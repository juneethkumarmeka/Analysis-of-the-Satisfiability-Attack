module basic_2500_25000_3000_50_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_1847,In_2270);
nand U1 (N_1,In_237,In_2403);
nand U2 (N_2,In_2098,In_1076);
and U3 (N_3,In_1670,In_83);
nor U4 (N_4,In_1703,In_2354);
nand U5 (N_5,In_1974,In_481);
or U6 (N_6,In_1660,In_1983);
and U7 (N_7,In_1508,In_1581);
nor U8 (N_8,In_2328,In_669);
nand U9 (N_9,In_912,In_2453);
nor U10 (N_10,In_2262,In_2035);
nor U11 (N_11,In_1385,In_545);
nor U12 (N_12,In_1635,In_255);
or U13 (N_13,In_247,In_324);
or U14 (N_14,In_1216,In_1415);
or U15 (N_15,In_777,In_102);
and U16 (N_16,In_2251,In_727);
nor U17 (N_17,In_1699,In_2303);
nand U18 (N_18,In_1715,In_2327);
nor U19 (N_19,In_1575,In_1356);
nand U20 (N_20,In_1763,In_1488);
nor U21 (N_21,In_1827,In_1350);
nor U22 (N_22,In_2061,In_2058);
nor U23 (N_23,In_2292,In_241);
and U24 (N_24,In_876,In_176);
and U25 (N_25,In_512,In_432);
nor U26 (N_26,In_128,In_2112);
nor U27 (N_27,In_1838,In_1769);
and U28 (N_28,In_2377,In_1275);
nand U29 (N_29,In_702,In_1897);
or U30 (N_30,In_736,In_1442);
and U31 (N_31,In_570,In_928);
or U32 (N_32,In_1549,In_1394);
and U33 (N_33,In_2359,In_1798);
and U34 (N_34,In_88,In_2461);
nand U35 (N_35,In_763,In_1485);
and U36 (N_36,In_1102,In_21);
nor U37 (N_37,In_349,In_1449);
nand U38 (N_38,In_323,In_1929);
nand U39 (N_39,In_1194,In_660);
nor U40 (N_40,In_1115,In_1105);
or U41 (N_41,In_1704,In_2466);
nor U42 (N_42,In_1396,In_1829);
nor U43 (N_43,In_231,In_528);
nand U44 (N_44,In_1122,In_1335);
nand U45 (N_45,In_1142,In_2233);
xnor U46 (N_46,In_869,In_2342);
xor U47 (N_47,In_801,In_540);
nor U48 (N_48,In_913,In_270);
and U49 (N_49,In_1724,In_534);
and U50 (N_50,In_41,In_1351);
or U51 (N_51,In_650,In_547);
nor U52 (N_52,In_1945,In_203);
or U53 (N_53,In_158,In_805);
nor U54 (N_54,In_2167,In_610);
nor U55 (N_55,In_2310,In_821);
nor U56 (N_56,In_1553,In_2029);
and U57 (N_57,In_1799,In_1792);
nand U58 (N_58,In_929,In_680);
and U59 (N_59,In_1578,In_2313);
xnor U60 (N_60,In_43,In_1013);
or U61 (N_61,In_963,In_2349);
or U62 (N_62,In_2030,In_2421);
nor U63 (N_63,In_1721,In_2041);
nand U64 (N_64,In_1251,In_1243);
and U65 (N_65,In_1873,In_1856);
and U66 (N_66,In_1674,In_403);
nor U67 (N_67,In_490,In_598);
nor U68 (N_68,In_542,In_1465);
or U69 (N_69,In_772,In_626);
nand U70 (N_70,In_2250,In_1949);
nand U71 (N_71,In_730,In_1622);
or U72 (N_72,In_1812,In_1828);
nand U73 (N_73,In_1035,In_1977);
or U74 (N_74,In_1229,In_1590);
or U75 (N_75,In_1080,In_877);
or U76 (N_76,In_1538,In_1679);
or U77 (N_77,In_1038,In_1073);
nand U78 (N_78,In_2192,In_134);
and U79 (N_79,In_68,In_1024);
nor U80 (N_80,In_1710,In_2415);
nand U81 (N_81,In_1061,In_180);
nand U82 (N_82,In_792,In_968);
and U83 (N_83,In_1678,In_2085);
nand U84 (N_84,In_605,In_604);
nor U85 (N_85,In_2200,In_1030);
and U86 (N_86,In_2395,In_58);
and U87 (N_87,In_1288,In_507);
or U88 (N_88,In_430,In_951);
or U89 (N_89,In_38,In_27);
and U90 (N_90,In_1614,In_165);
nand U91 (N_91,In_1492,In_249);
nor U92 (N_92,In_455,In_1595);
nand U93 (N_93,In_465,In_566);
nor U94 (N_94,In_1789,In_392);
xnor U95 (N_95,In_555,In_690);
and U96 (N_96,In_162,In_837);
and U97 (N_97,In_949,In_724);
and U98 (N_98,In_1259,In_1257);
or U99 (N_99,In_1777,In_1403);
or U100 (N_100,In_988,In_1392);
nor U101 (N_101,In_2459,In_1148);
nor U102 (N_102,In_1755,In_2215);
and U103 (N_103,In_750,In_1167);
nand U104 (N_104,In_1436,In_144);
or U105 (N_105,In_984,In_1957);
nand U106 (N_106,In_1365,In_1467);
nor U107 (N_107,In_1331,In_831);
nand U108 (N_108,In_1806,In_1540);
nor U109 (N_109,In_77,In_1564);
or U110 (N_110,In_674,In_862);
nand U111 (N_111,In_1069,In_819);
or U112 (N_112,In_2365,In_892);
nand U113 (N_113,In_227,In_256);
nand U114 (N_114,In_1489,In_1541);
xnor U115 (N_115,In_1127,In_1103);
or U116 (N_116,In_2477,In_1114);
nor U117 (N_117,In_338,In_2261);
xnor U118 (N_118,In_375,In_50);
and U119 (N_119,In_554,In_388);
nand U120 (N_120,In_520,In_1235);
or U121 (N_121,In_639,In_600);
nor U122 (N_122,In_1211,In_1072);
and U123 (N_123,In_1008,In_489);
and U124 (N_124,In_1079,In_1117);
and U125 (N_125,In_939,In_288);
nor U126 (N_126,In_1121,In_1547);
xor U127 (N_127,In_603,In_592);
nor U128 (N_128,In_720,In_2397);
nor U129 (N_129,In_1202,In_476);
or U130 (N_130,In_757,In_794);
nor U131 (N_131,In_1684,In_1800);
or U132 (N_132,In_1322,In_659);
and U133 (N_133,In_531,In_927);
or U134 (N_134,In_1656,In_836);
or U135 (N_135,In_1516,In_684);
xor U136 (N_136,In_2117,In_2394);
and U137 (N_137,In_2408,In_263);
nand U138 (N_138,In_78,In_1962);
or U139 (N_139,In_1807,In_1814);
nor U140 (N_140,In_1276,In_1645);
or U141 (N_141,In_596,In_1780);
and U142 (N_142,In_2267,In_411);
nor U143 (N_143,In_62,In_2148);
nand U144 (N_144,In_2027,In_133);
or U145 (N_145,In_2371,In_1874);
nor U146 (N_146,In_1401,In_1825);
xnor U147 (N_147,In_47,In_2175);
or U148 (N_148,In_1405,In_1757);
or U149 (N_149,In_1315,In_222);
nor U150 (N_150,In_1332,In_1817);
and U151 (N_151,In_1639,In_2176);
or U152 (N_152,In_1608,In_1661);
and U153 (N_153,In_441,In_1174);
and U154 (N_154,In_296,In_1867);
nand U155 (N_155,In_999,In_1698);
nand U156 (N_156,In_309,In_1846);
nand U157 (N_157,In_458,In_906);
or U158 (N_158,In_969,In_832);
nand U159 (N_159,In_56,In_1567);
nor U160 (N_160,In_1268,In_1004);
nand U161 (N_161,In_766,In_1985);
and U162 (N_162,In_808,In_1479);
nand U163 (N_163,In_2450,In_1176);
nor U164 (N_164,In_141,In_905);
nor U165 (N_165,In_1537,In_810);
nand U166 (N_166,In_632,In_813);
and U167 (N_167,In_1200,In_1425);
and U168 (N_168,In_223,In_1640);
and U169 (N_169,In_26,In_677);
nor U170 (N_170,In_30,In_2150);
and U171 (N_171,In_663,In_1033);
and U172 (N_172,In_2103,In_1533);
nand U173 (N_173,In_1697,In_1909);
nand U174 (N_174,In_1811,In_449);
nand U175 (N_175,In_491,In_494);
nand U176 (N_176,In_2014,In_2259);
nor U177 (N_177,In_2464,In_346);
or U178 (N_178,In_696,In_1470);
nand U179 (N_179,In_497,In_1961);
and U180 (N_180,In_2455,In_1976);
and U181 (N_181,In_1955,In_2384);
nor U182 (N_182,In_380,In_2067);
or U183 (N_183,In_967,In_602);
xnor U184 (N_184,In_53,In_2465);
and U185 (N_185,In_1217,In_1559);
nand U186 (N_186,In_2497,In_2146);
nand U187 (N_187,In_155,In_1823);
and U188 (N_188,In_437,In_1353);
nand U189 (N_189,In_1920,In_793);
or U190 (N_190,In_1053,In_880);
nand U191 (N_191,In_1071,In_1618);
nand U192 (N_192,In_1231,In_983);
or U193 (N_193,In_1098,In_1781);
or U194 (N_194,In_2158,In_893);
and U195 (N_195,In_1378,In_1190);
nand U196 (N_196,In_1839,In_820);
and U197 (N_197,In_2009,In_1313);
and U198 (N_198,In_482,In_1477);
nor U199 (N_199,In_1219,In_220);
or U200 (N_200,In_734,In_1865);
or U201 (N_201,In_814,In_2016);
or U202 (N_202,In_2232,In_2055);
or U203 (N_203,In_943,In_2319);
or U204 (N_204,In_302,In_2049);
or U205 (N_205,In_926,In_1292);
nor U206 (N_206,In_75,In_1001);
or U207 (N_207,In_2468,In_224);
or U208 (N_208,In_1334,In_2483);
nor U209 (N_209,In_888,In_151);
nand U210 (N_210,In_1233,In_1560);
or U211 (N_211,In_1527,In_2197);
nand U212 (N_212,In_958,In_1476);
or U213 (N_213,In_2171,In_806);
or U214 (N_214,In_1534,In_1308);
nand U215 (N_215,In_1499,In_1437);
or U216 (N_216,In_1579,In_2056);
nand U217 (N_217,In_1225,In_1768);
nand U218 (N_218,In_1066,In_2271);
xnor U219 (N_219,In_1043,In_633);
nand U220 (N_220,In_1017,In_1149);
and U221 (N_221,In_1990,In_167);
nor U222 (N_222,In_1152,In_1088);
nor U223 (N_223,In_258,In_1845);
nor U224 (N_224,In_889,In_1432);
and U225 (N_225,In_1742,In_1192);
nor U226 (N_226,In_2488,In_2025);
or U227 (N_227,In_2409,In_339);
or U228 (N_228,In_1993,In_1151);
and U229 (N_229,In_2454,In_890);
or U230 (N_230,In_101,In_285);
and U231 (N_231,In_901,In_828);
or U232 (N_232,In_1783,In_1862);
or U233 (N_233,In_1478,In_732);
and U234 (N_234,In_1486,In_93);
nand U235 (N_235,In_955,In_770);
nand U236 (N_236,In_2162,In_667);
xor U237 (N_237,In_1086,In_2333);
nand U238 (N_238,In_1170,In_817);
nor U239 (N_239,In_2368,In_1669);
or U240 (N_240,In_1959,In_401);
nand U241 (N_241,In_185,In_259);
nand U242 (N_242,In_2248,In_1878);
nor U243 (N_243,In_681,In_409);
or U244 (N_244,In_2063,In_1070);
or U245 (N_245,In_2425,In_737);
nor U246 (N_246,In_1228,In_1074);
xnor U247 (N_247,In_1852,In_662);
and U248 (N_248,In_530,In_846);
nand U249 (N_249,In_290,In_2194);
nand U250 (N_250,In_1239,In_1938);
and U251 (N_251,In_1441,In_1028);
nand U252 (N_252,In_1561,In_516);
and U253 (N_253,In_2124,In_1713);
nand U254 (N_254,In_1089,In_651);
and U255 (N_255,In_2140,In_1542);
and U256 (N_256,In_648,In_729);
or U257 (N_257,In_747,In_2152);
and U258 (N_258,In_1111,In_1397);
nor U259 (N_259,In_1842,In_2339);
nor U260 (N_260,In_1007,In_1469);
xnor U261 (N_261,In_1809,In_504);
nand U262 (N_262,In_2300,In_1002);
or U263 (N_263,In_2279,In_1455);
nand U264 (N_264,In_786,In_2411);
or U265 (N_265,In_18,In_138);
and U266 (N_266,In_2420,In_148);
and U267 (N_267,In_584,In_1501);
nor U268 (N_268,In_887,In_1997);
nand U269 (N_269,In_1637,In_2100);
nor U270 (N_270,In_2019,In_1594);
or U271 (N_271,In_2451,In_629);
xnor U272 (N_272,In_1910,In_1585);
nor U273 (N_273,In_2093,In_634);
and U274 (N_274,In_535,In_216);
or U275 (N_275,In_1487,In_576);
or U276 (N_276,In_433,In_553);
or U277 (N_277,In_904,In_1453);
and U278 (N_278,In_803,In_1510);
or U279 (N_279,In_2350,In_2096);
and U280 (N_280,In_936,In_2379);
nand U281 (N_281,In_587,In_331);
nor U282 (N_282,In_874,In_2037);
or U283 (N_283,In_400,In_1440);
and U284 (N_284,In_845,In_1868);
or U285 (N_285,In_2326,In_1081);
and U286 (N_286,In_95,In_1643);
and U287 (N_287,In_1328,In_2428);
nand U288 (N_288,In_1870,In_37);
nor U289 (N_289,In_2367,In_589);
or U290 (N_290,In_280,In_2137);
and U291 (N_291,In_1996,In_1876);
or U292 (N_292,In_1626,In_1324);
and U293 (N_293,In_475,In_563);
or U294 (N_294,In_1741,In_1031);
nor U295 (N_295,In_1925,In_1147);
nand U296 (N_296,In_1659,In_957);
and U297 (N_297,In_1109,In_2498);
or U298 (N_298,In_1050,In_1048);
nor U299 (N_299,In_881,In_1143);
nand U300 (N_300,In_1894,In_1490);
and U301 (N_301,In_2046,In_982);
and U302 (N_302,In_1671,In_1438);
nand U303 (N_303,In_1820,In_654);
nor U304 (N_304,In_24,In_1778);
or U305 (N_305,In_1141,In_1208);
nand U306 (N_306,In_172,In_1186);
nand U307 (N_307,In_454,In_485);
and U308 (N_308,In_1482,In_416);
nor U309 (N_309,In_170,In_2164);
and U310 (N_310,In_848,In_2213);
or U311 (N_311,In_562,In_2207);
nand U312 (N_312,In_1091,In_1927);
nor U313 (N_313,In_1067,In_1720);
or U314 (N_314,In_1238,In_2163);
and U315 (N_315,In_1956,In_80);
nand U316 (N_316,In_1157,In_1413);
nand U317 (N_317,In_2130,In_1722);
nor U318 (N_318,In_2238,In_1706);
xor U319 (N_319,In_518,In_627);
or U320 (N_320,In_410,In_1278);
nand U321 (N_321,In_2105,In_208);
or U322 (N_322,In_759,In_1859);
and U323 (N_323,In_2437,In_1832);
or U324 (N_324,In_1294,In_1646);
nor U325 (N_325,In_1756,In_97);
and U326 (N_326,In_1374,In_658);
nor U327 (N_327,In_2075,In_2043);
and U328 (N_328,In_179,In_2400);
nor U329 (N_329,In_2195,In_1253);
or U330 (N_330,In_1402,In_394);
and U331 (N_331,In_2011,In_1523);
or U332 (N_332,In_567,In_744);
nand U333 (N_333,In_436,In_1446);
nand U334 (N_334,In_2346,In_2042);
nor U335 (N_335,In_621,In_2434);
or U336 (N_336,In_2072,In_1279);
nor U337 (N_337,In_146,In_865);
and U338 (N_338,In_443,In_2241);
xnor U339 (N_339,In_2389,In_195);
nor U340 (N_340,In_29,In_2416);
xor U341 (N_341,In_108,In_71);
and U342 (N_342,In_1325,In_1901);
and U343 (N_343,In_2118,In_1759);
and U344 (N_344,In_98,In_201);
xor U345 (N_345,In_1796,In_70);
or U346 (N_346,In_265,In_593);
nor U347 (N_347,In_442,In_775);
and U348 (N_348,In_306,In_1039);
or U349 (N_349,In_1649,In_45);
nor U350 (N_350,In_468,In_1249);
nand U351 (N_351,In_63,In_2114);
or U352 (N_352,In_978,In_1158);
nor U353 (N_353,In_2495,In_384);
nand U354 (N_354,In_2357,In_966);
nand U355 (N_355,In_244,In_479);
nand U356 (N_356,In_2217,In_2083);
and U357 (N_357,In_767,In_184);
or U358 (N_358,In_735,In_1263);
nor U359 (N_359,In_48,In_1711);
or U360 (N_360,In_708,In_1299);
or U361 (N_361,In_1786,In_1558);
nor U362 (N_362,In_670,In_1339);
and U363 (N_363,In_2372,In_1444);
nand U364 (N_364,In_1199,In_515);
nand U365 (N_365,In_1171,In_412);
and U366 (N_366,In_1666,In_1361);
and U367 (N_367,In_645,In_875);
and U368 (N_368,In_1970,In_1252);
xor U369 (N_369,In_261,In_1146);
xnor U370 (N_370,In_2484,In_342);
nand U371 (N_371,In_87,In_156);
and U372 (N_372,In_334,In_2249);
nand U373 (N_373,In_1928,In_2191);
and U374 (N_374,In_352,In_234);
and U375 (N_375,In_120,In_2038);
or U376 (N_376,In_2022,In_1260);
nor U377 (N_377,In_1311,In_2006);
nor U378 (N_378,In_2291,In_390);
nand U379 (N_379,In_1400,In_1014);
and U380 (N_380,In_52,In_1978);
nand U381 (N_381,In_376,In_495);
and U382 (N_382,In_942,In_1960);
nand U383 (N_383,In_572,In_1518);
and U384 (N_384,In_34,In_478);
and U385 (N_385,In_675,In_1277);
nor U386 (N_386,In_370,In_1391);
and U387 (N_387,In_1304,In_2479);
nor U388 (N_388,In_1921,In_260);
and U389 (N_389,In_1907,In_1379);
or U390 (N_390,In_1557,In_1083);
nand U391 (N_391,In_106,In_886);
or U392 (N_392,In_991,In_2369);
and U393 (N_393,In_698,In_513);
nor U394 (N_394,In_90,In_1265);
or U395 (N_395,In_834,In_1535);
nand U396 (N_396,In_2401,In_818);
or U397 (N_397,In_2222,In_96);
or U398 (N_398,In_2321,In_1348);
or U399 (N_399,In_1886,In_1373);
nor U400 (N_400,In_1586,In_896);
and U401 (N_401,In_2390,In_419);
and U402 (N_402,In_868,In_2050);
or U403 (N_403,In_160,In_1389);
and U404 (N_404,In_2048,In_2269);
nor U405 (N_405,In_318,In_1184);
xor U406 (N_406,In_2094,In_2343);
xnor U407 (N_407,In_2265,In_312);
and U408 (N_408,In_861,In_2306);
or U409 (N_409,In_2398,In_1860);
or U410 (N_410,In_1676,In_1020);
nand U411 (N_411,In_1562,In_1879);
nand U412 (N_412,In_683,In_2101);
nor U413 (N_413,In_2051,In_413);
or U414 (N_414,In_1866,In_1688);
xnor U415 (N_415,In_1150,In_125);
nor U416 (N_416,In_1341,In_425);
or U417 (N_417,In_2255,In_225);
or U418 (N_418,In_283,In_788);
nor U419 (N_419,In_2438,In_161);
nand U420 (N_420,In_1367,In_699);
or U421 (N_421,In_1046,In_337);
nand U422 (N_422,In_2104,In_573);
and U423 (N_423,In_186,In_8);
nor U424 (N_424,In_1505,In_965);
nand U425 (N_425,In_439,In_758);
or U426 (N_426,In_1283,In_505);
or U427 (N_427,In_1887,In_1854);
nand U428 (N_428,In_2208,In_1108);
and U429 (N_429,In_712,In_2024);
and U430 (N_430,In_2108,In_1314);
and U431 (N_431,In_2302,In_492);
or U432 (N_432,In_776,In_835);
or U433 (N_433,In_560,In_1320);
nor U434 (N_434,In_311,In_1995);
or U435 (N_435,In_930,In_1398);
nand U436 (N_436,In_1498,In_2080);
nand U437 (N_437,In_107,In_840);
or U438 (N_438,In_2165,In_1693);
or U439 (N_439,In_1497,In_1185);
or U440 (N_440,In_2065,In_393);
nand U441 (N_441,In_2351,In_54);
and U442 (N_442,In_2402,In_333);
nor U443 (N_443,In_916,In_785);
and U444 (N_444,In_1620,In_1407);
and U445 (N_445,In_640,In_1681);
nand U446 (N_446,In_1802,In_1875);
or U447 (N_447,In_1291,In_1863);
nor U448 (N_448,In_1363,In_2166);
and U449 (N_449,In_453,In_2141);
or U450 (N_450,In_682,In_1125);
or U451 (N_451,In_2180,In_202);
or U452 (N_452,In_2422,In_351);
nand U453 (N_453,In_1045,In_543);
nand U454 (N_454,In_1946,In_1937);
and U455 (N_455,In_1491,In_2186);
or U456 (N_456,In_756,In_2337);
or U457 (N_457,In_1386,In_289);
xnor U458 (N_458,In_842,In_2266);
nand U459 (N_459,In_1691,In_2462);
nand U460 (N_460,In_365,In_517);
nand U461 (N_461,In_477,In_1484);
or U462 (N_462,In_1346,In_1329);
nor U463 (N_463,In_652,In_2135);
or U464 (N_464,In_60,In_1382);
and U465 (N_465,In_1164,In_40);
or U466 (N_466,In_565,In_625);
and U467 (N_467,In_1451,In_878);
nor U468 (N_468,In_1716,In_995);
nand U469 (N_469,In_1853,In_1627);
nand U470 (N_470,In_1986,In_1850);
and U471 (N_471,In_581,In_1175);
nor U472 (N_472,In_754,In_694);
or U473 (N_473,In_1040,In_1589);
nand U474 (N_474,In_1383,In_379);
or U475 (N_475,In_150,In_973);
or U476 (N_476,In_1784,In_812);
and U477 (N_477,In_85,In_2224);
nor U478 (N_478,In_666,In_2309);
and U479 (N_479,In_1326,In_1359);
nor U480 (N_480,In_2287,In_2297);
nor U481 (N_481,In_464,In_358);
and U482 (N_482,In_796,In_232);
nor U483 (N_483,In_686,In_1153);
and U484 (N_484,In_1087,In_1226);
or U485 (N_485,In_1668,In_807);
and U486 (N_486,In_1926,In_1187);
or U487 (N_487,In_175,In_304);
nor U488 (N_488,In_2414,In_200);
nor U489 (N_489,In_2318,In_325);
and U490 (N_490,In_1841,In_2023);
nand U491 (N_491,In_414,In_386);
nor U492 (N_492,In_250,In_743);
xor U493 (N_493,In_137,In_366);
or U494 (N_494,In_544,In_2332);
and U495 (N_495,In_779,In_2154);
xor U496 (N_496,In_1390,In_924);
nor U497 (N_497,In_1908,In_2078);
and U498 (N_498,In_166,In_1301);
nor U499 (N_499,In_76,In_2473);
and U500 (N_500,In_1023,In_2054);
or U501 (N_501,In_2044,N_269);
and U502 (N_502,In_32,In_2235);
xor U503 (N_503,In_2476,In_2139);
nand U504 (N_504,In_230,In_499);
nor U505 (N_505,In_327,In_2364);
nor U506 (N_506,In_2387,N_385);
nand U507 (N_507,In_804,In_1729);
nand U508 (N_508,N_213,In_211);
or U509 (N_509,N_196,N_251);
nand U510 (N_510,In_362,In_1520);
nand U511 (N_511,In_122,In_1592);
and U512 (N_512,In_2095,In_1064);
nor U513 (N_513,In_1290,In_2244);
nor U514 (N_514,In_268,In_2123);
and U515 (N_515,In_1059,In_2034);
or U516 (N_516,In_1922,In_1431);
nand U517 (N_517,N_7,N_266);
nand U518 (N_518,In_1135,In_1551);
nand U519 (N_519,In_700,In_2489);
nor U520 (N_520,N_43,In_1241);
and U521 (N_521,In_2375,In_614);
or U522 (N_522,In_305,In_2258);
and U523 (N_523,N_114,In_1269);
nor U524 (N_524,In_140,In_2405);
and U525 (N_525,In_2443,In_447);
and U526 (N_526,In_508,In_564);
nand U527 (N_527,N_227,In_833);
and U528 (N_528,In_858,N_300);
or U529 (N_529,In_456,In_1447);
nor U530 (N_530,In_980,N_499);
or U531 (N_531,N_231,In_1599);
nor U532 (N_532,In_117,In_2373);
and U533 (N_533,In_2340,In_2362);
and U534 (N_534,In_2155,In_1584);
nand U535 (N_535,In_1424,In_606);
nor U536 (N_536,In_500,In_187);
nor U537 (N_537,In_1026,In_1546);
and U538 (N_538,In_799,In_1761);
nor U539 (N_539,In_1813,In_1333);
nor U540 (N_540,In_1987,In_1966);
nor U541 (N_541,In_2491,In_1507);
or U542 (N_542,In_1460,In_509);
or U543 (N_543,In_1848,In_194);
and U544 (N_544,N_157,In_1858);
nand U545 (N_545,N_279,In_1494);
or U546 (N_546,N_482,In_826);
nor U547 (N_547,In_1988,In_1169);
and U548 (N_548,In_1298,In_1466);
and U549 (N_549,In_322,N_160);
nand U550 (N_550,In_977,In_2092);
or U551 (N_551,In_1924,In_89);
nor U552 (N_552,N_415,In_2177);
and U553 (N_553,In_1735,N_445);
and U554 (N_554,N_229,N_220);
nand U555 (N_555,N_424,N_302);
and U556 (N_556,N_26,In_790);
nor U557 (N_557,N_430,In_1734);
and U558 (N_558,In_769,N_249);
and U559 (N_559,N_493,In_1804);
or U560 (N_560,In_314,N_308);
and U561 (N_561,In_64,N_475);
or U562 (N_562,In_1738,In_1803);
nand U563 (N_563,In_2151,In_502);
and U564 (N_564,N_236,In_1791);
nor U565 (N_565,In_609,In_641);
and U566 (N_566,In_1022,In_1203);
and U567 (N_567,N_417,In_1287);
nor U568 (N_568,In_703,In_242);
nor U569 (N_569,In_1285,In_214);
xnor U570 (N_570,N_167,In_2008);
xor U571 (N_571,In_1439,N_234);
nand U572 (N_572,In_2018,In_463);
or U573 (N_573,N_473,In_1967);
nand U574 (N_574,In_1450,In_1282);
nand U575 (N_575,In_1113,In_157);
or U576 (N_576,In_1651,N_15);
nor U577 (N_577,N_88,In_1923);
or U578 (N_578,In_11,In_1000);
nand U579 (N_579,In_985,In_1036);
nor U580 (N_580,In_152,In_2047);
nand U581 (N_581,N_28,In_1418);
nor U582 (N_582,In_1819,In_1623);
and U583 (N_583,In_1018,In_191);
nor U584 (N_584,In_1736,N_70);
or U585 (N_585,N_248,In_922);
and U586 (N_586,In_340,N_54);
nor U587 (N_587,In_2231,In_335);
nand U588 (N_588,In_1349,In_590);
and U589 (N_589,N_259,In_2316);
nand U590 (N_590,In_1345,In_1273);
nand U591 (N_591,N_402,In_2431);
or U592 (N_592,N_384,In_2335);
nand U593 (N_593,N_450,N_342);
or U594 (N_594,In_1245,N_211);
and U595 (N_595,In_1588,In_2385);
xnor U596 (N_596,In_1834,N_389);
nand U597 (N_597,N_89,In_2345);
xor U598 (N_598,In_1213,N_148);
or U599 (N_599,In_431,N_138);
and U600 (N_600,N_357,In_278);
nor U601 (N_601,N_334,In_1221);
nor U602 (N_602,In_209,In_2234);
nand U603 (N_603,In_310,In_168);
and U604 (N_604,In_1015,In_326);
or U605 (N_605,N_490,In_1610);
or U606 (N_606,In_291,In_1471);
and U607 (N_607,In_1795,In_519);
or U608 (N_608,In_987,N_103);
nand U609 (N_609,N_288,In_1884);
or U610 (N_610,In_420,In_356);
or U611 (N_611,In_2138,In_1687);
and U612 (N_612,In_1468,In_1607);
or U613 (N_613,N_47,In_2156);
xor U614 (N_614,N_86,N_137);
nor U615 (N_615,In_183,N_143);
or U616 (N_616,In_1779,In_2446);
or U617 (N_617,In_1893,In_1227);
or U618 (N_618,In_2087,N_496);
nor U619 (N_619,In_961,In_435);
and U620 (N_620,In_1566,In_1888);
and U621 (N_621,In_1034,In_1864);
nand U622 (N_622,In_297,N_412);
or U623 (N_623,In_2144,N_378);
nand U624 (N_624,In_460,In_791);
or U625 (N_625,In_1935,N_49);
nand U626 (N_626,N_142,N_149);
or U627 (N_627,In_1092,In_1971);
and U628 (N_628,N_360,N_439);
and U629 (N_629,In_1555,In_328);
and U630 (N_630,In_2315,In_1675);
or U631 (N_631,In_1357,In_169);
nand U632 (N_632,In_2226,N_113);
nor U633 (N_633,In_271,N_171);
nor U634 (N_634,In_2301,In_1272);
nor U635 (N_635,N_257,In_2264);
or U636 (N_636,N_469,In_2374);
nor U637 (N_637,In_1406,In_2040);
or U638 (N_638,In_1565,In_219);
and U639 (N_639,N_313,In_1075);
xnor U640 (N_640,In_132,In_2472);
nor U641 (N_641,In_1376,In_923);
or U642 (N_642,In_784,In_882);
and U643 (N_643,N_147,N_75);
or U644 (N_644,In_533,In_1347);
nor U645 (N_645,In_1760,N_364);
or U646 (N_646,In_1496,In_2240);
nand U647 (N_647,In_1154,N_477);
nand U648 (N_648,In_721,In_1041);
and U649 (N_649,In_1270,In_1118);
or U650 (N_650,N_201,In_2329);
or U651 (N_651,In_124,In_1165);
and U652 (N_652,In_2071,N_173);
and U653 (N_653,In_613,N_436);
and U654 (N_654,In_171,In_1178);
nor U655 (N_655,In_72,In_707);
nand U656 (N_656,In_548,In_918);
nor U657 (N_657,N_193,N_395);
nor U658 (N_658,In_778,In_240);
nand U659 (N_659,In_1414,In_126);
nor U660 (N_660,N_440,In_899);
nand U661 (N_661,In_2228,In_1749);
nor U662 (N_662,In_1723,In_856);
or U663 (N_663,In_938,N_341);
nand U664 (N_664,In_1751,N_352);
nor U665 (N_665,In_1016,In_816);
xor U666 (N_666,In_264,In_2074);
or U667 (N_667,In_2366,In_1427);
or U668 (N_668,In_1330,In_1483);
and U669 (N_669,N_472,In_2452);
nand U670 (N_670,In_361,In_1826);
or U671 (N_671,In_701,N_354);
and U672 (N_672,In_28,N_125);
or U673 (N_673,N_416,In_2330);
nor U674 (N_674,In_1419,In_2485);
nand U675 (N_675,In_823,In_1172);
and U676 (N_676,In_2143,In_374);
nand U677 (N_677,N_126,N_467);
or U678 (N_678,N_146,In_1448);
nor U679 (N_679,N_197,In_1209);
or U680 (N_680,N_9,In_1388);
and U681 (N_681,In_921,In_1010);
nand U682 (N_682,In_1300,In_452);
nor U683 (N_683,In_1654,In_536);
or U684 (N_684,N_400,In_1625);
or U685 (N_685,N_221,In_695);
nand U686 (N_686,In_1522,In_205);
or U687 (N_687,In_44,In_1773);
nor U688 (N_688,In_2353,In_549);
nor U689 (N_689,In_1430,In_1650);
or U690 (N_690,In_2021,In_1719);
and U691 (N_691,In_1918,In_13);
xnor U692 (N_692,In_2142,N_144);
nor U693 (N_693,In_193,In_1412);
nor U694 (N_694,In_2089,N_83);
or U695 (N_695,In_0,N_30);
or U696 (N_696,In_900,In_1600);
nor U697 (N_697,N_176,N_332);
and U698 (N_698,In_809,In_599);
nand U699 (N_699,In_1702,In_749);
xor U700 (N_700,N_289,In_920);
nor U701 (N_701,In_867,In_438);
nand U702 (N_702,In_395,In_321);
nand U703 (N_703,In_2336,In_1094);
or U704 (N_704,In_493,In_2188);
or U705 (N_705,N_277,In_2407);
nand U706 (N_706,N_40,N_284);
nand U707 (N_707,In_2017,In_1503);
nand U708 (N_708,In_1543,N_299);
xnor U709 (N_709,In_1362,In_446);
nand U710 (N_710,In_733,In_113);
and U711 (N_711,In_1641,In_1824);
nor U712 (N_712,In_704,In_2086);
and U713 (N_713,N_317,In_539);
and U714 (N_714,N_460,In_2122);
nand U715 (N_715,In_1009,In_1242);
xnor U716 (N_716,In_1234,In_990);
nand U717 (N_717,In_1936,In_1998);
nor U718 (N_718,N_61,In_267);
and U719 (N_719,In_1753,In_2132);
nor U720 (N_720,N_438,In_1552);
nor U721 (N_721,In_765,In_1131);
and U722 (N_722,In_1583,N_242);
or U723 (N_723,In_871,In_872);
nand U724 (N_724,In_1504,In_2381);
nor U725 (N_725,N_60,In_841);
or U726 (N_726,In_1521,In_65);
and U727 (N_727,N_199,In_2439);
nor U728 (N_728,N_152,In_1342);
nor U729 (N_729,N_140,In_2284);
and U730 (N_730,N_457,N_177);
xnor U731 (N_731,In_636,N_254);
nor U732 (N_732,In_1730,N_79);
nor U733 (N_733,N_85,In_369);
xnor U734 (N_734,In_1062,N_121);
nor U735 (N_735,In_653,In_1601);
nor U736 (N_736,In_1569,In_474);
and U737 (N_737,In_915,N_208);
and U738 (N_738,In_514,In_1754);
and U739 (N_739,N_263,N_293);
or U740 (N_740,In_1980,In_1302);
nor U741 (N_741,In_1609,In_1340);
nand U742 (N_742,In_2290,In_1810);
nor U743 (N_743,In_2356,In_20);
or U744 (N_744,N_480,In_2392);
and U745 (N_745,In_1343,In_885);
nand U746 (N_746,In_276,N_492);
xor U747 (N_747,In_960,In_1463);
and U748 (N_748,In_1254,In_970);
and U749 (N_749,In_266,N_68);
nand U750 (N_750,In_81,N_390);
and U751 (N_751,N_362,N_403);
nand U752 (N_752,N_135,In_692);
nor U753 (N_753,In_484,In_2091);
nand U754 (N_754,In_1836,In_9);
and U755 (N_755,In_307,In_6);
nand U756 (N_756,In_739,In_486);
nor U757 (N_757,In_1354,N_96);
nand U758 (N_758,In_189,In_940);
or U759 (N_759,N_324,In_277);
or U760 (N_760,In_693,N_38);
nand U761 (N_761,N_14,In_714);
and U762 (N_762,In_1456,In_1078);
nor U763 (N_763,N_228,N_434);
and U764 (N_764,N_320,N_11);
and U765 (N_765,N_27,In_1642);
and U766 (N_766,In_2115,In_1709);
nor U767 (N_767,In_2432,In_691);
or U768 (N_768,In_2404,In_2129);
and U769 (N_769,In_1963,N_290);
nand U770 (N_770,In_199,N_178);
or U771 (N_771,N_1,N_192);
and U772 (N_772,In_2341,In_1964);
and U773 (N_773,In_1502,In_1305);
xor U774 (N_774,In_127,In_1410);
nor U775 (N_775,In_181,In_100);
or U776 (N_776,N_141,In_142);
xnor U777 (N_777,In_1653,N_419);
or U778 (N_778,In_470,In_1232);
nor U779 (N_779,In_1506,N_452);
nand U780 (N_780,In_57,In_1110);
or U781 (N_781,In_1903,In_1539);
or U782 (N_782,In_546,In_198);
nor U783 (N_783,In_2274,In_1054);
nand U784 (N_784,In_672,In_1128);
or U785 (N_785,N_94,In_1481);
xnor U786 (N_786,N_174,In_552);
and U787 (N_787,N_287,In_1612);
nor U788 (N_788,N_198,In_16);
nand U789 (N_789,In_273,In_948);
or U790 (N_790,N_92,N_58);
nor U791 (N_791,In_2257,In_355);
nand U792 (N_792,In_2070,In_173);
nor U793 (N_793,In_619,In_2220);
nor U794 (N_794,In_2444,In_1587);
nor U795 (N_795,In_1892,In_104);
and U796 (N_796,In_601,N_405);
or U797 (N_797,In_2467,N_350);
nand U798 (N_798,In_1683,N_478);
nand U799 (N_799,N_65,N_51);
nand U800 (N_800,In_2172,N_431);
nor U801 (N_801,In_2097,In_2120);
or U802 (N_802,In_92,In_396);
or U803 (N_803,In_1648,N_91);
nand U804 (N_804,N_207,N_19);
or U805 (N_805,In_1286,In_94);
or U806 (N_806,In_709,In_950);
nor U807 (N_807,N_312,In_2322);
nand U808 (N_808,In_1370,In_1740);
nor U809 (N_809,In_1421,In_1246);
and U810 (N_810,In_2174,In_1220);
nor U811 (N_811,In_33,In_1882);
or U812 (N_812,In_2221,In_706);
nor U813 (N_813,N_333,N_309);
or U814 (N_814,In_2225,In_1794);
or U815 (N_815,In_2268,N_463);
nand U816 (N_816,In_2079,N_338);
nor U817 (N_817,In_1531,N_261);
and U818 (N_818,In_2280,In_2410);
and U819 (N_819,N_245,In_385);
nand U820 (N_820,In_2486,In_1458);
nor U821 (N_821,In_1306,In_1605);
nor U822 (N_822,In_697,In_1849);
nor U823 (N_823,In_2157,In_1568);
nand U824 (N_824,N_194,In_2482);
or U825 (N_825,In_1764,In_450);
nor U826 (N_826,In_2160,In_301);
or U827 (N_827,In_558,N_344);
nor U828 (N_828,In_2278,In_1205);
nand U829 (N_829,In_1423,N_210);
xnor U830 (N_830,In_66,N_448);
nand U831 (N_831,In_2441,In_415);
and U832 (N_832,In_483,In_1638);
nor U833 (N_833,N_441,In_192);
nor U834 (N_834,N_73,In_1902);
or U835 (N_835,In_86,In_1417);
nand U836 (N_836,In_998,In_2281);
nor U837 (N_837,In_239,In_1725);
or U838 (N_838,N_163,In_2320);
nand U839 (N_839,In_1309,N_13);
nand U840 (N_840,In_212,N_315);
or U841 (N_841,In_1155,In_1454);
or U842 (N_842,In_2187,In_2153);
nor U843 (N_843,In_506,In_760);
nand U844 (N_844,In_1631,N_374);
nor U845 (N_845,N_124,In_1120);
nand U846 (N_846,In_2149,In_233);
or U847 (N_847,In_944,In_206);
and U848 (N_848,In_798,In_422);
nand U849 (N_849,In_2253,In_1563);
nand U850 (N_850,N_404,In_1785);
or U851 (N_851,In_153,In_1019);
or U852 (N_852,In_2109,N_348);
nor U853 (N_853,N_87,In_1106);
or U854 (N_854,N_329,In_1571);
and U855 (N_855,In_2286,N_33);
nor U856 (N_856,N_339,In_467);
or U857 (N_857,In_1593,In_408);
nand U858 (N_858,In_1011,In_668);
and U859 (N_859,In_119,In_1914);
nand U860 (N_860,In_139,In_661);
and U861 (N_861,N_435,In_1732);
xor U862 (N_862,In_624,In_1621);
and U863 (N_863,In_647,In_1616);
or U864 (N_864,In_1124,In_1191);
and U865 (N_865,In_406,In_2325);
and U866 (N_866,N_406,In_2338);
nor U867 (N_867,In_2386,N_123);
nand U868 (N_868,In_1934,N_184);
nand U869 (N_869,N_16,In_1821);
and U870 (N_870,In_1319,N_273);
nand U871 (N_871,In_1044,In_1689);
nand U872 (N_872,In_1274,N_285);
nor U873 (N_873,In_1765,N_485);
nor U874 (N_874,N_264,N_410);
or U875 (N_875,In_551,In_615);
nor U876 (N_876,N_372,In_857);
nor U877 (N_877,In_1060,In_1095);
nand U878 (N_878,In_1129,N_379);
and U879 (N_879,In_2412,In_382);
nor U880 (N_880,N_235,N_498);
and U881 (N_881,In_1360,In_716);
and U882 (N_882,In_299,N_465);
nand U883 (N_883,In_320,In_359);
and U884 (N_884,In_989,N_336);
and U885 (N_885,N_270,In_398);
or U886 (N_886,In_2113,In_236);
and U887 (N_887,In_1281,In_2277);
and U888 (N_888,In_2426,In_783);
and U889 (N_889,In_1215,N_53);
or U890 (N_890,N_116,In_262);
nand U891 (N_891,N_34,In_631);
and U892 (N_892,In_1179,In_2116);
nor U893 (N_893,In_1947,In_1883);
nand U894 (N_894,In_974,In_444);
nand U895 (N_895,N_247,In_1805);
nand U896 (N_896,In_860,N_337);
and U897 (N_897,In_1162,In_2159);
or U898 (N_898,In_1495,In_1989);
or U899 (N_899,N_456,N_319);
or U900 (N_900,In_2133,N_298);
nand U901 (N_901,In_1885,In_751);
nand U902 (N_902,In_103,In_740);
or U903 (N_903,In_843,In_1707);
nor U904 (N_904,In_722,In_738);
and U905 (N_905,In_360,N_459);
nand U906 (N_906,In_1197,N_189);
or U907 (N_907,In_1958,In_1634);
and U908 (N_908,N_226,In_1112);
nor U909 (N_909,N_139,In_1933);
nor U910 (N_910,In_1991,N_134);
nand U911 (N_911,N_275,In_1230);
nand U912 (N_912,In_145,In_1530);
nor U913 (N_913,In_891,In_1201);
and U914 (N_914,In_1377,In_2026);
or U915 (N_915,In_330,N_326);
and U916 (N_916,N_380,In_2068);
and U917 (N_917,In_2201,N_310);
or U918 (N_918,In_315,In_79);
nand U919 (N_919,In_909,In_679);
nor U920 (N_920,In_2299,N_470);
or U921 (N_921,N_218,In_336);
and U922 (N_922,N_427,In_731);
and U923 (N_923,In_2039,In_67);
and U924 (N_924,N_161,In_2456);
nor U925 (N_925,In_1090,In_2214);
or U926 (N_926,In_797,In_226);
nand U927 (N_927,N_396,In_423);
nand U928 (N_928,In_1183,In_782);
and U929 (N_929,In_1166,In_367);
or U930 (N_930,In_2481,In_424);
xor U931 (N_931,In_1029,In_1652);
or U932 (N_932,In_561,In_997);
nand U933 (N_933,In_591,In_1207);
or U934 (N_934,In_2406,In_1144);
nor U935 (N_935,In_1130,In_1435);
and U936 (N_936,N_117,In_1323);
and U937 (N_937,In_685,In_723);
or U938 (N_938,In_1705,In_2003);
nor U939 (N_939,In_2119,In_109);
and U940 (N_940,In_221,N_330);
nor U941 (N_941,In_1528,In_884);
nor U942 (N_942,In_91,In_69);
and U943 (N_943,N_45,N_433);
and U944 (N_944,In_188,In_1084);
and U945 (N_945,N_346,N_115);
and U946 (N_946,In_404,In_1603);
or U947 (N_947,N_278,In_1312);
and U948 (N_948,In_1411,N_486);
and U949 (N_949,N_215,In_2427);
nand U950 (N_950,In_855,In_2440);
and U951 (N_951,N_62,In_2032);
or U952 (N_952,In_417,In_1667);
nand U953 (N_953,In_2435,N_258);
or U954 (N_954,In_1250,N_345);
xnor U955 (N_955,In_2358,In_1051);
and U956 (N_956,In_1745,In_996);
nor U957 (N_957,In_741,In_2436);
nand U958 (N_958,In_1880,In_2183);
nand U959 (N_959,In_387,In_1942);
nand U960 (N_960,In_469,In_1948);
nor U961 (N_961,In_1517,In_2288);
nand U962 (N_962,N_195,In_2391);
and U963 (N_963,In_1840,N_119);
xnor U964 (N_964,In_1180,In_673);
nand U965 (N_965,N_271,In_897);
xnor U966 (N_966,In_718,N_484);
nand U967 (N_967,In_1965,In_2475);
nor U968 (N_968,In_1597,In_1012);
or U969 (N_969,In_2193,In_350);
and U970 (N_970,In_204,In_1236);
and U971 (N_971,In_538,N_214);
and U972 (N_972,In_580,N_291);
and U973 (N_973,In_863,N_373);
or U974 (N_974,In_254,In_300);
and U975 (N_975,In_2145,In_1057);
and U976 (N_976,In_762,In_628);
or U977 (N_977,N_358,In_1161);
and U978 (N_978,N_295,In_2308);
nor U979 (N_979,In_956,In_182);
or U980 (N_980,In_1525,In_2102);
nor U981 (N_981,N_181,In_2246);
or U982 (N_982,In_1911,In_1871);
nor U983 (N_983,N_187,N_488);
xor U984 (N_984,In_2413,In_597);
nor U985 (N_985,In_1744,In_112);
nand U986 (N_986,In_665,N_268);
and U987 (N_987,In_937,In_1472);
nor U988 (N_988,N_347,In_229);
nor U989 (N_989,N_164,In_2393);
or U990 (N_990,In_1628,In_1896);
or U991 (N_991,In_2305,In_1338);
nand U992 (N_992,In_1979,In_523);
nor U993 (N_993,N_386,In_163);
nand U994 (N_994,N_10,In_1371);
nor U995 (N_995,N_200,In_1818);
nor U996 (N_996,N_233,In_105);
nor U997 (N_997,In_1515,N_35);
xor U998 (N_998,In_2430,In_248);
and U999 (N_999,In_2490,In_49);
or U1000 (N_1000,N_753,In_678);
and U1001 (N_1001,In_1404,In_1284);
and U1002 (N_1002,In_620,In_2347);
and U1003 (N_1003,In_159,In_2239);
nand U1004 (N_1004,In_1047,N_687);
or U1005 (N_1005,N_937,In_2282);
nor U1006 (N_1006,N_5,N_230);
or U1007 (N_1007,N_801,N_425);
nand U1008 (N_1008,In_2045,In_2227);
nor U1009 (N_1009,N_694,In_859);
nand U1010 (N_1010,N_594,In_1182);
nand U1011 (N_1011,N_963,N_718);
nor U1012 (N_1012,In_1629,In_272);
nand U1013 (N_1013,In_1950,In_2423);
nand U1014 (N_1014,N_820,In_574);
and U1015 (N_1015,N_3,N_280);
nor U1016 (N_1016,N_602,In_671);
nor U1017 (N_1017,N_381,In_911);
and U1018 (N_1018,In_1380,N_172);
nor U1019 (N_1019,In_1368,In_2388);
nor U1020 (N_1020,N_204,N_369);
xnor U1021 (N_1021,In_623,In_164);
nor U1022 (N_1022,In_1372,In_617);
or U1023 (N_1023,N_614,N_790);
and U1024 (N_1024,In_2487,In_257);
and U1025 (N_1025,N_982,In_2396);
nor U1026 (N_1026,N_701,In_2289);
nor U1027 (N_1027,In_2417,In_2355);
or U1028 (N_1028,N_533,N_923);
or U1029 (N_1029,In_1835,In_1177);
nand U1030 (N_1030,In_894,N_796);
nor U1031 (N_1031,N_22,In_1509);
and U1032 (N_1032,N_742,N_978);
or U1033 (N_1033,N_569,N_515);
or U1034 (N_1034,In_883,In_459);
nor U1035 (N_1035,N_958,N_516);
and U1036 (N_1036,In_1677,In_149);
and U1037 (N_1037,In_418,N_365);
and U1038 (N_1038,In_174,In_952);
nand U1039 (N_1039,In_1766,In_1003);
or U1040 (N_1040,In_2210,N_999);
nand U1041 (N_1041,In_488,In_457);
nor U1042 (N_1042,N_570,N_894);
xnor U1043 (N_1043,N_175,N_575);
xnor U1044 (N_1044,In_1452,In_1969);
or U1045 (N_1045,N_992,In_2363);
nor U1046 (N_1046,N_778,In_1682);
nand U1047 (N_1047,In_1548,N_731);
or U1048 (N_1048,In_245,N_899);
or U1049 (N_1049,N_151,In_839);
or U1050 (N_1050,N_651,In_284);
nor U1051 (N_1051,In_687,N_661);
nand U1052 (N_1052,In_319,N_274);
nor U1053 (N_1053,In_1775,N_659);
xor U1054 (N_1054,In_719,N_821);
nor U1055 (N_1055,In_1767,N_993);
nor U1056 (N_1056,In_1223,N_669);
nand U1057 (N_1057,N_954,In_2492);
and U1058 (N_1058,In_19,N_443);
nand U1059 (N_1059,In_2066,In_1063);
and U1060 (N_1060,N_966,N_519);
nor U1061 (N_1061,In_116,N_451);
nand U1062 (N_1062,In_1256,In_1685);
nand U1063 (N_1063,N_327,N_853);
nand U1064 (N_1064,N_825,N_715);
or U1065 (N_1065,In_1104,In_992);
nor U1066 (N_1066,N_76,N_767);
and U1067 (N_1067,N_784,N_623);
nor U1068 (N_1068,In_1529,N_865);
nor U1069 (N_1069,N_716,N_688);
or U1070 (N_1070,In_503,N_684);
nand U1071 (N_1071,In_218,In_1464);
nor U1072 (N_1072,N_506,N_950);
nand U1073 (N_1073,In_7,N_513);
nand U1074 (N_1074,In_1787,In_2352);
or U1075 (N_1075,N_41,In_39);
nand U1076 (N_1076,N_863,N_785);
and U1077 (N_1077,In_1881,In_2059);
nand U1078 (N_1078,In_1973,N_601);
nor U1079 (N_1079,In_354,N_521);
or U1080 (N_1080,N_919,N_964);
and U1081 (N_1081,N_545,In_2382);
or U1082 (N_1082,In_979,In_2082);
and U1083 (N_1083,In_4,N_998);
and U1084 (N_1084,N_939,In_2478);
and U1085 (N_1085,N_36,In_2020);
nand U1086 (N_1086,In_2007,N_879);
nand U1087 (N_1087,N_185,In_332);
nand U1088 (N_1088,In_1445,N_655);
nor U1089 (N_1089,In_655,N_316);
nand U1090 (N_1090,N_50,In_2247);
and U1091 (N_1091,N_779,In_1591);
or U1092 (N_1092,N_813,In_2460);
nand U1093 (N_1093,N_696,N_675);
or U1094 (N_1094,In_2447,In_907);
nand U1095 (N_1095,In_525,In_656);
or U1096 (N_1096,In_2418,In_2344);
nor U1097 (N_1097,In_2260,N_892);
nor U1098 (N_1098,N_20,N_461);
nor U1099 (N_1099,In_2380,N_780);
nor U1100 (N_1100,N_133,In_557);
or U1101 (N_1101,N_241,N_552);
xor U1102 (N_1102,In_2296,In_1904);
or U1103 (N_1103,N_700,N_941);
or U1104 (N_1104,N_102,In_608);
nand U1105 (N_1105,N_107,In_473);
and U1106 (N_1106,In_827,In_1797);
xor U1107 (N_1107,In_1739,In_787);
or U1108 (N_1108,N_306,N_828);
and U1109 (N_1109,In_1042,In_864);
and U1110 (N_1110,In_1580,In_1366);
nand U1111 (N_1111,In_2147,N_949);
and U1112 (N_1112,N_729,N_885);
nand U1113 (N_1113,In_462,N_795);
nor U1114 (N_1114,N_281,N_896);
nor U1115 (N_1115,N_495,In_2134);
nor U1116 (N_1116,In_1913,In_2057);
nand U1117 (N_1117,In_2136,N_926);
or U1118 (N_1118,In_426,In_1247);
and U1119 (N_1119,In_377,In_1728);
nand U1120 (N_1120,N_479,N_548);
or U1121 (N_1121,In_1877,N_132);
and U1122 (N_1122,N_127,N_80);
or U1123 (N_1123,N_503,N_595);
or U1124 (N_1124,N_579,In_1900);
nor U1125 (N_1125,N_145,In_1097);
nand U1126 (N_1126,In_357,In_2031);
and U1127 (N_1127,N_838,In_287);
nand U1128 (N_1128,N_6,In_381);
and U1129 (N_1129,In_1992,N_957);
nor U1130 (N_1130,N_256,N_557);
nand U1131 (N_1131,In_1994,N_736);
and U1132 (N_1132,N_39,In_811);
and U1133 (N_1133,In_1999,N_895);
or U1134 (N_1134,In_371,In_1519);
or U1135 (N_1135,In_2383,N_619);
nor U1136 (N_1136,In_1574,N_845);
and U1137 (N_1137,N_807,N_650);
nand U1138 (N_1138,N_568,N_77);
or U1139 (N_1139,In_1393,In_1663);
or U1140 (N_1140,N_986,In_1891);
and U1141 (N_1141,In_962,N_282);
nor U1142 (N_1142,In_1196,In_1082);
or U1143 (N_1143,In_1816,N_740);
and U1144 (N_1144,N_423,In_1701);
and U1145 (N_1145,In_705,N_303);
or U1146 (N_1146,N_4,In_1536);
and U1147 (N_1147,In_2457,In_971);
or U1148 (N_1148,In_541,In_2073);
xnor U1149 (N_1149,In_1630,N_244);
nand U1150 (N_1150,N_830,In_25);
and U1151 (N_1151,N_524,In_1318);
nand U1152 (N_1152,N_771,In_1664);
or U1153 (N_1153,N_751,N_761);
or U1154 (N_1154,In_1145,In_1619);
nand U1155 (N_1155,In_1297,N_818);
and U1156 (N_1156,N_620,In_569);
nand U1157 (N_1157,N_349,In_1049);
nand U1158 (N_1158,In_946,In_59);
and U1159 (N_1159,In_1055,N_768);
or U1160 (N_1160,In_111,N_835);
and U1161 (N_1161,In_1596,N_565);
or U1162 (N_1162,In_844,N_224);
nor U1163 (N_1163,In_1545,In_795);
nor U1164 (N_1164,N_732,N_491);
nand U1165 (N_1165,N_179,N_869);
nor U1166 (N_1166,N_225,In_1459);
nor U1167 (N_1167,N_599,N_706);
or U1168 (N_1168,In_768,N_615);
and U1169 (N_1169,In_981,In_2376);
and U1170 (N_1170,N_558,N_632);
and U1171 (N_1171,In_1316,In_74);
nor U1172 (N_1172,In_1895,N_90);
nor U1173 (N_1173,In_537,In_851);
and U1174 (N_1174,In_755,N_605);
and U1175 (N_1175,In_1255,In_746);
nand U1176 (N_1176,N_900,N_411);
nand U1177 (N_1177,In_925,N_930);
nor U1178 (N_1178,In_207,In_2331);
and U1179 (N_1179,In_568,N_466);
nand U1180 (N_1180,In_622,N_681);
and U1181 (N_1181,In_1244,N_911);
nor U1182 (N_1182,N_66,N_929);
nor U1183 (N_1183,In_1544,In_1195);
nor U1184 (N_1184,In_1474,In_1717);
or U1185 (N_1185,N_223,N_877);
and U1186 (N_1186,N_432,N_549);
xnor U1187 (N_1187,In_2196,In_1611);
nor U1188 (N_1188,N_544,N_917);
and U1189 (N_1189,In_550,In_908);
or U1190 (N_1190,In_308,In_2052);
nor U1191 (N_1191,In_1173,N_756);
nand U1192 (N_1192,In_1428,N_78);
or U1193 (N_1193,In_2127,In_1982);
and U1194 (N_1194,In_579,In_2185);
nand U1195 (N_1195,In_1572,N_154);
nor U1196 (N_1196,In_1577,In_2360);
and U1197 (N_1197,In_771,N_678);
and U1198 (N_1198,N_202,N_876);
nor U1199 (N_1199,In_1006,N_833);
nand U1200 (N_1200,N_898,N_622);
and U1201 (N_1201,N_155,In_1168);
or U1202 (N_1202,In_286,N_984);
or U1203 (N_1203,In_1126,N_955);
nor U1204 (N_1204,N_959,N_680);
nand U1205 (N_1205,In_1188,In_480);
nand U1206 (N_1206,In_2256,In_1633);
nor U1207 (N_1207,N_286,In_2198);
and U1208 (N_1208,N_826,In_852);
nor U1209 (N_1209,In_2182,N_804);
or U1210 (N_1210,N_971,In_2471);
or U1211 (N_1211,N_359,In_1289);
nand U1212 (N_1212,N_960,In_129);
nor U1213 (N_1213,N_737,N_304);
nor U1214 (N_1214,In_1264,In_2110);
nor U1215 (N_1215,In_2499,In_2242);
or U1216 (N_1216,In_1321,In_2494);
and U1217 (N_1217,N_265,N_672);
or U1218 (N_1218,In_1224,N_840);
nor U1219 (N_1219,N_658,In_1941);
nor U1220 (N_1220,In_742,In_571);
nand U1221 (N_1221,In_1198,In_1762);
nand U1222 (N_1222,N_856,N_938);
and U1223 (N_1223,N_974,N_727);
nor U1224 (N_1224,In_114,N_777);
nor U1225 (N_1225,In_993,N_967);
or U1226 (N_1226,In_2273,In_130);
or U1227 (N_1227,In_2168,N_965);
and U1228 (N_1228,N_739,In_2314);
nand U1229 (N_1229,N_760,N_216);
nor U1230 (N_1230,N_250,In_2173);
and U1231 (N_1231,N_893,In_228);
nand U1232 (N_1232,N_21,N_464);
nor U1233 (N_1233,In_1526,In_2463);
nand U1234 (N_1234,N_84,In_2199);
and U1235 (N_1235,In_1733,In_1975);
nor U1236 (N_1236,In_1831,In_445);
nor U1237 (N_1237,In_931,N_307);
nand U1238 (N_1238,In_61,N_25);
nor U1239 (N_1239,N_714,N_497);
nor U1240 (N_1240,In_1336,In_1133);
or U1241 (N_1241,In_190,N_525);
and U1242 (N_1242,In_2179,In_373);
nor U1243 (N_1243,N_539,N_943);
and U1244 (N_1244,In_1119,In_1416);
and U1245 (N_1245,In_2004,N_375);
xor U1246 (N_1246,In_919,In_1662);
nor U1247 (N_1247,In_1381,In_1408);
nand U1248 (N_1248,N_587,In_1303);
or U1249 (N_1249,In_143,N_413);
or U1250 (N_1250,N_57,In_1714);
nor U1251 (N_1251,N_720,N_318);
or U1252 (N_1252,In_1750,N_945);
nand U1253 (N_1253,N_449,N_713);
or U1254 (N_1254,In_1822,In_1258);
and U1255 (N_1255,In_947,N_232);
or U1256 (N_1256,In_1857,In_2429);
and U1257 (N_1257,N_944,In_2053);
nand U1258 (N_1258,In_1905,N_382);
nor U1259 (N_1259,In_582,In_1);
and U1260 (N_1260,In_99,N_507);
and U1261 (N_1261,In_472,N_695);
nor U1262 (N_1262,In_1218,In_1204);
nand U1263 (N_1263,In_1123,N_563);
and U1264 (N_1264,In_131,N_916);
and U1265 (N_1265,In_1457,N_884);
and U1266 (N_1266,In_407,N_31);
nor U1267 (N_1267,N_934,In_428);
xor U1268 (N_1268,N_0,In_2298);
nor U1269 (N_1269,In_341,In_945);
or U1270 (N_1270,In_217,N_397);
or U1271 (N_1271,In_2111,In_298);
xnor U1272 (N_1272,N_639,In_51);
nor U1273 (N_1273,N_846,In_363);
nor U1274 (N_1274,N_867,In_1317);
nand U1275 (N_1275,N_653,N_504);
and U1276 (N_1276,N_755,N_769);
or U1277 (N_1277,In_2237,In_2126);
nand U1278 (N_1278,In_2169,N_522);
nor U1279 (N_1279,In_154,In_496);
or U1280 (N_1280,In_748,In_353);
or U1281 (N_1281,N_593,N_182);
nand U1282 (N_1282,N_994,In_471);
and U1283 (N_1283,N_108,In_2276);
xnor U1284 (N_1284,N_170,N_97);
nand U1285 (N_1285,In_2013,N_630);
or U1286 (N_1286,N_774,In_1426);
and U1287 (N_1287,In_1473,In_2252);
xor U1288 (N_1288,N_458,N_850);
or U1289 (N_1289,In_588,In_2218);
or U1290 (N_1290,N_387,In_829);
nor U1291 (N_1291,In_2088,N_843);
nor U1292 (N_1292,In_1261,In_2081);
nand U1293 (N_1293,In_215,N_870);
and U1294 (N_1294,N_559,N_946);
and U1295 (N_1295,N_985,In_1307);
nand U1296 (N_1296,In_1672,N_698);
nand U1297 (N_1297,In_17,In_2060);
nor U1298 (N_1298,N_738,In_630);
nand U1299 (N_1299,N_799,N_567);
nor U1300 (N_1300,N_162,N_810);
nand U1301 (N_1301,In_2285,In_292);
and U1302 (N_1302,In_343,N_775);
nor U1303 (N_1303,In_451,N_660);
nand U1304 (N_1304,In_253,N_328);
or U1305 (N_1305,N_902,In_2236);
and U1306 (N_1306,N_711,In_196);
nand U1307 (N_1307,N_890,N_98);
or U1308 (N_1308,In_2317,In_1266);
nor U1309 (N_1309,N_679,N_643);
or U1310 (N_1310,N_180,In_873);
and U1311 (N_1311,N_203,In_1514);
or U1312 (N_1312,In_2230,N_82);
or U1313 (N_1313,In_269,In_1429);
or U1314 (N_1314,In_1915,In_2);
nor U1315 (N_1315,N_81,N_331);
nor U1316 (N_1316,In_293,N_708);
and U1317 (N_1317,N_560,In_123);
nand U1318 (N_1318,In_238,N_562);
nor U1319 (N_1319,N_819,N_17);
nor U1320 (N_1320,In_1582,N_55);
and U1321 (N_1321,N_538,N_606);
nor U1322 (N_1322,N_150,N_356);
or U1323 (N_1323,In_935,In_903);
or U1324 (N_1324,N_762,In_1193);
nor U1325 (N_1325,N_812,N_629);
or U1326 (N_1326,In_1327,N_918);
or U1327 (N_1327,In_800,N_537);
nor U1328 (N_1328,In_1696,In_932);
and U1329 (N_1329,In_118,N_634);
nor U1330 (N_1330,N_690,N_165);
nor U1331 (N_1331,N_528,In_294);
and U1332 (N_1332,In_448,N_168);
or U1333 (N_1333,N_849,In_1005);
and U1334 (N_1334,N_882,In_854);
and U1335 (N_1335,In_710,N_508);
nand U1336 (N_1336,N_766,In_1673);
or U1337 (N_1337,In_866,In_1770);
or U1338 (N_1338,In_1375,In_1615);
or U1339 (N_1339,In_1513,In_1434);
nor U1340 (N_1340,In_2311,N_914);
and U1341 (N_1341,In_1746,In_1068);
or U1342 (N_1342,In_2442,N_426);
or U1343 (N_1343,N_101,N_578);
nand U1344 (N_1344,In_1512,In_2304);
nand U1345 (N_1345,N_829,N_648);
or U1346 (N_1346,N_717,In_1930);
and U1347 (N_1347,N_710,In_1384);
or U1348 (N_1348,N_995,N_219);
xnor U1349 (N_1349,N_398,N_633);
nor U1350 (N_1350,In_522,N_442);
and U1351 (N_1351,N_734,In_246);
and U1352 (N_1352,N_99,N_797);
or U1353 (N_1353,N_924,N_662);
nand U1354 (N_1354,In_618,N_907);
nor U1355 (N_1355,In_2445,In_1355);
nand U1356 (N_1356,In_2069,In_251);
nand U1357 (N_1357,In_2062,In_2181);
nand U1358 (N_1358,N_532,In_1906);
nand U1359 (N_1359,In_2334,In_1206);
nand U1360 (N_1360,In_1984,In_1037);
or U1361 (N_1361,In_688,In_2064);
and U1362 (N_1362,In_1939,N_95);
and U1363 (N_1363,In_1658,N_645);
nor U1364 (N_1364,N_546,N_340);
nand U1365 (N_1365,N_635,N_428);
xnor U1366 (N_1366,In_372,N_646);
nand U1367 (N_1367,In_838,N_597);
and U1368 (N_1368,N_921,N_968);
xor U1369 (N_1369,In_1271,N_724);
and U1370 (N_1370,In_1570,In_1647);
nand U1371 (N_1371,N_581,N_517);
and U1372 (N_1372,N_642,N_367);
or U1373 (N_1373,In_511,N_803);
nor U1374 (N_1374,N_129,In_2161);
or U1375 (N_1375,In_2076,N_590);
and U1376 (N_1376,N_598,In_774);
and U1377 (N_1377,In_2001,In_1830);
nor U1378 (N_1378,N_494,In_345);
nor U1379 (N_1379,In_1222,N_691);
nor U1380 (N_1380,N_972,N_961);
nor U1381 (N_1381,In_1692,N_2);
nor U1382 (N_1382,In_1613,In_1163);
nor U1383 (N_1383,In_461,In_524);
nand U1384 (N_1384,In_279,In_42);
nor U1385 (N_1385,In_1085,N_641);
and U1386 (N_1386,N_500,In_1052);
and U1387 (N_1387,N_24,In_849);
xnor U1388 (N_1388,N_566,In_1025);
nor U1389 (N_1389,In_1931,In_941);
nand U1390 (N_1390,In_2131,In_1712);
nor U1391 (N_1391,N_844,N_105);
nor U1392 (N_1392,In_2307,N_754);
nand U1393 (N_1393,In_1788,In_1093);
and U1394 (N_1394,N_130,N_321);
or U1395 (N_1395,N_18,In_2448);
nand U1396 (N_1396,In_646,N_63);
xor U1397 (N_1397,In_1056,In_1774);
xnor U1398 (N_1398,N_665,N_991);
nor U1399 (N_1399,N_422,N_977);
nand U1400 (N_1400,N_951,N_209);
and U1401 (N_1401,In_210,N_789);
nand U1402 (N_1402,In_825,In_728);
or U1403 (N_1403,In_2178,N_206);
nand U1404 (N_1404,In_1027,In_440);
nor U1405 (N_1405,N_842,N_540);
nand U1406 (N_1406,N_683,In_1556);
and U1407 (N_1407,N_613,In_1776);
nand U1408 (N_1408,In_1262,N_520);
and U1409 (N_1409,N_183,N_868);
nor U1410 (N_1410,In_1352,In_2275);
xnor U1411 (N_1411,In_1443,N_847);
nand U1412 (N_1412,N_947,N_536);
xor U1413 (N_1413,In_364,In_1160);
or U1414 (N_1414,N_322,In_1952);
and U1415 (N_1415,In_954,In_1972);
xor U1416 (N_1416,In_1737,N_535);
nor U1417 (N_1417,N_878,In_1758);
nand U1418 (N_1418,N_908,N_453);
and U1419 (N_1419,In_532,In_1771);
or U1420 (N_1420,N_741,In_2170);
and U1421 (N_1421,N_953,N_628);
or U1422 (N_1422,N_110,In_1032);
nand U1423 (N_1423,In_725,In_1296);
or U1424 (N_1424,In_498,In_815);
and U1425 (N_1425,N_343,N_915);
nor U1426 (N_1426,In_1159,In_847);
and U1427 (N_1427,N_292,N_610);
and U1428 (N_1428,In_466,In_1951);
or U1429 (N_1429,In_1944,N_393);
nand U1430 (N_1430,N_12,In_275);
and U1431 (N_1431,In_2190,In_850);
nand U1432 (N_1432,N_576,In_10);
nand U1433 (N_1433,N_276,N_542);
xor U1434 (N_1434,N_855,In_726);
or U1435 (N_1435,N_983,N_255);
and U1436 (N_1436,In_2323,N_699);
nor U1437 (N_1437,N_794,In_235);
nand U1438 (N_1438,In_1940,N_837);
xor U1439 (N_1439,In_2469,In_1855);
nand U1440 (N_1440,N_852,N_399);
nor U1441 (N_1441,N_806,N_388);
nor U1442 (N_1442,N_596,N_656);
nand U1443 (N_1443,N_839,N_166);
nor U1444 (N_1444,In_637,In_1096);
xnor U1445 (N_1445,In_313,N_580);
nand U1446 (N_1446,In_1657,N_834);
and U1447 (N_1447,N_783,N_534);
nand U1448 (N_1448,In_434,N_802);
or U1449 (N_1449,N_752,N_703);
and U1450 (N_1450,N_773,N_793);
nor U1451 (N_1451,N_913,N_67);
or U1452 (N_1452,In_1694,In_501);
nor U1453 (N_1453,In_147,N_747);
and U1454 (N_1454,N_922,In_529);
or U1455 (N_1455,In_649,N_956);
and U1456 (N_1456,In_2470,N_848);
nand U1457 (N_1457,N_191,N_745);
and U1458 (N_1458,In_824,N_750);
nor U1459 (N_1459,N_100,N_314);
nor U1460 (N_1460,In_1475,In_2493);
nor U1461 (N_1461,N_246,N_705);
nor U1462 (N_1462,In_2000,N_489);
nor U1463 (N_1463,In_972,In_2458);
nor U1464 (N_1464,N_743,In_898);
or U1465 (N_1465,N_23,N_817);
or U1466 (N_1466,In_2245,N_351);
nor U1467 (N_1467,In_556,N_370);
nor U1468 (N_1468,N_990,In_934);
nor U1469 (N_1469,In_2424,N_822);
or U1470 (N_1470,N_48,N_636);
nand U1471 (N_1471,In_2229,N_976);
nor U1472 (N_1472,N_721,N_649);
nor U1473 (N_1473,N_571,N_29);
and U1474 (N_1474,In_1680,In_2348);
or U1475 (N_1475,In_1077,N_730);
and U1476 (N_1476,In_1433,N_765);
and U1477 (N_1477,N_429,In_764);
and U1478 (N_1478,In_1134,N_421);
and U1479 (N_1479,In_316,N_928);
and U1480 (N_1480,In_397,N_728);
and U1481 (N_1481,In_1189,In_55);
and U1482 (N_1482,In_2433,N_37);
or U1483 (N_1483,In_329,In_1101);
and U1484 (N_1484,N_816,N_759);
or U1485 (N_1485,In_1107,In_1181);
or U1486 (N_1486,N_707,N_942);
or U1487 (N_1487,N_627,N_128);
nor U1488 (N_1488,N_874,N_611);
nor U1489 (N_1489,N_996,In_82);
and U1490 (N_1490,In_1917,In_1808);
nand U1491 (N_1491,N_392,In_676);
and U1492 (N_1492,In_1598,In_1644);
nor U1493 (N_1493,N_325,N_531);
xnor U1494 (N_1494,In_717,In_1708);
nand U1495 (N_1495,N_616,N_786);
nor U1496 (N_1496,In_2084,N_446);
and U1497 (N_1497,In_1655,N_866);
or U1498 (N_1498,N_625,N_677);
or U1499 (N_1499,N_296,In_2295);
nand U1500 (N_1500,In_1695,In_1624);
or U1501 (N_1501,N_664,N_682);
or U1502 (N_1502,N_805,N_1142);
nand U1503 (N_1503,N_1128,N_407);
nor U1504 (N_1504,N_541,N_1011);
and U1505 (N_1505,N_502,N_471);
nor U1506 (N_1506,N_746,In_976);
nand U1507 (N_1507,In_595,N_262);
nor U1508 (N_1508,N_1134,N_1090);
and U1509 (N_1509,N_1102,N_1362);
nand U1510 (N_1510,N_880,N_1395);
nor U1511 (N_1511,N_1496,N_1218);
nor U1512 (N_1512,N_454,N_1217);
nand U1513 (N_1513,In_2005,N_1020);
nor U1514 (N_1514,N_676,N_764);
nor U1515 (N_1515,In_1727,N_888);
nand U1516 (N_1516,N_64,In_1399);
nand U1517 (N_1517,N_704,N_1459);
or U1518 (N_1518,N_1368,N_1493);
and U1519 (N_1519,In_399,In_933);
nor U1520 (N_1520,N_260,N_1070);
and U1521 (N_1521,N_1146,In_959);
or U1522 (N_1522,N_1015,In_1058);
nor U1523 (N_1523,N_1222,In_745);
and U1524 (N_1524,In_2002,N_1159);
or U1525 (N_1525,N_772,N_1348);
nor U1526 (N_1526,N_1409,N_782);
or U1527 (N_1527,In_781,N_1155);
nor U1528 (N_1528,In_2028,In_2077);
nor U1529 (N_1529,N_1322,N_1356);
nand U1530 (N_1530,N_980,N_733);
and U1531 (N_1531,N_1037,In_1752);
or U1532 (N_1532,N_391,In_1493);
and U1533 (N_1533,N_1135,N_854);
or U1534 (N_1534,In_616,N_670);
or U1535 (N_1535,N_588,N_1027);
nand U1536 (N_1536,N_1446,N_353);
or U1537 (N_1537,N_222,In_1686);
or U1538 (N_1538,N_673,N_1068);
or U1539 (N_1539,N_638,N_1169);
or U1540 (N_1540,N_1125,N_758);
nand U1541 (N_1541,N_831,N_1019);
or U1542 (N_1542,N_904,In_575);
nor U1543 (N_1543,N_1482,In_853);
nand U1544 (N_1544,In_879,N_1269);
or U1545 (N_1545,In_427,N_1441);
nand U1546 (N_1546,N_1450,N_1399);
nor U1547 (N_1547,N_530,N_1061);
nand U1548 (N_1548,In_953,In_643);
or U1549 (N_1549,N_1248,N_674);
nor U1550 (N_1550,N_603,In_31);
and U1551 (N_1551,N_1282,N_476);
and U1552 (N_1552,In_5,N_626);
or U1553 (N_1553,N_920,N_1444);
nor U1554 (N_1554,In_303,N_1183);
nand U1555 (N_1555,N_1008,N_1145);
and U1556 (N_1556,In_2204,In_348);
and U1557 (N_1557,N_1491,N_1289);
or U1558 (N_1558,N_935,N_74);
and U1559 (N_1559,In_1100,N_1370);
nor U1560 (N_1560,N_44,N_1477);
nor U1561 (N_1561,N_1418,N_1460);
nand U1562 (N_1562,N_875,N_401);
or U1563 (N_1563,N_1420,N_726);
nor U1564 (N_1564,In_1782,N_1130);
or U1565 (N_1565,N_1413,N_1379);
or U1566 (N_1566,N_1445,N_1230);
nand U1567 (N_1567,N_1124,N_1288);
and U1568 (N_1568,N_1401,N_671);
or U1569 (N_1569,N_1198,N_243);
nand U1570 (N_1570,N_1039,In_2107);
or U1571 (N_1571,N_647,N_1171);
nor U1572 (N_1572,In_1912,N_1262);
and U1573 (N_1573,N_1344,In_421);
nand U1574 (N_1574,N_1285,N_1003);
xor U1575 (N_1575,N_749,In_2419);
and U1576 (N_1576,In_1801,N_505);
and U1577 (N_1577,N_1383,In_405);
nor U1578 (N_1578,N_1221,In_429);
or U1579 (N_1579,N_156,N_1347);
or U1580 (N_1580,N_585,N_1103);
and U1581 (N_1581,In_1748,N_1442);
or U1582 (N_1582,N_1333,N_1273);
or U1583 (N_1583,N_1311,N_1259);
nand U1584 (N_1584,N_1064,In_1837);
or U1585 (N_1585,N_1253,N_1371);
and U1586 (N_1586,N_1006,N_1082);
nor U1587 (N_1587,In_1772,In_2015);
or U1588 (N_1588,In_2254,N_118);
nor U1589 (N_1589,N_1021,In_1337);
and U1590 (N_1590,In_1815,N_912);
and U1591 (N_1591,N_1132,N_1012);
nand U1592 (N_1592,N_523,N_1091);
nand U1593 (N_1593,N_1213,N_1303);
nor U1594 (N_1594,N_1063,N_1224);
nand U1595 (N_1595,N_1234,N_1337);
and U1596 (N_1596,N_800,In_1532);
and U1597 (N_1597,N_1278,N_1291);
nor U1598 (N_1598,N_1170,N_1196);
or U1599 (N_1599,N_1349,N_1137);
nand U1600 (N_1600,N_608,N_861);
nor U1601 (N_1601,In_870,N_1261);
and U1602 (N_1602,N_1300,N_1480);
nor U1603 (N_1603,N_1054,In_789);
nand U1604 (N_1604,In_1726,In_1869);
or U1605 (N_1605,N_1484,N_1016);
or U1606 (N_1606,N_1425,N_814);
and U1607 (N_1607,N_217,N_1210);
or U1608 (N_1608,N_1351,In_1132);
nand U1609 (N_1609,N_1378,N_591);
nand U1610 (N_1610,N_1268,In_1981);
and U1611 (N_1611,N_1392,In_136);
and U1612 (N_1612,N_1452,In_2312);
or U1613 (N_1613,N_1394,N_1023);
nor U1614 (N_1614,N_212,In_1156);
xnor U1615 (N_1615,N_1240,In_642);
or U1616 (N_1616,N_253,In_822);
or U1617 (N_1617,N_612,N_363);
nor U1618 (N_1618,In_23,In_1422);
and U1619 (N_1619,N_1342,N_238);
nand U1620 (N_1620,In_713,N_186);
nand U1621 (N_1621,N_1229,N_188);
nand U1622 (N_1622,In_2010,N_543);
nor U1623 (N_1623,N_1270,In_487);
nor U1624 (N_1624,N_1398,N_1306);
nand U1625 (N_1625,In_1524,N_1168);
nand U1626 (N_1626,N_252,N_1405);
nand U1627 (N_1627,N_56,N_1161);
xnor U1628 (N_1628,N_1244,N_1166);
nand U1629 (N_1629,N_240,N_59);
nor U1630 (N_1630,N_962,N_1067);
and U1631 (N_1631,N_1226,N_1438);
nor U1632 (N_1632,N_609,In_594);
or U1633 (N_1633,In_1718,N_1298);
and U1634 (N_1634,N_906,N_1412);
or U1635 (N_1635,N_1297,In_3);
nor U1636 (N_1636,N_1353,N_1363);
and U1637 (N_1637,N_1180,N_1323);
or U1638 (N_1638,N_1302,In_638);
or U1639 (N_1639,N_547,N_886);
nand U1640 (N_1640,N_1390,N_1236);
and U1641 (N_1641,N_1443,N_1005);
and U1642 (N_1642,In_14,N_1108);
or U1643 (N_1643,N_501,N_1219);
and U1644 (N_1644,N_1369,N_841);
xnor U1645 (N_1645,N_1177,N_1263);
nor U1646 (N_1646,N_1029,In_644);
or U1647 (N_1647,N_1354,In_1550);
or U1648 (N_1648,In_391,N_512);
nor U1649 (N_1649,N_1173,In_521);
nand U1650 (N_1650,N_377,In_2128);
or U1651 (N_1651,N_1447,In_611);
nand U1652 (N_1652,N_809,N_1096);
nor U1653 (N_1653,N_1231,N_1000);
xor U1654 (N_1654,N_1305,In_197);
or U1655 (N_1655,N_1457,N_589);
nor U1656 (N_1656,N_1366,N_361);
nor U1657 (N_1657,N_1332,N_1265);
or U1658 (N_1658,N_770,N_1292);
or U1659 (N_1659,In_1240,N_1085);
and U1660 (N_1660,N_1455,In_1021);
or U1661 (N_1661,N_1163,N_1456);
or U1662 (N_1662,N_1220,N_887);
nor U1663 (N_1663,N_1463,N_1277);
nor U1664 (N_1664,N_1403,N_1275);
nor U1665 (N_1665,N_1098,In_964);
and U1666 (N_1666,In_110,In_2474);
nand U1667 (N_1667,N_857,N_1238);
nand U1668 (N_1668,N_1422,N_1164);
and U1669 (N_1669,In_402,N_1247);
nand U1670 (N_1670,N_1184,N_1185);
nand U1671 (N_1671,N_1228,N_1001);
nand U1672 (N_1672,N_586,In_802);
and U1673 (N_1673,In_1136,N_1343);
nand U1674 (N_1674,N_159,N_1089);
or U1675 (N_1675,N_903,N_1002);
nand U1676 (N_1676,N_1257,In_2216);
nand U1677 (N_1677,In_1364,In_1898);
and U1678 (N_1678,N_1312,N_1492);
and U1679 (N_1679,N_1280,N_1380);
or U1680 (N_1680,N_109,N_1421);
and U1681 (N_1681,N_1172,In_1212);
xnor U1682 (N_1682,N_1150,N_932);
or U1683 (N_1683,N_1267,N_1133);
or U1684 (N_1684,N_1118,N_1410);
and U1685 (N_1685,N_1359,N_509);
nor U1686 (N_1686,In_2189,N_529);
and U1687 (N_1687,N_891,N_1479);
or U1688 (N_1688,N_1320,N_131);
nor U1689 (N_1689,N_106,In_1700);
and U1690 (N_1690,N_1453,N_1175);
and U1691 (N_1691,N_1352,N_510);
or U1692 (N_1692,In_895,In_902);
and U1693 (N_1693,N_1487,N_1143);
and U1694 (N_1694,In_1790,In_135);
nor U1695 (N_1695,N_1301,N_297);
and U1696 (N_1696,In_1420,N_1427);
nand U1697 (N_1697,N_1385,In_1511);
and U1698 (N_1698,N_1065,N_640);
and U1699 (N_1699,N_693,N_1497);
or U1700 (N_1700,N_1110,N_1283);
nand U1701 (N_1701,In_2099,N_1088);
nor U1702 (N_1702,N_1041,N_735);
nand U1703 (N_1703,N_975,N_408);
or U1704 (N_1704,N_1367,N_1440);
nand U1705 (N_1705,In_1369,N_283);
nand U1706 (N_1706,N_1052,N_973);
nand U1707 (N_1707,In_583,N_8);
or U1708 (N_1708,In_1844,N_1047);
nand U1709 (N_1709,N_1148,In_917);
nor U1710 (N_1710,N_1470,N_936);
or U1711 (N_1711,N_1407,N_551);
nand U1712 (N_1712,N_1123,In_1861);
nor U1713 (N_1713,N_1151,N_637);
or U1714 (N_1714,N_1424,In_281);
xnor U1715 (N_1715,N_1149,N_1328);
or U1716 (N_1716,N_394,N_1464);
and U1717 (N_1717,N_1308,N_1435);
nand U1718 (N_1718,N_1038,N_1364);
and U1719 (N_1719,N_905,N_1216);
nand U1720 (N_1720,N_618,In_2361);
or U1721 (N_1721,N_1458,N_1246);
or U1722 (N_1722,In_1409,N_1433);
or U1723 (N_1723,In_2206,In_368);
and U1724 (N_1724,N_881,N_527);
and U1725 (N_1725,In_1731,N_1397);
nand U1726 (N_1726,N_668,N_1190);
and U1727 (N_1727,N_873,N_600);
or U1728 (N_1728,N_1056,N_1072);
or U1729 (N_1729,N_1111,N_1053);
nor U1730 (N_1730,N_414,N_1271);
and U1731 (N_1731,N_1254,N_592);
or U1732 (N_1732,N_1121,In_2272);
or U1733 (N_1733,N_1239,N_1062);
and U1734 (N_1734,In_2243,N_574);
nand U1735 (N_1735,In_1602,In_2209);
or U1736 (N_1736,N_1049,N_948);
or U1737 (N_1737,N_1360,In_282);
or U1738 (N_1738,In_2184,N_72);
nand U1739 (N_1739,In_1833,In_2090);
or U1740 (N_1740,N_1461,N_554);
and U1741 (N_1741,N_1416,N_1017);
nand U1742 (N_1742,N_1051,In_252);
nor U1743 (N_1743,N_1279,N_689);
nor U1744 (N_1744,In_2212,In_15);
nand U1745 (N_1745,N_1154,N_1030);
nand U1746 (N_1746,N_860,In_1280);
nor U1747 (N_1747,In_986,In_1295);
or U1748 (N_1748,In_2036,N_1035);
or U1749 (N_1749,N_697,N_686);
and U1750 (N_1750,N_1423,N_1167);
or U1751 (N_1751,N_1473,N_572);
nor U1752 (N_1752,N_1429,In_1932);
nand U1753 (N_1753,N_1084,N_1287);
nand U1754 (N_1754,N_1260,N_1310);
nand U1755 (N_1755,N_561,N_725);
and U1756 (N_1756,N_871,N_1309);
and U1757 (N_1757,N_1028,In_1480);
or U1758 (N_1758,N_1316,N_1372);
and U1759 (N_1759,N_1406,N_462);
and U1760 (N_1760,N_1044,N_1034);
or U1761 (N_1761,In_389,N_1093);
or U1762 (N_1762,N_1242,N_631);
nor U1763 (N_1763,N_1045,N_1437);
or U1764 (N_1764,In_84,N_1074);
xor U1765 (N_1765,N_1060,N_1189);
nor U1766 (N_1766,In_1310,N_1162);
or U1767 (N_1767,N_1144,N_1494);
and U1768 (N_1768,N_366,N_1252);
nand U1769 (N_1769,N_1434,In_1690);
or U1770 (N_1770,N_692,In_2211);
or U1771 (N_1771,N_617,In_2125);
or U1772 (N_1772,N_1223,N_112);
nor U1773 (N_1773,N_1451,N_355);
nand U1774 (N_1774,N_1488,N_1119);
nor U1775 (N_1775,In_178,N_1036);
or U1776 (N_1776,N_582,In_635);
nor U1777 (N_1777,N_931,N_1073);
nand U1778 (N_1778,N_120,N_239);
nor U1779 (N_1779,N_1138,N_1249);
nand U1780 (N_1780,In_1617,N_1448);
nor U1781 (N_1781,N_719,N_556);
nor U1782 (N_1782,N_901,N_1331);
or U1783 (N_1783,N_1326,N_1340);
and U1784 (N_1784,N_69,N_1317);
and U1785 (N_1785,N_1382,N_1040);
or U1786 (N_1786,In_1395,N_1436);
or U1787 (N_1787,N_511,N_93);
and U1788 (N_1788,N_925,N_1043);
and U1789 (N_1789,N_836,In_1248);
nor U1790 (N_1790,N_757,N_573);
xor U1791 (N_1791,In_773,N_1207);
nor U1792 (N_1792,N_1211,N_455);
nor U1793 (N_1793,N_1059,N_305);
and U1794 (N_1794,N_1215,N_1243);
nor U1795 (N_1795,In_1943,N_1078);
nor U1796 (N_1796,N_1046,N_1208);
or U1797 (N_1797,In_274,N_526);
or U1798 (N_1798,N_1467,In_2294);
xnor U1799 (N_1799,In_1604,N_702);
or U1800 (N_1800,N_553,In_1606);
nor U1801 (N_1801,N_1293,N_1469);
nand U1802 (N_1802,In_2399,N_1387);
or U1803 (N_1803,N_1097,In_1890);
nor U1804 (N_1804,N_1139,N_1389);
or U1805 (N_1805,In_295,N_1314);
or U1806 (N_1806,N_1076,N_1321);
nand U1807 (N_1807,N_1099,N_1115);
nand U1808 (N_1808,N_1081,N_1299);
or U1809 (N_1809,N_1087,In_657);
nand U1810 (N_1810,N_883,N_1071);
nand U1811 (N_1811,N_791,In_1899);
nand U1812 (N_1812,In_1138,N_1258);
and U1813 (N_1813,N_1255,N_909);
nor U1814 (N_1814,N_811,In_1573);
or U1815 (N_1815,N_1205,In_1636);
and U1816 (N_1816,N_474,N_1199);
xnor U1817 (N_1817,N_979,N_798);
and U1818 (N_1818,N_564,N_1375);
and U1819 (N_1819,N_1495,In_780);
nor U1820 (N_1820,N_1462,N_763);
nor U1821 (N_1821,N_1122,N_1430);
nand U1822 (N_1822,N_1010,N_1276);
nand U1823 (N_1823,In_378,In_1344);
or U1824 (N_1824,N_153,N_781);
nor U1825 (N_1825,N_1319,N_1113);
or U1826 (N_1826,N_1318,N_1489);
xor U1827 (N_1827,N_1201,In_2203);
and U1828 (N_1828,In_1843,N_205);
or U1829 (N_1829,In_1140,In_1214);
nor U1830 (N_1830,N_1106,In_510);
nand U1831 (N_1831,N_1004,N_1157);
and U1832 (N_1832,N_722,N_1414);
or U1833 (N_1833,N_301,N_481);
nor U1834 (N_1834,N_815,N_1295);
nand U1835 (N_1835,N_1404,In_578);
and U1836 (N_1836,N_1411,N_644);
or U1837 (N_1837,In_213,In_1554);
nand U1838 (N_1838,In_753,N_1195);
nor U1839 (N_1839,In_1461,N_1120);
and U1840 (N_1840,N_654,N_1095);
nand U1841 (N_1841,N_1066,N_1153);
and U1842 (N_1842,N_1290,N_685);
and U1843 (N_1843,In_612,N_1109);
or U1844 (N_1844,N_1313,In_1953);
nand U1845 (N_1845,N_1481,N_607);
nand U1846 (N_1846,N_604,N_859);
nand U1847 (N_1847,N_1077,N_1086);
and U1848 (N_1848,In_1116,N_46);
and U1849 (N_1849,N_376,N_1428);
nand U1850 (N_1850,In_1851,In_1968);
nand U1851 (N_1851,N_1485,N_1187);
or U1852 (N_1852,In_914,N_1232);
or U1853 (N_1853,N_1104,N_1325);
or U1854 (N_1854,N_1140,N_823);
xnor U1855 (N_1855,N_1182,N_970);
and U1856 (N_1856,N_1376,In_527);
nor U1857 (N_1857,N_709,N_1454);
nand U1858 (N_1858,In_2263,N_1136);
nand U1859 (N_1859,In_2378,N_335);
nand U1860 (N_1860,N_1057,N_910);
nor U1861 (N_1861,N_158,N_1202);
and U1862 (N_1862,N_1327,In_1916);
nand U1863 (N_1863,N_1388,N_824);
or U1864 (N_1864,In_2324,N_122);
or U1865 (N_1865,N_988,N_483);
and U1866 (N_1866,N_969,N_1338);
nor U1867 (N_1867,In_177,N_1432);
or U1868 (N_1868,N_1200,N_487);
nand U1869 (N_1869,N_1237,N_1474);
nor U1870 (N_1870,N_32,In_1099);
xor U1871 (N_1871,In_761,In_526);
or U1872 (N_1872,N_1013,In_12);
nand U1873 (N_1873,N_294,N_788);
and U1874 (N_1874,N_1296,N_748);
nor U1875 (N_1875,N_1192,In_1919);
and U1876 (N_1876,In_752,N_1274);
nand U1877 (N_1877,N_1374,N_1475);
nand U1878 (N_1878,In_121,In_1632);
nand U1879 (N_1879,N_657,N_1324);
or U1880 (N_1880,In_2223,N_927);
nand U1881 (N_1881,N_42,N_787);
and U1882 (N_1882,N_1486,N_1188);
xnor U1883 (N_1883,In_344,In_1576);
and U1884 (N_1884,N_514,N_1336);
or U1885 (N_1885,N_1339,N_1471);
or U1886 (N_1886,In_994,N_418);
and U1887 (N_1887,N_1032,N_550);
and U1888 (N_1888,N_1100,N_1384);
and U1889 (N_1889,In_2449,N_1417);
or U1890 (N_1890,In_2106,N_1281);
nand U1891 (N_1891,N_1284,N_555);
and U1892 (N_1892,In_910,N_1055);
and U1893 (N_1893,N_1483,N_1105);
nor U1894 (N_1894,In_1793,In_1872);
or U1895 (N_1895,N_1026,In_73);
or U1896 (N_1896,N_1402,N_104);
nand U1897 (N_1897,N_71,N_1014);
nor U1898 (N_1898,N_1152,N_1024);
and U1899 (N_1899,N_1341,N_1250);
or U1900 (N_1900,N_1355,In_317);
and U1901 (N_1901,N_267,N_1101);
and U1902 (N_1902,N_1181,N_1465);
nor U1903 (N_1903,N_1126,N_1478);
and U1904 (N_1904,N_1358,N_1009);
nor U1905 (N_1905,N_621,N_237);
nand U1906 (N_1906,N_997,In_2033);
or U1907 (N_1907,N_624,N_827);
nand U1908 (N_1908,N_1490,N_1080);
nor U1909 (N_1909,N_518,N_1408);
xnor U1910 (N_1910,N_1373,N_1160);
nand U1911 (N_1911,In_607,N_1345);
nand U1912 (N_1912,In_689,In_1139);
and U1913 (N_1913,N_1092,In_35);
and U1914 (N_1914,N_723,N_447);
or U1915 (N_1915,N_52,N_1191);
and U1916 (N_1916,N_577,N_311);
nor U1917 (N_1917,N_1468,N_666);
nand U1918 (N_1918,N_1304,In_2496);
and U1919 (N_1919,N_1307,N_409);
or U1920 (N_1920,N_169,In_46);
nor U1921 (N_1921,N_1156,N_1251);
xor U1922 (N_1922,N_663,N_323);
or U1923 (N_1923,N_1472,N_1186);
and U1924 (N_1924,N_1204,N_1083);
nor U1925 (N_1925,In_664,N_1022);
and U1926 (N_1926,N_808,N_1212);
nor U1927 (N_1927,N_1206,In_1500);
or U1928 (N_1928,In_830,N_1179);
and U1929 (N_1929,N_1391,In_1387);
and U1930 (N_1930,N_1129,In_1293);
nor U1931 (N_1931,N_851,N_1264);
and U1932 (N_1932,N_1225,In_2293);
and U1933 (N_1933,In_2480,N_1116);
or U1934 (N_1934,N_1147,N_1079);
nor U1935 (N_1935,N_1393,N_712);
and U1936 (N_1936,N_136,N_1386);
nand U1937 (N_1937,In_2283,N_1272);
or U1938 (N_1938,N_437,In_347);
and U1939 (N_1939,N_1178,In_1210);
or U1940 (N_1940,In_115,N_1365);
nor U1941 (N_1941,N_468,N_989);
nor U1942 (N_1942,N_1315,N_1499);
nand U1943 (N_1943,N_1419,N_1018);
and U1944 (N_1944,N_981,N_1396);
or U1945 (N_1945,N_1256,N_1127);
nor U1946 (N_1946,N_1266,N_368);
and U1947 (N_1947,N_444,N_1334);
and U1948 (N_1948,N_1131,N_1203);
or U1949 (N_1949,In_1954,N_832);
or U1950 (N_1950,In_1267,In_1065);
nor U1951 (N_1951,N_1117,In_1747);
nor U1952 (N_1952,N_111,In_1358);
nor U1953 (N_1953,N_1439,N_1350);
nand U1954 (N_1954,N_1031,In_711);
nand U1955 (N_1955,N_652,N_1050);
nor U1956 (N_1956,In_22,N_1058);
and U1957 (N_1957,N_1069,N_862);
nand U1958 (N_1958,N_1114,N_1233);
nand U1959 (N_1959,In_559,In_2219);
nand U1960 (N_1960,N_1165,In_586);
nand U1961 (N_1961,N_371,N_1176);
and U1962 (N_1962,N_667,In_36);
nor U1963 (N_1963,N_383,In_1889);
nor U1964 (N_1964,N_776,In_585);
nor U1965 (N_1965,N_1042,N_889);
nand U1966 (N_1966,N_933,N_420);
nand U1967 (N_1967,N_1294,N_1235);
or U1968 (N_1968,N_1335,In_2205);
nor U1969 (N_1969,N_1381,In_1462);
and U1970 (N_1970,N_190,N_1209);
and U1971 (N_1971,In_975,N_1048);
and U1972 (N_1972,In_577,N_897);
nor U1973 (N_1973,In_715,N_1415);
and U1974 (N_1974,In_243,N_584);
or U1975 (N_1975,N_1286,N_272);
or U1976 (N_1976,N_1400,N_940);
and U1977 (N_1977,N_1158,N_1141);
nand U1978 (N_1978,N_583,In_383);
or U1979 (N_1979,N_1241,In_2202);
and U1980 (N_1980,In_1665,N_1466);
and U1981 (N_1981,N_987,N_1361);
or U1982 (N_1982,N_1174,N_858);
nor U1983 (N_1983,N_1214,In_2370);
nor U1984 (N_1984,N_1193,N_1426);
or U1985 (N_1985,N_1330,In_2121);
nand U1986 (N_1986,N_1357,N_1449);
and U1987 (N_1987,N_1431,N_1112);
nor U1988 (N_1988,N_1007,N_872);
or U1989 (N_1989,N_1075,In_1237);
and U1990 (N_1990,N_1377,N_1107);
nor U1991 (N_1991,N_1194,N_952);
or U1992 (N_1992,N_1245,N_1329);
and U1993 (N_1993,N_1033,In_1137);
nor U1994 (N_1994,N_1476,N_1094);
nor U1995 (N_1995,N_1197,N_792);
nor U1996 (N_1996,In_2012,In_1743);
xor U1997 (N_1997,N_864,N_1346);
nand U1998 (N_1998,N_1025,N_744);
nor U1999 (N_1999,N_1227,N_1498);
and U2000 (N_2000,N_1515,N_1625);
nor U2001 (N_2001,N_1561,N_1681);
nand U2002 (N_2002,N_1851,N_1546);
nor U2003 (N_2003,N_1655,N_1976);
or U2004 (N_2004,N_1646,N_1910);
and U2005 (N_2005,N_1500,N_1771);
nor U2006 (N_2006,N_1652,N_1760);
nor U2007 (N_2007,N_1885,N_1815);
nor U2008 (N_2008,N_1817,N_1977);
nor U2009 (N_2009,N_1841,N_1565);
or U2010 (N_2010,N_1856,N_1537);
and U2011 (N_2011,N_1979,N_1833);
nor U2012 (N_2012,N_1878,N_1837);
nand U2013 (N_2013,N_1677,N_1658);
nor U2014 (N_2014,N_1890,N_1603);
nor U2015 (N_2015,N_1644,N_1587);
and U2016 (N_2016,N_1715,N_1968);
nor U2017 (N_2017,N_1525,N_1987);
and U2018 (N_2018,N_1539,N_1960);
nand U2019 (N_2019,N_1531,N_1673);
nand U2020 (N_2020,N_1674,N_1584);
nor U2021 (N_2021,N_1519,N_1970);
and U2022 (N_2022,N_1688,N_1527);
and U2023 (N_2023,N_1796,N_1710);
nand U2024 (N_2024,N_1764,N_1689);
nor U2025 (N_2025,N_1854,N_1605);
or U2026 (N_2026,N_1941,N_1859);
or U2027 (N_2027,N_1812,N_1575);
nand U2028 (N_2028,N_1819,N_1834);
and U2029 (N_2029,N_1538,N_1744);
nor U2030 (N_2030,N_1807,N_1732);
nor U2031 (N_2031,N_1653,N_1876);
nand U2032 (N_2032,N_1926,N_1782);
and U2033 (N_2033,N_1905,N_1717);
and U2034 (N_2034,N_1591,N_1863);
nor U2035 (N_2035,N_1982,N_1946);
and U2036 (N_2036,N_1684,N_1903);
nor U2037 (N_2037,N_1618,N_1844);
nor U2038 (N_2038,N_1777,N_1708);
nor U2039 (N_2039,N_1639,N_1517);
nand U2040 (N_2040,N_1852,N_1778);
and U2041 (N_2041,N_1745,N_1628);
nand U2042 (N_2042,N_1767,N_1985);
and U2043 (N_2043,N_1925,N_1911);
nor U2044 (N_2044,N_1692,N_1509);
and U2045 (N_2045,N_1614,N_1608);
nor U2046 (N_2046,N_1757,N_1523);
xnor U2047 (N_2047,N_1576,N_1578);
nor U2048 (N_2048,N_1849,N_1973);
nor U2049 (N_2049,N_1897,N_1747);
or U2050 (N_2050,N_1836,N_1709);
nand U2051 (N_2051,N_1786,N_1621);
and U2052 (N_2052,N_1893,N_1814);
nor U2053 (N_2053,N_1555,N_1889);
and U2054 (N_2054,N_1508,N_1549);
nand U2055 (N_2055,N_1753,N_1999);
or U2056 (N_2056,N_1927,N_1759);
nor U2057 (N_2057,N_1702,N_1716);
nand U2058 (N_2058,N_1797,N_1739);
nor U2059 (N_2059,N_1627,N_1540);
nand U2060 (N_2060,N_1723,N_1742);
or U2061 (N_2061,N_1533,N_1630);
or U2062 (N_2062,N_1511,N_1912);
and U2063 (N_2063,N_1522,N_1776);
nor U2064 (N_2064,N_1743,N_1660);
and U2065 (N_2065,N_1866,N_1676);
or U2066 (N_2066,N_1512,N_1920);
or U2067 (N_2067,N_1956,N_1789);
and U2068 (N_2068,N_1507,N_1774);
nand U2069 (N_2069,N_1929,N_1592);
or U2070 (N_2070,N_1953,N_1899);
nor U2071 (N_2071,N_1731,N_1824);
nor U2072 (N_2072,N_1727,N_1867);
nand U2073 (N_2073,N_1637,N_1619);
and U2074 (N_2074,N_1733,N_1762);
nand U2075 (N_2075,N_1884,N_1922);
or U2076 (N_2076,N_1827,N_1808);
or U2077 (N_2077,N_1810,N_1791);
nor U2078 (N_2078,N_1597,N_1700);
nor U2079 (N_2079,N_1823,N_1612);
nand U2080 (N_2080,N_1635,N_1934);
xnor U2081 (N_2081,N_1928,N_1643);
nand U2082 (N_2082,N_1773,N_1853);
or U2083 (N_2083,N_1580,N_1756);
nor U2084 (N_2084,N_1626,N_1736);
and U2085 (N_2085,N_1790,N_1992);
or U2086 (N_2086,N_1931,N_1633);
or U2087 (N_2087,N_1570,N_1919);
and U2088 (N_2088,N_1785,N_1502);
or U2089 (N_2089,N_1556,N_1935);
nand U2090 (N_2090,N_1962,N_1991);
nand U2091 (N_2091,N_1750,N_1940);
or U2092 (N_2092,N_1983,N_1703);
nor U2093 (N_2093,N_1887,N_1942);
nand U2094 (N_2094,N_1847,N_1712);
nand U2095 (N_2095,N_1559,N_1665);
or U2096 (N_2096,N_1908,N_1802);
or U2097 (N_2097,N_1650,N_1959);
nor U2098 (N_2098,N_1954,N_1645);
nand U2099 (N_2099,N_1877,N_1557);
or U2100 (N_2100,N_1938,N_1879);
nand U2101 (N_2101,N_1583,N_1640);
or U2102 (N_2102,N_1800,N_1670);
or U2103 (N_2103,N_1901,N_1861);
or U2104 (N_2104,N_1825,N_1662);
nor U2105 (N_2105,N_1921,N_1696);
xor U2106 (N_2106,N_1683,N_1520);
nand U2107 (N_2107,N_1726,N_1846);
nor U2108 (N_2108,N_1564,N_1839);
or U2109 (N_2109,N_1820,N_1933);
and U2110 (N_2110,N_1634,N_1536);
nor U2111 (N_2111,N_1506,N_1947);
and U2112 (N_2112,N_1661,N_1799);
and U2113 (N_2113,N_1951,N_1704);
xnor U2114 (N_2114,N_1963,N_1737);
nor U2115 (N_2115,N_1687,N_1685);
and U2116 (N_2116,N_1809,N_1813);
or U2117 (N_2117,N_1598,N_1740);
nor U2118 (N_2118,N_1686,N_1532);
nor U2119 (N_2119,N_1524,N_1943);
and U2120 (N_2120,N_1986,N_1895);
nor U2121 (N_2121,N_1599,N_1569);
and U2122 (N_2122,N_1838,N_1504);
or U2123 (N_2123,N_1832,N_1923);
nor U2124 (N_2124,N_1600,N_1924);
nor U2125 (N_2125,N_1930,N_1850);
xnor U2126 (N_2126,N_1858,N_1748);
and U2127 (N_2127,N_1896,N_1794);
nor U2128 (N_2128,N_1892,N_1752);
nor U2129 (N_2129,N_1544,N_1535);
and U2130 (N_2130,N_1988,N_1651);
nand U2131 (N_2131,N_1718,N_1705);
nand U2132 (N_2132,N_1937,N_1840);
and U2133 (N_2133,N_1965,N_1811);
nand U2134 (N_2134,N_1521,N_1730);
nor U2135 (N_2135,N_1711,N_1554);
nand U2136 (N_2136,N_1870,N_1695);
or U2137 (N_2137,N_1843,N_1969);
xor U2138 (N_2138,N_1596,N_1957);
nor U2139 (N_2139,N_1678,N_1551);
and U2140 (N_2140,N_1784,N_1798);
and U2141 (N_2141,N_1936,N_1697);
nor U2142 (N_2142,N_1528,N_1952);
nand U2143 (N_2143,N_1542,N_1898);
nor U2144 (N_2144,N_1914,N_1913);
or U2145 (N_2145,N_1585,N_1775);
nand U2146 (N_2146,N_1981,N_1666);
or U2147 (N_2147,N_1588,N_1735);
nand U2148 (N_2148,N_1829,N_1980);
nand U2149 (N_2149,N_1719,N_1579);
nand U2150 (N_2150,N_1706,N_1505);
xnor U2151 (N_2151,N_1624,N_1803);
and U2152 (N_2152,N_1958,N_1616);
and U2153 (N_2153,N_1868,N_1615);
or U2154 (N_2154,N_1516,N_1875);
and U2155 (N_2155,N_1606,N_1882);
and U2156 (N_2156,N_1806,N_1869);
nand U2157 (N_2157,N_1904,N_1560);
and U2158 (N_2158,N_1932,N_1978);
nand U2159 (N_2159,N_1558,N_1553);
nor U2160 (N_2160,N_1656,N_1530);
nor U2161 (N_2161,N_1566,N_1996);
or U2162 (N_2162,N_1694,N_1667);
nor U2163 (N_2163,N_1581,N_1971);
nand U2164 (N_2164,N_1779,N_1550);
and U2165 (N_2165,N_1792,N_1826);
nand U2166 (N_2166,N_1769,N_1984);
nand U2167 (N_2167,N_1573,N_1816);
nor U2168 (N_2168,N_1891,N_1801);
or U2169 (N_2169,N_1623,N_1543);
nand U2170 (N_2170,N_1765,N_1842);
and U2171 (N_2171,N_1641,N_1602);
or U2172 (N_2172,N_1620,N_1669);
nand U2173 (N_2173,N_1648,N_1572);
and U2174 (N_2174,N_1755,N_1691);
and U2175 (N_2175,N_1995,N_1944);
nand U2176 (N_2176,N_1874,N_1793);
or U2177 (N_2177,N_1741,N_1763);
nand U2178 (N_2178,N_1865,N_1541);
nand U2179 (N_2179,N_1664,N_1918);
nor U2180 (N_2180,N_1994,N_1534);
xnor U2181 (N_2181,N_1967,N_1857);
and U2182 (N_2182,N_1754,N_1698);
and U2183 (N_2183,N_1781,N_1855);
or U2184 (N_2184,N_1894,N_1835);
or U2185 (N_2185,N_1631,N_1900);
or U2186 (N_2186,N_1780,N_1993);
nand U2187 (N_2187,N_1513,N_1582);
nor U2188 (N_2188,N_1610,N_1638);
nand U2189 (N_2189,N_1647,N_1873);
and U2190 (N_2190,N_1848,N_1595);
nor U2191 (N_2191,N_1872,N_1975);
nand U2192 (N_2192,N_1888,N_1883);
nand U2193 (N_2193,N_1663,N_1768);
and U2194 (N_2194,N_1672,N_1998);
or U2195 (N_2195,N_1804,N_1636);
nor U2196 (N_2196,N_1679,N_1675);
nor U2197 (N_2197,N_1568,N_1787);
or U2198 (N_2198,N_1964,N_1734);
nor U2199 (N_2199,N_1728,N_1654);
nand U2200 (N_2200,N_1722,N_1671);
or U2201 (N_2201,N_1862,N_1552);
and U2202 (N_2202,N_1713,N_1966);
and U2203 (N_2203,N_1701,N_1590);
and U2204 (N_2204,N_1860,N_1818);
or U2205 (N_2205,N_1707,N_1529);
xnor U2206 (N_2206,N_1830,N_1822);
or U2207 (N_2207,N_1906,N_1586);
nor U2208 (N_2208,N_1939,N_1788);
and U2209 (N_2209,N_1567,N_1749);
nand U2210 (N_2210,N_1761,N_1772);
and U2211 (N_2211,N_1563,N_1547);
nand U2212 (N_2212,N_1548,N_1622);
nor U2213 (N_2213,N_1725,N_1668);
nand U2214 (N_2214,N_1501,N_1657);
nor U2215 (N_2215,N_1972,N_1693);
or U2216 (N_2216,N_1770,N_1907);
nor U2217 (N_2217,N_1997,N_1649);
or U2218 (N_2218,N_1659,N_1989);
nor U2219 (N_2219,N_1699,N_1514);
nor U2220 (N_2220,N_1738,N_1594);
and U2221 (N_2221,N_1974,N_1593);
nor U2222 (N_2222,N_1682,N_1950);
nor U2223 (N_2223,N_1629,N_1909);
and U2224 (N_2224,N_1917,N_1915);
or U2225 (N_2225,N_1613,N_1571);
or U2226 (N_2226,N_1945,N_1611);
xor U2227 (N_2227,N_1783,N_1751);
nand U2228 (N_2228,N_1721,N_1729);
nor U2229 (N_2229,N_1990,N_1845);
and U2230 (N_2230,N_1805,N_1881);
nand U2231 (N_2231,N_1574,N_1545);
or U2232 (N_2232,N_1766,N_1577);
nor U2233 (N_2233,N_1503,N_1871);
and U2234 (N_2234,N_1526,N_1632);
and U2235 (N_2235,N_1916,N_1831);
and U2236 (N_2236,N_1961,N_1902);
and U2237 (N_2237,N_1680,N_1720);
nand U2238 (N_2238,N_1758,N_1518);
or U2239 (N_2239,N_1724,N_1880);
nand U2240 (N_2240,N_1886,N_1949);
and U2241 (N_2241,N_1562,N_1604);
nand U2242 (N_2242,N_1955,N_1609);
and U2243 (N_2243,N_1795,N_1642);
nand U2244 (N_2244,N_1510,N_1607);
nand U2245 (N_2245,N_1948,N_1821);
nor U2246 (N_2246,N_1714,N_1601);
and U2247 (N_2247,N_1864,N_1690);
nand U2248 (N_2248,N_1617,N_1589);
nor U2249 (N_2249,N_1746,N_1828);
or U2250 (N_2250,N_1537,N_1683);
and U2251 (N_2251,N_1877,N_1941);
nand U2252 (N_2252,N_1550,N_1807);
or U2253 (N_2253,N_1960,N_1584);
or U2254 (N_2254,N_1917,N_1593);
nand U2255 (N_2255,N_1849,N_1999);
or U2256 (N_2256,N_1750,N_1515);
and U2257 (N_2257,N_1585,N_1991);
and U2258 (N_2258,N_1560,N_1980);
nor U2259 (N_2259,N_1876,N_1979);
and U2260 (N_2260,N_1582,N_1969);
nor U2261 (N_2261,N_1884,N_1902);
and U2262 (N_2262,N_1903,N_1638);
nor U2263 (N_2263,N_1650,N_1971);
nand U2264 (N_2264,N_1668,N_1720);
or U2265 (N_2265,N_1588,N_1833);
or U2266 (N_2266,N_1889,N_1732);
nand U2267 (N_2267,N_1621,N_1805);
and U2268 (N_2268,N_1596,N_1903);
and U2269 (N_2269,N_1606,N_1663);
and U2270 (N_2270,N_1674,N_1921);
nor U2271 (N_2271,N_1701,N_1779);
or U2272 (N_2272,N_1923,N_1620);
nand U2273 (N_2273,N_1990,N_1933);
nand U2274 (N_2274,N_1837,N_1890);
nand U2275 (N_2275,N_1704,N_1917);
and U2276 (N_2276,N_1547,N_1543);
nor U2277 (N_2277,N_1962,N_1595);
or U2278 (N_2278,N_1694,N_1576);
nand U2279 (N_2279,N_1573,N_1552);
xnor U2280 (N_2280,N_1962,N_1531);
or U2281 (N_2281,N_1886,N_1659);
or U2282 (N_2282,N_1913,N_1824);
or U2283 (N_2283,N_1577,N_1659);
or U2284 (N_2284,N_1999,N_1875);
nor U2285 (N_2285,N_1763,N_1533);
or U2286 (N_2286,N_1775,N_1833);
and U2287 (N_2287,N_1850,N_1973);
or U2288 (N_2288,N_1860,N_1628);
nand U2289 (N_2289,N_1618,N_1624);
nand U2290 (N_2290,N_1549,N_1978);
and U2291 (N_2291,N_1853,N_1744);
or U2292 (N_2292,N_1929,N_1875);
nor U2293 (N_2293,N_1521,N_1778);
and U2294 (N_2294,N_1934,N_1590);
nor U2295 (N_2295,N_1874,N_1829);
or U2296 (N_2296,N_1903,N_1715);
nand U2297 (N_2297,N_1757,N_1537);
xnor U2298 (N_2298,N_1704,N_1875);
or U2299 (N_2299,N_1545,N_1749);
or U2300 (N_2300,N_1819,N_1917);
and U2301 (N_2301,N_1621,N_1888);
and U2302 (N_2302,N_1743,N_1893);
nor U2303 (N_2303,N_1888,N_1720);
and U2304 (N_2304,N_1833,N_1888);
and U2305 (N_2305,N_1722,N_1533);
nand U2306 (N_2306,N_1559,N_1942);
and U2307 (N_2307,N_1611,N_1995);
nor U2308 (N_2308,N_1935,N_1973);
nand U2309 (N_2309,N_1547,N_1631);
nor U2310 (N_2310,N_1582,N_1583);
or U2311 (N_2311,N_1958,N_1576);
or U2312 (N_2312,N_1589,N_1527);
nor U2313 (N_2313,N_1993,N_1844);
or U2314 (N_2314,N_1705,N_1548);
nand U2315 (N_2315,N_1846,N_1518);
nor U2316 (N_2316,N_1656,N_1983);
or U2317 (N_2317,N_1844,N_1990);
or U2318 (N_2318,N_1696,N_1854);
or U2319 (N_2319,N_1821,N_1844);
nand U2320 (N_2320,N_1581,N_1769);
and U2321 (N_2321,N_1579,N_1901);
nor U2322 (N_2322,N_1567,N_1965);
nor U2323 (N_2323,N_1741,N_1695);
and U2324 (N_2324,N_1758,N_1733);
nor U2325 (N_2325,N_1618,N_1801);
or U2326 (N_2326,N_1778,N_1685);
or U2327 (N_2327,N_1513,N_1870);
nor U2328 (N_2328,N_1777,N_1949);
nand U2329 (N_2329,N_1825,N_1638);
nand U2330 (N_2330,N_1557,N_1749);
nor U2331 (N_2331,N_1718,N_1695);
nor U2332 (N_2332,N_1658,N_1755);
and U2333 (N_2333,N_1562,N_1610);
nor U2334 (N_2334,N_1753,N_1673);
and U2335 (N_2335,N_1998,N_1745);
nor U2336 (N_2336,N_1809,N_1920);
and U2337 (N_2337,N_1736,N_1968);
nand U2338 (N_2338,N_1940,N_1622);
nor U2339 (N_2339,N_1717,N_1659);
or U2340 (N_2340,N_1553,N_1515);
or U2341 (N_2341,N_1952,N_1612);
and U2342 (N_2342,N_1710,N_1681);
or U2343 (N_2343,N_1886,N_1752);
nand U2344 (N_2344,N_1616,N_1570);
or U2345 (N_2345,N_1532,N_1521);
nor U2346 (N_2346,N_1963,N_1513);
or U2347 (N_2347,N_1595,N_1741);
and U2348 (N_2348,N_1886,N_1830);
or U2349 (N_2349,N_1513,N_1923);
xor U2350 (N_2350,N_1886,N_1981);
nand U2351 (N_2351,N_1926,N_1600);
nor U2352 (N_2352,N_1594,N_1946);
nand U2353 (N_2353,N_1994,N_1619);
or U2354 (N_2354,N_1764,N_1532);
nor U2355 (N_2355,N_1804,N_1875);
nand U2356 (N_2356,N_1943,N_1701);
and U2357 (N_2357,N_1976,N_1576);
nor U2358 (N_2358,N_1759,N_1675);
and U2359 (N_2359,N_1618,N_1625);
nand U2360 (N_2360,N_1947,N_1580);
nor U2361 (N_2361,N_1893,N_1596);
nand U2362 (N_2362,N_1854,N_1693);
and U2363 (N_2363,N_1751,N_1862);
nand U2364 (N_2364,N_1604,N_1623);
nand U2365 (N_2365,N_1895,N_1612);
nand U2366 (N_2366,N_1742,N_1612);
nor U2367 (N_2367,N_1669,N_1914);
nor U2368 (N_2368,N_1624,N_1982);
nor U2369 (N_2369,N_1743,N_1776);
or U2370 (N_2370,N_1996,N_1976);
and U2371 (N_2371,N_1724,N_1646);
and U2372 (N_2372,N_1674,N_1899);
nor U2373 (N_2373,N_1818,N_1663);
or U2374 (N_2374,N_1819,N_1951);
and U2375 (N_2375,N_1516,N_1606);
and U2376 (N_2376,N_1886,N_1892);
and U2377 (N_2377,N_1943,N_1541);
nor U2378 (N_2378,N_1795,N_1682);
xnor U2379 (N_2379,N_1949,N_1841);
nand U2380 (N_2380,N_1569,N_1807);
or U2381 (N_2381,N_1651,N_1942);
and U2382 (N_2382,N_1871,N_1508);
nor U2383 (N_2383,N_1741,N_1532);
or U2384 (N_2384,N_1838,N_1637);
or U2385 (N_2385,N_1743,N_1636);
nand U2386 (N_2386,N_1623,N_1827);
and U2387 (N_2387,N_1840,N_1656);
nand U2388 (N_2388,N_1742,N_1682);
nand U2389 (N_2389,N_1566,N_1764);
nand U2390 (N_2390,N_1520,N_1579);
xor U2391 (N_2391,N_1529,N_1652);
or U2392 (N_2392,N_1986,N_1564);
and U2393 (N_2393,N_1943,N_1818);
nand U2394 (N_2394,N_1845,N_1873);
nor U2395 (N_2395,N_1559,N_1733);
nand U2396 (N_2396,N_1806,N_1606);
nand U2397 (N_2397,N_1958,N_1774);
nand U2398 (N_2398,N_1541,N_1736);
and U2399 (N_2399,N_1968,N_1899);
or U2400 (N_2400,N_1637,N_1693);
xnor U2401 (N_2401,N_1952,N_1692);
or U2402 (N_2402,N_1769,N_1820);
or U2403 (N_2403,N_1828,N_1585);
and U2404 (N_2404,N_1605,N_1901);
or U2405 (N_2405,N_1947,N_1794);
nand U2406 (N_2406,N_1605,N_1921);
nand U2407 (N_2407,N_1656,N_1881);
and U2408 (N_2408,N_1848,N_1741);
or U2409 (N_2409,N_1532,N_1877);
nand U2410 (N_2410,N_1882,N_1632);
and U2411 (N_2411,N_1624,N_1605);
or U2412 (N_2412,N_1763,N_1773);
nand U2413 (N_2413,N_1613,N_1762);
nand U2414 (N_2414,N_1578,N_1501);
nor U2415 (N_2415,N_1759,N_1920);
nor U2416 (N_2416,N_1966,N_1736);
and U2417 (N_2417,N_1510,N_1719);
nand U2418 (N_2418,N_1568,N_1504);
and U2419 (N_2419,N_1899,N_1881);
nand U2420 (N_2420,N_1926,N_1591);
or U2421 (N_2421,N_1605,N_1729);
and U2422 (N_2422,N_1798,N_1928);
nor U2423 (N_2423,N_1914,N_1873);
and U2424 (N_2424,N_1743,N_1915);
or U2425 (N_2425,N_1607,N_1504);
and U2426 (N_2426,N_1794,N_1659);
nor U2427 (N_2427,N_1752,N_1707);
or U2428 (N_2428,N_1755,N_1574);
nor U2429 (N_2429,N_1641,N_1576);
or U2430 (N_2430,N_1724,N_1961);
and U2431 (N_2431,N_1602,N_1998);
and U2432 (N_2432,N_1722,N_1931);
or U2433 (N_2433,N_1798,N_1516);
nand U2434 (N_2434,N_1944,N_1595);
and U2435 (N_2435,N_1986,N_1559);
or U2436 (N_2436,N_1541,N_1503);
or U2437 (N_2437,N_1816,N_1681);
nor U2438 (N_2438,N_1881,N_1770);
and U2439 (N_2439,N_1501,N_1734);
nand U2440 (N_2440,N_1572,N_1850);
nor U2441 (N_2441,N_1859,N_1977);
nand U2442 (N_2442,N_1994,N_1848);
and U2443 (N_2443,N_1721,N_1686);
and U2444 (N_2444,N_1734,N_1507);
nor U2445 (N_2445,N_1675,N_1686);
nor U2446 (N_2446,N_1931,N_1576);
nor U2447 (N_2447,N_1954,N_1605);
nor U2448 (N_2448,N_1948,N_1825);
and U2449 (N_2449,N_1852,N_1981);
or U2450 (N_2450,N_1716,N_1749);
nor U2451 (N_2451,N_1803,N_1981);
or U2452 (N_2452,N_1613,N_1977);
xnor U2453 (N_2453,N_1898,N_1648);
and U2454 (N_2454,N_1878,N_1661);
nor U2455 (N_2455,N_1708,N_1762);
nor U2456 (N_2456,N_1890,N_1554);
nor U2457 (N_2457,N_1743,N_1549);
and U2458 (N_2458,N_1561,N_1821);
nand U2459 (N_2459,N_1945,N_1573);
and U2460 (N_2460,N_1652,N_1903);
and U2461 (N_2461,N_1813,N_1598);
nand U2462 (N_2462,N_1604,N_1542);
or U2463 (N_2463,N_1579,N_1671);
and U2464 (N_2464,N_1603,N_1907);
or U2465 (N_2465,N_1658,N_1874);
nand U2466 (N_2466,N_1623,N_1796);
or U2467 (N_2467,N_1560,N_1656);
nand U2468 (N_2468,N_1950,N_1573);
nor U2469 (N_2469,N_1764,N_1907);
and U2470 (N_2470,N_1715,N_1518);
nand U2471 (N_2471,N_1940,N_1509);
and U2472 (N_2472,N_1795,N_1513);
nand U2473 (N_2473,N_1525,N_1794);
and U2474 (N_2474,N_1983,N_1852);
and U2475 (N_2475,N_1542,N_1581);
nand U2476 (N_2476,N_1844,N_1675);
and U2477 (N_2477,N_1573,N_1988);
xor U2478 (N_2478,N_1987,N_1759);
nor U2479 (N_2479,N_1930,N_1958);
or U2480 (N_2480,N_1925,N_1626);
nor U2481 (N_2481,N_1586,N_1830);
and U2482 (N_2482,N_1720,N_1677);
nor U2483 (N_2483,N_1505,N_1924);
and U2484 (N_2484,N_1741,N_1938);
and U2485 (N_2485,N_1675,N_1649);
nand U2486 (N_2486,N_1537,N_1988);
nor U2487 (N_2487,N_1708,N_1686);
nor U2488 (N_2488,N_1785,N_1851);
and U2489 (N_2489,N_1997,N_1868);
nor U2490 (N_2490,N_1885,N_1846);
nand U2491 (N_2491,N_1823,N_1967);
nor U2492 (N_2492,N_1503,N_1548);
or U2493 (N_2493,N_1782,N_1788);
nand U2494 (N_2494,N_1685,N_1518);
xor U2495 (N_2495,N_1565,N_1599);
nand U2496 (N_2496,N_1757,N_1545);
nor U2497 (N_2497,N_1649,N_1927);
or U2498 (N_2498,N_1526,N_1651);
or U2499 (N_2499,N_1969,N_1739);
or U2500 (N_2500,N_2165,N_2335);
nor U2501 (N_2501,N_2462,N_2179);
and U2502 (N_2502,N_2433,N_2065);
nor U2503 (N_2503,N_2375,N_2098);
nor U2504 (N_2504,N_2155,N_2312);
and U2505 (N_2505,N_2429,N_2002);
or U2506 (N_2506,N_2170,N_2351);
nor U2507 (N_2507,N_2217,N_2446);
or U2508 (N_2508,N_2035,N_2085);
nor U2509 (N_2509,N_2323,N_2099);
and U2510 (N_2510,N_2338,N_2075);
nand U2511 (N_2511,N_2344,N_2223);
and U2512 (N_2512,N_2396,N_2040);
or U2513 (N_2513,N_2291,N_2203);
nand U2514 (N_2514,N_2271,N_2381);
nand U2515 (N_2515,N_2314,N_2473);
nand U2516 (N_2516,N_2192,N_2359);
nor U2517 (N_2517,N_2290,N_2043);
and U2518 (N_2518,N_2215,N_2311);
nand U2519 (N_2519,N_2218,N_2293);
and U2520 (N_2520,N_2250,N_2464);
xor U2521 (N_2521,N_2106,N_2425);
or U2522 (N_2522,N_2116,N_2133);
nand U2523 (N_2523,N_2339,N_2229);
nand U2524 (N_2524,N_2354,N_2317);
or U2525 (N_2525,N_2048,N_2360);
nor U2526 (N_2526,N_2493,N_2350);
or U2527 (N_2527,N_2292,N_2301);
and U2528 (N_2528,N_2104,N_2006);
and U2529 (N_2529,N_2141,N_2492);
or U2530 (N_2530,N_2295,N_2285);
nor U2531 (N_2531,N_2255,N_2274);
and U2532 (N_2532,N_2091,N_2368);
or U2533 (N_2533,N_2448,N_2276);
nor U2534 (N_2534,N_2157,N_2431);
nand U2535 (N_2535,N_2299,N_2022);
xor U2536 (N_2536,N_2406,N_2036);
nor U2537 (N_2537,N_2298,N_2168);
or U2538 (N_2538,N_2222,N_2069);
or U2539 (N_2539,N_2162,N_2310);
and U2540 (N_2540,N_2054,N_2173);
nand U2541 (N_2541,N_2348,N_2485);
nand U2542 (N_2542,N_2171,N_2051);
or U2543 (N_2543,N_2181,N_2233);
or U2544 (N_2544,N_2038,N_2214);
and U2545 (N_2545,N_2352,N_2023);
xor U2546 (N_2546,N_2014,N_2343);
nor U2547 (N_2547,N_2392,N_2417);
nand U2548 (N_2548,N_2187,N_2019);
nor U2549 (N_2549,N_2001,N_2449);
and U2550 (N_2550,N_2264,N_2411);
or U2551 (N_2551,N_2282,N_2435);
nor U2552 (N_2552,N_2163,N_2126);
nand U2553 (N_2553,N_2076,N_2458);
nor U2554 (N_2554,N_2196,N_2058);
nand U2555 (N_2555,N_2231,N_2367);
nor U2556 (N_2556,N_2101,N_2119);
nand U2557 (N_2557,N_2167,N_2062);
and U2558 (N_2558,N_2305,N_2444);
and U2559 (N_2559,N_2018,N_2258);
nand U2560 (N_2560,N_2487,N_2379);
and U2561 (N_2561,N_2150,N_2269);
or U2562 (N_2562,N_2390,N_2287);
and U2563 (N_2563,N_2248,N_2220);
and U2564 (N_2564,N_2304,N_2486);
nor U2565 (N_2565,N_2089,N_2064);
or U2566 (N_2566,N_2245,N_2188);
nor U2567 (N_2567,N_2052,N_2407);
nor U2568 (N_2568,N_2147,N_2034);
or U2569 (N_2569,N_2041,N_2373);
or U2570 (N_2570,N_2415,N_2465);
or U2571 (N_2571,N_2260,N_2160);
and U2572 (N_2572,N_2388,N_2357);
or U2573 (N_2573,N_2088,N_2049);
and U2574 (N_2574,N_2183,N_2194);
or U2575 (N_2575,N_2427,N_2240);
nor U2576 (N_2576,N_2084,N_2327);
and U2577 (N_2577,N_2494,N_2152);
and U2578 (N_2578,N_2056,N_2334);
nor U2579 (N_2579,N_2208,N_2073);
and U2580 (N_2580,N_2130,N_2166);
nand U2581 (N_2581,N_2237,N_2221);
nand U2582 (N_2582,N_2008,N_2438);
nand U2583 (N_2583,N_2137,N_2477);
or U2584 (N_2584,N_2238,N_2140);
or U2585 (N_2585,N_2322,N_2093);
nor U2586 (N_2586,N_2016,N_2441);
and U2587 (N_2587,N_2185,N_2262);
nand U2588 (N_2588,N_2450,N_2083);
nor U2589 (N_2589,N_2309,N_2315);
or U2590 (N_2590,N_2398,N_2384);
and U2591 (N_2591,N_2371,N_2046);
nand U2592 (N_2592,N_2151,N_2060);
nor U2593 (N_2593,N_2055,N_2186);
or U2594 (N_2594,N_2000,N_2125);
and U2595 (N_2595,N_2200,N_2112);
and U2596 (N_2596,N_2161,N_2190);
nor U2597 (N_2597,N_2419,N_2401);
nor U2598 (N_2598,N_2294,N_2275);
or U2599 (N_2599,N_2436,N_2078);
nor U2600 (N_2600,N_2347,N_2471);
nand U2601 (N_2601,N_2103,N_2337);
or U2602 (N_2602,N_2109,N_2189);
and U2603 (N_2603,N_2184,N_2176);
or U2604 (N_2604,N_2121,N_2489);
nor U2605 (N_2605,N_2482,N_2479);
nor U2606 (N_2606,N_2329,N_2445);
or U2607 (N_2607,N_2107,N_2086);
or U2608 (N_2608,N_2077,N_2164);
or U2609 (N_2609,N_2118,N_2281);
nor U2610 (N_2610,N_2355,N_2136);
nand U2611 (N_2611,N_2267,N_2191);
nand U2612 (N_2612,N_2251,N_2097);
and U2613 (N_2613,N_2270,N_2346);
nand U2614 (N_2614,N_2306,N_2113);
xnor U2615 (N_2615,N_2363,N_2122);
nor U2616 (N_2616,N_2138,N_2135);
and U2617 (N_2617,N_2483,N_2402);
nand U2618 (N_2618,N_2059,N_2497);
nand U2619 (N_2619,N_2100,N_2132);
nor U2620 (N_2620,N_2128,N_2365);
or U2621 (N_2621,N_2047,N_2289);
nor U2622 (N_2622,N_2480,N_2143);
or U2623 (N_2623,N_2239,N_2385);
and U2624 (N_2624,N_2094,N_2488);
nand U2625 (N_2625,N_2228,N_2131);
or U2626 (N_2626,N_2403,N_2030);
nor U2627 (N_2627,N_2111,N_2453);
and U2628 (N_2628,N_2216,N_2028);
nor U2629 (N_2629,N_2272,N_2263);
nand U2630 (N_2630,N_2284,N_2484);
nand U2631 (N_2631,N_2230,N_2108);
nor U2632 (N_2632,N_2358,N_2080);
nand U2633 (N_2633,N_2297,N_2300);
nand U2634 (N_2634,N_2349,N_2095);
nor U2635 (N_2635,N_2026,N_2376);
or U2636 (N_2636,N_2235,N_2345);
nand U2637 (N_2637,N_2273,N_2495);
and U2638 (N_2638,N_2268,N_2090);
nor U2639 (N_2639,N_2257,N_2017);
nor U2640 (N_2640,N_2400,N_2209);
and U2641 (N_2641,N_2279,N_2259);
or U2642 (N_2642,N_2120,N_2256);
nor U2643 (N_2643,N_2197,N_2288);
nand U2644 (N_2644,N_2456,N_2387);
or U2645 (N_2645,N_2244,N_2336);
or U2646 (N_2646,N_2474,N_2283);
or U2647 (N_2647,N_2148,N_2124);
nand U2648 (N_2648,N_2443,N_2333);
or U2649 (N_2649,N_2020,N_2081);
and U2650 (N_2650,N_2468,N_2455);
or U2651 (N_2651,N_2249,N_2174);
nand U2652 (N_2652,N_2280,N_2423);
nand U2653 (N_2653,N_2286,N_2370);
and U2654 (N_2654,N_2204,N_2442);
nor U2655 (N_2655,N_2012,N_2405);
and U2656 (N_2656,N_2408,N_2416);
nor U2657 (N_2657,N_2071,N_2011);
and U2658 (N_2658,N_2117,N_2478);
nand U2659 (N_2659,N_2045,N_2127);
and U2660 (N_2660,N_2394,N_2198);
nand U2661 (N_2661,N_2154,N_2397);
or U2662 (N_2662,N_2361,N_2341);
nor U2663 (N_2663,N_2496,N_2180);
nor U2664 (N_2664,N_2374,N_2451);
and U2665 (N_2665,N_2261,N_2469);
nand U2666 (N_2666,N_2470,N_2007);
or U2667 (N_2667,N_2153,N_2457);
or U2668 (N_2668,N_2211,N_2421);
nor U2669 (N_2669,N_2378,N_2145);
nand U2670 (N_2670,N_2102,N_2205);
or U2671 (N_2671,N_2364,N_2362);
nor U2672 (N_2672,N_2342,N_2226);
and U2673 (N_2673,N_2061,N_2475);
and U2674 (N_2674,N_2463,N_2372);
nor U2675 (N_2675,N_2383,N_2236);
and U2676 (N_2676,N_2472,N_2193);
nand U2677 (N_2677,N_2243,N_2439);
or U2678 (N_2678,N_2146,N_2032);
nor U2679 (N_2679,N_2206,N_2074);
or U2680 (N_2680,N_2201,N_2325);
or U2681 (N_2681,N_2027,N_2393);
nand U2682 (N_2682,N_2447,N_2159);
or U2683 (N_2683,N_2498,N_2009);
xor U2684 (N_2684,N_2420,N_2114);
nand U2685 (N_2685,N_2178,N_2144);
nor U2686 (N_2686,N_2015,N_2067);
or U2687 (N_2687,N_2210,N_2066);
or U2688 (N_2688,N_2324,N_2366);
or U2689 (N_2689,N_2404,N_2319);
or U2690 (N_2690,N_2182,N_2328);
nand U2691 (N_2691,N_2434,N_2021);
and U2692 (N_2692,N_2332,N_2195);
and U2693 (N_2693,N_2172,N_2050);
nor U2694 (N_2694,N_2321,N_2278);
and U2695 (N_2695,N_2252,N_2013);
nor U2696 (N_2696,N_2242,N_2369);
or U2697 (N_2697,N_2105,N_2440);
or U2698 (N_2698,N_2079,N_2010);
and U2699 (N_2699,N_2156,N_2481);
and U2700 (N_2700,N_2005,N_2031);
nor U2701 (N_2701,N_2042,N_2207);
and U2702 (N_2702,N_2296,N_2377);
nor U2703 (N_2703,N_2072,N_2414);
and U2704 (N_2704,N_2382,N_2142);
nand U2705 (N_2705,N_2212,N_2320);
nor U2706 (N_2706,N_2491,N_2063);
nor U2707 (N_2707,N_2307,N_2330);
nand U2708 (N_2708,N_2318,N_2467);
nor U2709 (N_2709,N_2277,N_2302);
or U2710 (N_2710,N_2308,N_2432);
nand U2711 (N_2711,N_2424,N_2039);
or U2712 (N_2712,N_2158,N_2202);
and U2713 (N_2713,N_2460,N_2004);
nor U2714 (N_2714,N_2316,N_2123);
nor U2715 (N_2715,N_2037,N_2082);
and U2716 (N_2716,N_2254,N_2070);
or U2717 (N_2717,N_2428,N_2227);
nor U2718 (N_2718,N_2380,N_2092);
and U2719 (N_2719,N_2356,N_2331);
or U2720 (N_2720,N_2115,N_2025);
nand U2721 (N_2721,N_2461,N_2303);
nor U2722 (N_2722,N_2024,N_2234);
nand U2723 (N_2723,N_2241,N_2175);
or U2724 (N_2724,N_2232,N_2437);
and U2725 (N_2725,N_2246,N_2033);
and U2726 (N_2726,N_2454,N_2213);
nor U2727 (N_2727,N_2110,N_2499);
or U2728 (N_2728,N_2057,N_2044);
nor U2729 (N_2729,N_2265,N_2422);
or U2730 (N_2730,N_2068,N_2219);
nand U2731 (N_2731,N_2413,N_2253);
or U2732 (N_2732,N_2096,N_2386);
nand U2733 (N_2733,N_2129,N_2169);
nor U2734 (N_2734,N_2389,N_2029);
nand U2735 (N_2735,N_2326,N_2452);
or U2736 (N_2736,N_2412,N_2466);
xor U2737 (N_2737,N_2459,N_2225);
and U2738 (N_2738,N_2224,N_2395);
and U2739 (N_2739,N_2340,N_2410);
nor U2740 (N_2740,N_2418,N_2409);
nand U2741 (N_2741,N_2313,N_2139);
xor U2742 (N_2742,N_2430,N_2391);
nor U2743 (N_2743,N_2199,N_2003);
nand U2744 (N_2744,N_2490,N_2177);
nand U2745 (N_2745,N_2476,N_2053);
nand U2746 (N_2746,N_2266,N_2247);
xnor U2747 (N_2747,N_2353,N_2426);
nor U2748 (N_2748,N_2149,N_2134);
nand U2749 (N_2749,N_2399,N_2087);
and U2750 (N_2750,N_2092,N_2220);
or U2751 (N_2751,N_2353,N_2107);
nand U2752 (N_2752,N_2209,N_2342);
or U2753 (N_2753,N_2043,N_2086);
and U2754 (N_2754,N_2422,N_2104);
or U2755 (N_2755,N_2040,N_2053);
or U2756 (N_2756,N_2136,N_2278);
or U2757 (N_2757,N_2456,N_2463);
nor U2758 (N_2758,N_2301,N_2131);
nor U2759 (N_2759,N_2311,N_2493);
and U2760 (N_2760,N_2320,N_2203);
and U2761 (N_2761,N_2010,N_2186);
nand U2762 (N_2762,N_2065,N_2365);
or U2763 (N_2763,N_2184,N_2277);
nor U2764 (N_2764,N_2283,N_2207);
nand U2765 (N_2765,N_2478,N_2057);
and U2766 (N_2766,N_2351,N_2302);
or U2767 (N_2767,N_2023,N_2165);
or U2768 (N_2768,N_2414,N_2485);
or U2769 (N_2769,N_2269,N_2138);
or U2770 (N_2770,N_2366,N_2290);
nand U2771 (N_2771,N_2318,N_2371);
nor U2772 (N_2772,N_2101,N_2153);
nand U2773 (N_2773,N_2232,N_2466);
nand U2774 (N_2774,N_2088,N_2109);
xor U2775 (N_2775,N_2133,N_2207);
nor U2776 (N_2776,N_2069,N_2358);
nor U2777 (N_2777,N_2084,N_2301);
or U2778 (N_2778,N_2289,N_2251);
nand U2779 (N_2779,N_2260,N_2453);
nor U2780 (N_2780,N_2216,N_2365);
or U2781 (N_2781,N_2378,N_2498);
and U2782 (N_2782,N_2194,N_2099);
nand U2783 (N_2783,N_2323,N_2113);
and U2784 (N_2784,N_2381,N_2031);
nor U2785 (N_2785,N_2133,N_2473);
nor U2786 (N_2786,N_2390,N_2286);
and U2787 (N_2787,N_2149,N_2493);
or U2788 (N_2788,N_2135,N_2355);
or U2789 (N_2789,N_2066,N_2376);
nor U2790 (N_2790,N_2064,N_2049);
nand U2791 (N_2791,N_2042,N_2005);
nor U2792 (N_2792,N_2116,N_2375);
nand U2793 (N_2793,N_2108,N_2354);
xnor U2794 (N_2794,N_2051,N_2429);
and U2795 (N_2795,N_2245,N_2358);
nor U2796 (N_2796,N_2022,N_2353);
nand U2797 (N_2797,N_2115,N_2244);
nand U2798 (N_2798,N_2348,N_2327);
nor U2799 (N_2799,N_2332,N_2461);
nor U2800 (N_2800,N_2198,N_2281);
and U2801 (N_2801,N_2259,N_2397);
or U2802 (N_2802,N_2232,N_2216);
nand U2803 (N_2803,N_2024,N_2209);
or U2804 (N_2804,N_2282,N_2462);
or U2805 (N_2805,N_2131,N_2166);
and U2806 (N_2806,N_2026,N_2161);
and U2807 (N_2807,N_2332,N_2000);
nand U2808 (N_2808,N_2444,N_2175);
or U2809 (N_2809,N_2063,N_2081);
nand U2810 (N_2810,N_2004,N_2356);
or U2811 (N_2811,N_2377,N_2495);
xnor U2812 (N_2812,N_2427,N_2476);
nand U2813 (N_2813,N_2253,N_2377);
or U2814 (N_2814,N_2144,N_2413);
xor U2815 (N_2815,N_2342,N_2184);
or U2816 (N_2816,N_2059,N_2459);
nand U2817 (N_2817,N_2203,N_2410);
nor U2818 (N_2818,N_2443,N_2083);
and U2819 (N_2819,N_2185,N_2322);
or U2820 (N_2820,N_2031,N_2064);
nand U2821 (N_2821,N_2296,N_2009);
and U2822 (N_2822,N_2152,N_2000);
nor U2823 (N_2823,N_2270,N_2209);
or U2824 (N_2824,N_2275,N_2101);
nand U2825 (N_2825,N_2067,N_2238);
nand U2826 (N_2826,N_2386,N_2038);
nor U2827 (N_2827,N_2138,N_2168);
nor U2828 (N_2828,N_2090,N_2196);
and U2829 (N_2829,N_2361,N_2232);
or U2830 (N_2830,N_2059,N_2148);
nor U2831 (N_2831,N_2341,N_2345);
or U2832 (N_2832,N_2233,N_2176);
nand U2833 (N_2833,N_2475,N_2375);
and U2834 (N_2834,N_2321,N_2271);
or U2835 (N_2835,N_2475,N_2136);
nor U2836 (N_2836,N_2346,N_2122);
nand U2837 (N_2837,N_2425,N_2396);
nor U2838 (N_2838,N_2218,N_2363);
and U2839 (N_2839,N_2442,N_2429);
and U2840 (N_2840,N_2275,N_2442);
nor U2841 (N_2841,N_2198,N_2086);
and U2842 (N_2842,N_2089,N_2347);
and U2843 (N_2843,N_2009,N_2255);
nor U2844 (N_2844,N_2357,N_2365);
and U2845 (N_2845,N_2236,N_2310);
nor U2846 (N_2846,N_2157,N_2115);
and U2847 (N_2847,N_2257,N_2052);
nand U2848 (N_2848,N_2304,N_2020);
nand U2849 (N_2849,N_2339,N_2223);
nor U2850 (N_2850,N_2003,N_2117);
nor U2851 (N_2851,N_2358,N_2141);
or U2852 (N_2852,N_2092,N_2281);
nor U2853 (N_2853,N_2109,N_2091);
nand U2854 (N_2854,N_2321,N_2352);
nand U2855 (N_2855,N_2332,N_2026);
nand U2856 (N_2856,N_2147,N_2134);
or U2857 (N_2857,N_2373,N_2074);
and U2858 (N_2858,N_2349,N_2140);
nor U2859 (N_2859,N_2264,N_2131);
or U2860 (N_2860,N_2196,N_2494);
nand U2861 (N_2861,N_2225,N_2132);
or U2862 (N_2862,N_2236,N_2020);
nor U2863 (N_2863,N_2151,N_2152);
and U2864 (N_2864,N_2390,N_2050);
nor U2865 (N_2865,N_2383,N_2244);
nor U2866 (N_2866,N_2421,N_2084);
nor U2867 (N_2867,N_2005,N_2399);
and U2868 (N_2868,N_2079,N_2353);
nor U2869 (N_2869,N_2258,N_2041);
and U2870 (N_2870,N_2248,N_2121);
nor U2871 (N_2871,N_2258,N_2194);
nand U2872 (N_2872,N_2086,N_2312);
nor U2873 (N_2873,N_2235,N_2426);
or U2874 (N_2874,N_2434,N_2089);
or U2875 (N_2875,N_2048,N_2447);
nand U2876 (N_2876,N_2215,N_2222);
and U2877 (N_2877,N_2312,N_2184);
nand U2878 (N_2878,N_2386,N_2204);
and U2879 (N_2879,N_2079,N_2113);
nand U2880 (N_2880,N_2055,N_2116);
nand U2881 (N_2881,N_2352,N_2086);
or U2882 (N_2882,N_2420,N_2346);
nand U2883 (N_2883,N_2210,N_2146);
or U2884 (N_2884,N_2329,N_2060);
and U2885 (N_2885,N_2472,N_2112);
nor U2886 (N_2886,N_2076,N_2116);
or U2887 (N_2887,N_2073,N_2150);
and U2888 (N_2888,N_2166,N_2081);
nand U2889 (N_2889,N_2240,N_2486);
nand U2890 (N_2890,N_2424,N_2284);
or U2891 (N_2891,N_2054,N_2363);
nand U2892 (N_2892,N_2406,N_2016);
nand U2893 (N_2893,N_2405,N_2427);
nor U2894 (N_2894,N_2011,N_2424);
and U2895 (N_2895,N_2281,N_2426);
or U2896 (N_2896,N_2483,N_2148);
nand U2897 (N_2897,N_2226,N_2044);
nor U2898 (N_2898,N_2311,N_2011);
or U2899 (N_2899,N_2160,N_2154);
or U2900 (N_2900,N_2049,N_2377);
and U2901 (N_2901,N_2014,N_2195);
or U2902 (N_2902,N_2253,N_2075);
nand U2903 (N_2903,N_2042,N_2002);
or U2904 (N_2904,N_2357,N_2292);
nand U2905 (N_2905,N_2134,N_2046);
or U2906 (N_2906,N_2057,N_2078);
nand U2907 (N_2907,N_2042,N_2097);
nand U2908 (N_2908,N_2130,N_2115);
nand U2909 (N_2909,N_2414,N_2361);
nand U2910 (N_2910,N_2126,N_2054);
nor U2911 (N_2911,N_2248,N_2146);
nor U2912 (N_2912,N_2483,N_2197);
nand U2913 (N_2913,N_2009,N_2492);
or U2914 (N_2914,N_2263,N_2208);
and U2915 (N_2915,N_2284,N_2199);
and U2916 (N_2916,N_2191,N_2491);
nor U2917 (N_2917,N_2495,N_2222);
and U2918 (N_2918,N_2140,N_2155);
or U2919 (N_2919,N_2377,N_2341);
and U2920 (N_2920,N_2312,N_2393);
or U2921 (N_2921,N_2193,N_2246);
or U2922 (N_2922,N_2374,N_2278);
nand U2923 (N_2923,N_2063,N_2268);
or U2924 (N_2924,N_2448,N_2211);
and U2925 (N_2925,N_2323,N_2355);
and U2926 (N_2926,N_2183,N_2094);
and U2927 (N_2927,N_2468,N_2076);
and U2928 (N_2928,N_2498,N_2061);
xnor U2929 (N_2929,N_2364,N_2267);
or U2930 (N_2930,N_2453,N_2208);
nor U2931 (N_2931,N_2312,N_2201);
nor U2932 (N_2932,N_2204,N_2420);
nand U2933 (N_2933,N_2304,N_2448);
nand U2934 (N_2934,N_2187,N_2154);
and U2935 (N_2935,N_2297,N_2239);
nor U2936 (N_2936,N_2123,N_2276);
nand U2937 (N_2937,N_2249,N_2011);
nand U2938 (N_2938,N_2418,N_2473);
nor U2939 (N_2939,N_2224,N_2316);
nand U2940 (N_2940,N_2114,N_2277);
nand U2941 (N_2941,N_2472,N_2488);
and U2942 (N_2942,N_2139,N_2246);
or U2943 (N_2943,N_2334,N_2403);
and U2944 (N_2944,N_2228,N_2321);
nor U2945 (N_2945,N_2359,N_2369);
or U2946 (N_2946,N_2116,N_2456);
and U2947 (N_2947,N_2013,N_2247);
and U2948 (N_2948,N_2490,N_2167);
and U2949 (N_2949,N_2026,N_2104);
and U2950 (N_2950,N_2171,N_2260);
nand U2951 (N_2951,N_2281,N_2124);
nand U2952 (N_2952,N_2097,N_2423);
and U2953 (N_2953,N_2451,N_2191);
and U2954 (N_2954,N_2439,N_2052);
and U2955 (N_2955,N_2465,N_2012);
or U2956 (N_2956,N_2045,N_2199);
or U2957 (N_2957,N_2275,N_2322);
and U2958 (N_2958,N_2337,N_2037);
nand U2959 (N_2959,N_2407,N_2210);
and U2960 (N_2960,N_2166,N_2163);
or U2961 (N_2961,N_2000,N_2477);
nor U2962 (N_2962,N_2180,N_2062);
or U2963 (N_2963,N_2169,N_2176);
nand U2964 (N_2964,N_2133,N_2202);
or U2965 (N_2965,N_2004,N_2468);
and U2966 (N_2966,N_2306,N_2214);
nor U2967 (N_2967,N_2289,N_2339);
nand U2968 (N_2968,N_2355,N_2326);
nand U2969 (N_2969,N_2050,N_2474);
nand U2970 (N_2970,N_2116,N_2432);
nand U2971 (N_2971,N_2125,N_2348);
nor U2972 (N_2972,N_2444,N_2388);
and U2973 (N_2973,N_2292,N_2278);
nor U2974 (N_2974,N_2213,N_2180);
and U2975 (N_2975,N_2475,N_2108);
and U2976 (N_2976,N_2458,N_2096);
nand U2977 (N_2977,N_2358,N_2490);
or U2978 (N_2978,N_2209,N_2045);
nand U2979 (N_2979,N_2105,N_2321);
nor U2980 (N_2980,N_2001,N_2244);
and U2981 (N_2981,N_2475,N_2465);
or U2982 (N_2982,N_2382,N_2201);
or U2983 (N_2983,N_2498,N_2114);
and U2984 (N_2984,N_2468,N_2473);
and U2985 (N_2985,N_2231,N_2309);
and U2986 (N_2986,N_2340,N_2384);
nor U2987 (N_2987,N_2434,N_2199);
and U2988 (N_2988,N_2099,N_2087);
and U2989 (N_2989,N_2216,N_2291);
and U2990 (N_2990,N_2315,N_2270);
xor U2991 (N_2991,N_2068,N_2074);
or U2992 (N_2992,N_2232,N_2099);
or U2993 (N_2993,N_2479,N_2312);
nor U2994 (N_2994,N_2479,N_2380);
nor U2995 (N_2995,N_2397,N_2451);
and U2996 (N_2996,N_2491,N_2226);
and U2997 (N_2997,N_2217,N_2344);
or U2998 (N_2998,N_2230,N_2394);
and U2999 (N_2999,N_2010,N_2000);
or U3000 (N_3000,N_2822,N_2693);
nand U3001 (N_3001,N_2887,N_2780);
nor U3002 (N_3002,N_2866,N_2662);
nor U3003 (N_3003,N_2984,N_2606);
and U3004 (N_3004,N_2621,N_2827);
or U3005 (N_3005,N_2572,N_2775);
nor U3006 (N_3006,N_2604,N_2973);
and U3007 (N_3007,N_2510,N_2627);
and U3008 (N_3008,N_2824,N_2936);
nor U3009 (N_3009,N_2565,N_2514);
or U3010 (N_3010,N_2798,N_2669);
or U3011 (N_3011,N_2533,N_2578);
nand U3012 (N_3012,N_2964,N_2707);
nor U3013 (N_3013,N_2779,N_2992);
or U3014 (N_3014,N_2969,N_2714);
or U3015 (N_3015,N_2790,N_2966);
nor U3016 (N_3016,N_2848,N_2724);
and U3017 (N_3017,N_2738,N_2642);
nor U3018 (N_3018,N_2588,N_2586);
and U3019 (N_3019,N_2647,N_2654);
and U3020 (N_3020,N_2573,N_2876);
or U3021 (N_3021,N_2659,N_2894);
and U3022 (N_3022,N_2551,N_2907);
xnor U3023 (N_3023,N_2997,N_2879);
nand U3024 (N_3024,N_2751,N_2532);
and U3025 (N_3025,N_2545,N_2835);
or U3026 (N_3026,N_2759,N_2765);
or U3027 (N_3027,N_2701,N_2526);
nand U3028 (N_3028,N_2793,N_2819);
xor U3029 (N_3029,N_2600,N_2683);
or U3030 (N_3030,N_2708,N_2908);
nand U3031 (N_3031,N_2797,N_2843);
nand U3032 (N_3032,N_2762,N_2921);
and U3033 (N_3033,N_2943,N_2684);
and U3034 (N_3034,N_2981,N_2933);
nor U3035 (N_3035,N_2605,N_2672);
nor U3036 (N_3036,N_2729,N_2541);
and U3037 (N_3037,N_2858,N_2952);
and U3038 (N_3038,N_2886,N_2567);
nor U3039 (N_3039,N_2633,N_2601);
xor U3040 (N_3040,N_2677,N_2910);
and U3041 (N_3041,N_2881,N_2599);
nor U3042 (N_3042,N_2776,N_2769);
or U3043 (N_3043,N_2616,N_2562);
xor U3044 (N_3044,N_2975,N_2632);
or U3045 (N_3045,N_2717,N_2715);
and U3046 (N_3046,N_2517,N_2882);
nand U3047 (N_3047,N_2788,N_2688);
nor U3048 (N_3048,N_2681,N_2813);
or U3049 (N_3049,N_2970,N_2608);
and U3050 (N_3050,N_2505,N_2877);
nor U3051 (N_3051,N_2689,N_2953);
and U3052 (N_3052,N_2694,N_2983);
or U3053 (N_3053,N_2513,N_2682);
nand U3054 (N_3054,N_2752,N_2963);
nor U3055 (N_3055,N_2611,N_2718);
or U3056 (N_3056,N_2965,N_2893);
nand U3057 (N_3057,N_2686,N_2516);
or U3058 (N_3058,N_2916,N_2512);
and U3059 (N_3059,N_2617,N_2940);
nand U3060 (N_3060,N_2732,N_2840);
and U3061 (N_3061,N_2704,N_2546);
or U3062 (N_3062,N_2740,N_2998);
or U3063 (N_3063,N_2622,N_2706);
nand U3064 (N_3064,N_2656,N_2530);
or U3065 (N_3065,N_2919,N_2868);
or U3066 (N_3066,N_2875,N_2579);
and U3067 (N_3067,N_2698,N_2584);
and U3068 (N_3068,N_2671,N_2990);
nor U3069 (N_3069,N_2988,N_2781);
or U3070 (N_3070,N_2703,N_2630);
and U3071 (N_3071,N_2959,N_2709);
or U3072 (N_3072,N_2861,N_2917);
and U3073 (N_3073,N_2628,N_2869);
or U3074 (N_3074,N_2838,N_2763);
nand U3075 (N_3075,N_2854,N_2646);
or U3076 (N_3076,N_2576,N_2577);
nor U3077 (N_3077,N_2673,N_2692);
and U3078 (N_3078,N_2663,N_2949);
nand U3079 (N_3079,N_2528,N_2644);
nor U3080 (N_3080,N_2836,N_2734);
nand U3081 (N_3081,N_2980,N_2537);
nor U3082 (N_3082,N_2592,N_2913);
nand U3083 (N_3083,N_2851,N_2634);
nor U3084 (N_3084,N_2653,N_2817);
xor U3085 (N_3085,N_2782,N_2666);
nand U3086 (N_3086,N_2620,N_2764);
nor U3087 (N_3087,N_2503,N_2748);
nand U3088 (N_3088,N_2711,N_2539);
or U3089 (N_3089,N_2956,N_2810);
nand U3090 (N_3090,N_2538,N_2597);
or U3091 (N_3091,N_2705,N_2585);
nand U3092 (N_3092,N_2852,N_2839);
and U3093 (N_3093,N_2501,N_2638);
nor U3094 (N_3094,N_2504,N_2543);
or U3095 (N_3095,N_2747,N_2667);
nor U3096 (N_3096,N_2926,N_2939);
and U3097 (N_3097,N_2741,N_2796);
and U3098 (N_3098,N_2590,N_2687);
nor U3099 (N_3099,N_2668,N_2697);
nor U3100 (N_3100,N_2960,N_2880);
nand U3101 (N_3101,N_2772,N_2986);
and U3102 (N_3102,N_2589,N_2758);
nor U3103 (N_3103,N_2791,N_2806);
nand U3104 (N_3104,N_2976,N_2550);
nand U3105 (N_3105,N_2524,N_2625);
or U3106 (N_3106,N_2954,N_2955);
or U3107 (N_3107,N_2925,N_2598);
and U3108 (N_3108,N_2898,N_2957);
nor U3109 (N_3109,N_2691,N_2613);
nand U3110 (N_3110,N_2815,N_2520);
nand U3111 (N_3111,N_2911,N_2730);
or U3112 (N_3112,N_2830,N_2857);
nand U3113 (N_3113,N_2811,N_2942);
nand U3114 (N_3114,N_2623,N_2721);
nor U3115 (N_3115,N_2612,N_2859);
nand U3116 (N_3116,N_2902,N_2581);
or U3117 (N_3117,N_2792,N_2658);
or U3118 (N_3118,N_2996,N_2794);
or U3119 (N_3119,N_2664,N_2795);
nor U3120 (N_3120,N_2944,N_2582);
nor U3121 (N_3121,N_2770,N_2999);
nor U3122 (N_3122,N_2750,N_2856);
and U3123 (N_3123,N_2789,N_2555);
nand U3124 (N_3124,N_2676,N_2923);
nor U3125 (N_3125,N_2831,N_2544);
nand U3126 (N_3126,N_2873,N_2728);
or U3127 (N_3127,N_2833,N_2665);
and U3128 (N_3128,N_2725,N_2872);
nand U3129 (N_3129,N_2523,N_2896);
or U3130 (N_3130,N_2920,N_2746);
nand U3131 (N_3131,N_2828,N_2778);
or U3132 (N_3132,N_2784,N_2593);
nand U3133 (N_3133,N_2652,N_2771);
nor U3134 (N_3134,N_2823,N_2821);
or U3135 (N_3135,N_2609,N_2648);
and U3136 (N_3136,N_2534,N_2727);
and U3137 (N_3137,N_2945,N_2846);
nor U3138 (N_3138,N_2834,N_2549);
nand U3139 (N_3139,N_2660,N_2842);
and U3140 (N_3140,N_2767,N_2863);
nand U3141 (N_3141,N_2649,N_2837);
and U3142 (N_3142,N_2874,N_2571);
nand U3143 (N_3143,N_2812,N_2774);
or U3144 (N_3144,N_2744,N_2962);
or U3145 (N_3145,N_2749,N_2733);
nor U3146 (N_3146,N_2826,N_2560);
nor U3147 (N_3147,N_2756,N_2761);
or U3148 (N_3148,N_2971,N_2888);
and U3149 (N_3149,N_2643,N_2700);
or U3150 (N_3150,N_2801,N_2878);
and U3151 (N_3151,N_2935,N_2624);
or U3152 (N_3152,N_2864,N_2900);
nor U3153 (N_3153,N_2603,N_2760);
xnor U3154 (N_3154,N_2675,N_2518);
nor U3155 (N_3155,N_2540,N_2702);
or U3156 (N_3156,N_2909,N_2557);
nand U3157 (N_3157,N_2987,N_2853);
or U3158 (N_3158,N_2574,N_2766);
or U3159 (N_3159,N_2651,N_2891);
or U3160 (N_3160,N_2950,N_2841);
nor U3161 (N_3161,N_2757,N_2696);
nand U3162 (N_3162,N_2948,N_2884);
xor U3163 (N_3163,N_2650,N_2977);
or U3164 (N_3164,N_2614,N_2575);
nand U3165 (N_3165,N_2777,N_2629);
nor U3166 (N_3166,N_2928,N_2993);
nor U3167 (N_3167,N_2890,N_2972);
or U3168 (N_3168,N_2580,N_2832);
and U3169 (N_3169,N_2636,N_2802);
nor U3170 (N_3170,N_2610,N_2979);
or U3171 (N_3171,N_2800,N_2712);
nor U3172 (N_3172,N_2500,N_2937);
nand U3173 (N_3173,N_2912,N_2755);
nand U3174 (N_3174,N_2547,N_2994);
nor U3175 (N_3175,N_2525,N_2602);
xor U3176 (N_3176,N_2906,N_2559);
nor U3177 (N_3177,N_2968,N_2903);
nor U3178 (N_3178,N_2849,N_2786);
and U3179 (N_3179,N_2904,N_2548);
or U3180 (N_3180,N_2938,N_2787);
and U3181 (N_3181,N_2768,N_2922);
nand U3182 (N_3182,N_2871,N_2930);
nor U3183 (N_3183,N_2670,N_2515);
or U3184 (N_3184,N_2946,N_2743);
nand U3185 (N_3185,N_2635,N_2985);
and U3186 (N_3186,N_2640,N_2974);
and U3187 (N_3187,N_2596,N_2554);
nand U3188 (N_3188,N_2542,N_2915);
nor U3189 (N_3189,N_2690,N_2508);
nand U3190 (N_3190,N_2901,N_2958);
xnor U3191 (N_3191,N_2947,N_2511);
nor U3192 (N_3192,N_2850,N_2737);
or U3193 (N_3193,N_2587,N_2674);
and U3194 (N_3194,N_2726,N_2637);
nor U3195 (N_3195,N_2521,N_2951);
or U3196 (N_3196,N_2695,N_2914);
nor U3197 (N_3197,N_2867,N_2566);
xor U3198 (N_3198,N_2570,N_2657);
and U3199 (N_3199,N_2556,N_2989);
and U3200 (N_3200,N_2929,N_2753);
and U3201 (N_3201,N_2527,N_2594);
and U3202 (N_3202,N_2641,N_2655);
nor U3203 (N_3203,N_2558,N_2805);
and U3204 (N_3204,N_2631,N_2889);
or U3205 (N_3205,N_2803,N_2961);
nor U3206 (N_3206,N_2924,N_2897);
and U3207 (N_3207,N_2885,N_2722);
nand U3208 (N_3208,N_2710,N_2529);
nand U3209 (N_3209,N_2742,N_2731);
or U3210 (N_3210,N_2595,N_2844);
and U3211 (N_3211,N_2568,N_2591);
nor U3212 (N_3212,N_2807,N_2847);
nand U3213 (N_3213,N_2745,N_2799);
and U3214 (N_3214,N_2618,N_2995);
nor U3215 (N_3215,N_2991,N_2583);
nor U3216 (N_3216,N_2509,N_2845);
nand U3217 (N_3217,N_2619,N_2895);
and U3218 (N_3218,N_2536,N_2561);
and U3219 (N_3219,N_2716,N_2685);
and U3220 (N_3220,N_2535,N_2720);
nand U3221 (N_3221,N_2931,N_2818);
and U3222 (N_3222,N_2804,N_2552);
nor U3223 (N_3223,N_2860,N_2899);
nand U3224 (N_3224,N_2607,N_2569);
or U3225 (N_3225,N_2892,N_2564);
nand U3226 (N_3226,N_2754,N_2699);
nand U3227 (N_3227,N_2553,N_2865);
nor U3228 (N_3228,N_2918,N_2723);
nand U3229 (N_3229,N_2645,N_2967);
or U3230 (N_3230,N_2679,N_2661);
or U3231 (N_3231,N_2883,N_2626);
and U3232 (N_3232,N_2982,N_2531);
nand U3233 (N_3233,N_2808,N_2825);
and U3234 (N_3234,N_2809,N_2978);
and U3235 (N_3235,N_2563,N_2736);
nor U3236 (N_3236,N_2862,N_2829);
or U3237 (N_3237,N_2739,N_2502);
nor U3238 (N_3238,N_2507,N_2735);
nand U3239 (N_3239,N_2506,N_2680);
nor U3240 (N_3240,N_2713,N_2934);
nand U3241 (N_3241,N_2519,N_2855);
nor U3242 (N_3242,N_2785,N_2941);
nor U3243 (N_3243,N_2522,N_2870);
nand U3244 (N_3244,N_2905,N_2820);
and U3245 (N_3245,N_2773,N_2639);
or U3246 (N_3246,N_2816,N_2932);
and U3247 (N_3247,N_2783,N_2615);
nor U3248 (N_3248,N_2678,N_2814);
and U3249 (N_3249,N_2927,N_2719);
nand U3250 (N_3250,N_2892,N_2847);
xor U3251 (N_3251,N_2584,N_2714);
or U3252 (N_3252,N_2876,N_2818);
and U3253 (N_3253,N_2741,N_2688);
nor U3254 (N_3254,N_2967,N_2733);
nand U3255 (N_3255,N_2833,N_2550);
nand U3256 (N_3256,N_2559,N_2582);
or U3257 (N_3257,N_2759,N_2831);
and U3258 (N_3258,N_2761,N_2971);
nand U3259 (N_3259,N_2675,N_2715);
and U3260 (N_3260,N_2533,N_2827);
nor U3261 (N_3261,N_2668,N_2844);
nor U3262 (N_3262,N_2889,N_2629);
or U3263 (N_3263,N_2515,N_2961);
nand U3264 (N_3264,N_2598,N_2809);
or U3265 (N_3265,N_2827,N_2542);
and U3266 (N_3266,N_2537,N_2874);
or U3267 (N_3267,N_2576,N_2848);
or U3268 (N_3268,N_2579,N_2559);
and U3269 (N_3269,N_2992,N_2692);
or U3270 (N_3270,N_2866,N_2564);
nor U3271 (N_3271,N_2899,N_2517);
nand U3272 (N_3272,N_2606,N_2937);
nor U3273 (N_3273,N_2921,N_2675);
and U3274 (N_3274,N_2838,N_2652);
nor U3275 (N_3275,N_2504,N_2801);
nand U3276 (N_3276,N_2509,N_2547);
nand U3277 (N_3277,N_2582,N_2759);
xor U3278 (N_3278,N_2898,N_2576);
nor U3279 (N_3279,N_2979,N_2650);
and U3280 (N_3280,N_2641,N_2830);
nor U3281 (N_3281,N_2614,N_2936);
and U3282 (N_3282,N_2733,N_2633);
nor U3283 (N_3283,N_2834,N_2554);
nand U3284 (N_3284,N_2945,N_2749);
or U3285 (N_3285,N_2628,N_2730);
and U3286 (N_3286,N_2522,N_2976);
xor U3287 (N_3287,N_2684,N_2882);
nand U3288 (N_3288,N_2660,N_2931);
nor U3289 (N_3289,N_2937,N_2593);
nand U3290 (N_3290,N_2525,N_2687);
nand U3291 (N_3291,N_2744,N_2930);
nand U3292 (N_3292,N_2778,N_2573);
and U3293 (N_3293,N_2595,N_2840);
or U3294 (N_3294,N_2860,N_2837);
nand U3295 (N_3295,N_2918,N_2830);
nand U3296 (N_3296,N_2724,N_2506);
nand U3297 (N_3297,N_2736,N_2940);
nand U3298 (N_3298,N_2702,N_2784);
or U3299 (N_3299,N_2790,N_2899);
and U3300 (N_3300,N_2624,N_2610);
or U3301 (N_3301,N_2949,N_2808);
nand U3302 (N_3302,N_2563,N_2993);
nor U3303 (N_3303,N_2514,N_2881);
and U3304 (N_3304,N_2527,N_2692);
nor U3305 (N_3305,N_2993,N_2921);
nor U3306 (N_3306,N_2647,N_2910);
nor U3307 (N_3307,N_2925,N_2724);
nand U3308 (N_3308,N_2625,N_2580);
nor U3309 (N_3309,N_2739,N_2516);
and U3310 (N_3310,N_2971,N_2877);
or U3311 (N_3311,N_2918,N_2798);
and U3312 (N_3312,N_2887,N_2738);
and U3313 (N_3313,N_2548,N_2856);
nor U3314 (N_3314,N_2988,N_2582);
nand U3315 (N_3315,N_2916,N_2586);
nand U3316 (N_3316,N_2590,N_2838);
and U3317 (N_3317,N_2748,N_2919);
nand U3318 (N_3318,N_2667,N_2724);
and U3319 (N_3319,N_2552,N_2824);
nor U3320 (N_3320,N_2606,N_2796);
or U3321 (N_3321,N_2722,N_2811);
xnor U3322 (N_3322,N_2695,N_2902);
nor U3323 (N_3323,N_2558,N_2769);
nand U3324 (N_3324,N_2873,N_2550);
nand U3325 (N_3325,N_2775,N_2647);
nand U3326 (N_3326,N_2628,N_2971);
nand U3327 (N_3327,N_2975,N_2950);
or U3328 (N_3328,N_2523,N_2517);
nor U3329 (N_3329,N_2633,N_2960);
nand U3330 (N_3330,N_2892,N_2816);
nor U3331 (N_3331,N_2815,N_2626);
and U3332 (N_3332,N_2880,N_2843);
and U3333 (N_3333,N_2533,N_2691);
nand U3334 (N_3334,N_2566,N_2983);
nor U3335 (N_3335,N_2828,N_2736);
nor U3336 (N_3336,N_2820,N_2696);
xnor U3337 (N_3337,N_2885,N_2720);
nor U3338 (N_3338,N_2991,N_2593);
and U3339 (N_3339,N_2931,N_2809);
nor U3340 (N_3340,N_2988,N_2895);
nor U3341 (N_3341,N_2892,N_2906);
or U3342 (N_3342,N_2569,N_2839);
and U3343 (N_3343,N_2649,N_2852);
nor U3344 (N_3344,N_2581,N_2785);
nand U3345 (N_3345,N_2996,N_2745);
or U3346 (N_3346,N_2980,N_2801);
nor U3347 (N_3347,N_2761,N_2526);
nor U3348 (N_3348,N_2506,N_2683);
or U3349 (N_3349,N_2582,N_2951);
nand U3350 (N_3350,N_2882,N_2791);
or U3351 (N_3351,N_2546,N_2786);
nand U3352 (N_3352,N_2829,N_2506);
nand U3353 (N_3353,N_2948,N_2666);
or U3354 (N_3354,N_2569,N_2665);
nor U3355 (N_3355,N_2617,N_2563);
nor U3356 (N_3356,N_2933,N_2757);
and U3357 (N_3357,N_2893,N_2657);
or U3358 (N_3358,N_2798,N_2832);
nand U3359 (N_3359,N_2808,N_2938);
nand U3360 (N_3360,N_2993,N_2653);
nand U3361 (N_3361,N_2681,N_2639);
xnor U3362 (N_3362,N_2695,N_2807);
nand U3363 (N_3363,N_2671,N_2541);
and U3364 (N_3364,N_2634,N_2509);
and U3365 (N_3365,N_2742,N_2894);
xor U3366 (N_3366,N_2894,N_2508);
or U3367 (N_3367,N_2693,N_2607);
or U3368 (N_3368,N_2673,N_2722);
nand U3369 (N_3369,N_2641,N_2612);
or U3370 (N_3370,N_2550,N_2544);
and U3371 (N_3371,N_2951,N_2855);
or U3372 (N_3372,N_2656,N_2674);
nor U3373 (N_3373,N_2647,N_2921);
and U3374 (N_3374,N_2548,N_2596);
nand U3375 (N_3375,N_2750,N_2658);
nor U3376 (N_3376,N_2543,N_2635);
or U3377 (N_3377,N_2752,N_2718);
and U3378 (N_3378,N_2761,N_2880);
nand U3379 (N_3379,N_2812,N_2993);
and U3380 (N_3380,N_2825,N_2975);
nor U3381 (N_3381,N_2843,N_2748);
nor U3382 (N_3382,N_2686,N_2786);
nand U3383 (N_3383,N_2923,N_2559);
nand U3384 (N_3384,N_2745,N_2987);
nand U3385 (N_3385,N_2580,N_2683);
and U3386 (N_3386,N_2793,N_2589);
nor U3387 (N_3387,N_2583,N_2763);
nor U3388 (N_3388,N_2628,N_2798);
and U3389 (N_3389,N_2502,N_2730);
xnor U3390 (N_3390,N_2502,N_2719);
nor U3391 (N_3391,N_2816,N_2634);
nand U3392 (N_3392,N_2628,N_2537);
nand U3393 (N_3393,N_2720,N_2614);
nor U3394 (N_3394,N_2768,N_2853);
nor U3395 (N_3395,N_2667,N_2973);
and U3396 (N_3396,N_2802,N_2905);
and U3397 (N_3397,N_2966,N_2849);
and U3398 (N_3398,N_2964,N_2712);
nand U3399 (N_3399,N_2920,N_2750);
xnor U3400 (N_3400,N_2698,N_2948);
nor U3401 (N_3401,N_2892,N_2986);
or U3402 (N_3402,N_2810,N_2728);
nand U3403 (N_3403,N_2770,N_2522);
and U3404 (N_3404,N_2943,N_2672);
and U3405 (N_3405,N_2889,N_2857);
nand U3406 (N_3406,N_2997,N_2827);
nand U3407 (N_3407,N_2654,N_2714);
nand U3408 (N_3408,N_2532,N_2829);
and U3409 (N_3409,N_2639,N_2581);
or U3410 (N_3410,N_2591,N_2665);
and U3411 (N_3411,N_2637,N_2526);
nand U3412 (N_3412,N_2922,N_2946);
or U3413 (N_3413,N_2503,N_2687);
nand U3414 (N_3414,N_2958,N_2825);
nor U3415 (N_3415,N_2777,N_2557);
nand U3416 (N_3416,N_2932,N_2711);
xnor U3417 (N_3417,N_2685,N_2578);
or U3418 (N_3418,N_2770,N_2838);
nor U3419 (N_3419,N_2713,N_2521);
and U3420 (N_3420,N_2569,N_2832);
or U3421 (N_3421,N_2902,N_2719);
or U3422 (N_3422,N_2990,N_2524);
nand U3423 (N_3423,N_2955,N_2826);
nand U3424 (N_3424,N_2832,N_2740);
and U3425 (N_3425,N_2606,N_2547);
and U3426 (N_3426,N_2784,N_2922);
or U3427 (N_3427,N_2701,N_2573);
nor U3428 (N_3428,N_2668,N_2758);
nor U3429 (N_3429,N_2560,N_2745);
and U3430 (N_3430,N_2982,N_2979);
or U3431 (N_3431,N_2900,N_2940);
or U3432 (N_3432,N_2829,N_2569);
or U3433 (N_3433,N_2794,N_2970);
nor U3434 (N_3434,N_2907,N_2953);
nand U3435 (N_3435,N_2616,N_2581);
nor U3436 (N_3436,N_2914,N_2923);
nand U3437 (N_3437,N_2547,N_2678);
nand U3438 (N_3438,N_2798,N_2837);
or U3439 (N_3439,N_2620,N_2979);
nor U3440 (N_3440,N_2552,N_2762);
nor U3441 (N_3441,N_2937,N_2654);
nand U3442 (N_3442,N_2940,N_2655);
nand U3443 (N_3443,N_2629,N_2518);
nor U3444 (N_3444,N_2833,N_2548);
nor U3445 (N_3445,N_2692,N_2896);
nor U3446 (N_3446,N_2647,N_2708);
nor U3447 (N_3447,N_2906,N_2608);
nor U3448 (N_3448,N_2533,N_2603);
nand U3449 (N_3449,N_2903,N_2753);
nor U3450 (N_3450,N_2585,N_2703);
or U3451 (N_3451,N_2646,N_2968);
nand U3452 (N_3452,N_2506,N_2971);
nand U3453 (N_3453,N_2769,N_2744);
and U3454 (N_3454,N_2709,N_2592);
or U3455 (N_3455,N_2923,N_2683);
or U3456 (N_3456,N_2851,N_2861);
nand U3457 (N_3457,N_2604,N_2649);
or U3458 (N_3458,N_2964,N_2652);
or U3459 (N_3459,N_2957,N_2535);
nor U3460 (N_3460,N_2805,N_2871);
or U3461 (N_3461,N_2828,N_2827);
or U3462 (N_3462,N_2992,N_2985);
nand U3463 (N_3463,N_2716,N_2648);
and U3464 (N_3464,N_2629,N_2501);
nand U3465 (N_3465,N_2841,N_2914);
nor U3466 (N_3466,N_2627,N_2764);
nor U3467 (N_3467,N_2931,N_2975);
nor U3468 (N_3468,N_2550,N_2514);
or U3469 (N_3469,N_2942,N_2851);
xor U3470 (N_3470,N_2844,N_2741);
and U3471 (N_3471,N_2902,N_2613);
and U3472 (N_3472,N_2528,N_2521);
or U3473 (N_3473,N_2974,N_2630);
and U3474 (N_3474,N_2759,N_2805);
or U3475 (N_3475,N_2823,N_2581);
xor U3476 (N_3476,N_2866,N_2502);
or U3477 (N_3477,N_2987,N_2899);
or U3478 (N_3478,N_2874,N_2834);
and U3479 (N_3479,N_2521,N_2678);
and U3480 (N_3480,N_2796,N_2747);
nor U3481 (N_3481,N_2633,N_2703);
and U3482 (N_3482,N_2653,N_2982);
and U3483 (N_3483,N_2739,N_2580);
nand U3484 (N_3484,N_2787,N_2657);
or U3485 (N_3485,N_2795,N_2575);
and U3486 (N_3486,N_2757,N_2603);
and U3487 (N_3487,N_2639,N_2846);
nand U3488 (N_3488,N_2650,N_2695);
nor U3489 (N_3489,N_2556,N_2912);
and U3490 (N_3490,N_2910,N_2643);
nand U3491 (N_3491,N_2955,N_2924);
nor U3492 (N_3492,N_2737,N_2710);
nor U3493 (N_3493,N_2696,N_2985);
nand U3494 (N_3494,N_2710,N_2562);
and U3495 (N_3495,N_2806,N_2569);
nor U3496 (N_3496,N_2520,N_2601);
nor U3497 (N_3497,N_2546,N_2814);
and U3498 (N_3498,N_2951,N_2826);
nor U3499 (N_3499,N_2626,N_2573);
or U3500 (N_3500,N_3045,N_3305);
xor U3501 (N_3501,N_3337,N_3031);
and U3502 (N_3502,N_3028,N_3355);
or U3503 (N_3503,N_3482,N_3233);
or U3504 (N_3504,N_3067,N_3412);
nor U3505 (N_3505,N_3144,N_3261);
nand U3506 (N_3506,N_3078,N_3154);
nand U3507 (N_3507,N_3300,N_3225);
and U3508 (N_3508,N_3285,N_3170);
and U3509 (N_3509,N_3242,N_3119);
nand U3510 (N_3510,N_3431,N_3231);
nand U3511 (N_3511,N_3486,N_3432);
and U3512 (N_3512,N_3060,N_3008);
and U3513 (N_3513,N_3322,N_3309);
nor U3514 (N_3514,N_3160,N_3320);
xnor U3515 (N_3515,N_3422,N_3338);
nand U3516 (N_3516,N_3084,N_3376);
or U3517 (N_3517,N_3459,N_3414);
nor U3518 (N_3518,N_3162,N_3130);
and U3519 (N_3519,N_3037,N_3014);
or U3520 (N_3520,N_3229,N_3265);
and U3521 (N_3521,N_3110,N_3105);
nand U3522 (N_3522,N_3380,N_3100);
and U3523 (N_3523,N_3319,N_3394);
nor U3524 (N_3524,N_3442,N_3142);
or U3525 (N_3525,N_3013,N_3150);
nor U3526 (N_3526,N_3097,N_3001);
nor U3527 (N_3527,N_3308,N_3342);
nor U3528 (N_3528,N_3088,N_3054);
nand U3529 (N_3529,N_3195,N_3369);
and U3530 (N_3530,N_3306,N_3435);
or U3531 (N_3531,N_3359,N_3258);
nor U3532 (N_3532,N_3217,N_3147);
and U3533 (N_3533,N_3096,N_3057);
nor U3534 (N_3534,N_3377,N_3026);
nand U3535 (N_3535,N_3458,N_3248);
nor U3536 (N_3536,N_3244,N_3087);
nor U3537 (N_3537,N_3047,N_3395);
or U3538 (N_3538,N_3043,N_3348);
and U3539 (N_3539,N_3234,N_3210);
or U3540 (N_3540,N_3325,N_3099);
nor U3541 (N_3541,N_3135,N_3176);
nor U3542 (N_3542,N_3102,N_3205);
or U3543 (N_3543,N_3161,N_3282);
and U3544 (N_3544,N_3221,N_3403);
and U3545 (N_3545,N_3200,N_3232);
nor U3546 (N_3546,N_3071,N_3438);
nand U3547 (N_3547,N_3303,N_3490);
or U3548 (N_3548,N_3464,N_3451);
nand U3549 (N_3549,N_3035,N_3434);
xor U3550 (N_3550,N_3273,N_3391);
nor U3551 (N_3551,N_3137,N_3297);
nor U3552 (N_3552,N_3418,N_3456);
and U3553 (N_3553,N_3321,N_3447);
nand U3554 (N_3554,N_3362,N_3336);
or U3555 (N_3555,N_3034,N_3347);
and U3556 (N_3556,N_3404,N_3151);
nand U3557 (N_3557,N_3240,N_3016);
nor U3558 (N_3558,N_3264,N_3344);
and U3559 (N_3559,N_3296,N_3201);
nand U3560 (N_3560,N_3367,N_3477);
or U3561 (N_3561,N_3196,N_3385);
or U3562 (N_3562,N_3211,N_3283);
nand U3563 (N_3563,N_3222,N_3169);
nand U3564 (N_3564,N_3123,N_3198);
and U3565 (N_3565,N_3167,N_3061);
nand U3566 (N_3566,N_3266,N_3298);
and U3567 (N_3567,N_3117,N_3461);
and U3568 (N_3568,N_3474,N_3327);
nand U3569 (N_3569,N_3081,N_3386);
and U3570 (N_3570,N_3304,N_3440);
nand U3571 (N_3571,N_3236,N_3106);
xnor U3572 (N_3572,N_3289,N_3357);
xor U3573 (N_3573,N_3223,N_3335);
and U3574 (N_3574,N_3029,N_3245);
nor U3575 (N_3575,N_3324,N_3062);
or U3576 (N_3576,N_3463,N_3288);
nor U3577 (N_3577,N_3468,N_3098);
or U3578 (N_3578,N_3277,N_3146);
and U3579 (N_3579,N_3382,N_3295);
nor U3580 (N_3580,N_3317,N_3156);
and U3581 (N_3581,N_3000,N_3024);
nand U3582 (N_3582,N_3488,N_3199);
nor U3583 (N_3583,N_3493,N_3360);
nor U3584 (N_3584,N_3393,N_3247);
nand U3585 (N_3585,N_3122,N_3272);
and U3586 (N_3586,N_3290,N_3495);
nand U3587 (N_3587,N_3301,N_3187);
xnor U3588 (N_3588,N_3249,N_3185);
nor U3589 (N_3589,N_3085,N_3333);
nor U3590 (N_3590,N_3019,N_3094);
nand U3591 (N_3591,N_3433,N_3454);
nand U3592 (N_3592,N_3375,N_3471);
nand U3593 (N_3593,N_3082,N_3326);
or U3594 (N_3594,N_3239,N_3421);
and U3595 (N_3595,N_3113,N_3152);
or U3596 (N_3596,N_3025,N_3483);
and U3597 (N_3597,N_3165,N_3402);
nand U3598 (N_3598,N_3315,N_3473);
nand U3599 (N_3599,N_3109,N_3379);
nand U3600 (N_3600,N_3383,N_3095);
nor U3601 (N_3601,N_3115,N_3332);
or U3602 (N_3602,N_3466,N_3120);
nor U3603 (N_3603,N_3059,N_3188);
or U3604 (N_3604,N_3193,N_3489);
nor U3605 (N_3605,N_3033,N_3416);
nand U3606 (N_3606,N_3207,N_3191);
nand U3607 (N_3607,N_3441,N_3075);
and U3608 (N_3608,N_3184,N_3055);
and U3609 (N_3609,N_3230,N_3125);
nor U3610 (N_3610,N_3006,N_3243);
and U3611 (N_3611,N_3140,N_3168);
and U3612 (N_3612,N_3250,N_3036);
nand U3613 (N_3613,N_3323,N_3172);
or U3614 (N_3614,N_3491,N_3093);
or U3615 (N_3615,N_3330,N_3164);
nor U3616 (N_3616,N_3133,N_3018);
or U3617 (N_3617,N_3259,N_3280);
nand U3618 (N_3618,N_3462,N_3453);
or U3619 (N_3619,N_3287,N_3420);
nor U3620 (N_3620,N_3126,N_3370);
or U3621 (N_3621,N_3053,N_3050);
nand U3622 (N_3622,N_3499,N_3279);
or U3623 (N_3623,N_3238,N_3148);
nand U3624 (N_3624,N_3138,N_3291);
and U3625 (N_3625,N_3032,N_3423);
nand U3626 (N_3626,N_3051,N_3262);
and U3627 (N_3627,N_3350,N_3074);
nor U3628 (N_3628,N_3202,N_3400);
or U3629 (N_3629,N_3389,N_3443);
nand U3630 (N_3630,N_3153,N_3455);
nor U3631 (N_3631,N_3334,N_3346);
or U3632 (N_3632,N_3341,N_3424);
xnor U3633 (N_3633,N_3178,N_3166);
and U3634 (N_3634,N_3478,N_3343);
and U3635 (N_3635,N_3470,N_3437);
nand U3636 (N_3636,N_3003,N_3173);
or U3637 (N_3637,N_3163,N_3048);
and U3638 (N_3638,N_3182,N_3409);
nand U3639 (N_3639,N_3020,N_3373);
nand U3640 (N_3640,N_3214,N_3398);
xnor U3641 (N_3641,N_3132,N_3040);
nand U3642 (N_3642,N_3446,N_3010);
nand U3643 (N_3643,N_3378,N_3179);
nand U3644 (N_3644,N_3406,N_3030);
and U3645 (N_3645,N_3263,N_3044);
nor U3646 (N_3646,N_3310,N_3318);
nand U3647 (N_3647,N_3425,N_3022);
and U3648 (N_3648,N_3415,N_3215);
nor U3649 (N_3649,N_3253,N_3209);
and U3650 (N_3650,N_3267,N_3103);
nor U3651 (N_3651,N_3364,N_3313);
and U3652 (N_3652,N_3387,N_3015);
and U3653 (N_3653,N_3136,N_3427);
nand U3654 (N_3654,N_3257,N_3203);
nand U3655 (N_3655,N_3080,N_3371);
nor U3656 (N_3656,N_3246,N_3481);
or U3657 (N_3657,N_3017,N_3066);
nor U3658 (N_3658,N_3197,N_3065);
and U3659 (N_3659,N_3177,N_3396);
nand U3660 (N_3660,N_3274,N_3311);
and U3661 (N_3661,N_3316,N_3129);
nor U3662 (N_3662,N_3307,N_3208);
nor U3663 (N_3663,N_3235,N_3042);
nor U3664 (N_3664,N_3108,N_3049);
and U3665 (N_3665,N_3340,N_3388);
nor U3666 (N_3666,N_3284,N_3460);
or U3667 (N_3667,N_3293,N_3157);
nor U3668 (N_3668,N_3005,N_3363);
and U3669 (N_3669,N_3116,N_3011);
nand U3670 (N_3670,N_3226,N_3063);
nor U3671 (N_3671,N_3374,N_3021);
or U3672 (N_3672,N_3128,N_3410);
nor U3673 (N_3673,N_3183,N_3012);
and U3674 (N_3674,N_3218,N_3448);
nand U3675 (N_3675,N_3083,N_3092);
nand U3676 (N_3676,N_3487,N_3352);
nand U3677 (N_3677,N_3181,N_3328);
nand U3678 (N_3678,N_3407,N_3299);
nand U3679 (N_3679,N_3417,N_3254);
and U3680 (N_3680,N_3155,N_3227);
nor U3681 (N_3681,N_3439,N_3397);
nand U3682 (N_3682,N_3220,N_3428);
nand U3683 (N_3683,N_3213,N_3159);
nor U3684 (N_3684,N_3046,N_3294);
and U3685 (N_3685,N_3484,N_3292);
and U3686 (N_3686,N_3390,N_3175);
and U3687 (N_3687,N_3212,N_3426);
and U3688 (N_3688,N_3286,N_3312);
or U3689 (N_3689,N_3276,N_3145);
and U3690 (N_3690,N_3121,N_3469);
nand U3691 (N_3691,N_3452,N_3450);
nor U3692 (N_3692,N_3480,N_3068);
and U3693 (N_3693,N_3275,N_3064);
and U3694 (N_3694,N_3381,N_3131);
nor U3695 (N_3695,N_3118,N_3039);
and U3696 (N_3696,N_3497,N_3445);
nor U3697 (N_3697,N_3171,N_3091);
xor U3698 (N_3698,N_3009,N_3436);
or U3699 (N_3699,N_3358,N_3216);
nor U3700 (N_3700,N_3219,N_3408);
or U3701 (N_3701,N_3281,N_3090);
nor U3702 (N_3702,N_3401,N_3127);
and U3703 (N_3703,N_3457,N_3339);
and U3704 (N_3704,N_3302,N_3314);
nand U3705 (N_3705,N_3430,N_3124);
nand U3706 (N_3706,N_3349,N_3411);
and U3707 (N_3707,N_3268,N_3354);
and U3708 (N_3708,N_3134,N_3413);
xor U3709 (N_3709,N_3076,N_3023);
or U3710 (N_3710,N_3190,N_3189);
and U3711 (N_3711,N_3429,N_3072);
and U3712 (N_3712,N_3351,N_3372);
and U3713 (N_3713,N_3052,N_3069);
nor U3714 (N_3714,N_3331,N_3077);
xnor U3715 (N_3715,N_3419,N_3492);
or U3716 (N_3716,N_3206,N_3158);
nand U3717 (N_3717,N_3485,N_3365);
and U3718 (N_3718,N_3027,N_3255);
or U3719 (N_3719,N_3141,N_3149);
and U3720 (N_3720,N_3476,N_3260);
nor U3721 (N_3721,N_3467,N_3104);
and U3722 (N_3722,N_3058,N_3007);
or U3723 (N_3723,N_3139,N_3101);
nor U3724 (N_3724,N_3089,N_3405);
nand U3725 (N_3725,N_3112,N_3228);
and U3726 (N_3726,N_3038,N_3465);
and U3727 (N_3727,N_3498,N_3496);
or U3728 (N_3728,N_3269,N_3194);
xnor U3729 (N_3729,N_3143,N_3356);
and U3730 (N_3730,N_3392,N_3079);
nor U3731 (N_3731,N_3086,N_3366);
or U3732 (N_3732,N_3270,N_3114);
nand U3733 (N_3733,N_3251,N_3271);
and U3734 (N_3734,N_3174,N_3329);
or U3735 (N_3735,N_3041,N_3192);
or U3736 (N_3736,N_3353,N_3361);
and U3737 (N_3737,N_3107,N_3368);
and U3738 (N_3738,N_3241,N_3494);
nor U3739 (N_3739,N_3224,N_3180);
nand U3740 (N_3740,N_3449,N_3111);
or U3741 (N_3741,N_3073,N_3384);
and U3742 (N_3742,N_3256,N_3252);
and U3743 (N_3743,N_3444,N_3070);
nor U3744 (N_3744,N_3472,N_3237);
nor U3745 (N_3745,N_3056,N_3399);
and U3746 (N_3746,N_3475,N_3278);
xnor U3747 (N_3747,N_3479,N_3004);
nand U3748 (N_3748,N_3002,N_3186);
nor U3749 (N_3749,N_3204,N_3345);
and U3750 (N_3750,N_3372,N_3225);
nand U3751 (N_3751,N_3157,N_3364);
nand U3752 (N_3752,N_3315,N_3467);
or U3753 (N_3753,N_3369,N_3333);
or U3754 (N_3754,N_3219,N_3130);
or U3755 (N_3755,N_3235,N_3212);
nand U3756 (N_3756,N_3135,N_3443);
and U3757 (N_3757,N_3264,N_3372);
or U3758 (N_3758,N_3182,N_3346);
nor U3759 (N_3759,N_3143,N_3491);
or U3760 (N_3760,N_3076,N_3064);
and U3761 (N_3761,N_3333,N_3387);
or U3762 (N_3762,N_3433,N_3104);
nor U3763 (N_3763,N_3198,N_3000);
nand U3764 (N_3764,N_3146,N_3135);
or U3765 (N_3765,N_3440,N_3035);
nand U3766 (N_3766,N_3402,N_3292);
or U3767 (N_3767,N_3295,N_3229);
or U3768 (N_3768,N_3045,N_3009);
and U3769 (N_3769,N_3193,N_3043);
nand U3770 (N_3770,N_3022,N_3003);
or U3771 (N_3771,N_3376,N_3333);
or U3772 (N_3772,N_3476,N_3473);
nand U3773 (N_3773,N_3009,N_3394);
nor U3774 (N_3774,N_3264,N_3243);
nor U3775 (N_3775,N_3350,N_3333);
nand U3776 (N_3776,N_3204,N_3282);
nor U3777 (N_3777,N_3391,N_3146);
nand U3778 (N_3778,N_3104,N_3332);
nor U3779 (N_3779,N_3425,N_3016);
or U3780 (N_3780,N_3428,N_3452);
nor U3781 (N_3781,N_3360,N_3475);
and U3782 (N_3782,N_3282,N_3392);
or U3783 (N_3783,N_3492,N_3301);
nor U3784 (N_3784,N_3397,N_3322);
and U3785 (N_3785,N_3488,N_3042);
nand U3786 (N_3786,N_3348,N_3284);
nor U3787 (N_3787,N_3390,N_3403);
and U3788 (N_3788,N_3498,N_3385);
and U3789 (N_3789,N_3101,N_3242);
nor U3790 (N_3790,N_3295,N_3034);
and U3791 (N_3791,N_3086,N_3289);
and U3792 (N_3792,N_3093,N_3225);
or U3793 (N_3793,N_3450,N_3004);
nand U3794 (N_3794,N_3032,N_3285);
and U3795 (N_3795,N_3160,N_3392);
nor U3796 (N_3796,N_3464,N_3219);
nor U3797 (N_3797,N_3258,N_3094);
nor U3798 (N_3798,N_3252,N_3481);
nor U3799 (N_3799,N_3165,N_3149);
or U3800 (N_3800,N_3379,N_3074);
or U3801 (N_3801,N_3001,N_3310);
nand U3802 (N_3802,N_3071,N_3437);
and U3803 (N_3803,N_3254,N_3460);
nor U3804 (N_3804,N_3054,N_3087);
or U3805 (N_3805,N_3181,N_3450);
and U3806 (N_3806,N_3162,N_3143);
and U3807 (N_3807,N_3032,N_3354);
or U3808 (N_3808,N_3261,N_3106);
and U3809 (N_3809,N_3434,N_3204);
xnor U3810 (N_3810,N_3130,N_3059);
or U3811 (N_3811,N_3230,N_3069);
nor U3812 (N_3812,N_3123,N_3449);
xor U3813 (N_3813,N_3189,N_3354);
or U3814 (N_3814,N_3050,N_3283);
nand U3815 (N_3815,N_3153,N_3404);
nand U3816 (N_3816,N_3465,N_3078);
or U3817 (N_3817,N_3217,N_3496);
and U3818 (N_3818,N_3132,N_3098);
nand U3819 (N_3819,N_3217,N_3268);
nand U3820 (N_3820,N_3120,N_3186);
or U3821 (N_3821,N_3358,N_3215);
nor U3822 (N_3822,N_3060,N_3067);
and U3823 (N_3823,N_3353,N_3339);
and U3824 (N_3824,N_3082,N_3066);
and U3825 (N_3825,N_3099,N_3481);
xnor U3826 (N_3826,N_3040,N_3174);
or U3827 (N_3827,N_3134,N_3321);
nand U3828 (N_3828,N_3439,N_3047);
nor U3829 (N_3829,N_3002,N_3433);
nand U3830 (N_3830,N_3279,N_3059);
or U3831 (N_3831,N_3238,N_3004);
and U3832 (N_3832,N_3349,N_3144);
nor U3833 (N_3833,N_3486,N_3261);
nor U3834 (N_3834,N_3066,N_3459);
and U3835 (N_3835,N_3067,N_3020);
and U3836 (N_3836,N_3148,N_3167);
or U3837 (N_3837,N_3385,N_3481);
and U3838 (N_3838,N_3279,N_3259);
and U3839 (N_3839,N_3441,N_3091);
nor U3840 (N_3840,N_3495,N_3175);
nor U3841 (N_3841,N_3355,N_3104);
and U3842 (N_3842,N_3213,N_3090);
nor U3843 (N_3843,N_3261,N_3364);
nand U3844 (N_3844,N_3292,N_3235);
and U3845 (N_3845,N_3478,N_3337);
and U3846 (N_3846,N_3334,N_3001);
and U3847 (N_3847,N_3257,N_3397);
or U3848 (N_3848,N_3328,N_3415);
nor U3849 (N_3849,N_3137,N_3140);
or U3850 (N_3850,N_3281,N_3070);
and U3851 (N_3851,N_3130,N_3235);
or U3852 (N_3852,N_3443,N_3437);
or U3853 (N_3853,N_3194,N_3442);
or U3854 (N_3854,N_3203,N_3455);
and U3855 (N_3855,N_3363,N_3250);
nor U3856 (N_3856,N_3481,N_3287);
or U3857 (N_3857,N_3312,N_3301);
or U3858 (N_3858,N_3222,N_3116);
or U3859 (N_3859,N_3167,N_3229);
nor U3860 (N_3860,N_3374,N_3205);
or U3861 (N_3861,N_3425,N_3177);
or U3862 (N_3862,N_3010,N_3076);
and U3863 (N_3863,N_3383,N_3433);
or U3864 (N_3864,N_3487,N_3095);
or U3865 (N_3865,N_3129,N_3231);
nand U3866 (N_3866,N_3303,N_3041);
or U3867 (N_3867,N_3470,N_3332);
or U3868 (N_3868,N_3009,N_3054);
nand U3869 (N_3869,N_3054,N_3211);
or U3870 (N_3870,N_3097,N_3432);
and U3871 (N_3871,N_3220,N_3025);
and U3872 (N_3872,N_3081,N_3257);
or U3873 (N_3873,N_3023,N_3164);
or U3874 (N_3874,N_3279,N_3422);
nor U3875 (N_3875,N_3016,N_3190);
nor U3876 (N_3876,N_3136,N_3046);
and U3877 (N_3877,N_3103,N_3230);
xnor U3878 (N_3878,N_3156,N_3181);
xor U3879 (N_3879,N_3068,N_3218);
nor U3880 (N_3880,N_3083,N_3288);
and U3881 (N_3881,N_3230,N_3107);
or U3882 (N_3882,N_3230,N_3261);
nand U3883 (N_3883,N_3125,N_3426);
or U3884 (N_3884,N_3107,N_3236);
nor U3885 (N_3885,N_3041,N_3153);
nand U3886 (N_3886,N_3218,N_3003);
xor U3887 (N_3887,N_3448,N_3388);
or U3888 (N_3888,N_3197,N_3311);
and U3889 (N_3889,N_3249,N_3173);
nor U3890 (N_3890,N_3296,N_3317);
nand U3891 (N_3891,N_3190,N_3366);
and U3892 (N_3892,N_3314,N_3244);
nor U3893 (N_3893,N_3231,N_3133);
and U3894 (N_3894,N_3142,N_3070);
and U3895 (N_3895,N_3033,N_3316);
or U3896 (N_3896,N_3463,N_3167);
or U3897 (N_3897,N_3412,N_3330);
and U3898 (N_3898,N_3384,N_3089);
or U3899 (N_3899,N_3048,N_3041);
or U3900 (N_3900,N_3027,N_3440);
and U3901 (N_3901,N_3065,N_3184);
and U3902 (N_3902,N_3494,N_3014);
and U3903 (N_3903,N_3274,N_3352);
nor U3904 (N_3904,N_3235,N_3314);
or U3905 (N_3905,N_3315,N_3476);
and U3906 (N_3906,N_3205,N_3270);
or U3907 (N_3907,N_3058,N_3389);
and U3908 (N_3908,N_3279,N_3403);
nand U3909 (N_3909,N_3283,N_3048);
and U3910 (N_3910,N_3269,N_3041);
or U3911 (N_3911,N_3014,N_3004);
and U3912 (N_3912,N_3448,N_3045);
nor U3913 (N_3913,N_3465,N_3214);
and U3914 (N_3914,N_3322,N_3487);
nand U3915 (N_3915,N_3021,N_3257);
nand U3916 (N_3916,N_3151,N_3201);
and U3917 (N_3917,N_3326,N_3040);
nor U3918 (N_3918,N_3302,N_3030);
nor U3919 (N_3919,N_3044,N_3436);
and U3920 (N_3920,N_3193,N_3094);
xor U3921 (N_3921,N_3276,N_3361);
nand U3922 (N_3922,N_3321,N_3200);
and U3923 (N_3923,N_3053,N_3216);
or U3924 (N_3924,N_3334,N_3418);
nand U3925 (N_3925,N_3248,N_3273);
nand U3926 (N_3926,N_3088,N_3128);
and U3927 (N_3927,N_3259,N_3416);
and U3928 (N_3928,N_3237,N_3125);
or U3929 (N_3929,N_3029,N_3487);
nand U3930 (N_3930,N_3254,N_3122);
or U3931 (N_3931,N_3034,N_3055);
and U3932 (N_3932,N_3075,N_3187);
nor U3933 (N_3933,N_3219,N_3283);
or U3934 (N_3934,N_3006,N_3100);
nand U3935 (N_3935,N_3057,N_3414);
nand U3936 (N_3936,N_3471,N_3034);
xor U3937 (N_3937,N_3217,N_3263);
nor U3938 (N_3938,N_3211,N_3412);
nor U3939 (N_3939,N_3261,N_3465);
nor U3940 (N_3940,N_3096,N_3380);
nor U3941 (N_3941,N_3354,N_3491);
and U3942 (N_3942,N_3225,N_3114);
nor U3943 (N_3943,N_3236,N_3276);
nor U3944 (N_3944,N_3413,N_3312);
nand U3945 (N_3945,N_3094,N_3475);
xor U3946 (N_3946,N_3194,N_3210);
nand U3947 (N_3947,N_3348,N_3080);
nand U3948 (N_3948,N_3351,N_3259);
or U3949 (N_3949,N_3165,N_3466);
nor U3950 (N_3950,N_3153,N_3145);
nand U3951 (N_3951,N_3401,N_3429);
nor U3952 (N_3952,N_3291,N_3416);
or U3953 (N_3953,N_3269,N_3198);
or U3954 (N_3954,N_3478,N_3467);
nor U3955 (N_3955,N_3245,N_3186);
nor U3956 (N_3956,N_3416,N_3437);
nand U3957 (N_3957,N_3022,N_3327);
nor U3958 (N_3958,N_3355,N_3388);
nor U3959 (N_3959,N_3312,N_3124);
nand U3960 (N_3960,N_3322,N_3066);
nor U3961 (N_3961,N_3211,N_3358);
nand U3962 (N_3962,N_3477,N_3174);
and U3963 (N_3963,N_3209,N_3027);
nor U3964 (N_3964,N_3396,N_3479);
nor U3965 (N_3965,N_3176,N_3017);
nand U3966 (N_3966,N_3057,N_3314);
nand U3967 (N_3967,N_3102,N_3240);
or U3968 (N_3968,N_3046,N_3225);
and U3969 (N_3969,N_3156,N_3479);
and U3970 (N_3970,N_3340,N_3494);
nand U3971 (N_3971,N_3146,N_3309);
or U3972 (N_3972,N_3221,N_3300);
nand U3973 (N_3973,N_3088,N_3179);
nor U3974 (N_3974,N_3191,N_3211);
or U3975 (N_3975,N_3461,N_3194);
and U3976 (N_3976,N_3202,N_3453);
nor U3977 (N_3977,N_3072,N_3466);
or U3978 (N_3978,N_3335,N_3302);
or U3979 (N_3979,N_3173,N_3453);
or U3980 (N_3980,N_3048,N_3157);
and U3981 (N_3981,N_3289,N_3309);
nand U3982 (N_3982,N_3052,N_3147);
or U3983 (N_3983,N_3447,N_3047);
or U3984 (N_3984,N_3257,N_3126);
nand U3985 (N_3985,N_3471,N_3439);
and U3986 (N_3986,N_3471,N_3157);
nor U3987 (N_3987,N_3004,N_3080);
and U3988 (N_3988,N_3002,N_3379);
and U3989 (N_3989,N_3047,N_3118);
nor U3990 (N_3990,N_3498,N_3229);
nand U3991 (N_3991,N_3118,N_3198);
nor U3992 (N_3992,N_3092,N_3069);
nand U3993 (N_3993,N_3184,N_3026);
xnor U3994 (N_3994,N_3214,N_3329);
nand U3995 (N_3995,N_3198,N_3142);
and U3996 (N_3996,N_3112,N_3291);
nand U3997 (N_3997,N_3167,N_3206);
or U3998 (N_3998,N_3140,N_3240);
and U3999 (N_3999,N_3255,N_3032);
or U4000 (N_4000,N_3755,N_3996);
and U4001 (N_4001,N_3806,N_3533);
or U4002 (N_4002,N_3890,N_3546);
nand U4003 (N_4003,N_3782,N_3685);
nor U4004 (N_4004,N_3560,N_3976);
and U4005 (N_4005,N_3690,N_3787);
nor U4006 (N_4006,N_3828,N_3503);
nor U4007 (N_4007,N_3762,N_3720);
xor U4008 (N_4008,N_3670,N_3711);
and U4009 (N_4009,N_3633,N_3748);
and U4010 (N_4010,N_3651,N_3741);
nand U4011 (N_4011,N_3545,N_3613);
nand U4012 (N_4012,N_3944,N_3884);
nand U4013 (N_4013,N_3561,N_3550);
or U4014 (N_4014,N_3570,N_3522);
nand U4015 (N_4015,N_3639,N_3568);
and U4016 (N_4016,N_3852,N_3802);
nor U4017 (N_4017,N_3640,N_3812);
nor U4018 (N_4018,N_3962,N_3899);
or U4019 (N_4019,N_3593,N_3977);
xor U4020 (N_4020,N_3587,N_3527);
or U4021 (N_4021,N_3657,N_3742);
xor U4022 (N_4022,N_3644,N_3847);
and U4023 (N_4023,N_3672,N_3577);
or U4024 (N_4024,N_3653,N_3511);
nor U4025 (N_4025,N_3776,N_3796);
nand U4026 (N_4026,N_3871,N_3572);
nor U4027 (N_4027,N_3951,N_3600);
or U4028 (N_4028,N_3895,N_3662);
nor U4029 (N_4029,N_3681,N_3874);
or U4030 (N_4030,N_3746,N_3514);
nand U4031 (N_4031,N_3795,N_3980);
and U4032 (N_4032,N_3810,N_3821);
or U4033 (N_4033,N_3630,N_3800);
nor U4034 (N_4034,N_3961,N_3612);
xnor U4035 (N_4035,N_3887,N_3908);
or U4036 (N_4036,N_3739,N_3982);
or U4037 (N_4037,N_3872,N_3752);
nor U4038 (N_4038,N_3837,N_3931);
nand U4039 (N_4039,N_3615,N_3637);
or U4040 (N_4040,N_3913,N_3942);
nor U4041 (N_4041,N_3766,N_3967);
and U4042 (N_4042,N_3710,N_3716);
nand U4043 (N_4043,N_3801,N_3906);
and U4044 (N_4044,N_3547,N_3697);
nand U4045 (N_4045,N_3731,N_3502);
or U4046 (N_4046,N_3754,N_3616);
or U4047 (N_4047,N_3656,N_3713);
and U4048 (N_4048,N_3963,N_3728);
and U4049 (N_4049,N_3636,N_3599);
or U4050 (N_4050,N_3531,N_3719);
nor U4051 (N_4051,N_3680,N_3687);
nand U4052 (N_4052,N_3509,N_3729);
or U4053 (N_4053,N_3888,N_3970);
nand U4054 (N_4054,N_3679,N_3540);
nand U4055 (N_4055,N_3751,N_3870);
nor U4056 (N_4056,N_3506,N_3992);
nand U4057 (N_4057,N_3715,N_3936);
nor U4058 (N_4058,N_3948,N_3964);
or U4059 (N_4059,N_3902,N_3829);
and U4060 (N_4060,N_3983,N_3535);
and U4061 (N_4061,N_3595,N_3559);
nor U4062 (N_4062,N_3608,N_3543);
nand U4063 (N_4063,N_3738,N_3641);
and U4064 (N_4064,N_3834,N_3537);
or U4065 (N_4065,N_3933,N_3573);
nor U4066 (N_4066,N_3648,N_3596);
nand U4067 (N_4067,N_3767,N_3512);
or U4068 (N_4068,N_3588,N_3822);
and U4069 (N_4069,N_3794,N_3844);
and U4070 (N_4070,N_3501,N_3551);
nor U4071 (N_4071,N_3989,N_3517);
or U4072 (N_4072,N_3959,N_3924);
nand U4073 (N_4073,N_3791,N_3571);
nor U4074 (N_4074,N_3905,N_3622);
or U4075 (N_4075,N_3869,N_3859);
nor U4076 (N_4076,N_3629,N_3659);
and U4077 (N_4077,N_3873,N_3921);
nor U4078 (N_4078,N_3603,N_3865);
nor U4079 (N_4079,N_3567,N_3709);
or U4080 (N_4080,N_3826,N_3749);
or U4081 (N_4081,N_3526,N_3886);
nand U4082 (N_4082,N_3584,N_3623);
and U4083 (N_4083,N_3860,N_3943);
nor U4084 (N_4084,N_3733,N_3744);
nor U4085 (N_4085,N_3785,N_3957);
and U4086 (N_4086,N_3638,N_3987);
or U4087 (N_4087,N_3703,N_3524);
nand U4088 (N_4088,N_3513,N_3553);
nand U4089 (N_4089,N_3912,N_3777);
nor U4090 (N_4090,N_3893,N_3532);
nor U4091 (N_4091,N_3705,N_3909);
and U4092 (N_4092,N_3876,N_3698);
nand U4093 (N_4093,N_3722,N_3863);
and U4094 (N_4094,N_3625,N_3712);
and U4095 (N_4095,N_3566,N_3799);
or U4096 (N_4096,N_3730,N_3889);
or U4097 (N_4097,N_3652,N_3790);
or U4098 (N_4098,N_3804,N_3508);
and U4099 (N_4099,N_3918,N_3922);
and U4100 (N_4100,N_3634,N_3986);
or U4101 (N_4101,N_3792,N_3530);
nand U4102 (N_4102,N_3669,N_3862);
or U4103 (N_4103,N_3718,N_3786);
nand U4104 (N_4104,N_3984,N_3952);
nor U4105 (N_4105,N_3580,N_3507);
or U4106 (N_4106,N_3949,N_3660);
nor U4107 (N_4107,N_3617,N_3997);
nand U4108 (N_4108,N_3556,N_3856);
and U4109 (N_4109,N_3814,N_3529);
and U4110 (N_4110,N_3735,N_3937);
or U4111 (N_4111,N_3611,N_3689);
and U4112 (N_4112,N_3896,N_3939);
or U4113 (N_4113,N_3867,N_3940);
or U4114 (N_4114,N_3528,N_3857);
nand U4115 (N_4115,N_3973,N_3702);
or U4116 (N_4116,N_3538,N_3745);
and U4117 (N_4117,N_3548,N_3974);
nand U4118 (N_4118,N_3650,N_3759);
xor U4119 (N_4119,N_3793,N_3819);
and U4120 (N_4120,N_3988,N_3975);
nor U4121 (N_4121,N_3851,N_3695);
nand U4122 (N_4122,N_3621,N_3704);
or U4123 (N_4123,N_3858,N_3645);
nand U4124 (N_4124,N_3985,N_3558);
nand U4125 (N_4125,N_3534,N_3825);
nor U4126 (N_4126,N_3555,N_3809);
or U4127 (N_4127,N_3781,N_3756);
or U4128 (N_4128,N_3753,N_3654);
and U4129 (N_4129,N_3866,N_3520);
or U4130 (N_4130,N_3758,N_3945);
nand U4131 (N_4131,N_3504,N_3946);
or U4132 (N_4132,N_3700,N_3552);
or U4133 (N_4133,N_3882,N_3549);
and U4134 (N_4134,N_3598,N_3678);
nor U4135 (N_4135,N_3877,N_3590);
and U4136 (N_4136,N_3916,N_3891);
and U4137 (N_4137,N_3525,N_3676);
nand U4138 (N_4138,N_3830,N_3544);
and U4139 (N_4139,N_3723,N_3671);
or U4140 (N_4140,N_3663,N_3823);
nand U4141 (N_4141,N_3848,N_3591);
nor U4142 (N_4142,N_3892,N_3764);
or U4143 (N_4143,N_3798,N_3521);
or U4144 (N_4144,N_3979,N_3808);
or U4145 (N_4145,N_3618,N_3696);
or U4146 (N_4146,N_3881,N_3803);
nor U4147 (N_4147,N_3838,N_3845);
nand U4148 (N_4148,N_3515,N_3635);
or U4149 (N_4149,N_3727,N_3563);
nand U4150 (N_4150,N_3624,N_3628);
xnor U4151 (N_4151,N_3778,N_3647);
and U4152 (N_4152,N_3914,N_3861);
nor U4153 (N_4153,N_3763,N_3953);
or U4154 (N_4154,N_3765,N_3594);
nand U4155 (N_4155,N_3771,N_3941);
nand U4156 (N_4156,N_3947,N_3868);
nor U4157 (N_4157,N_3592,N_3578);
and U4158 (N_4158,N_3954,N_3614);
nand U4159 (N_4159,N_3911,N_3717);
and U4160 (N_4160,N_3775,N_3740);
and U4161 (N_4161,N_3993,N_3875);
or U4162 (N_4162,N_3539,N_3842);
nor U4163 (N_4163,N_3688,N_3677);
nor U4164 (N_4164,N_3646,N_3724);
or U4165 (N_4165,N_3649,N_3925);
nand U4166 (N_4166,N_3897,N_3562);
or U4167 (N_4167,N_3510,N_3894);
xor U4168 (N_4168,N_3674,N_3699);
nand U4169 (N_4169,N_3994,N_3789);
xor U4170 (N_4170,N_3926,N_3965);
and U4171 (N_4171,N_3841,N_3706);
xnor U4172 (N_4172,N_3816,N_3850);
or U4173 (N_4173,N_3835,N_3518);
nor U4174 (N_4174,N_3589,N_3505);
and U4175 (N_4175,N_3643,N_3516);
nand U4176 (N_4176,N_3920,N_3928);
nor U4177 (N_4177,N_3901,N_3541);
nor U4178 (N_4178,N_3607,N_3606);
or U4179 (N_4179,N_3779,N_3938);
and U4180 (N_4180,N_3668,N_3569);
nor U4181 (N_4181,N_3631,N_3864);
and U4182 (N_4182,N_3966,N_3813);
and U4183 (N_4183,N_3923,N_3581);
nor U4184 (N_4184,N_3770,N_3536);
nor U4185 (N_4185,N_3575,N_3900);
nand U4186 (N_4186,N_3743,N_3831);
nand U4187 (N_4187,N_3610,N_3772);
nand U4188 (N_4188,N_3788,N_3574);
or U4189 (N_4189,N_3692,N_3878);
nand U4190 (N_4190,N_3855,N_3978);
nor U4191 (N_4191,N_3990,N_3910);
nand U4192 (N_4192,N_3708,N_3691);
and U4193 (N_4193,N_3734,N_3684);
and U4194 (N_4194,N_3661,N_3955);
and U4195 (N_4195,N_3999,N_3626);
or U4196 (N_4196,N_3693,N_3620);
or U4197 (N_4197,N_3880,N_3673);
or U4198 (N_4198,N_3956,N_3736);
nor U4199 (N_4199,N_3998,N_3919);
nor U4200 (N_4200,N_3805,N_3972);
or U4201 (N_4201,N_3666,N_3917);
nor U4202 (N_4202,N_3686,N_3619);
and U4203 (N_4203,N_3557,N_3784);
or U4204 (N_4204,N_3971,N_3773);
and U4205 (N_4205,N_3694,N_3760);
and U4206 (N_4206,N_3769,N_3846);
or U4207 (N_4207,N_3683,N_3833);
nor U4208 (N_4208,N_3929,N_3854);
nand U4209 (N_4209,N_3583,N_3597);
nand U4210 (N_4210,N_3602,N_3658);
xnor U4211 (N_4211,N_3500,N_3627);
nand U4212 (N_4212,N_3609,N_3832);
or U4213 (N_4213,N_3721,N_3519);
nand U4214 (N_4214,N_3675,N_3667);
xor U4215 (N_4215,N_3737,N_3601);
or U4216 (N_4216,N_3582,N_3995);
and U4217 (N_4217,N_3907,N_3843);
nand U4218 (N_4218,N_3579,N_3840);
and U4219 (N_4219,N_3780,N_3932);
nor U4220 (N_4220,N_3565,N_3818);
or U4221 (N_4221,N_3958,N_3576);
and U4222 (N_4222,N_3968,N_3768);
nand U4223 (N_4223,N_3757,N_3585);
nor U4224 (N_4224,N_3927,N_3898);
and U4225 (N_4225,N_3827,N_3849);
nor U4226 (N_4226,N_3824,N_3836);
nor U4227 (N_4227,N_3915,N_3934);
nor U4228 (N_4228,N_3783,N_3732);
nor U4229 (N_4229,N_3554,N_3839);
or U4230 (N_4230,N_3586,N_3811);
nor U4231 (N_4231,N_3714,N_3991);
nor U4232 (N_4232,N_3707,N_3950);
or U4233 (N_4233,N_3807,N_3817);
or U4234 (N_4234,N_3665,N_3747);
and U4235 (N_4235,N_3642,N_3969);
nor U4236 (N_4236,N_3930,N_3981);
and U4237 (N_4237,N_3815,N_3883);
nand U4238 (N_4238,N_3904,N_3604);
or U4239 (N_4239,N_3655,N_3885);
and U4240 (N_4240,N_3774,N_3750);
nand U4241 (N_4241,N_3761,N_3725);
or U4242 (N_4242,N_3853,N_3797);
nor U4243 (N_4243,N_3820,N_3935);
nand U4244 (N_4244,N_3632,N_3701);
nor U4245 (N_4245,N_3542,N_3903);
nand U4246 (N_4246,N_3879,N_3682);
and U4247 (N_4247,N_3726,N_3960);
nor U4248 (N_4248,N_3664,N_3564);
nand U4249 (N_4249,N_3605,N_3523);
or U4250 (N_4250,N_3538,N_3946);
nor U4251 (N_4251,N_3527,N_3734);
and U4252 (N_4252,N_3649,N_3511);
nand U4253 (N_4253,N_3772,N_3650);
nand U4254 (N_4254,N_3779,N_3911);
nor U4255 (N_4255,N_3870,N_3656);
and U4256 (N_4256,N_3732,N_3939);
or U4257 (N_4257,N_3512,N_3957);
nor U4258 (N_4258,N_3623,N_3557);
or U4259 (N_4259,N_3833,N_3935);
nor U4260 (N_4260,N_3592,N_3697);
and U4261 (N_4261,N_3886,N_3869);
and U4262 (N_4262,N_3887,N_3672);
nand U4263 (N_4263,N_3900,N_3517);
nand U4264 (N_4264,N_3791,N_3734);
nand U4265 (N_4265,N_3571,N_3549);
nand U4266 (N_4266,N_3566,N_3745);
nor U4267 (N_4267,N_3985,N_3797);
nor U4268 (N_4268,N_3751,N_3658);
nor U4269 (N_4269,N_3851,N_3898);
nor U4270 (N_4270,N_3793,N_3936);
and U4271 (N_4271,N_3535,N_3914);
nand U4272 (N_4272,N_3507,N_3987);
or U4273 (N_4273,N_3880,N_3763);
or U4274 (N_4274,N_3791,N_3591);
or U4275 (N_4275,N_3814,N_3941);
xor U4276 (N_4276,N_3730,N_3643);
and U4277 (N_4277,N_3523,N_3958);
nor U4278 (N_4278,N_3948,N_3594);
nor U4279 (N_4279,N_3583,N_3755);
nor U4280 (N_4280,N_3968,N_3834);
or U4281 (N_4281,N_3563,N_3717);
and U4282 (N_4282,N_3973,N_3960);
or U4283 (N_4283,N_3974,N_3721);
nor U4284 (N_4284,N_3864,N_3870);
or U4285 (N_4285,N_3627,N_3871);
or U4286 (N_4286,N_3752,N_3964);
or U4287 (N_4287,N_3546,N_3855);
nor U4288 (N_4288,N_3675,N_3872);
and U4289 (N_4289,N_3812,N_3661);
and U4290 (N_4290,N_3870,N_3935);
nor U4291 (N_4291,N_3708,N_3716);
or U4292 (N_4292,N_3636,N_3680);
and U4293 (N_4293,N_3832,N_3810);
nand U4294 (N_4294,N_3583,N_3651);
and U4295 (N_4295,N_3891,N_3513);
and U4296 (N_4296,N_3948,N_3805);
and U4297 (N_4297,N_3614,N_3871);
xor U4298 (N_4298,N_3829,N_3730);
nor U4299 (N_4299,N_3674,N_3868);
or U4300 (N_4300,N_3611,N_3620);
and U4301 (N_4301,N_3703,N_3627);
and U4302 (N_4302,N_3615,N_3936);
and U4303 (N_4303,N_3910,N_3605);
or U4304 (N_4304,N_3659,N_3563);
and U4305 (N_4305,N_3535,N_3840);
nor U4306 (N_4306,N_3935,N_3644);
nor U4307 (N_4307,N_3557,N_3533);
and U4308 (N_4308,N_3855,N_3901);
nor U4309 (N_4309,N_3993,N_3573);
and U4310 (N_4310,N_3512,N_3898);
xor U4311 (N_4311,N_3930,N_3677);
nand U4312 (N_4312,N_3982,N_3519);
nor U4313 (N_4313,N_3966,N_3604);
nor U4314 (N_4314,N_3701,N_3795);
nor U4315 (N_4315,N_3775,N_3768);
or U4316 (N_4316,N_3952,N_3641);
or U4317 (N_4317,N_3501,N_3623);
or U4318 (N_4318,N_3782,N_3715);
nor U4319 (N_4319,N_3578,N_3502);
or U4320 (N_4320,N_3676,N_3563);
or U4321 (N_4321,N_3624,N_3529);
and U4322 (N_4322,N_3943,N_3911);
xnor U4323 (N_4323,N_3955,N_3660);
or U4324 (N_4324,N_3654,N_3539);
nor U4325 (N_4325,N_3790,N_3816);
and U4326 (N_4326,N_3697,N_3939);
and U4327 (N_4327,N_3676,N_3978);
nand U4328 (N_4328,N_3981,N_3547);
and U4329 (N_4329,N_3882,N_3602);
or U4330 (N_4330,N_3998,N_3738);
nand U4331 (N_4331,N_3552,N_3716);
nor U4332 (N_4332,N_3587,N_3976);
nor U4333 (N_4333,N_3520,N_3914);
and U4334 (N_4334,N_3594,N_3968);
or U4335 (N_4335,N_3787,N_3752);
and U4336 (N_4336,N_3578,N_3614);
or U4337 (N_4337,N_3773,N_3895);
nor U4338 (N_4338,N_3829,N_3781);
and U4339 (N_4339,N_3768,N_3955);
or U4340 (N_4340,N_3813,N_3563);
nor U4341 (N_4341,N_3778,N_3539);
nand U4342 (N_4342,N_3667,N_3883);
nand U4343 (N_4343,N_3560,N_3763);
nor U4344 (N_4344,N_3717,N_3568);
nand U4345 (N_4345,N_3501,N_3753);
xor U4346 (N_4346,N_3658,N_3588);
or U4347 (N_4347,N_3801,N_3526);
nand U4348 (N_4348,N_3988,N_3815);
or U4349 (N_4349,N_3917,N_3843);
and U4350 (N_4350,N_3969,N_3780);
nand U4351 (N_4351,N_3668,N_3605);
nor U4352 (N_4352,N_3971,N_3540);
or U4353 (N_4353,N_3718,N_3876);
nor U4354 (N_4354,N_3790,N_3546);
or U4355 (N_4355,N_3947,N_3994);
or U4356 (N_4356,N_3725,N_3825);
or U4357 (N_4357,N_3543,N_3601);
nor U4358 (N_4358,N_3979,N_3713);
or U4359 (N_4359,N_3730,N_3806);
nand U4360 (N_4360,N_3944,N_3841);
xor U4361 (N_4361,N_3904,N_3909);
or U4362 (N_4362,N_3876,N_3907);
or U4363 (N_4363,N_3928,N_3676);
and U4364 (N_4364,N_3675,N_3593);
nand U4365 (N_4365,N_3995,N_3549);
nor U4366 (N_4366,N_3802,N_3636);
or U4367 (N_4367,N_3993,N_3566);
and U4368 (N_4368,N_3558,N_3893);
and U4369 (N_4369,N_3793,N_3917);
or U4370 (N_4370,N_3851,N_3609);
and U4371 (N_4371,N_3607,N_3974);
and U4372 (N_4372,N_3724,N_3893);
nor U4373 (N_4373,N_3524,N_3589);
and U4374 (N_4374,N_3993,N_3771);
nand U4375 (N_4375,N_3707,N_3850);
or U4376 (N_4376,N_3544,N_3781);
nor U4377 (N_4377,N_3675,N_3905);
nor U4378 (N_4378,N_3995,N_3771);
xnor U4379 (N_4379,N_3912,N_3670);
nor U4380 (N_4380,N_3948,N_3635);
or U4381 (N_4381,N_3955,N_3709);
or U4382 (N_4382,N_3921,N_3999);
or U4383 (N_4383,N_3804,N_3757);
or U4384 (N_4384,N_3530,N_3578);
xor U4385 (N_4385,N_3973,N_3559);
xnor U4386 (N_4386,N_3629,N_3792);
or U4387 (N_4387,N_3789,N_3889);
xnor U4388 (N_4388,N_3507,N_3514);
nand U4389 (N_4389,N_3543,N_3856);
nand U4390 (N_4390,N_3765,N_3759);
and U4391 (N_4391,N_3654,N_3512);
or U4392 (N_4392,N_3864,N_3670);
and U4393 (N_4393,N_3653,N_3694);
nand U4394 (N_4394,N_3928,N_3549);
and U4395 (N_4395,N_3653,N_3506);
and U4396 (N_4396,N_3927,N_3526);
nand U4397 (N_4397,N_3941,N_3849);
nor U4398 (N_4398,N_3740,N_3921);
nor U4399 (N_4399,N_3727,N_3906);
and U4400 (N_4400,N_3934,N_3734);
and U4401 (N_4401,N_3944,N_3706);
or U4402 (N_4402,N_3554,N_3643);
or U4403 (N_4403,N_3957,N_3586);
or U4404 (N_4404,N_3565,N_3647);
nor U4405 (N_4405,N_3891,N_3580);
or U4406 (N_4406,N_3965,N_3610);
nand U4407 (N_4407,N_3591,N_3554);
or U4408 (N_4408,N_3813,N_3981);
nor U4409 (N_4409,N_3745,N_3768);
nand U4410 (N_4410,N_3976,N_3540);
nor U4411 (N_4411,N_3833,N_3787);
or U4412 (N_4412,N_3933,N_3657);
and U4413 (N_4413,N_3879,N_3889);
and U4414 (N_4414,N_3763,N_3551);
xor U4415 (N_4415,N_3590,N_3598);
nor U4416 (N_4416,N_3866,N_3610);
nand U4417 (N_4417,N_3926,N_3948);
xnor U4418 (N_4418,N_3662,N_3926);
nand U4419 (N_4419,N_3843,N_3946);
nor U4420 (N_4420,N_3546,N_3934);
or U4421 (N_4421,N_3622,N_3673);
nand U4422 (N_4422,N_3608,N_3954);
nor U4423 (N_4423,N_3500,N_3651);
or U4424 (N_4424,N_3990,N_3787);
or U4425 (N_4425,N_3741,N_3501);
and U4426 (N_4426,N_3861,N_3946);
or U4427 (N_4427,N_3898,N_3989);
nor U4428 (N_4428,N_3827,N_3563);
nand U4429 (N_4429,N_3907,N_3851);
or U4430 (N_4430,N_3573,N_3564);
nand U4431 (N_4431,N_3533,N_3931);
nand U4432 (N_4432,N_3677,N_3518);
nor U4433 (N_4433,N_3636,N_3804);
nor U4434 (N_4434,N_3773,N_3721);
xnor U4435 (N_4435,N_3877,N_3981);
or U4436 (N_4436,N_3656,N_3720);
nand U4437 (N_4437,N_3948,N_3842);
and U4438 (N_4438,N_3592,N_3649);
xnor U4439 (N_4439,N_3959,N_3652);
nand U4440 (N_4440,N_3518,N_3537);
nand U4441 (N_4441,N_3631,N_3912);
and U4442 (N_4442,N_3727,N_3981);
xor U4443 (N_4443,N_3889,N_3937);
nor U4444 (N_4444,N_3825,N_3678);
or U4445 (N_4445,N_3570,N_3874);
and U4446 (N_4446,N_3647,N_3643);
nand U4447 (N_4447,N_3701,N_3716);
nand U4448 (N_4448,N_3905,N_3851);
or U4449 (N_4449,N_3963,N_3758);
or U4450 (N_4450,N_3509,N_3727);
and U4451 (N_4451,N_3962,N_3519);
nor U4452 (N_4452,N_3996,N_3611);
nand U4453 (N_4453,N_3891,N_3886);
nor U4454 (N_4454,N_3836,N_3989);
and U4455 (N_4455,N_3667,N_3616);
and U4456 (N_4456,N_3688,N_3820);
or U4457 (N_4457,N_3821,N_3761);
nor U4458 (N_4458,N_3770,N_3771);
nor U4459 (N_4459,N_3820,N_3906);
or U4460 (N_4460,N_3788,N_3682);
or U4461 (N_4461,N_3944,N_3816);
nor U4462 (N_4462,N_3604,N_3959);
or U4463 (N_4463,N_3561,N_3855);
nand U4464 (N_4464,N_3549,N_3500);
nor U4465 (N_4465,N_3667,N_3908);
xnor U4466 (N_4466,N_3718,N_3590);
nand U4467 (N_4467,N_3996,N_3942);
nand U4468 (N_4468,N_3605,N_3988);
and U4469 (N_4469,N_3715,N_3773);
nand U4470 (N_4470,N_3834,N_3964);
nand U4471 (N_4471,N_3628,N_3870);
or U4472 (N_4472,N_3540,N_3718);
or U4473 (N_4473,N_3861,N_3726);
and U4474 (N_4474,N_3811,N_3781);
nor U4475 (N_4475,N_3941,N_3969);
and U4476 (N_4476,N_3754,N_3518);
xnor U4477 (N_4477,N_3726,N_3696);
nand U4478 (N_4478,N_3715,N_3974);
nor U4479 (N_4479,N_3681,N_3573);
and U4480 (N_4480,N_3862,N_3666);
or U4481 (N_4481,N_3729,N_3870);
nand U4482 (N_4482,N_3659,N_3671);
and U4483 (N_4483,N_3662,N_3827);
or U4484 (N_4484,N_3953,N_3695);
nor U4485 (N_4485,N_3931,N_3725);
nor U4486 (N_4486,N_3875,N_3808);
and U4487 (N_4487,N_3785,N_3862);
or U4488 (N_4488,N_3825,N_3961);
and U4489 (N_4489,N_3699,N_3632);
nand U4490 (N_4490,N_3923,N_3995);
nor U4491 (N_4491,N_3869,N_3624);
nand U4492 (N_4492,N_3623,N_3568);
nand U4493 (N_4493,N_3535,N_3647);
xor U4494 (N_4494,N_3596,N_3597);
or U4495 (N_4495,N_3795,N_3913);
or U4496 (N_4496,N_3568,N_3855);
nor U4497 (N_4497,N_3658,N_3739);
nor U4498 (N_4498,N_3623,N_3928);
or U4499 (N_4499,N_3665,N_3577);
or U4500 (N_4500,N_4327,N_4142);
or U4501 (N_4501,N_4357,N_4394);
nand U4502 (N_4502,N_4300,N_4307);
nor U4503 (N_4503,N_4365,N_4100);
and U4504 (N_4504,N_4465,N_4147);
and U4505 (N_4505,N_4039,N_4472);
or U4506 (N_4506,N_4242,N_4305);
or U4507 (N_4507,N_4024,N_4036);
nor U4508 (N_4508,N_4167,N_4027);
or U4509 (N_4509,N_4238,N_4051);
nand U4510 (N_4510,N_4445,N_4169);
nor U4511 (N_4511,N_4494,N_4450);
and U4512 (N_4512,N_4399,N_4135);
nand U4513 (N_4513,N_4134,N_4206);
and U4514 (N_4514,N_4186,N_4273);
nor U4515 (N_4515,N_4468,N_4294);
or U4516 (N_4516,N_4432,N_4409);
or U4517 (N_4517,N_4210,N_4408);
or U4518 (N_4518,N_4261,N_4175);
xnor U4519 (N_4519,N_4265,N_4412);
and U4520 (N_4520,N_4433,N_4339);
and U4521 (N_4521,N_4092,N_4011);
nand U4522 (N_4522,N_4462,N_4106);
nand U4523 (N_4523,N_4352,N_4032);
nand U4524 (N_4524,N_4444,N_4488);
xnor U4525 (N_4525,N_4292,N_4376);
nor U4526 (N_4526,N_4221,N_4340);
and U4527 (N_4527,N_4386,N_4043);
nand U4528 (N_4528,N_4013,N_4089);
or U4529 (N_4529,N_4150,N_4296);
and U4530 (N_4530,N_4220,N_4298);
nor U4531 (N_4531,N_4470,N_4196);
and U4532 (N_4532,N_4304,N_4390);
and U4533 (N_4533,N_4231,N_4377);
and U4534 (N_4534,N_4277,N_4184);
nor U4535 (N_4535,N_4228,N_4197);
nand U4536 (N_4536,N_4463,N_4435);
and U4537 (N_4537,N_4002,N_4424);
or U4538 (N_4538,N_4306,N_4192);
nand U4539 (N_4539,N_4170,N_4455);
nand U4540 (N_4540,N_4404,N_4118);
or U4541 (N_4541,N_4317,N_4268);
nor U4542 (N_4542,N_4152,N_4278);
nand U4543 (N_4543,N_4474,N_4022);
and U4544 (N_4544,N_4393,N_4359);
or U4545 (N_4545,N_4178,N_4497);
and U4546 (N_4546,N_4103,N_4166);
or U4547 (N_4547,N_4379,N_4145);
xor U4548 (N_4548,N_4094,N_4258);
nand U4549 (N_4549,N_4388,N_4498);
or U4550 (N_4550,N_4337,N_4213);
nor U4551 (N_4551,N_4283,N_4074);
or U4552 (N_4552,N_4256,N_4185);
and U4553 (N_4553,N_4173,N_4097);
and U4554 (N_4554,N_4476,N_4417);
nor U4555 (N_4555,N_4234,N_4284);
nor U4556 (N_4556,N_4368,N_4452);
and U4557 (N_4557,N_4236,N_4132);
and U4558 (N_4558,N_4275,N_4453);
nor U4559 (N_4559,N_4397,N_4403);
nand U4560 (N_4560,N_4044,N_4461);
nand U4561 (N_4561,N_4299,N_4082);
nand U4562 (N_4562,N_4285,N_4354);
and U4563 (N_4563,N_4454,N_4373);
and U4564 (N_4564,N_4230,N_4343);
xor U4565 (N_4565,N_4021,N_4114);
and U4566 (N_4566,N_4158,N_4018);
or U4567 (N_4567,N_4102,N_4301);
or U4568 (N_4568,N_4112,N_4211);
nand U4569 (N_4569,N_4257,N_4437);
nand U4570 (N_4570,N_4070,N_4405);
nand U4571 (N_4571,N_4010,N_4068);
and U4572 (N_4572,N_4180,N_4053);
nor U4573 (N_4573,N_4322,N_4204);
nor U4574 (N_4574,N_4338,N_4413);
nor U4575 (N_4575,N_4163,N_4364);
nor U4576 (N_4576,N_4076,N_4382);
nand U4577 (N_4577,N_4218,N_4289);
nand U4578 (N_4578,N_4168,N_4090);
nand U4579 (N_4579,N_4355,N_4270);
nor U4580 (N_4580,N_4119,N_4083);
or U4581 (N_4581,N_4223,N_4492);
and U4582 (N_4582,N_4235,N_4224);
or U4583 (N_4583,N_4179,N_4443);
or U4584 (N_4584,N_4334,N_4477);
or U4585 (N_4585,N_4323,N_4155);
nand U4586 (N_4586,N_4123,N_4378);
xor U4587 (N_4587,N_4269,N_4203);
nand U4588 (N_4588,N_4007,N_4342);
nor U4589 (N_4589,N_4266,N_4049);
or U4590 (N_4590,N_4212,N_4191);
or U4591 (N_4591,N_4064,N_4050);
and U4592 (N_4592,N_4005,N_4457);
and U4593 (N_4593,N_4017,N_4183);
nor U4594 (N_4594,N_4136,N_4411);
and U4595 (N_4595,N_4225,N_4216);
or U4596 (N_4596,N_4128,N_4120);
xnor U4597 (N_4597,N_4441,N_4481);
and U4598 (N_4598,N_4440,N_4396);
nand U4599 (N_4599,N_4161,N_4019);
nand U4600 (N_4600,N_4320,N_4372);
nor U4601 (N_4601,N_4260,N_4062);
and U4602 (N_4602,N_4137,N_4237);
and U4603 (N_4603,N_4088,N_4389);
nor U4604 (N_4604,N_4483,N_4016);
nor U4605 (N_4605,N_4420,N_4366);
xor U4606 (N_4606,N_4263,N_4034);
and U4607 (N_4607,N_4316,N_4029);
nor U4608 (N_4608,N_4113,N_4217);
and U4609 (N_4609,N_4361,N_4060);
or U4610 (N_4610,N_4375,N_4302);
nor U4611 (N_4611,N_4402,N_4310);
and U4612 (N_4612,N_4456,N_4008);
and U4613 (N_4613,N_4015,N_4276);
or U4614 (N_4614,N_4482,N_4189);
and U4615 (N_4615,N_4434,N_4030);
and U4616 (N_4616,N_4144,N_4140);
and U4617 (N_4617,N_4287,N_4367);
and U4618 (N_4618,N_4233,N_4293);
nand U4619 (N_4619,N_4421,N_4148);
nand U4620 (N_4620,N_4071,N_4344);
nand U4621 (N_4621,N_4124,N_4351);
nor U4622 (N_4622,N_4250,N_4303);
nand U4623 (N_4623,N_4117,N_4057);
and U4624 (N_4624,N_4133,N_4448);
nand U4625 (N_4625,N_4232,N_4254);
nand U4626 (N_4626,N_4395,N_4406);
nand U4627 (N_4627,N_4190,N_4297);
and U4628 (N_4628,N_4165,N_4077);
nor U4629 (N_4629,N_4146,N_4127);
and U4630 (N_4630,N_4108,N_4193);
and U4631 (N_4631,N_4398,N_4227);
or U4632 (N_4632,N_4346,N_4069);
nor U4633 (N_4633,N_4176,N_4247);
nand U4634 (N_4634,N_4122,N_4380);
or U4635 (N_4635,N_4329,N_4073);
and U4636 (N_4636,N_4348,N_4429);
and U4637 (N_4637,N_4360,N_4243);
nand U4638 (N_4638,N_4141,N_4047);
nor U4639 (N_4639,N_4086,N_4349);
and U4640 (N_4640,N_4309,N_4286);
or U4641 (N_4641,N_4037,N_4075);
or U4642 (N_4642,N_4072,N_4369);
or U4643 (N_4643,N_4332,N_4259);
or U4644 (N_4644,N_4109,N_4362);
or U4645 (N_4645,N_4489,N_4249);
nor U4646 (N_4646,N_4290,N_4171);
nand U4647 (N_4647,N_4341,N_4356);
xor U4648 (N_4648,N_4115,N_4104);
nand U4649 (N_4649,N_4330,N_4451);
and U4650 (N_4650,N_4000,N_4449);
and U4651 (N_4651,N_4479,N_4241);
nand U4652 (N_4652,N_4387,N_4004);
xnor U4653 (N_4653,N_4058,N_4181);
or U4654 (N_4654,N_4222,N_4093);
nor U4655 (N_4655,N_4281,N_4484);
nand U4656 (N_4656,N_4023,N_4110);
and U4657 (N_4657,N_4084,N_4208);
nor U4658 (N_4658,N_4052,N_4045);
nor U4659 (N_4659,N_4464,N_4426);
and U4660 (N_4660,N_4080,N_4499);
and U4661 (N_4661,N_4478,N_4055);
nand U4662 (N_4662,N_4061,N_4467);
and U4663 (N_4663,N_4198,N_4153);
nor U4664 (N_4664,N_4458,N_4214);
or U4665 (N_4665,N_4098,N_4475);
or U4666 (N_4666,N_4157,N_4031);
nand U4667 (N_4667,N_4188,N_4264);
or U4668 (N_4668,N_4079,N_4495);
and U4669 (N_4669,N_4430,N_4318);
or U4670 (N_4670,N_4333,N_4091);
nand U4671 (N_4671,N_4251,N_4207);
or U4672 (N_4672,N_4442,N_4126);
nand U4673 (N_4673,N_4374,N_4026);
and U4674 (N_4674,N_4130,N_4226);
nor U4675 (N_4675,N_4295,N_4014);
nor U4676 (N_4676,N_4446,N_4182);
nand U4677 (N_4677,N_4081,N_4428);
xnor U4678 (N_4678,N_4383,N_4324);
nor U4679 (N_4679,N_4202,N_4172);
nand U4680 (N_4680,N_4245,N_4418);
nand U4681 (N_4681,N_4407,N_4469);
nand U4682 (N_4682,N_4491,N_4255);
nand U4683 (N_4683,N_4056,N_4336);
nor U4684 (N_4684,N_4358,N_4156);
nor U4685 (N_4685,N_4422,N_4248);
or U4686 (N_4686,N_4078,N_4125);
and U4687 (N_4687,N_4414,N_4066);
nor U4688 (N_4688,N_4347,N_4003);
and U4689 (N_4689,N_4447,N_4041);
nand U4690 (N_4690,N_4138,N_4240);
nand U4691 (N_4691,N_4028,N_4262);
and U4692 (N_4692,N_4459,N_4466);
nor U4693 (N_4693,N_4438,N_4490);
nand U4694 (N_4694,N_4042,N_4328);
xor U4695 (N_4695,N_4040,N_4215);
nand U4696 (N_4696,N_4012,N_4205);
and U4697 (N_4697,N_4154,N_4035);
nor U4698 (N_4698,N_4020,N_4496);
xnor U4699 (N_4699,N_4063,N_4177);
and U4700 (N_4700,N_4111,N_4423);
nand U4701 (N_4701,N_4195,N_4326);
or U4702 (N_4702,N_4436,N_4485);
nor U4703 (N_4703,N_4335,N_4151);
and U4704 (N_4704,N_4252,N_4385);
nand U4705 (N_4705,N_4291,N_4280);
xnor U4706 (N_4706,N_4282,N_4279);
and U4707 (N_4707,N_4159,N_4149);
and U4708 (N_4708,N_4486,N_4054);
nor U4709 (N_4709,N_4087,N_4308);
or U4710 (N_4710,N_4219,N_4439);
and U4711 (N_4711,N_4415,N_4370);
nor U4712 (N_4712,N_4384,N_4099);
and U4713 (N_4713,N_4239,N_4229);
or U4714 (N_4714,N_4431,N_4187);
and U4715 (N_4715,N_4174,N_4162);
or U4716 (N_4716,N_4325,N_4312);
nor U4717 (N_4717,N_4311,N_4038);
nor U4718 (N_4718,N_4143,N_4116);
nor U4719 (N_4719,N_4121,N_4067);
nor U4720 (N_4720,N_4160,N_4096);
nor U4721 (N_4721,N_4314,N_4272);
nor U4722 (N_4722,N_4139,N_4046);
or U4723 (N_4723,N_4001,N_4105);
nand U4724 (N_4724,N_4345,N_4493);
and U4725 (N_4725,N_4401,N_4381);
nand U4726 (N_4726,N_4209,N_4487);
nand U4727 (N_4727,N_4048,N_4025);
or U4728 (N_4728,N_4033,N_4410);
and U4729 (N_4729,N_4244,N_4471);
or U4730 (N_4730,N_4331,N_4253);
nor U4731 (N_4731,N_4059,N_4427);
or U4732 (N_4732,N_4391,N_4480);
xor U4733 (N_4733,N_4164,N_4363);
nand U4734 (N_4734,N_4419,N_4416);
xor U4735 (N_4735,N_4095,N_4425);
or U4736 (N_4736,N_4246,N_4288);
nand U4737 (N_4737,N_4194,N_4460);
nor U4738 (N_4738,N_4371,N_4199);
nand U4739 (N_4739,N_4200,N_4006);
or U4740 (N_4740,N_4353,N_4315);
nor U4741 (N_4741,N_4267,N_4321);
nor U4742 (N_4742,N_4392,N_4065);
nor U4743 (N_4743,N_4085,N_4473);
nor U4744 (N_4744,N_4101,N_4129);
xnor U4745 (N_4745,N_4400,N_4274);
nor U4746 (N_4746,N_4271,N_4319);
and U4747 (N_4747,N_4009,N_4201);
nand U4748 (N_4748,N_4131,N_4313);
or U4749 (N_4749,N_4107,N_4350);
or U4750 (N_4750,N_4258,N_4047);
or U4751 (N_4751,N_4383,N_4309);
nor U4752 (N_4752,N_4360,N_4392);
nand U4753 (N_4753,N_4087,N_4206);
nand U4754 (N_4754,N_4026,N_4499);
and U4755 (N_4755,N_4123,N_4433);
or U4756 (N_4756,N_4416,N_4236);
nand U4757 (N_4757,N_4460,N_4369);
nor U4758 (N_4758,N_4465,N_4023);
and U4759 (N_4759,N_4209,N_4402);
nand U4760 (N_4760,N_4270,N_4278);
nand U4761 (N_4761,N_4055,N_4079);
nor U4762 (N_4762,N_4287,N_4008);
and U4763 (N_4763,N_4086,N_4484);
nand U4764 (N_4764,N_4381,N_4198);
and U4765 (N_4765,N_4152,N_4117);
xor U4766 (N_4766,N_4273,N_4030);
and U4767 (N_4767,N_4130,N_4198);
and U4768 (N_4768,N_4352,N_4268);
or U4769 (N_4769,N_4355,N_4228);
and U4770 (N_4770,N_4234,N_4183);
and U4771 (N_4771,N_4377,N_4233);
nor U4772 (N_4772,N_4148,N_4108);
nor U4773 (N_4773,N_4339,N_4239);
and U4774 (N_4774,N_4023,N_4161);
or U4775 (N_4775,N_4139,N_4300);
xor U4776 (N_4776,N_4463,N_4199);
xnor U4777 (N_4777,N_4216,N_4313);
nor U4778 (N_4778,N_4301,N_4076);
or U4779 (N_4779,N_4078,N_4471);
nor U4780 (N_4780,N_4223,N_4161);
and U4781 (N_4781,N_4246,N_4149);
or U4782 (N_4782,N_4320,N_4464);
nand U4783 (N_4783,N_4263,N_4415);
nor U4784 (N_4784,N_4048,N_4155);
nor U4785 (N_4785,N_4223,N_4145);
nand U4786 (N_4786,N_4337,N_4246);
nor U4787 (N_4787,N_4378,N_4392);
and U4788 (N_4788,N_4079,N_4091);
or U4789 (N_4789,N_4328,N_4446);
nand U4790 (N_4790,N_4303,N_4099);
nand U4791 (N_4791,N_4340,N_4431);
or U4792 (N_4792,N_4196,N_4240);
and U4793 (N_4793,N_4082,N_4109);
or U4794 (N_4794,N_4297,N_4290);
nand U4795 (N_4795,N_4039,N_4450);
or U4796 (N_4796,N_4429,N_4118);
nand U4797 (N_4797,N_4100,N_4444);
nand U4798 (N_4798,N_4247,N_4114);
or U4799 (N_4799,N_4158,N_4418);
nand U4800 (N_4800,N_4150,N_4451);
and U4801 (N_4801,N_4263,N_4373);
or U4802 (N_4802,N_4136,N_4498);
or U4803 (N_4803,N_4402,N_4464);
nor U4804 (N_4804,N_4380,N_4411);
or U4805 (N_4805,N_4375,N_4170);
nand U4806 (N_4806,N_4049,N_4345);
nor U4807 (N_4807,N_4348,N_4301);
nor U4808 (N_4808,N_4027,N_4113);
nand U4809 (N_4809,N_4013,N_4380);
and U4810 (N_4810,N_4219,N_4447);
or U4811 (N_4811,N_4489,N_4140);
nand U4812 (N_4812,N_4247,N_4156);
nand U4813 (N_4813,N_4167,N_4213);
xnor U4814 (N_4814,N_4005,N_4073);
or U4815 (N_4815,N_4302,N_4400);
and U4816 (N_4816,N_4454,N_4246);
nand U4817 (N_4817,N_4054,N_4056);
and U4818 (N_4818,N_4329,N_4021);
or U4819 (N_4819,N_4374,N_4009);
nand U4820 (N_4820,N_4060,N_4013);
nor U4821 (N_4821,N_4123,N_4015);
or U4822 (N_4822,N_4109,N_4494);
and U4823 (N_4823,N_4306,N_4254);
or U4824 (N_4824,N_4374,N_4044);
xnor U4825 (N_4825,N_4123,N_4106);
and U4826 (N_4826,N_4045,N_4409);
nand U4827 (N_4827,N_4132,N_4413);
and U4828 (N_4828,N_4359,N_4422);
nor U4829 (N_4829,N_4114,N_4362);
and U4830 (N_4830,N_4244,N_4227);
nor U4831 (N_4831,N_4264,N_4437);
and U4832 (N_4832,N_4468,N_4134);
nor U4833 (N_4833,N_4046,N_4413);
and U4834 (N_4834,N_4176,N_4411);
and U4835 (N_4835,N_4161,N_4375);
nand U4836 (N_4836,N_4231,N_4107);
nor U4837 (N_4837,N_4240,N_4028);
nor U4838 (N_4838,N_4147,N_4167);
nand U4839 (N_4839,N_4195,N_4469);
and U4840 (N_4840,N_4452,N_4211);
or U4841 (N_4841,N_4149,N_4134);
or U4842 (N_4842,N_4451,N_4147);
nor U4843 (N_4843,N_4056,N_4427);
nor U4844 (N_4844,N_4015,N_4132);
nand U4845 (N_4845,N_4101,N_4471);
nand U4846 (N_4846,N_4255,N_4231);
and U4847 (N_4847,N_4085,N_4063);
and U4848 (N_4848,N_4494,N_4043);
nand U4849 (N_4849,N_4166,N_4442);
nor U4850 (N_4850,N_4122,N_4386);
nand U4851 (N_4851,N_4014,N_4403);
or U4852 (N_4852,N_4324,N_4231);
or U4853 (N_4853,N_4090,N_4363);
and U4854 (N_4854,N_4462,N_4119);
or U4855 (N_4855,N_4371,N_4253);
and U4856 (N_4856,N_4243,N_4016);
and U4857 (N_4857,N_4309,N_4194);
nor U4858 (N_4858,N_4326,N_4051);
and U4859 (N_4859,N_4165,N_4243);
nor U4860 (N_4860,N_4306,N_4173);
nor U4861 (N_4861,N_4249,N_4051);
and U4862 (N_4862,N_4015,N_4094);
or U4863 (N_4863,N_4183,N_4333);
nor U4864 (N_4864,N_4137,N_4177);
nor U4865 (N_4865,N_4346,N_4134);
nor U4866 (N_4866,N_4072,N_4225);
and U4867 (N_4867,N_4220,N_4030);
nand U4868 (N_4868,N_4119,N_4227);
and U4869 (N_4869,N_4241,N_4153);
and U4870 (N_4870,N_4329,N_4014);
or U4871 (N_4871,N_4151,N_4323);
nor U4872 (N_4872,N_4084,N_4355);
nor U4873 (N_4873,N_4465,N_4296);
and U4874 (N_4874,N_4414,N_4208);
nor U4875 (N_4875,N_4215,N_4412);
nand U4876 (N_4876,N_4348,N_4201);
nor U4877 (N_4877,N_4231,N_4408);
and U4878 (N_4878,N_4429,N_4198);
nor U4879 (N_4879,N_4108,N_4404);
nand U4880 (N_4880,N_4192,N_4024);
nand U4881 (N_4881,N_4055,N_4024);
nor U4882 (N_4882,N_4158,N_4265);
or U4883 (N_4883,N_4097,N_4123);
and U4884 (N_4884,N_4487,N_4393);
nor U4885 (N_4885,N_4492,N_4080);
or U4886 (N_4886,N_4329,N_4307);
nand U4887 (N_4887,N_4192,N_4221);
nand U4888 (N_4888,N_4491,N_4405);
or U4889 (N_4889,N_4180,N_4430);
nand U4890 (N_4890,N_4430,N_4423);
or U4891 (N_4891,N_4149,N_4351);
or U4892 (N_4892,N_4321,N_4388);
nor U4893 (N_4893,N_4049,N_4166);
or U4894 (N_4894,N_4419,N_4216);
or U4895 (N_4895,N_4067,N_4355);
nor U4896 (N_4896,N_4195,N_4378);
and U4897 (N_4897,N_4441,N_4267);
nor U4898 (N_4898,N_4356,N_4488);
and U4899 (N_4899,N_4462,N_4179);
nor U4900 (N_4900,N_4352,N_4366);
and U4901 (N_4901,N_4214,N_4254);
or U4902 (N_4902,N_4240,N_4386);
nand U4903 (N_4903,N_4351,N_4284);
nor U4904 (N_4904,N_4297,N_4065);
or U4905 (N_4905,N_4198,N_4152);
nor U4906 (N_4906,N_4059,N_4338);
nor U4907 (N_4907,N_4150,N_4185);
nor U4908 (N_4908,N_4379,N_4037);
nor U4909 (N_4909,N_4350,N_4179);
nor U4910 (N_4910,N_4145,N_4052);
or U4911 (N_4911,N_4102,N_4275);
or U4912 (N_4912,N_4187,N_4441);
nor U4913 (N_4913,N_4382,N_4374);
or U4914 (N_4914,N_4037,N_4378);
nor U4915 (N_4915,N_4407,N_4379);
and U4916 (N_4916,N_4460,N_4488);
nor U4917 (N_4917,N_4483,N_4161);
and U4918 (N_4918,N_4203,N_4382);
nand U4919 (N_4919,N_4375,N_4127);
nand U4920 (N_4920,N_4194,N_4335);
or U4921 (N_4921,N_4429,N_4143);
or U4922 (N_4922,N_4410,N_4383);
nor U4923 (N_4923,N_4460,N_4467);
and U4924 (N_4924,N_4095,N_4337);
nor U4925 (N_4925,N_4439,N_4351);
nor U4926 (N_4926,N_4377,N_4436);
and U4927 (N_4927,N_4292,N_4491);
and U4928 (N_4928,N_4486,N_4460);
nor U4929 (N_4929,N_4070,N_4491);
or U4930 (N_4930,N_4098,N_4179);
and U4931 (N_4931,N_4087,N_4288);
nor U4932 (N_4932,N_4169,N_4187);
or U4933 (N_4933,N_4112,N_4184);
nor U4934 (N_4934,N_4282,N_4231);
or U4935 (N_4935,N_4169,N_4197);
nand U4936 (N_4936,N_4018,N_4196);
nand U4937 (N_4937,N_4228,N_4261);
nor U4938 (N_4938,N_4125,N_4374);
nor U4939 (N_4939,N_4480,N_4222);
nor U4940 (N_4940,N_4393,N_4406);
and U4941 (N_4941,N_4342,N_4038);
nand U4942 (N_4942,N_4088,N_4121);
nand U4943 (N_4943,N_4293,N_4016);
nand U4944 (N_4944,N_4012,N_4175);
or U4945 (N_4945,N_4068,N_4352);
nor U4946 (N_4946,N_4002,N_4071);
or U4947 (N_4947,N_4185,N_4048);
nand U4948 (N_4948,N_4109,N_4478);
nand U4949 (N_4949,N_4101,N_4023);
or U4950 (N_4950,N_4281,N_4044);
or U4951 (N_4951,N_4334,N_4021);
nor U4952 (N_4952,N_4248,N_4129);
or U4953 (N_4953,N_4278,N_4154);
or U4954 (N_4954,N_4371,N_4421);
nand U4955 (N_4955,N_4039,N_4458);
or U4956 (N_4956,N_4494,N_4400);
and U4957 (N_4957,N_4118,N_4170);
or U4958 (N_4958,N_4324,N_4161);
nand U4959 (N_4959,N_4231,N_4240);
nor U4960 (N_4960,N_4404,N_4277);
or U4961 (N_4961,N_4331,N_4149);
or U4962 (N_4962,N_4312,N_4410);
and U4963 (N_4963,N_4310,N_4087);
nand U4964 (N_4964,N_4071,N_4495);
nand U4965 (N_4965,N_4162,N_4064);
nor U4966 (N_4966,N_4353,N_4450);
nand U4967 (N_4967,N_4135,N_4369);
or U4968 (N_4968,N_4037,N_4128);
nor U4969 (N_4969,N_4337,N_4038);
nand U4970 (N_4970,N_4332,N_4173);
nand U4971 (N_4971,N_4490,N_4184);
and U4972 (N_4972,N_4488,N_4161);
and U4973 (N_4973,N_4410,N_4105);
or U4974 (N_4974,N_4330,N_4447);
nand U4975 (N_4975,N_4013,N_4384);
nand U4976 (N_4976,N_4449,N_4048);
nor U4977 (N_4977,N_4383,N_4170);
nor U4978 (N_4978,N_4148,N_4124);
and U4979 (N_4979,N_4458,N_4383);
nor U4980 (N_4980,N_4499,N_4329);
xnor U4981 (N_4981,N_4308,N_4093);
xor U4982 (N_4982,N_4411,N_4043);
or U4983 (N_4983,N_4118,N_4123);
and U4984 (N_4984,N_4399,N_4369);
nor U4985 (N_4985,N_4303,N_4235);
and U4986 (N_4986,N_4011,N_4086);
and U4987 (N_4987,N_4356,N_4057);
and U4988 (N_4988,N_4432,N_4237);
or U4989 (N_4989,N_4100,N_4326);
nand U4990 (N_4990,N_4332,N_4138);
xor U4991 (N_4991,N_4368,N_4416);
xor U4992 (N_4992,N_4103,N_4076);
or U4993 (N_4993,N_4247,N_4059);
or U4994 (N_4994,N_4037,N_4219);
or U4995 (N_4995,N_4311,N_4335);
or U4996 (N_4996,N_4178,N_4315);
or U4997 (N_4997,N_4189,N_4108);
nor U4998 (N_4998,N_4236,N_4145);
nor U4999 (N_4999,N_4047,N_4469);
and U5000 (N_5000,N_4670,N_4994);
nand U5001 (N_5001,N_4616,N_4795);
or U5002 (N_5002,N_4708,N_4625);
and U5003 (N_5003,N_4837,N_4594);
and U5004 (N_5004,N_4714,N_4979);
nand U5005 (N_5005,N_4789,N_4623);
xor U5006 (N_5006,N_4915,N_4820);
and U5007 (N_5007,N_4744,N_4530);
and U5008 (N_5008,N_4908,N_4515);
nand U5009 (N_5009,N_4788,N_4597);
nor U5010 (N_5010,N_4936,N_4856);
nand U5011 (N_5011,N_4800,N_4751);
nor U5012 (N_5012,N_4956,N_4650);
and U5013 (N_5013,N_4907,N_4719);
or U5014 (N_5014,N_4881,N_4707);
or U5015 (N_5015,N_4859,N_4666);
nand U5016 (N_5016,N_4521,N_4763);
and U5017 (N_5017,N_4713,N_4639);
nand U5018 (N_5018,N_4547,N_4601);
nor U5019 (N_5019,N_4502,N_4848);
nor U5020 (N_5020,N_4618,N_4636);
nor U5021 (N_5021,N_4775,N_4823);
nand U5022 (N_5022,N_4892,N_4501);
or U5023 (N_5023,N_4790,N_4894);
nor U5024 (N_5024,N_4786,N_4920);
nor U5025 (N_5025,N_4741,N_4614);
xnor U5026 (N_5026,N_4993,N_4922);
nor U5027 (N_5027,N_4628,N_4943);
nor U5028 (N_5028,N_4762,N_4661);
or U5029 (N_5029,N_4598,N_4975);
and U5030 (N_5030,N_4629,N_4553);
nor U5031 (N_5031,N_4978,N_4822);
nand U5032 (N_5032,N_4632,N_4529);
or U5033 (N_5033,N_4753,N_4561);
and U5034 (N_5034,N_4702,N_4906);
nand U5035 (N_5035,N_4738,N_4566);
nand U5036 (N_5036,N_4635,N_4701);
nor U5037 (N_5037,N_4532,N_4793);
and U5038 (N_5038,N_4752,N_4615);
nor U5039 (N_5039,N_4571,N_4682);
and U5040 (N_5040,N_4876,N_4551);
and U5041 (N_5041,N_4930,N_4893);
nor U5042 (N_5042,N_4658,N_4986);
nor U5043 (N_5043,N_4603,N_4558);
xnor U5044 (N_5044,N_4729,N_4630);
or U5045 (N_5045,N_4510,N_4836);
nand U5046 (N_5046,N_4890,N_4649);
nor U5047 (N_5047,N_4883,N_4989);
nor U5048 (N_5048,N_4850,N_4518);
and U5049 (N_5049,N_4681,N_4912);
nand U5050 (N_5050,N_4727,N_4677);
or U5051 (N_5051,N_4562,N_4589);
or U5052 (N_5052,N_4815,N_4716);
xnor U5053 (N_5053,N_4575,N_4634);
nor U5054 (N_5054,N_4605,N_4891);
or U5055 (N_5055,N_4965,N_4916);
and U5056 (N_5056,N_4969,N_4572);
nor U5057 (N_5057,N_4731,N_4573);
nand U5058 (N_5058,N_4869,N_4750);
nand U5059 (N_5059,N_4770,N_4759);
nor U5060 (N_5060,N_4540,N_4581);
and U5061 (N_5061,N_4543,N_4875);
or U5062 (N_5062,N_4609,N_4673);
nor U5063 (N_5063,N_4611,N_4717);
nand U5064 (N_5064,N_4726,N_4797);
nor U5065 (N_5065,N_4966,N_4809);
xnor U5066 (N_5066,N_4805,N_4944);
or U5067 (N_5067,N_4816,N_4980);
and U5068 (N_5068,N_4653,N_4604);
nand U5069 (N_5069,N_4686,N_4842);
or U5070 (N_5070,N_4991,N_4870);
nand U5071 (N_5071,N_4830,N_4563);
nor U5072 (N_5072,N_4997,N_4517);
and U5073 (N_5073,N_4503,N_4829);
nor U5074 (N_5074,N_4919,N_4570);
or U5075 (N_5075,N_4949,N_4678);
and U5076 (N_5076,N_4568,N_4801);
and U5077 (N_5077,N_4525,N_4508);
xor U5078 (N_5078,N_4835,N_4987);
nor U5079 (N_5079,N_4813,N_4712);
or U5080 (N_5080,N_4841,N_4735);
and U5081 (N_5081,N_4971,N_4780);
or U5082 (N_5082,N_4692,N_4698);
nand U5083 (N_5083,N_4847,N_4659);
or U5084 (N_5084,N_4700,N_4642);
or U5085 (N_5085,N_4621,N_4703);
and U5086 (N_5086,N_4882,N_4757);
or U5087 (N_5087,N_4819,N_4524);
and U5088 (N_5088,N_4742,N_4582);
nor U5089 (N_5089,N_4917,N_4981);
nand U5090 (N_5090,N_4544,N_4537);
nor U5091 (N_5091,N_4855,N_4669);
and U5092 (N_5092,N_4909,N_4596);
nor U5093 (N_5093,N_4705,N_4808);
and U5094 (N_5094,N_4671,N_4760);
nand U5095 (N_5095,N_4542,N_4580);
nand U5096 (N_5096,N_4846,N_4948);
or U5097 (N_5097,N_4940,N_4730);
or U5098 (N_5098,N_4693,N_4843);
nand U5099 (N_5099,N_4565,N_4814);
xnor U5100 (N_5100,N_4683,N_4668);
nand U5101 (N_5101,N_4811,N_4807);
or U5102 (N_5102,N_4810,N_4884);
nand U5103 (N_5103,N_4945,N_4783);
or U5104 (N_5104,N_4592,N_4583);
or U5105 (N_5105,N_4796,N_4584);
or U5106 (N_5106,N_4874,N_4858);
and U5107 (N_5107,N_4506,N_4739);
nand U5108 (N_5108,N_4862,N_4748);
nor U5109 (N_5109,N_4754,N_4576);
nand U5110 (N_5110,N_4867,N_4844);
nor U5111 (N_5111,N_4655,N_4756);
nor U5112 (N_5112,N_4764,N_4734);
nand U5113 (N_5113,N_4999,N_4990);
nor U5114 (N_5114,N_4868,N_4888);
nand U5115 (N_5115,N_4982,N_4526);
nand U5116 (N_5116,N_4560,N_4732);
and U5117 (N_5117,N_4545,N_4695);
or U5118 (N_5118,N_4769,N_4672);
and U5119 (N_5119,N_4901,N_4685);
xnor U5120 (N_5120,N_4918,N_4527);
or U5121 (N_5121,N_4593,N_4952);
and U5122 (N_5122,N_4896,N_4995);
or U5123 (N_5123,N_4520,N_4765);
xor U5124 (N_5124,N_4513,N_4897);
nor U5125 (N_5125,N_4531,N_4652);
and U5126 (N_5126,N_4758,N_4784);
nor U5127 (N_5127,N_4976,N_4736);
nand U5128 (N_5128,N_4647,N_4791);
or U5129 (N_5129,N_4509,N_4657);
nor U5130 (N_5130,N_4617,N_4984);
nor U5131 (N_5131,N_4746,N_4539);
and U5132 (N_5132,N_4626,N_4961);
nand U5133 (N_5133,N_4559,N_4675);
or U5134 (N_5134,N_4691,N_4660);
and U5135 (N_5135,N_4610,N_4690);
or U5136 (N_5136,N_4864,N_4887);
or U5137 (N_5137,N_4722,N_4684);
and U5138 (N_5138,N_4885,N_4939);
or U5139 (N_5139,N_4970,N_4895);
nand U5140 (N_5140,N_4812,N_4903);
and U5141 (N_5141,N_4904,N_4724);
and U5142 (N_5142,N_4654,N_4640);
nand U5143 (N_5143,N_4960,N_4926);
nand U5144 (N_5144,N_4612,N_4767);
nand U5145 (N_5145,N_4803,N_4607);
nand U5146 (N_5146,N_4638,N_4555);
and U5147 (N_5147,N_4927,N_4694);
or U5148 (N_5148,N_4535,N_4799);
and U5149 (N_5149,N_4689,N_4905);
or U5150 (N_5150,N_4931,N_4878);
nor U5151 (N_5151,N_4857,N_4910);
nor U5152 (N_5152,N_4785,N_4959);
nand U5153 (N_5153,N_4512,N_4646);
nand U5154 (N_5154,N_4834,N_4504);
nor U5155 (N_5155,N_4911,N_4967);
nand U5156 (N_5156,N_4955,N_4998);
and U5157 (N_5157,N_4947,N_4935);
xnor U5158 (N_5158,N_4633,N_4929);
nor U5159 (N_5159,N_4921,N_4941);
nand U5160 (N_5160,N_4877,N_4715);
and U5161 (N_5161,N_4833,N_4585);
and U5162 (N_5162,N_4866,N_4889);
nor U5163 (N_5163,N_4900,N_4740);
or U5164 (N_5164,N_4554,N_4879);
nand U5165 (N_5165,N_4773,N_4516);
nor U5166 (N_5166,N_4772,N_4950);
nor U5167 (N_5167,N_4792,N_4588);
nor U5168 (N_5168,N_4914,N_4974);
or U5169 (N_5169,N_4579,N_4600);
and U5170 (N_5170,N_4505,N_4865);
and U5171 (N_5171,N_4818,N_4778);
or U5172 (N_5172,N_4802,N_4552);
xor U5173 (N_5173,N_4641,N_4577);
nor U5174 (N_5174,N_4861,N_4608);
nor U5175 (N_5175,N_4710,N_4711);
nand U5176 (N_5176,N_4840,N_4849);
nand U5177 (N_5177,N_4590,N_4680);
nand U5178 (N_5178,N_4992,N_4806);
nand U5179 (N_5179,N_4964,N_4522);
nor U5180 (N_5180,N_4624,N_4873);
nor U5181 (N_5181,N_4782,N_4733);
nor U5182 (N_5182,N_4794,N_4776);
nor U5183 (N_5183,N_4962,N_4709);
and U5184 (N_5184,N_4913,N_4942);
and U5185 (N_5185,N_4871,N_4953);
or U5186 (N_5186,N_4854,N_4860);
and U5187 (N_5187,N_4667,N_4988);
nor U5188 (N_5188,N_4872,N_4523);
or U5189 (N_5189,N_4839,N_4851);
nor U5190 (N_5190,N_4637,N_4721);
nor U5191 (N_5191,N_4899,N_4595);
or U5192 (N_5192,N_4826,N_4804);
or U5193 (N_5193,N_4766,N_4602);
nor U5194 (N_5194,N_4599,N_4699);
and U5195 (N_5195,N_4928,N_4587);
and U5196 (N_5196,N_4737,N_4845);
and U5197 (N_5197,N_4863,N_4674);
nand U5198 (N_5198,N_4781,N_4688);
or U5199 (N_5199,N_4696,N_4706);
nand U5200 (N_5200,N_4679,N_4643);
nor U5201 (N_5201,N_4852,N_4951);
xor U5202 (N_5202,N_4968,N_4687);
or U5203 (N_5203,N_4645,N_4656);
or U5204 (N_5204,N_4983,N_4723);
and U5205 (N_5205,N_4676,N_4924);
nand U5206 (N_5206,N_4880,N_4923);
xor U5207 (N_5207,N_4534,N_4768);
nand U5208 (N_5208,N_4821,N_4591);
or U5209 (N_5209,N_4946,N_4662);
nor U5210 (N_5210,N_4771,N_4550);
nand U5211 (N_5211,N_4720,N_4925);
and U5212 (N_5212,N_4564,N_4958);
or U5213 (N_5213,N_4831,N_4761);
and U5214 (N_5214,N_4957,N_4697);
nor U5215 (N_5215,N_4567,N_4937);
or U5216 (N_5216,N_4934,N_4832);
or U5217 (N_5217,N_4824,N_4549);
nand U5218 (N_5218,N_4500,N_4644);
nand U5219 (N_5219,N_4725,N_4973);
and U5220 (N_5220,N_4798,N_4541);
or U5221 (N_5221,N_4665,N_4507);
nand U5222 (N_5222,N_4619,N_4546);
or U5223 (N_5223,N_4886,N_4779);
nor U5224 (N_5224,N_4996,N_4774);
and U5225 (N_5225,N_4648,N_4743);
or U5226 (N_5226,N_4972,N_4745);
and U5227 (N_5227,N_4606,N_4627);
nand U5228 (N_5228,N_4519,N_4985);
nand U5229 (N_5229,N_4574,N_4569);
or U5230 (N_5230,N_4511,N_4578);
nor U5231 (N_5231,N_4663,N_4536);
nor U5232 (N_5232,N_4718,N_4977);
or U5233 (N_5233,N_4817,N_4777);
and U5234 (N_5234,N_4613,N_4514);
and U5235 (N_5235,N_4749,N_4853);
and U5236 (N_5236,N_4932,N_4938);
nand U5237 (N_5237,N_4828,N_4664);
or U5238 (N_5238,N_4827,N_4557);
nor U5239 (N_5239,N_4954,N_4898);
and U5240 (N_5240,N_4548,N_4533);
nand U5241 (N_5241,N_4620,N_4556);
and U5242 (N_5242,N_4902,N_4586);
nand U5243 (N_5243,N_4631,N_4728);
nand U5244 (N_5244,N_4538,N_4838);
nor U5245 (N_5245,N_4755,N_4528);
or U5246 (N_5246,N_4825,N_4704);
nor U5247 (N_5247,N_4933,N_4622);
nor U5248 (N_5248,N_4747,N_4651);
nor U5249 (N_5249,N_4787,N_4963);
and U5250 (N_5250,N_4537,N_4893);
nor U5251 (N_5251,N_4778,N_4988);
nand U5252 (N_5252,N_4750,N_4639);
or U5253 (N_5253,N_4863,N_4506);
and U5254 (N_5254,N_4704,N_4554);
and U5255 (N_5255,N_4739,N_4718);
or U5256 (N_5256,N_4638,N_4642);
nand U5257 (N_5257,N_4782,N_4854);
nand U5258 (N_5258,N_4922,N_4861);
or U5259 (N_5259,N_4647,N_4508);
or U5260 (N_5260,N_4510,N_4957);
and U5261 (N_5261,N_4783,N_4587);
nor U5262 (N_5262,N_4619,N_4514);
or U5263 (N_5263,N_4571,N_4741);
nand U5264 (N_5264,N_4746,N_4737);
nor U5265 (N_5265,N_4521,N_4685);
xor U5266 (N_5266,N_4519,N_4958);
nand U5267 (N_5267,N_4934,N_4882);
xnor U5268 (N_5268,N_4696,N_4734);
nor U5269 (N_5269,N_4600,N_4926);
and U5270 (N_5270,N_4952,N_4607);
nand U5271 (N_5271,N_4992,N_4651);
nor U5272 (N_5272,N_4727,N_4956);
and U5273 (N_5273,N_4608,N_4853);
or U5274 (N_5274,N_4639,N_4643);
and U5275 (N_5275,N_4748,N_4510);
and U5276 (N_5276,N_4509,N_4649);
or U5277 (N_5277,N_4822,N_4976);
and U5278 (N_5278,N_4519,N_4556);
nand U5279 (N_5279,N_4892,N_4904);
or U5280 (N_5280,N_4568,N_4627);
or U5281 (N_5281,N_4944,N_4899);
or U5282 (N_5282,N_4664,N_4804);
nor U5283 (N_5283,N_4958,N_4921);
nand U5284 (N_5284,N_4981,N_4727);
nor U5285 (N_5285,N_4525,N_4719);
nor U5286 (N_5286,N_4733,N_4942);
or U5287 (N_5287,N_4611,N_4989);
nand U5288 (N_5288,N_4814,N_4799);
and U5289 (N_5289,N_4892,N_4792);
nand U5290 (N_5290,N_4593,N_4920);
xnor U5291 (N_5291,N_4953,N_4548);
or U5292 (N_5292,N_4987,N_4800);
or U5293 (N_5293,N_4875,N_4863);
nor U5294 (N_5294,N_4549,N_4800);
and U5295 (N_5295,N_4577,N_4824);
nor U5296 (N_5296,N_4921,N_4982);
nand U5297 (N_5297,N_4628,N_4529);
or U5298 (N_5298,N_4894,N_4900);
or U5299 (N_5299,N_4842,N_4818);
and U5300 (N_5300,N_4667,N_4953);
nand U5301 (N_5301,N_4589,N_4676);
and U5302 (N_5302,N_4719,N_4820);
or U5303 (N_5303,N_4829,N_4523);
nand U5304 (N_5304,N_4709,N_4922);
nor U5305 (N_5305,N_4631,N_4815);
or U5306 (N_5306,N_4850,N_4811);
nor U5307 (N_5307,N_4666,N_4955);
or U5308 (N_5308,N_4695,N_4577);
nand U5309 (N_5309,N_4540,N_4805);
nor U5310 (N_5310,N_4581,N_4956);
and U5311 (N_5311,N_4654,N_4823);
and U5312 (N_5312,N_4963,N_4768);
nor U5313 (N_5313,N_4803,N_4552);
and U5314 (N_5314,N_4962,N_4940);
or U5315 (N_5315,N_4555,N_4593);
nor U5316 (N_5316,N_4790,N_4770);
or U5317 (N_5317,N_4977,N_4571);
nor U5318 (N_5318,N_4581,N_4534);
nor U5319 (N_5319,N_4840,N_4796);
and U5320 (N_5320,N_4502,N_4582);
nand U5321 (N_5321,N_4746,N_4844);
nand U5322 (N_5322,N_4621,N_4826);
nand U5323 (N_5323,N_4919,N_4629);
nand U5324 (N_5324,N_4831,N_4976);
or U5325 (N_5325,N_4562,N_4888);
nor U5326 (N_5326,N_4788,N_4817);
nand U5327 (N_5327,N_4521,N_4627);
and U5328 (N_5328,N_4663,N_4807);
nand U5329 (N_5329,N_4768,N_4984);
and U5330 (N_5330,N_4733,N_4743);
nor U5331 (N_5331,N_4540,N_4967);
xnor U5332 (N_5332,N_4766,N_4904);
nor U5333 (N_5333,N_4582,N_4865);
nor U5334 (N_5334,N_4799,N_4899);
and U5335 (N_5335,N_4644,N_4636);
and U5336 (N_5336,N_4685,N_4774);
nand U5337 (N_5337,N_4754,N_4777);
and U5338 (N_5338,N_4771,N_4622);
nand U5339 (N_5339,N_4760,N_4931);
nand U5340 (N_5340,N_4925,N_4894);
nand U5341 (N_5341,N_4882,N_4777);
nor U5342 (N_5342,N_4685,N_4844);
nor U5343 (N_5343,N_4749,N_4768);
nand U5344 (N_5344,N_4776,N_4969);
or U5345 (N_5345,N_4943,N_4823);
nor U5346 (N_5346,N_4539,N_4837);
nor U5347 (N_5347,N_4888,N_4845);
nor U5348 (N_5348,N_4625,N_4966);
or U5349 (N_5349,N_4672,N_4863);
or U5350 (N_5350,N_4910,N_4611);
nand U5351 (N_5351,N_4502,N_4866);
nand U5352 (N_5352,N_4643,N_4910);
or U5353 (N_5353,N_4741,N_4856);
nor U5354 (N_5354,N_4760,N_4785);
and U5355 (N_5355,N_4818,N_4997);
nand U5356 (N_5356,N_4851,N_4848);
nor U5357 (N_5357,N_4747,N_4902);
nand U5358 (N_5358,N_4791,N_4792);
nand U5359 (N_5359,N_4846,N_4703);
or U5360 (N_5360,N_4958,N_4622);
nor U5361 (N_5361,N_4945,N_4623);
nor U5362 (N_5362,N_4556,N_4964);
nand U5363 (N_5363,N_4710,N_4940);
or U5364 (N_5364,N_4922,N_4551);
nor U5365 (N_5365,N_4865,N_4938);
nor U5366 (N_5366,N_4749,N_4829);
or U5367 (N_5367,N_4787,N_4832);
or U5368 (N_5368,N_4659,N_4831);
nor U5369 (N_5369,N_4850,N_4865);
nor U5370 (N_5370,N_4935,N_4828);
nand U5371 (N_5371,N_4975,N_4906);
nand U5372 (N_5372,N_4859,N_4920);
and U5373 (N_5373,N_4645,N_4598);
nor U5374 (N_5374,N_4756,N_4760);
or U5375 (N_5375,N_4910,N_4833);
nor U5376 (N_5376,N_4881,N_4878);
or U5377 (N_5377,N_4663,N_4566);
or U5378 (N_5378,N_4529,N_4987);
nor U5379 (N_5379,N_4906,N_4661);
and U5380 (N_5380,N_4709,N_4905);
nor U5381 (N_5381,N_4703,N_4827);
nand U5382 (N_5382,N_4689,N_4645);
nor U5383 (N_5383,N_4530,N_4753);
and U5384 (N_5384,N_4616,N_4571);
nor U5385 (N_5385,N_4605,N_4680);
xor U5386 (N_5386,N_4771,N_4539);
and U5387 (N_5387,N_4565,N_4556);
and U5388 (N_5388,N_4548,N_4529);
or U5389 (N_5389,N_4531,N_4947);
and U5390 (N_5390,N_4934,N_4635);
nor U5391 (N_5391,N_4910,N_4993);
xnor U5392 (N_5392,N_4852,N_4945);
nand U5393 (N_5393,N_4587,N_4745);
nand U5394 (N_5394,N_4732,N_4593);
nor U5395 (N_5395,N_4796,N_4593);
nand U5396 (N_5396,N_4726,N_4810);
nand U5397 (N_5397,N_4567,N_4678);
and U5398 (N_5398,N_4603,N_4632);
or U5399 (N_5399,N_4827,N_4767);
nor U5400 (N_5400,N_4851,N_4568);
and U5401 (N_5401,N_4905,N_4575);
nand U5402 (N_5402,N_4587,N_4998);
nor U5403 (N_5403,N_4677,N_4944);
nor U5404 (N_5404,N_4845,N_4791);
or U5405 (N_5405,N_4644,N_4637);
or U5406 (N_5406,N_4745,N_4955);
xor U5407 (N_5407,N_4502,N_4685);
nor U5408 (N_5408,N_4729,N_4981);
xnor U5409 (N_5409,N_4855,N_4992);
nand U5410 (N_5410,N_4646,N_4890);
or U5411 (N_5411,N_4883,N_4776);
nand U5412 (N_5412,N_4639,N_4823);
nand U5413 (N_5413,N_4648,N_4803);
or U5414 (N_5414,N_4948,N_4909);
nand U5415 (N_5415,N_4871,N_4703);
nand U5416 (N_5416,N_4932,N_4502);
and U5417 (N_5417,N_4800,N_4779);
or U5418 (N_5418,N_4552,N_4706);
xor U5419 (N_5419,N_4835,N_4753);
xor U5420 (N_5420,N_4805,N_4916);
or U5421 (N_5421,N_4951,N_4903);
or U5422 (N_5422,N_4843,N_4890);
and U5423 (N_5423,N_4610,N_4679);
and U5424 (N_5424,N_4762,N_4544);
nand U5425 (N_5425,N_4834,N_4563);
or U5426 (N_5426,N_4805,N_4567);
nand U5427 (N_5427,N_4731,N_4572);
nor U5428 (N_5428,N_4715,N_4787);
xor U5429 (N_5429,N_4606,N_4777);
nand U5430 (N_5430,N_4972,N_4529);
nand U5431 (N_5431,N_4509,N_4613);
and U5432 (N_5432,N_4805,N_4832);
nand U5433 (N_5433,N_4568,N_4547);
and U5434 (N_5434,N_4712,N_4935);
nor U5435 (N_5435,N_4767,N_4747);
or U5436 (N_5436,N_4654,N_4701);
nor U5437 (N_5437,N_4603,N_4586);
nor U5438 (N_5438,N_4653,N_4940);
or U5439 (N_5439,N_4709,N_4582);
nand U5440 (N_5440,N_4500,N_4622);
nand U5441 (N_5441,N_4529,N_4768);
or U5442 (N_5442,N_4849,N_4603);
nor U5443 (N_5443,N_4672,N_4732);
or U5444 (N_5444,N_4971,N_4635);
or U5445 (N_5445,N_4688,N_4660);
nand U5446 (N_5446,N_4811,N_4869);
and U5447 (N_5447,N_4803,N_4831);
nand U5448 (N_5448,N_4818,N_4977);
nor U5449 (N_5449,N_4617,N_4768);
and U5450 (N_5450,N_4899,N_4932);
nand U5451 (N_5451,N_4879,N_4804);
and U5452 (N_5452,N_4558,N_4589);
or U5453 (N_5453,N_4816,N_4817);
or U5454 (N_5454,N_4787,N_4916);
xnor U5455 (N_5455,N_4872,N_4538);
nand U5456 (N_5456,N_4895,N_4712);
and U5457 (N_5457,N_4820,N_4909);
nor U5458 (N_5458,N_4750,N_4792);
or U5459 (N_5459,N_4682,N_4804);
or U5460 (N_5460,N_4882,N_4869);
and U5461 (N_5461,N_4798,N_4646);
or U5462 (N_5462,N_4922,N_4637);
or U5463 (N_5463,N_4539,N_4759);
nor U5464 (N_5464,N_4546,N_4914);
or U5465 (N_5465,N_4938,N_4811);
and U5466 (N_5466,N_4750,N_4891);
nor U5467 (N_5467,N_4645,N_4922);
and U5468 (N_5468,N_4544,N_4855);
or U5469 (N_5469,N_4755,N_4823);
or U5470 (N_5470,N_4698,N_4831);
or U5471 (N_5471,N_4674,N_4756);
nand U5472 (N_5472,N_4501,N_4855);
and U5473 (N_5473,N_4673,N_4579);
nand U5474 (N_5474,N_4770,N_4661);
nand U5475 (N_5475,N_4800,N_4613);
or U5476 (N_5476,N_4652,N_4787);
nor U5477 (N_5477,N_4699,N_4978);
and U5478 (N_5478,N_4715,N_4785);
nor U5479 (N_5479,N_4629,N_4669);
xnor U5480 (N_5480,N_4837,N_4844);
or U5481 (N_5481,N_4621,N_4961);
or U5482 (N_5482,N_4521,N_4910);
nor U5483 (N_5483,N_4902,N_4749);
and U5484 (N_5484,N_4900,N_4636);
and U5485 (N_5485,N_4729,N_4612);
and U5486 (N_5486,N_4845,N_4531);
xor U5487 (N_5487,N_4623,N_4516);
xnor U5488 (N_5488,N_4618,N_4660);
nand U5489 (N_5489,N_4793,N_4829);
nand U5490 (N_5490,N_4846,N_4907);
nand U5491 (N_5491,N_4692,N_4773);
nor U5492 (N_5492,N_4880,N_4740);
nand U5493 (N_5493,N_4712,N_4577);
nand U5494 (N_5494,N_4663,N_4886);
nand U5495 (N_5495,N_4693,N_4839);
and U5496 (N_5496,N_4934,N_4831);
nor U5497 (N_5497,N_4769,N_4995);
or U5498 (N_5498,N_4763,N_4731);
nand U5499 (N_5499,N_4594,N_4792);
and U5500 (N_5500,N_5427,N_5151);
nand U5501 (N_5501,N_5159,N_5443);
nor U5502 (N_5502,N_5267,N_5055);
and U5503 (N_5503,N_5147,N_5431);
and U5504 (N_5504,N_5009,N_5010);
and U5505 (N_5505,N_5488,N_5471);
nand U5506 (N_5506,N_5350,N_5412);
nand U5507 (N_5507,N_5453,N_5014);
or U5508 (N_5508,N_5152,N_5142);
or U5509 (N_5509,N_5302,N_5292);
and U5510 (N_5510,N_5325,N_5202);
nor U5511 (N_5511,N_5176,N_5163);
nor U5512 (N_5512,N_5063,N_5253);
and U5513 (N_5513,N_5106,N_5269);
or U5514 (N_5514,N_5383,N_5463);
and U5515 (N_5515,N_5333,N_5149);
and U5516 (N_5516,N_5284,N_5005);
or U5517 (N_5517,N_5229,N_5354);
nor U5518 (N_5518,N_5286,N_5217);
nor U5519 (N_5519,N_5037,N_5456);
or U5520 (N_5520,N_5128,N_5296);
nand U5521 (N_5521,N_5061,N_5119);
or U5522 (N_5522,N_5421,N_5281);
nand U5523 (N_5523,N_5068,N_5365);
nand U5524 (N_5524,N_5209,N_5023);
or U5525 (N_5525,N_5204,N_5411);
nor U5526 (N_5526,N_5091,N_5348);
or U5527 (N_5527,N_5392,N_5353);
xor U5528 (N_5528,N_5417,N_5024);
and U5529 (N_5529,N_5072,N_5025);
nor U5530 (N_5530,N_5377,N_5442);
and U5531 (N_5531,N_5356,N_5224);
or U5532 (N_5532,N_5195,N_5329);
nand U5533 (N_5533,N_5225,N_5248);
and U5534 (N_5534,N_5324,N_5002);
or U5535 (N_5535,N_5041,N_5309);
xor U5536 (N_5536,N_5180,N_5045);
nand U5537 (N_5537,N_5315,N_5227);
xnor U5538 (N_5538,N_5008,N_5319);
or U5539 (N_5539,N_5215,N_5028);
or U5540 (N_5540,N_5337,N_5207);
or U5541 (N_5541,N_5059,N_5481);
and U5542 (N_5542,N_5379,N_5385);
nor U5543 (N_5543,N_5439,N_5485);
and U5544 (N_5544,N_5219,N_5054);
or U5545 (N_5545,N_5369,N_5484);
and U5546 (N_5546,N_5079,N_5170);
and U5547 (N_5547,N_5285,N_5032);
nand U5548 (N_5548,N_5083,N_5130);
or U5549 (N_5549,N_5346,N_5342);
or U5550 (N_5550,N_5373,N_5251);
or U5551 (N_5551,N_5073,N_5069);
and U5552 (N_5552,N_5468,N_5496);
or U5553 (N_5553,N_5189,N_5276);
or U5554 (N_5554,N_5165,N_5361);
or U5555 (N_5555,N_5378,N_5179);
and U5556 (N_5556,N_5199,N_5455);
and U5557 (N_5557,N_5287,N_5234);
and U5558 (N_5558,N_5164,N_5338);
nand U5559 (N_5559,N_5418,N_5306);
and U5560 (N_5560,N_5092,N_5283);
or U5561 (N_5561,N_5186,N_5425);
nand U5562 (N_5562,N_5031,N_5039);
nor U5563 (N_5563,N_5133,N_5101);
or U5564 (N_5564,N_5310,N_5080);
nor U5565 (N_5565,N_5398,N_5191);
or U5566 (N_5566,N_5071,N_5479);
nor U5567 (N_5567,N_5146,N_5026);
nor U5568 (N_5568,N_5150,N_5428);
and U5569 (N_5569,N_5019,N_5016);
or U5570 (N_5570,N_5331,N_5095);
nand U5571 (N_5571,N_5438,N_5339);
and U5572 (N_5572,N_5279,N_5345);
nor U5573 (N_5573,N_5047,N_5465);
and U5574 (N_5574,N_5247,N_5249);
and U5575 (N_5575,N_5052,N_5185);
nand U5576 (N_5576,N_5211,N_5067);
nand U5577 (N_5577,N_5498,N_5275);
or U5578 (N_5578,N_5006,N_5178);
and U5579 (N_5579,N_5405,N_5305);
or U5580 (N_5580,N_5136,N_5493);
and U5581 (N_5581,N_5492,N_5018);
nor U5582 (N_5582,N_5115,N_5138);
or U5583 (N_5583,N_5413,N_5486);
nand U5584 (N_5584,N_5237,N_5386);
and U5585 (N_5585,N_5436,N_5460);
nand U5586 (N_5586,N_5260,N_5221);
or U5587 (N_5587,N_5371,N_5196);
nand U5588 (N_5588,N_5020,N_5289);
and U5589 (N_5589,N_5173,N_5190);
nand U5590 (N_5590,N_5034,N_5074);
or U5591 (N_5591,N_5084,N_5473);
nor U5592 (N_5592,N_5222,N_5408);
nand U5593 (N_5593,N_5332,N_5394);
or U5594 (N_5594,N_5096,N_5352);
nand U5595 (N_5595,N_5452,N_5192);
or U5596 (N_5596,N_5304,N_5022);
nand U5597 (N_5597,N_5391,N_5334);
or U5598 (N_5598,N_5193,N_5044);
nand U5599 (N_5599,N_5000,N_5432);
and U5600 (N_5600,N_5087,N_5001);
and U5601 (N_5601,N_5297,N_5499);
and U5602 (N_5602,N_5349,N_5291);
nand U5603 (N_5603,N_5467,N_5184);
and U5604 (N_5604,N_5321,N_5375);
nor U5605 (N_5605,N_5316,N_5104);
nor U5606 (N_5606,N_5478,N_5343);
or U5607 (N_5607,N_5301,N_5447);
nand U5608 (N_5608,N_5200,N_5030);
nand U5609 (N_5609,N_5144,N_5490);
nand U5610 (N_5610,N_5230,N_5078);
nor U5611 (N_5611,N_5434,N_5457);
and U5612 (N_5612,N_5308,N_5422);
or U5613 (N_5613,N_5414,N_5216);
and U5614 (N_5614,N_5435,N_5395);
xnor U5615 (N_5615,N_5111,N_5218);
or U5616 (N_5616,N_5317,N_5363);
nand U5617 (N_5617,N_5158,N_5433);
and U5618 (N_5618,N_5359,N_5131);
nor U5619 (N_5619,N_5497,N_5208);
or U5620 (N_5620,N_5077,N_5407);
or U5621 (N_5621,N_5271,N_5042);
nand U5622 (N_5622,N_5265,N_5241);
and U5623 (N_5623,N_5326,N_5154);
or U5624 (N_5624,N_5261,N_5036);
nor U5625 (N_5625,N_5420,N_5277);
nand U5626 (N_5626,N_5451,N_5127);
and U5627 (N_5627,N_5172,N_5288);
and U5628 (N_5628,N_5233,N_5226);
and U5629 (N_5629,N_5058,N_5043);
or U5630 (N_5630,N_5065,N_5303);
or U5631 (N_5631,N_5480,N_5344);
nand U5632 (N_5632,N_5116,N_5290);
nor U5633 (N_5633,N_5174,N_5476);
nor U5634 (N_5634,N_5125,N_5475);
nor U5635 (N_5635,N_5187,N_5168);
or U5636 (N_5636,N_5491,N_5089);
and U5637 (N_5637,N_5238,N_5135);
and U5638 (N_5638,N_5293,N_5424);
or U5639 (N_5639,N_5007,N_5099);
or U5640 (N_5640,N_5462,N_5155);
or U5641 (N_5641,N_5409,N_5390);
xor U5642 (N_5642,N_5143,N_5198);
and U5643 (N_5643,N_5017,N_5206);
or U5644 (N_5644,N_5210,N_5214);
nand U5645 (N_5645,N_5157,N_5094);
nor U5646 (N_5646,N_5445,N_5254);
or U5647 (N_5647,N_5410,N_5416);
nand U5648 (N_5648,N_5160,N_5235);
or U5649 (N_5649,N_5278,N_5320);
or U5650 (N_5650,N_5323,N_5300);
nand U5651 (N_5651,N_5062,N_5013);
and U5652 (N_5652,N_5360,N_5403);
nor U5653 (N_5653,N_5366,N_5312);
nand U5654 (N_5654,N_5162,N_5169);
nor U5655 (N_5655,N_5437,N_5213);
or U5656 (N_5656,N_5057,N_5470);
nor U5657 (N_5657,N_5440,N_5181);
and U5658 (N_5658,N_5085,N_5256);
nand U5659 (N_5659,N_5220,N_5401);
nand U5660 (N_5660,N_5134,N_5141);
nor U5661 (N_5661,N_5194,N_5129);
and U5662 (N_5662,N_5376,N_5011);
or U5663 (N_5663,N_5108,N_5252);
and U5664 (N_5664,N_5123,N_5228);
nand U5665 (N_5665,N_5171,N_5430);
or U5666 (N_5666,N_5464,N_5050);
nand U5667 (N_5667,N_5311,N_5029);
or U5668 (N_5668,N_5120,N_5419);
and U5669 (N_5669,N_5081,N_5448);
nand U5670 (N_5670,N_5429,N_5066);
nor U5671 (N_5671,N_5474,N_5015);
xor U5672 (N_5672,N_5027,N_5082);
nand U5673 (N_5673,N_5070,N_5075);
or U5674 (N_5674,N_5482,N_5076);
nor U5675 (N_5675,N_5355,N_5167);
or U5676 (N_5676,N_5231,N_5166);
nand U5677 (N_5677,N_5175,N_5212);
nor U5678 (N_5678,N_5381,N_5100);
or U5679 (N_5679,N_5327,N_5380);
nand U5680 (N_5680,N_5335,N_5357);
and U5681 (N_5681,N_5270,N_5124);
or U5682 (N_5682,N_5203,N_5090);
nand U5683 (N_5683,N_5459,N_5280);
or U5684 (N_5684,N_5415,N_5258);
or U5685 (N_5685,N_5046,N_5243);
nand U5686 (N_5686,N_5003,N_5012);
or U5687 (N_5687,N_5040,N_5097);
and U5688 (N_5688,N_5004,N_5188);
nor U5689 (N_5689,N_5384,N_5367);
nand U5690 (N_5690,N_5259,N_5400);
or U5691 (N_5691,N_5139,N_5368);
nand U5692 (N_5692,N_5223,N_5295);
and U5693 (N_5693,N_5033,N_5268);
nor U5694 (N_5694,N_5035,N_5298);
nor U5695 (N_5695,N_5201,N_5406);
nand U5696 (N_5696,N_5402,N_5318);
nor U5697 (N_5697,N_5093,N_5105);
nor U5698 (N_5698,N_5145,N_5107);
or U5699 (N_5699,N_5262,N_5274);
nand U5700 (N_5700,N_5053,N_5264);
nand U5701 (N_5701,N_5049,N_5336);
and U5702 (N_5702,N_5487,N_5494);
or U5703 (N_5703,N_5399,N_5404);
or U5704 (N_5704,N_5244,N_5454);
and U5705 (N_5705,N_5477,N_5382);
nor U5706 (N_5706,N_5372,N_5118);
nand U5707 (N_5707,N_5362,N_5132);
nand U5708 (N_5708,N_5250,N_5266);
nor U5709 (N_5709,N_5060,N_5197);
or U5710 (N_5710,N_5396,N_5472);
or U5711 (N_5711,N_5177,N_5364);
and U5712 (N_5712,N_5441,N_5088);
xnor U5713 (N_5713,N_5246,N_5126);
nor U5714 (N_5714,N_5112,N_5347);
or U5715 (N_5715,N_5450,N_5183);
or U5716 (N_5716,N_5466,N_5423);
nor U5717 (N_5717,N_5117,N_5294);
nor U5718 (N_5718,N_5370,N_5140);
or U5719 (N_5719,N_5389,N_5449);
and U5720 (N_5720,N_5148,N_5240);
nor U5721 (N_5721,N_5205,N_5358);
nand U5722 (N_5722,N_5495,N_5299);
and U5723 (N_5723,N_5374,N_5489);
nand U5724 (N_5724,N_5110,N_5257);
nand U5725 (N_5725,N_5102,N_5388);
nand U5726 (N_5726,N_5182,N_5340);
or U5727 (N_5727,N_5313,N_5113);
or U5728 (N_5728,N_5137,N_5387);
and U5729 (N_5729,N_5341,N_5397);
or U5730 (N_5730,N_5056,N_5446);
nor U5731 (N_5731,N_5236,N_5328);
or U5732 (N_5732,N_5314,N_5461);
nand U5733 (N_5733,N_5263,N_5121);
nand U5734 (N_5734,N_5048,N_5239);
nand U5735 (N_5735,N_5156,N_5255);
nand U5736 (N_5736,N_5122,N_5086);
nand U5737 (N_5737,N_5426,N_5161);
nor U5738 (N_5738,N_5098,N_5109);
nor U5739 (N_5739,N_5351,N_5232);
or U5740 (N_5740,N_5242,N_5245);
nor U5741 (N_5741,N_5444,N_5458);
or U5742 (N_5742,N_5064,N_5393);
nand U5743 (N_5743,N_5330,N_5153);
or U5744 (N_5744,N_5051,N_5282);
and U5745 (N_5745,N_5307,N_5483);
and U5746 (N_5746,N_5021,N_5103);
nor U5747 (N_5747,N_5114,N_5273);
and U5748 (N_5748,N_5038,N_5322);
and U5749 (N_5749,N_5469,N_5272);
nand U5750 (N_5750,N_5095,N_5395);
nor U5751 (N_5751,N_5240,N_5138);
and U5752 (N_5752,N_5221,N_5061);
nand U5753 (N_5753,N_5146,N_5179);
nor U5754 (N_5754,N_5164,N_5281);
and U5755 (N_5755,N_5110,N_5057);
nor U5756 (N_5756,N_5215,N_5418);
or U5757 (N_5757,N_5161,N_5121);
nand U5758 (N_5758,N_5216,N_5044);
or U5759 (N_5759,N_5007,N_5450);
nand U5760 (N_5760,N_5019,N_5030);
nand U5761 (N_5761,N_5126,N_5105);
or U5762 (N_5762,N_5217,N_5386);
or U5763 (N_5763,N_5393,N_5454);
nand U5764 (N_5764,N_5415,N_5073);
and U5765 (N_5765,N_5315,N_5440);
or U5766 (N_5766,N_5498,N_5224);
and U5767 (N_5767,N_5243,N_5063);
nand U5768 (N_5768,N_5225,N_5127);
nand U5769 (N_5769,N_5283,N_5352);
nand U5770 (N_5770,N_5058,N_5081);
or U5771 (N_5771,N_5188,N_5307);
or U5772 (N_5772,N_5336,N_5368);
or U5773 (N_5773,N_5063,N_5397);
and U5774 (N_5774,N_5377,N_5274);
or U5775 (N_5775,N_5454,N_5368);
and U5776 (N_5776,N_5355,N_5087);
and U5777 (N_5777,N_5294,N_5482);
nand U5778 (N_5778,N_5155,N_5309);
and U5779 (N_5779,N_5391,N_5180);
and U5780 (N_5780,N_5431,N_5020);
nand U5781 (N_5781,N_5421,N_5465);
and U5782 (N_5782,N_5407,N_5078);
or U5783 (N_5783,N_5422,N_5025);
or U5784 (N_5784,N_5434,N_5115);
nand U5785 (N_5785,N_5125,N_5191);
or U5786 (N_5786,N_5058,N_5389);
and U5787 (N_5787,N_5498,N_5420);
or U5788 (N_5788,N_5128,N_5343);
or U5789 (N_5789,N_5427,N_5360);
and U5790 (N_5790,N_5388,N_5464);
or U5791 (N_5791,N_5197,N_5236);
or U5792 (N_5792,N_5413,N_5150);
nor U5793 (N_5793,N_5401,N_5496);
nand U5794 (N_5794,N_5323,N_5371);
or U5795 (N_5795,N_5008,N_5368);
or U5796 (N_5796,N_5266,N_5249);
and U5797 (N_5797,N_5157,N_5484);
nand U5798 (N_5798,N_5097,N_5416);
nor U5799 (N_5799,N_5158,N_5282);
and U5800 (N_5800,N_5170,N_5297);
or U5801 (N_5801,N_5039,N_5304);
nor U5802 (N_5802,N_5281,N_5335);
nand U5803 (N_5803,N_5107,N_5392);
nand U5804 (N_5804,N_5309,N_5460);
and U5805 (N_5805,N_5475,N_5285);
and U5806 (N_5806,N_5081,N_5461);
nor U5807 (N_5807,N_5395,N_5027);
or U5808 (N_5808,N_5498,N_5132);
nor U5809 (N_5809,N_5038,N_5434);
or U5810 (N_5810,N_5068,N_5488);
and U5811 (N_5811,N_5155,N_5356);
nor U5812 (N_5812,N_5066,N_5100);
or U5813 (N_5813,N_5020,N_5287);
or U5814 (N_5814,N_5494,N_5060);
nor U5815 (N_5815,N_5268,N_5077);
and U5816 (N_5816,N_5286,N_5177);
or U5817 (N_5817,N_5429,N_5439);
nand U5818 (N_5818,N_5387,N_5293);
nor U5819 (N_5819,N_5345,N_5036);
and U5820 (N_5820,N_5432,N_5264);
or U5821 (N_5821,N_5272,N_5101);
or U5822 (N_5822,N_5324,N_5194);
nand U5823 (N_5823,N_5339,N_5478);
nor U5824 (N_5824,N_5440,N_5157);
or U5825 (N_5825,N_5199,N_5484);
or U5826 (N_5826,N_5200,N_5155);
nor U5827 (N_5827,N_5388,N_5161);
or U5828 (N_5828,N_5133,N_5013);
and U5829 (N_5829,N_5180,N_5079);
nor U5830 (N_5830,N_5471,N_5348);
nand U5831 (N_5831,N_5001,N_5390);
nand U5832 (N_5832,N_5496,N_5291);
nand U5833 (N_5833,N_5286,N_5245);
nand U5834 (N_5834,N_5073,N_5182);
nor U5835 (N_5835,N_5215,N_5404);
nand U5836 (N_5836,N_5332,N_5406);
and U5837 (N_5837,N_5463,N_5373);
or U5838 (N_5838,N_5102,N_5313);
or U5839 (N_5839,N_5398,N_5016);
and U5840 (N_5840,N_5361,N_5150);
nand U5841 (N_5841,N_5286,N_5142);
nand U5842 (N_5842,N_5226,N_5136);
and U5843 (N_5843,N_5236,N_5490);
nand U5844 (N_5844,N_5021,N_5434);
nor U5845 (N_5845,N_5012,N_5436);
xnor U5846 (N_5846,N_5088,N_5141);
nand U5847 (N_5847,N_5010,N_5013);
or U5848 (N_5848,N_5347,N_5114);
nor U5849 (N_5849,N_5101,N_5368);
and U5850 (N_5850,N_5256,N_5015);
or U5851 (N_5851,N_5431,N_5289);
nand U5852 (N_5852,N_5374,N_5243);
and U5853 (N_5853,N_5458,N_5286);
or U5854 (N_5854,N_5195,N_5412);
nand U5855 (N_5855,N_5281,N_5380);
nor U5856 (N_5856,N_5443,N_5173);
or U5857 (N_5857,N_5248,N_5378);
nor U5858 (N_5858,N_5497,N_5320);
xor U5859 (N_5859,N_5300,N_5384);
nor U5860 (N_5860,N_5423,N_5379);
or U5861 (N_5861,N_5329,N_5357);
and U5862 (N_5862,N_5317,N_5257);
or U5863 (N_5863,N_5148,N_5434);
nor U5864 (N_5864,N_5460,N_5496);
nand U5865 (N_5865,N_5472,N_5225);
and U5866 (N_5866,N_5129,N_5120);
nand U5867 (N_5867,N_5277,N_5407);
or U5868 (N_5868,N_5484,N_5349);
nand U5869 (N_5869,N_5481,N_5387);
and U5870 (N_5870,N_5076,N_5067);
nor U5871 (N_5871,N_5395,N_5349);
and U5872 (N_5872,N_5150,N_5358);
or U5873 (N_5873,N_5108,N_5206);
and U5874 (N_5874,N_5494,N_5379);
or U5875 (N_5875,N_5333,N_5021);
or U5876 (N_5876,N_5031,N_5310);
and U5877 (N_5877,N_5424,N_5491);
nor U5878 (N_5878,N_5241,N_5268);
and U5879 (N_5879,N_5475,N_5451);
nand U5880 (N_5880,N_5208,N_5112);
and U5881 (N_5881,N_5138,N_5463);
nor U5882 (N_5882,N_5136,N_5437);
nand U5883 (N_5883,N_5384,N_5202);
nor U5884 (N_5884,N_5058,N_5234);
nand U5885 (N_5885,N_5217,N_5080);
nand U5886 (N_5886,N_5479,N_5070);
and U5887 (N_5887,N_5456,N_5094);
or U5888 (N_5888,N_5131,N_5331);
or U5889 (N_5889,N_5231,N_5240);
and U5890 (N_5890,N_5218,N_5235);
nand U5891 (N_5891,N_5344,N_5387);
or U5892 (N_5892,N_5249,N_5260);
or U5893 (N_5893,N_5395,N_5028);
nand U5894 (N_5894,N_5022,N_5377);
nor U5895 (N_5895,N_5443,N_5091);
or U5896 (N_5896,N_5218,N_5156);
nor U5897 (N_5897,N_5332,N_5104);
nand U5898 (N_5898,N_5175,N_5065);
nand U5899 (N_5899,N_5310,N_5414);
and U5900 (N_5900,N_5465,N_5393);
nand U5901 (N_5901,N_5406,N_5238);
or U5902 (N_5902,N_5394,N_5461);
nand U5903 (N_5903,N_5442,N_5119);
or U5904 (N_5904,N_5053,N_5259);
nor U5905 (N_5905,N_5431,N_5052);
nand U5906 (N_5906,N_5107,N_5196);
nand U5907 (N_5907,N_5144,N_5197);
and U5908 (N_5908,N_5203,N_5152);
and U5909 (N_5909,N_5174,N_5441);
nor U5910 (N_5910,N_5286,N_5042);
nor U5911 (N_5911,N_5352,N_5325);
or U5912 (N_5912,N_5358,N_5311);
nand U5913 (N_5913,N_5068,N_5227);
or U5914 (N_5914,N_5400,N_5084);
xor U5915 (N_5915,N_5318,N_5153);
nand U5916 (N_5916,N_5276,N_5464);
nor U5917 (N_5917,N_5409,N_5154);
nand U5918 (N_5918,N_5179,N_5152);
and U5919 (N_5919,N_5092,N_5051);
nor U5920 (N_5920,N_5017,N_5398);
and U5921 (N_5921,N_5167,N_5216);
or U5922 (N_5922,N_5341,N_5398);
nor U5923 (N_5923,N_5407,N_5336);
or U5924 (N_5924,N_5001,N_5060);
or U5925 (N_5925,N_5226,N_5461);
nor U5926 (N_5926,N_5032,N_5408);
and U5927 (N_5927,N_5327,N_5162);
and U5928 (N_5928,N_5125,N_5304);
nor U5929 (N_5929,N_5092,N_5343);
nor U5930 (N_5930,N_5342,N_5409);
or U5931 (N_5931,N_5396,N_5357);
nand U5932 (N_5932,N_5380,N_5272);
nor U5933 (N_5933,N_5487,N_5475);
and U5934 (N_5934,N_5364,N_5372);
and U5935 (N_5935,N_5341,N_5213);
nand U5936 (N_5936,N_5497,N_5431);
nand U5937 (N_5937,N_5483,N_5024);
nor U5938 (N_5938,N_5326,N_5003);
or U5939 (N_5939,N_5278,N_5309);
nand U5940 (N_5940,N_5072,N_5364);
nor U5941 (N_5941,N_5233,N_5495);
or U5942 (N_5942,N_5244,N_5370);
nor U5943 (N_5943,N_5002,N_5495);
nand U5944 (N_5944,N_5499,N_5467);
nand U5945 (N_5945,N_5015,N_5458);
and U5946 (N_5946,N_5446,N_5121);
or U5947 (N_5947,N_5498,N_5120);
and U5948 (N_5948,N_5305,N_5397);
xnor U5949 (N_5949,N_5286,N_5188);
nor U5950 (N_5950,N_5401,N_5225);
nand U5951 (N_5951,N_5277,N_5310);
or U5952 (N_5952,N_5282,N_5319);
or U5953 (N_5953,N_5028,N_5135);
nand U5954 (N_5954,N_5115,N_5156);
or U5955 (N_5955,N_5199,N_5009);
nor U5956 (N_5956,N_5383,N_5022);
nand U5957 (N_5957,N_5143,N_5363);
nand U5958 (N_5958,N_5279,N_5264);
nor U5959 (N_5959,N_5223,N_5435);
nor U5960 (N_5960,N_5431,N_5179);
and U5961 (N_5961,N_5488,N_5322);
or U5962 (N_5962,N_5331,N_5319);
nand U5963 (N_5963,N_5383,N_5330);
nand U5964 (N_5964,N_5145,N_5359);
nand U5965 (N_5965,N_5105,N_5434);
nor U5966 (N_5966,N_5259,N_5323);
nand U5967 (N_5967,N_5259,N_5478);
or U5968 (N_5968,N_5098,N_5052);
and U5969 (N_5969,N_5174,N_5044);
xnor U5970 (N_5970,N_5277,N_5487);
nor U5971 (N_5971,N_5026,N_5415);
nor U5972 (N_5972,N_5377,N_5285);
nor U5973 (N_5973,N_5401,N_5049);
nor U5974 (N_5974,N_5027,N_5336);
or U5975 (N_5975,N_5235,N_5149);
or U5976 (N_5976,N_5132,N_5443);
nand U5977 (N_5977,N_5338,N_5010);
nand U5978 (N_5978,N_5410,N_5205);
or U5979 (N_5979,N_5229,N_5042);
and U5980 (N_5980,N_5472,N_5163);
nand U5981 (N_5981,N_5321,N_5274);
nand U5982 (N_5982,N_5273,N_5077);
and U5983 (N_5983,N_5384,N_5304);
nor U5984 (N_5984,N_5364,N_5474);
nand U5985 (N_5985,N_5213,N_5495);
nor U5986 (N_5986,N_5173,N_5419);
nor U5987 (N_5987,N_5143,N_5059);
or U5988 (N_5988,N_5298,N_5329);
nand U5989 (N_5989,N_5028,N_5047);
nand U5990 (N_5990,N_5257,N_5469);
and U5991 (N_5991,N_5484,N_5307);
and U5992 (N_5992,N_5360,N_5063);
or U5993 (N_5993,N_5013,N_5293);
or U5994 (N_5994,N_5020,N_5177);
nand U5995 (N_5995,N_5415,N_5274);
nand U5996 (N_5996,N_5492,N_5464);
or U5997 (N_5997,N_5119,N_5121);
and U5998 (N_5998,N_5456,N_5419);
and U5999 (N_5999,N_5337,N_5043);
and U6000 (N_6000,N_5795,N_5656);
nor U6001 (N_6001,N_5705,N_5612);
or U6002 (N_6002,N_5765,N_5584);
nand U6003 (N_6003,N_5918,N_5972);
nand U6004 (N_6004,N_5936,N_5619);
nor U6005 (N_6005,N_5877,N_5812);
or U6006 (N_6006,N_5846,N_5794);
and U6007 (N_6007,N_5997,N_5807);
and U6008 (N_6008,N_5767,N_5579);
or U6009 (N_6009,N_5746,N_5681);
nor U6010 (N_6010,N_5992,N_5930);
nand U6011 (N_6011,N_5554,N_5676);
nand U6012 (N_6012,N_5551,N_5655);
and U6013 (N_6013,N_5915,N_5647);
and U6014 (N_6014,N_5650,N_5710);
nand U6015 (N_6015,N_5751,N_5924);
nand U6016 (N_6016,N_5802,N_5974);
or U6017 (N_6017,N_5788,N_5805);
nand U6018 (N_6018,N_5525,N_5881);
and U6019 (N_6019,N_5943,N_5882);
or U6020 (N_6020,N_5633,N_5904);
nor U6021 (N_6021,N_5591,N_5847);
nand U6022 (N_6022,N_5916,N_5913);
or U6023 (N_6023,N_5862,N_5500);
or U6024 (N_6024,N_5585,N_5900);
and U6025 (N_6025,N_5820,N_5885);
or U6026 (N_6026,N_5986,N_5575);
and U6027 (N_6027,N_5609,N_5892);
or U6028 (N_6028,N_5798,N_5828);
or U6029 (N_6029,N_5880,N_5898);
and U6030 (N_6030,N_5757,N_5561);
and U6031 (N_6031,N_5824,N_5671);
nor U6032 (N_6032,N_5637,N_5782);
and U6033 (N_6033,N_5535,N_5590);
or U6034 (N_6034,N_5929,N_5822);
nor U6035 (N_6035,N_5715,N_5772);
or U6036 (N_6036,N_5960,N_5917);
nor U6037 (N_6037,N_5578,N_5537);
and U6038 (N_6038,N_5555,N_5611);
nor U6039 (N_6039,N_5963,N_5534);
or U6040 (N_6040,N_5965,N_5839);
xor U6041 (N_6041,N_5810,N_5544);
or U6042 (N_6042,N_5704,N_5566);
or U6043 (N_6043,N_5513,N_5693);
nand U6044 (N_6044,N_5865,N_5691);
nor U6045 (N_6045,N_5879,N_5982);
nand U6046 (N_6046,N_5632,N_5686);
nor U6047 (N_6047,N_5902,N_5922);
or U6048 (N_6048,N_5750,N_5533);
nand U6049 (N_6049,N_5556,N_5803);
nor U6050 (N_6050,N_5653,N_5981);
nand U6051 (N_6051,N_5737,N_5593);
and U6052 (N_6052,N_5791,N_5515);
or U6053 (N_6053,N_5783,N_5840);
or U6054 (N_6054,N_5914,N_5861);
and U6055 (N_6055,N_5849,N_5665);
nand U6056 (N_6056,N_5595,N_5835);
nand U6057 (N_6057,N_5996,N_5573);
xor U6058 (N_6058,N_5945,N_5511);
nand U6059 (N_6059,N_5729,N_5934);
nor U6060 (N_6060,N_5638,N_5541);
and U6061 (N_6061,N_5850,N_5958);
nor U6062 (N_6062,N_5658,N_5649);
nor U6063 (N_6063,N_5939,N_5713);
or U6064 (N_6064,N_5733,N_5826);
nand U6065 (N_6065,N_5680,N_5539);
and U6066 (N_6066,N_5626,N_5778);
and U6067 (N_6067,N_5829,N_5779);
nand U6068 (N_6068,N_5896,N_5644);
nor U6069 (N_6069,N_5955,N_5505);
nor U6070 (N_6070,N_5718,N_5780);
and U6071 (N_6071,N_5999,N_5545);
and U6072 (N_6072,N_5871,N_5838);
nand U6073 (N_6073,N_5538,N_5908);
nor U6074 (N_6074,N_5530,N_5621);
or U6075 (N_6075,N_5640,N_5600);
nand U6076 (N_6076,N_5953,N_5635);
nor U6077 (N_6077,N_5690,N_5893);
and U6078 (N_6078,N_5589,N_5601);
nor U6079 (N_6079,N_5948,N_5689);
and U6080 (N_6080,N_5518,N_5954);
nand U6081 (N_6081,N_5502,N_5927);
or U6082 (N_6082,N_5773,N_5740);
xnor U6083 (N_6083,N_5598,N_5570);
nor U6084 (N_6084,N_5753,N_5856);
or U6085 (N_6085,N_5703,N_5832);
or U6086 (N_6086,N_5800,N_5764);
or U6087 (N_6087,N_5911,N_5969);
and U6088 (N_6088,N_5756,N_5508);
and U6089 (N_6089,N_5947,N_5866);
or U6090 (N_6090,N_5894,N_5966);
and U6091 (N_6091,N_5909,N_5771);
nor U6092 (N_6092,N_5546,N_5588);
or U6093 (N_6093,N_5868,N_5859);
or U6094 (N_6094,N_5967,N_5891);
and U6095 (N_6095,N_5864,N_5991);
or U6096 (N_6096,N_5989,N_5701);
or U6097 (N_6097,N_5957,N_5639);
nand U6098 (N_6098,N_5606,N_5651);
nor U6099 (N_6099,N_5770,N_5547);
and U6100 (N_6100,N_5670,N_5851);
nand U6101 (N_6101,N_5987,N_5792);
nor U6102 (N_6102,N_5521,N_5559);
nand U6103 (N_6103,N_5652,N_5597);
and U6104 (N_6104,N_5532,N_5769);
and U6105 (N_6105,N_5608,N_5744);
nand U6106 (N_6106,N_5677,N_5522);
or U6107 (N_6107,N_5825,N_5636);
and U6108 (N_6108,N_5925,N_5980);
or U6109 (N_6109,N_5979,N_5776);
or U6110 (N_6110,N_5735,N_5631);
xor U6111 (N_6111,N_5815,N_5952);
or U6112 (N_6112,N_5749,N_5899);
and U6113 (N_6113,N_5666,N_5845);
nor U6114 (N_6114,N_5994,N_5628);
nand U6115 (N_6115,N_5577,N_5971);
or U6116 (N_6116,N_5560,N_5562);
nand U6117 (N_6117,N_5620,N_5873);
and U6118 (N_6118,N_5875,N_5622);
and U6119 (N_6119,N_5901,N_5962);
or U6120 (N_6120,N_5724,N_5853);
nor U6121 (N_6121,N_5514,N_5748);
or U6122 (N_6122,N_5625,N_5602);
nand U6123 (N_6123,N_5563,N_5932);
or U6124 (N_6124,N_5811,N_5884);
and U6125 (N_6125,N_5732,N_5926);
or U6126 (N_6126,N_5543,N_5920);
nand U6127 (N_6127,N_5833,N_5692);
nand U6128 (N_6128,N_5777,N_5694);
and U6129 (N_6129,N_5906,N_5503);
nor U6130 (N_6130,N_5801,N_5886);
nor U6131 (N_6131,N_5728,N_5940);
and U6132 (N_6132,N_5709,N_5526);
nand U6133 (N_6133,N_5870,N_5695);
and U6134 (N_6134,N_5552,N_5574);
nor U6135 (N_6135,N_5928,N_5984);
nand U6136 (N_6136,N_5998,N_5507);
nand U6137 (N_6137,N_5531,N_5572);
and U6138 (N_6138,N_5854,N_5604);
nand U6139 (N_6139,N_5978,N_5642);
nor U6140 (N_6140,N_5617,N_5697);
and U6141 (N_6141,N_5938,N_5645);
nand U6142 (N_6142,N_5506,N_5641);
and U6143 (N_6143,N_5726,N_5941);
and U6144 (N_6144,N_5942,N_5752);
and U6145 (N_6145,N_5781,N_5834);
and U6146 (N_6146,N_5582,N_5565);
nor U6147 (N_6147,N_5897,N_5657);
and U6148 (N_6148,N_5919,N_5592);
xnor U6149 (N_6149,N_5564,N_5687);
and U6150 (N_6150,N_5512,N_5624);
xnor U6151 (N_6151,N_5736,N_5599);
or U6152 (N_6152,N_5809,N_5576);
nor U6153 (N_6153,N_5813,N_5707);
nor U6154 (N_6154,N_5977,N_5661);
xnor U6155 (N_6155,N_5842,N_5869);
and U6156 (N_6156,N_5643,N_5634);
nand U6157 (N_6157,N_5571,N_5614);
and U6158 (N_6158,N_5890,N_5678);
nand U6159 (N_6159,N_5723,N_5983);
nand U6160 (N_6160,N_5883,N_5933);
or U6161 (N_6161,N_5876,N_5731);
nand U6162 (N_6162,N_5509,N_5747);
nand U6163 (N_6163,N_5527,N_5821);
and U6164 (N_6164,N_5654,N_5907);
nand U6165 (N_6165,N_5895,N_5730);
nand U6166 (N_6166,N_5517,N_5667);
and U6167 (N_6167,N_5787,N_5717);
nor U6168 (N_6168,N_5540,N_5855);
or U6169 (N_6169,N_5827,N_5831);
and U6170 (N_6170,N_5581,N_5720);
nor U6171 (N_6171,N_5596,N_5674);
nand U6172 (N_6172,N_5951,N_5519);
nand U6173 (N_6173,N_5536,N_5973);
and U6174 (N_6174,N_5557,N_5580);
nor U6175 (N_6175,N_5975,N_5745);
nand U6176 (N_6176,N_5630,N_5623);
and U6177 (N_6177,N_5520,N_5528);
nand U6178 (N_6178,N_5775,N_5889);
and U6179 (N_6179,N_5714,N_5949);
or U6180 (N_6180,N_5524,N_5660);
nand U6181 (N_6181,N_5672,N_5629);
or U6182 (N_6182,N_5607,N_5841);
or U6183 (N_6183,N_5793,N_5766);
or U6184 (N_6184,N_5727,N_5857);
or U6185 (N_6185,N_5796,N_5558);
and U6186 (N_6186,N_5808,N_5569);
nand U6187 (N_6187,N_5743,N_5610);
and U6188 (N_6188,N_5529,N_5830);
nor U6189 (N_6189,N_5843,N_5874);
and U6190 (N_6190,N_5931,N_5734);
nand U6191 (N_6191,N_5935,N_5615);
and U6192 (N_6192,N_5944,N_5848);
and U6193 (N_6193,N_5719,N_5836);
or U6194 (N_6194,N_5618,N_5587);
nor U6195 (N_6195,N_5860,N_5993);
nor U6196 (N_6196,N_5613,N_5648);
nand U6197 (N_6197,N_5804,N_5668);
nor U6198 (N_6198,N_5970,N_5685);
and U6199 (N_6199,N_5568,N_5878);
or U6200 (N_6200,N_5905,N_5698);
nor U6201 (N_6201,N_5669,N_5675);
nor U6202 (N_6202,N_5664,N_5959);
nand U6203 (N_6203,N_5863,N_5852);
or U6204 (N_6204,N_5768,N_5706);
or U6205 (N_6205,N_5721,N_5659);
or U6206 (N_6206,N_5837,N_5683);
and U6207 (N_6207,N_5627,N_5504);
and U6208 (N_6208,N_5819,N_5708);
and U6209 (N_6209,N_5550,N_5988);
nand U6210 (N_6210,N_5567,N_5759);
nand U6211 (N_6211,N_5964,N_5616);
xor U6212 (N_6212,N_5646,N_5682);
and U6213 (N_6213,N_5956,N_5976);
or U6214 (N_6214,N_5739,N_5789);
nand U6215 (N_6215,N_5797,N_5679);
and U6216 (N_6216,N_5761,N_5968);
or U6217 (N_6217,N_5758,N_5760);
nand U6218 (N_6218,N_5662,N_5818);
or U6219 (N_6219,N_5742,N_5741);
and U6220 (N_6220,N_5696,N_5823);
or U6221 (N_6221,N_5688,N_5946);
nand U6222 (N_6222,N_5814,N_5784);
and U6223 (N_6223,N_5785,N_5790);
nor U6224 (N_6224,N_5887,N_5910);
or U6225 (N_6225,N_5702,N_5763);
nand U6226 (N_6226,N_5921,N_5716);
nor U6227 (N_6227,N_5995,N_5725);
nor U6228 (N_6228,N_5950,N_5548);
or U6229 (N_6229,N_5786,N_5516);
and U6230 (N_6230,N_5923,N_5699);
nand U6231 (N_6231,N_5523,N_5553);
nand U6232 (N_6232,N_5937,N_5586);
or U6233 (N_6233,N_5990,N_5700);
nor U6234 (N_6234,N_5799,N_5712);
and U6235 (N_6235,N_5806,N_5912);
nor U6236 (N_6236,N_5603,N_5985);
nor U6237 (N_6237,N_5858,N_5762);
nor U6238 (N_6238,N_5754,N_5844);
xor U6239 (N_6239,N_5711,N_5684);
and U6240 (N_6240,N_5501,N_5755);
or U6241 (N_6241,N_5594,N_5722);
nor U6242 (N_6242,N_5888,N_5903);
or U6243 (N_6243,N_5663,N_5583);
or U6244 (N_6244,N_5961,N_5738);
nor U6245 (N_6245,N_5510,N_5872);
and U6246 (N_6246,N_5867,N_5673);
nor U6247 (N_6247,N_5549,N_5816);
and U6248 (N_6248,N_5817,N_5605);
nand U6249 (N_6249,N_5542,N_5774);
nor U6250 (N_6250,N_5859,N_5647);
and U6251 (N_6251,N_5973,N_5956);
nor U6252 (N_6252,N_5639,N_5882);
nand U6253 (N_6253,N_5547,N_5550);
nor U6254 (N_6254,N_5893,N_5819);
xnor U6255 (N_6255,N_5907,N_5990);
nor U6256 (N_6256,N_5700,N_5764);
nand U6257 (N_6257,N_5552,N_5793);
and U6258 (N_6258,N_5816,N_5903);
nand U6259 (N_6259,N_5856,N_5857);
nand U6260 (N_6260,N_5986,N_5609);
nand U6261 (N_6261,N_5766,N_5942);
nand U6262 (N_6262,N_5767,N_5688);
nor U6263 (N_6263,N_5666,N_5789);
nand U6264 (N_6264,N_5988,N_5917);
nor U6265 (N_6265,N_5706,N_5669);
or U6266 (N_6266,N_5952,N_5505);
and U6267 (N_6267,N_5964,N_5732);
or U6268 (N_6268,N_5942,N_5673);
and U6269 (N_6269,N_5759,N_5842);
nand U6270 (N_6270,N_5623,N_5558);
nand U6271 (N_6271,N_5927,N_5564);
nor U6272 (N_6272,N_5961,N_5745);
or U6273 (N_6273,N_5628,N_5668);
and U6274 (N_6274,N_5719,N_5980);
nand U6275 (N_6275,N_5641,N_5696);
or U6276 (N_6276,N_5788,N_5629);
or U6277 (N_6277,N_5639,N_5702);
nand U6278 (N_6278,N_5562,N_5928);
or U6279 (N_6279,N_5562,N_5738);
nand U6280 (N_6280,N_5626,N_5994);
or U6281 (N_6281,N_5551,N_5823);
nand U6282 (N_6282,N_5895,N_5894);
and U6283 (N_6283,N_5700,N_5656);
and U6284 (N_6284,N_5998,N_5586);
or U6285 (N_6285,N_5715,N_5988);
nor U6286 (N_6286,N_5696,N_5754);
nand U6287 (N_6287,N_5851,N_5890);
or U6288 (N_6288,N_5518,N_5872);
and U6289 (N_6289,N_5522,N_5839);
nand U6290 (N_6290,N_5737,N_5639);
and U6291 (N_6291,N_5850,N_5771);
xnor U6292 (N_6292,N_5749,N_5568);
nand U6293 (N_6293,N_5636,N_5742);
or U6294 (N_6294,N_5661,N_5966);
and U6295 (N_6295,N_5584,N_5787);
nand U6296 (N_6296,N_5515,N_5806);
nand U6297 (N_6297,N_5873,N_5885);
or U6298 (N_6298,N_5792,N_5861);
nor U6299 (N_6299,N_5520,N_5747);
or U6300 (N_6300,N_5678,N_5807);
or U6301 (N_6301,N_5614,N_5669);
nor U6302 (N_6302,N_5925,N_5805);
or U6303 (N_6303,N_5793,N_5901);
nand U6304 (N_6304,N_5887,N_5684);
nor U6305 (N_6305,N_5532,N_5707);
and U6306 (N_6306,N_5665,N_5743);
or U6307 (N_6307,N_5856,N_5812);
or U6308 (N_6308,N_5842,N_5672);
and U6309 (N_6309,N_5655,N_5717);
and U6310 (N_6310,N_5756,N_5724);
nor U6311 (N_6311,N_5799,N_5745);
xor U6312 (N_6312,N_5620,N_5948);
nand U6313 (N_6313,N_5982,N_5539);
nand U6314 (N_6314,N_5655,N_5721);
nand U6315 (N_6315,N_5551,N_5915);
nand U6316 (N_6316,N_5659,N_5794);
and U6317 (N_6317,N_5632,N_5909);
nor U6318 (N_6318,N_5777,N_5820);
nand U6319 (N_6319,N_5572,N_5613);
nand U6320 (N_6320,N_5750,N_5986);
or U6321 (N_6321,N_5569,N_5904);
or U6322 (N_6322,N_5518,N_5810);
or U6323 (N_6323,N_5772,N_5644);
and U6324 (N_6324,N_5773,N_5657);
nand U6325 (N_6325,N_5582,N_5510);
nor U6326 (N_6326,N_5692,N_5890);
nand U6327 (N_6327,N_5865,N_5552);
and U6328 (N_6328,N_5971,N_5749);
and U6329 (N_6329,N_5681,N_5515);
or U6330 (N_6330,N_5506,N_5744);
and U6331 (N_6331,N_5914,N_5612);
nor U6332 (N_6332,N_5990,N_5848);
nand U6333 (N_6333,N_5877,N_5933);
nand U6334 (N_6334,N_5600,N_5845);
nand U6335 (N_6335,N_5831,N_5894);
and U6336 (N_6336,N_5876,N_5600);
nor U6337 (N_6337,N_5672,N_5866);
nor U6338 (N_6338,N_5833,N_5835);
or U6339 (N_6339,N_5914,N_5539);
or U6340 (N_6340,N_5868,N_5820);
nand U6341 (N_6341,N_5663,N_5773);
nand U6342 (N_6342,N_5707,N_5663);
nand U6343 (N_6343,N_5926,N_5631);
nand U6344 (N_6344,N_5541,N_5917);
and U6345 (N_6345,N_5611,N_5614);
or U6346 (N_6346,N_5920,N_5600);
nand U6347 (N_6347,N_5933,N_5834);
and U6348 (N_6348,N_5925,N_5971);
and U6349 (N_6349,N_5871,N_5807);
nand U6350 (N_6350,N_5507,N_5595);
nand U6351 (N_6351,N_5587,N_5743);
and U6352 (N_6352,N_5541,N_5655);
and U6353 (N_6353,N_5722,N_5696);
nor U6354 (N_6354,N_5591,N_5711);
or U6355 (N_6355,N_5508,N_5884);
nand U6356 (N_6356,N_5929,N_5933);
or U6357 (N_6357,N_5891,N_5618);
nand U6358 (N_6358,N_5823,N_5745);
nand U6359 (N_6359,N_5943,N_5551);
or U6360 (N_6360,N_5617,N_5891);
nand U6361 (N_6361,N_5839,N_5845);
and U6362 (N_6362,N_5569,N_5800);
and U6363 (N_6363,N_5543,N_5914);
or U6364 (N_6364,N_5990,N_5806);
nand U6365 (N_6365,N_5586,N_5955);
nand U6366 (N_6366,N_5555,N_5561);
and U6367 (N_6367,N_5872,N_5878);
and U6368 (N_6368,N_5844,N_5947);
nor U6369 (N_6369,N_5955,N_5841);
or U6370 (N_6370,N_5866,N_5506);
nand U6371 (N_6371,N_5811,N_5958);
nor U6372 (N_6372,N_5876,N_5942);
nor U6373 (N_6373,N_5945,N_5793);
or U6374 (N_6374,N_5671,N_5776);
and U6375 (N_6375,N_5982,N_5810);
and U6376 (N_6376,N_5588,N_5761);
or U6377 (N_6377,N_5630,N_5943);
and U6378 (N_6378,N_5861,N_5595);
and U6379 (N_6379,N_5837,N_5861);
or U6380 (N_6380,N_5568,N_5655);
and U6381 (N_6381,N_5768,N_5638);
and U6382 (N_6382,N_5834,N_5582);
or U6383 (N_6383,N_5855,N_5952);
nand U6384 (N_6384,N_5992,N_5548);
and U6385 (N_6385,N_5658,N_5983);
nand U6386 (N_6386,N_5726,N_5546);
or U6387 (N_6387,N_5777,N_5592);
and U6388 (N_6388,N_5745,N_5808);
or U6389 (N_6389,N_5721,N_5855);
and U6390 (N_6390,N_5571,N_5766);
or U6391 (N_6391,N_5786,N_5539);
and U6392 (N_6392,N_5635,N_5535);
or U6393 (N_6393,N_5988,N_5860);
xor U6394 (N_6394,N_5663,N_5944);
nand U6395 (N_6395,N_5835,N_5757);
or U6396 (N_6396,N_5976,N_5768);
nand U6397 (N_6397,N_5763,N_5977);
and U6398 (N_6398,N_5854,N_5670);
nor U6399 (N_6399,N_5649,N_5936);
nor U6400 (N_6400,N_5996,N_5770);
nand U6401 (N_6401,N_5679,N_5873);
and U6402 (N_6402,N_5958,N_5505);
nand U6403 (N_6403,N_5644,N_5630);
nor U6404 (N_6404,N_5711,N_5996);
and U6405 (N_6405,N_5919,N_5536);
nand U6406 (N_6406,N_5565,N_5508);
nor U6407 (N_6407,N_5814,N_5583);
nand U6408 (N_6408,N_5841,N_5970);
nor U6409 (N_6409,N_5613,N_5560);
nor U6410 (N_6410,N_5965,N_5969);
and U6411 (N_6411,N_5552,N_5594);
nand U6412 (N_6412,N_5988,N_5511);
nor U6413 (N_6413,N_5832,N_5554);
nor U6414 (N_6414,N_5740,N_5849);
or U6415 (N_6415,N_5768,N_5913);
and U6416 (N_6416,N_5996,N_5951);
nand U6417 (N_6417,N_5587,N_5871);
xnor U6418 (N_6418,N_5616,N_5640);
or U6419 (N_6419,N_5751,N_5637);
or U6420 (N_6420,N_5675,N_5752);
and U6421 (N_6421,N_5603,N_5553);
nand U6422 (N_6422,N_5964,N_5885);
nor U6423 (N_6423,N_5964,N_5809);
nand U6424 (N_6424,N_5583,N_5623);
or U6425 (N_6425,N_5970,N_5631);
nor U6426 (N_6426,N_5985,N_5504);
nand U6427 (N_6427,N_5592,N_5798);
or U6428 (N_6428,N_5846,N_5919);
nand U6429 (N_6429,N_5550,N_5611);
nor U6430 (N_6430,N_5553,N_5635);
nand U6431 (N_6431,N_5970,N_5966);
nand U6432 (N_6432,N_5920,N_5535);
and U6433 (N_6433,N_5537,N_5671);
nand U6434 (N_6434,N_5608,N_5951);
and U6435 (N_6435,N_5871,N_5667);
nand U6436 (N_6436,N_5925,N_5872);
nor U6437 (N_6437,N_5806,N_5519);
nor U6438 (N_6438,N_5839,N_5826);
nor U6439 (N_6439,N_5694,N_5868);
or U6440 (N_6440,N_5633,N_5833);
and U6441 (N_6441,N_5919,N_5970);
nor U6442 (N_6442,N_5612,N_5678);
nand U6443 (N_6443,N_5514,N_5795);
or U6444 (N_6444,N_5648,N_5600);
nor U6445 (N_6445,N_5904,N_5799);
or U6446 (N_6446,N_5941,N_5754);
nand U6447 (N_6447,N_5766,N_5928);
or U6448 (N_6448,N_5762,N_5655);
nand U6449 (N_6449,N_5760,N_5651);
or U6450 (N_6450,N_5695,N_5518);
nand U6451 (N_6451,N_5836,N_5767);
or U6452 (N_6452,N_5564,N_5811);
or U6453 (N_6453,N_5992,N_5707);
nor U6454 (N_6454,N_5546,N_5811);
and U6455 (N_6455,N_5688,N_5712);
and U6456 (N_6456,N_5940,N_5921);
nor U6457 (N_6457,N_5686,N_5688);
and U6458 (N_6458,N_5533,N_5696);
and U6459 (N_6459,N_5716,N_5917);
or U6460 (N_6460,N_5751,N_5859);
nand U6461 (N_6461,N_5696,N_5747);
nand U6462 (N_6462,N_5737,N_5861);
nor U6463 (N_6463,N_5931,N_5815);
or U6464 (N_6464,N_5869,N_5891);
or U6465 (N_6465,N_5803,N_5921);
and U6466 (N_6466,N_5582,N_5964);
nor U6467 (N_6467,N_5743,N_5908);
and U6468 (N_6468,N_5736,N_5622);
and U6469 (N_6469,N_5726,N_5744);
or U6470 (N_6470,N_5653,N_5962);
or U6471 (N_6471,N_5903,N_5665);
or U6472 (N_6472,N_5694,N_5523);
and U6473 (N_6473,N_5920,N_5944);
and U6474 (N_6474,N_5736,N_5760);
and U6475 (N_6475,N_5589,N_5557);
nand U6476 (N_6476,N_5960,N_5580);
or U6477 (N_6477,N_5653,N_5783);
xnor U6478 (N_6478,N_5506,N_5720);
nor U6479 (N_6479,N_5703,N_5649);
and U6480 (N_6480,N_5672,N_5549);
or U6481 (N_6481,N_5889,N_5559);
or U6482 (N_6482,N_5756,N_5894);
and U6483 (N_6483,N_5651,N_5924);
nand U6484 (N_6484,N_5933,N_5870);
and U6485 (N_6485,N_5725,N_5935);
xor U6486 (N_6486,N_5992,N_5817);
nor U6487 (N_6487,N_5774,N_5918);
and U6488 (N_6488,N_5821,N_5738);
nor U6489 (N_6489,N_5550,N_5653);
and U6490 (N_6490,N_5923,N_5873);
nor U6491 (N_6491,N_5826,N_5816);
nor U6492 (N_6492,N_5906,N_5644);
or U6493 (N_6493,N_5869,N_5555);
or U6494 (N_6494,N_5571,N_5928);
and U6495 (N_6495,N_5835,N_5596);
or U6496 (N_6496,N_5791,N_5769);
nand U6497 (N_6497,N_5771,N_5887);
or U6498 (N_6498,N_5526,N_5979);
nand U6499 (N_6499,N_5630,N_5746);
xor U6500 (N_6500,N_6083,N_6413);
nor U6501 (N_6501,N_6493,N_6310);
nor U6502 (N_6502,N_6367,N_6060);
nor U6503 (N_6503,N_6406,N_6027);
nor U6504 (N_6504,N_6264,N_6096);
and U6505 (N_6505,N_6260,N_6022);
and U6506 (N_6506,N_6097,N_6474);
nor U6507 (N_6507,N_6462,N_6444);
or U6508 (N_6508,N_6357,N_6349);
nor U6509 (N_6509,N_6385,N_6318);
nand U6510 (N_6510,N_6194,N_6322);
nor U6511 (N_6511,N_6377,N_6336);
nor U6512 (N_6512,N_6240,N_6425);
nand U6513 (N_6513,N_6200,N_6272);
nand U6514 (N_6514,N_6472,N_6375);
nor U6515 (N_6515,N_6205,N_6086);
nand U6516 (N_6516,N_6064,N_6118);
or U6517 (N_6517,N_6355,N_6207);
nand U6518 (N_6518,N_6422,N_6286);
or U6519 (N_6519,N_6008,N_6091);
and U6520 (N_6520,N_6259,N_6285);
and U6521 (N_6521,N_6266,N_6085);
nand U6522 (N_6522,N_6049,N_6360);
nor U6523 (N_6523,N_6499,N_6089);
nor U6524 (N_6524,N_6056,N_6024);
xor U6525 (N_6525,N_6078,N_6195);
nand U6526 (N_6526,N_6456,N_6072);
nor U6527 (N_6527,N_6485,N_6244);
nor U6528 (N_6528,N_6410,N_6235);
or U6529 (N_6529,N_6013,N_6404);
nor U6530 (N_6530,N_6368,N_6210);
nor U6531 (N_6531,N_6304,N_6009);
and U6532 (N_6532,N_6137,N_6476);
nand U6533 (N_6533,N_6341,N_6003);
nor U6534 (N_6534,N_6370,N_6247);
nor U6535 (N_6535,N_6397,N_6016);
and U6536 (N_6536,N_6364,N_6356);
nand U6537 (N_6537,N_6265,N_6035);
and U6538 (N_6538,N_6081,N_6284);
and U6539 (N_6539,N_6411,N_6111);
or U6540 (N_6540,N_6074,N_6290);
nand U6541 (N_6541,N_6116,N_6495);
or U6542 (N_6542,N_6449,N_6090);
or U6543 (N_6543,N_6252,N_6028);
and U6544 (N_6544,N_6112,N_6012);
or U6545 (N_6545,N_6131,N_6047);
or U6546 (N_6546,N_6312,N_6154);
or U6547 (N_6547,N_6156,N_6458);
and U6548 (N_6548,N_6026,N_6299);
nand U6549 (N_6549,N_6044,N_6316);
nand U6550 (N_6550,N_6359,N_6424);
nor U6551 (N_6551,N_6269,N_6196);
or U6552 (N_6552,N_6189,N_6101);
or U6553 (N_6553,N_6007,N_6239);
or U6554 (N_6554,N_6295,N_6158);
nand U6555 (N_6555,N_6435,N_6021);
nand U6556 (N_6556,N_6457,N_6015);
nor U6557 (N_6557,N_6416,N_6080);
nor U6558 (N_6558,N_6045,N_6324);
nand U6559 (N_6559,N_6020,N_6484);
nor U6560 (N_6560,N_6236,N_6464);
and U6561 (N_6561,N_6376,N_6139);
nor U6562 (N_6562,N_6143,N_6395);
nor U6563 (N_6563,N_6400,N_6128);
nor U6564 (N_6564,N_6306,N_6215);
or U6565 (N_6565,N_6394,N_6005);
nand U6566 (N_6566,N_6063,N_6423);
nor U6567 (N_6567,N_6327,N_6165);
or U6568 (N_6568,N_6268,N_6415);
nor U6569 (N_6569,N_6030,N_6103);
xor U6570 (N_6570,N_6100,N_6427);
or U6571 (N_6571,N_6408,N_6159);
nand U6572 (N_6572,N_6463,N_6490);
and U6573 (N_6573,N_6167,N_6480);
nor U6574 (N_6574,N_6294,N_6088);
or U6575 (N_6575,N_6492,N_6419);
and U6576 (N_6576,N_6323,N_6203);
and U6577 (N_6577,N_6213,N_6498);
nor U6578 (N_6578,N_6114,N_6270);
or U6579 (N_6579,N_6230,N_6308);
nand U6580 (N_6580,N_6439,N_6076);
nand U6581 (N_6581,N_6126,N_6038);
and U6582 (N_6582,N_6187,N_6202);
nor U6583 (N_6583,N_6055,N_6447);
nor U6584 (N_6584,N_6105,N_6084);
nand U6585 (N_6585,N_6381,N_6362);
or U6586 (N_6586,N_6333,N_6298);
and U6587 (N_6587,N_6421,N_6099);
and U6588 (N_6588,N_6221,N_6451);
nand U6589 (N_6589,N_6352,N_6384);
nand U6590 (N_6590,N_6460,N_6188);
and U6591 (N_6591,N_6066,N_6329);
nand U6592 (N_6592,N_6296,N_6023);
nand U6593 (N_6593,N_6162,N_6151);
nand U6594 (N_6594,N_6051,N_6275);
and U6595 (N_6595,N_6130,N_6067);
and U6596 (N_6596,N_6147,N_6233);
and U6597 (N_6597,N_6366,N_6095);
nand U6598 (N_6598,N_6283,N_6305);
nand U6599 (N_6599,N_6133,N_6040);
and U6600 (N_6600,N_6109,N_6288);
or U6601 (N_6601,N_6497,N_6053);
and U6602 (N_6602,N_6245,N_6071);
or U6603 (N_6603,N_6330,N_6321);
and U6604 (N_6604,N_6319,N_6328);
nand U6605 (N_6605,N_6034,N_6436);
and U6606 (N_6606,N_6190,N_6405);
or U6607 (N_6607,N_6466,N_6250);
or U6608 (N_6608,N_6036,N_6301);
or U6609 (N_6609,N_6032,N_6052);
or U6610 (N_6610,N_6050,N_6471);
nand U6611 (N_6611,N_6127,N_6093);
or U6612 (N_6612,N_6382,N_6371);
xor U6613 (N_6613,N_6217,N_6365);
nand U6614 (N_6614,N_6082,N_6280);
or U6615 (N_6615,N_6448,N_6238);
nor U6616 (N_6616,N_6231,N_6123);
and U6617 (N_6617,N_6345,N_6418);
nor U6618 (N_6618,N_6465,N_6059);
or U6619 (N_6619,N_6380,N_6004);
nor U6620 (N_6620,N_6006,N_6428);
nor U6621 (N_6621,N_6120,N_6054);
nor U6622 (N_6622,N_6379,N_6242);
nand U6623 (N_6623,N_6019,N_6197);
nor U6624 (N_6624,N_6479,N_6234);
nand U6625 (N_6625,N_6430,N_6145);
or U6626 (N_6626,N_6115,N_6223);
nor U6627 (N_6627,N_6338,N_6262);
and U6628 (N_6628,N_6303,N_6104);
xor U6629 (N_6629,N_6191,N_6271);
or U6630 (N_6630,N_6174,N_6075);
nand U6631 (N_6631,N_6206,N_6258);
nor U6632 (N_6632,N_6369,N_6496);
or U6633 (N_6633,N_6398,N_6176);
and U6634 (N_6634,N_6315,N_6273);
nor U6635 (N_6635,N_6237,N_6353);
nor U6636 (N_6636,N_6113,N_6487);
nand U6637 (N_6637,N_6168,N_6442);
xor U6638 (N_6638,N_6478,N_6136);
or U6639 (N_6639,N_6486,N_6274);
and U6640 (N_6640,N_6256,N_6431);
xor U6641 (N_6641,N_6440,N_6092);
and U6642 (N_6642,N_6140,N_6261);
xor U6643 (N_6643,N_6445,N_6106);
nor U6644 (N_6644,N_6443,N_6039);
or U6645 (N_6645,N_6177,N_6372);
nand U6646 (N_6646,N_6175,N_6263);
nor U6647 (N_6647,N_6342,N_6317);
nor U6648 (N_6648,N_6402,N_6166);
and U6649 (N_6649,N_6332,N_6161);
nor U6650 (N_6650,N_6392,N_6433);
nand U6651 (N_6651,N_6470,N_6426);
and U6652 (N_6652,N_6212,N_6383);
nor U6653 (N_6653,N_6201,N_6184);
or U6654 (N_6654,N_6488,N_6029);
nand U6655 (N_6655,N_6361,N_6253);
nor U6656 (N_6656,N_6193,N_6011);
nand U6657 (N_6657,N_6218,N_6347);
or U6658 (N_6658,N_6125,N_6157);
nor U6659 (N_6659,N_6152,N_6287);
nor U6660 (N_6660,N_6208,N_6388);
or U6661 (N_6661,N_6469,N_6142);
nor U6662 (N_6662,N_6414,N_6452);
and U6663 (N_6663,N_6307,N_6468);
and U6664 (N_6664,N_6409,N_6246);
and U6665 (N_6665,N_6216,N_6222);
and U6666 (N_6666,N_6354,N_6390);
and U6667 (N_6667,N_6094,N_6396);
and U6668 (N_6668,N_6249,N_6041);
or U6669 (N_6669,N_6257,N_6220);
or U6670 (N_6670,N_6098,N_6185);
nor U6671 (N_6671,N_6477,N_6062);
nor U6672 (N_6672,N_6279,N_6079);
or U6673 (N_6673,N_6037,N_6155);
or U6674 (N_6674,N_6199,N_6344);
or U6675 (N_6675,N_6311,N_6134);
and U6676 (N_6676,N_6399,N_6135);
nor U6677 (N_6677,N_6241,N_6070);
nor U6678 (N_6678,N_6122,N_6232);
nand U6679 (N_6679,N_6254,N_6068);
or U6680 (N_6680,N_6282,N_6225);
nor U6681 (N_6681,N_6348,N_6378);
and U6682 (N_6682,N_6292,N_6180);
nor U6683 (N_6683,N_6373,N_6407);
or U6684 (N_6684,N_6073,N_6450);
nor U6685 (N_6685,N_6467,N_6334);
or U6686 (N_6686,N_6343,N_6033);
or U6687 (N_6687,N_6281,N_6461);
nand U6688 (N_6688,N_6335,N_6224);
nor U6689 (N_6689,N_6192,N_6417);
and U6690 (N_6690,N_6297,N_6031);
nand U6691 (N_6691,N_6255,N_6391);
or U6692 (N_6692,N_6001,N_6179);
nand U6693 (N_6693,N_6267,N_6017);
nor U6694 (N_6694,N_6339,N_6313);
and U6695 (N_6695,N_6058,N_6403);
nor U6696 (N_6696,N_6204,N_6132);
or U6697 (N_6697,N_6401,N_6107);
or U6698 (N_6698,N_6077,N_6289);
nor U6699 (N_6699,N_6446,N_6214);
or U6700 (N_6700,N_6164,N_6172);
nand U6701 (N_6701,N_6434,N_6482);
nor U6702 (N_6702,N_6481,N_6069);
and U6703 (N_6703,N_6248,N_6432);
and U6704 (N_6704,N_6186,N_6173);
and U6705 (N_6705,N_6129,N_6002);
or U6706 (N_6706,N_6043,N_6102);
and U6707 (N_6707,N_6211,N_6320);
nand U6708 (N_6708,N_6489,N_6491);
nor U6709 (N_6709,N_6119,N_6420);
and U6710 (N_6710,N_6293,N_6243);
or U6711 (N_6711,N_6087,N_6014);
or U6712 (N_6712,N_6146,N_6229);
nor U6713 (N_6713,N_6277,N_6374);
and U6714 (N_6714,N_6170,N_6325);
nor U6715 (N_6715,N_6441,N_6025);
nand U6716 (N_6716,N_6065,N_6459);
nor U6717 (N_6717,N_6429,N_6473);
nand U6718 (N_6718,N_6163,N_6010);
or U6719 (N_6719,N_6150,N_6278);
or U6720 (N_6720,N_6178,N_6314);
nor U6721 (N_6721,N_6181,N_6302);
nor U6722 (N_6722,N_6363,N_6160);
or U6723 (N_6723,N_6454,N_6331);
and U6724 (N_6724,N_6386,N_6227);
nor U6725 (N_6725,N_6455,N_6124);
nand U6726 (N_6726,N_6437,N_6183);
or U6727 (N_6727,N_6300,N_6121);
or U6728 (N_6728,N_6198,N_6018);
or U6729 (N_6729,N_6048,N_6309);
and U6730 (N_6730,N_6219,N_6389);
nand U6731 (N_6731,N_6494,N_6117);
nand U6732 (N_6732,N_6046,N_6483);
nor U6733 (N_6733,N_6182,N_6340);
or U6734 (N_6734,N_6350,N_6337);
and U6735 (N_6735,N_6291,N_6138);
nand U6736 (N_6736,N_6141,N_6276);
or U6737 (N_6737,N_6346,N_6453);
and U6738 (N_6738,N_6209,N_6438);
and U6739 (N_6739,N_6169,N_6042);
nand U6740 (N_6740,N_6000,N_6351);
nand U6741 (N_6741,N_6110,N_6387);
nand U6742 (N_6742,N_6148,N_6475);
or U6743 (N_6743,N_6057,N_6144);
nor U6744 (N_6744,N_6171,N_6061);
and U6745 (N_6745,N_6153,N_6412);
nand U6746 (N_6746,N_6228,N_6149);
and U6747 (N_6747,N_6108,N_6251);
nand U6748 (N_6748,N_6393,N_6326);
or U6749 (N_6749,N_6358,N_6226);
or U6750 (N_6750,N_6452,N_6172);
nand U6751 (N_6751,N_6038,N_6432);
nor U6752 (N_6752,N_6412,N_6401);
or U6753 (N_6753,N_6323,N_6111);
nand U6754 (N_6754,N_6471,N_6118);
or U6755 (N_6755,N_6086,N_6342);
or U6756 (N_6756,N_6381,N_6103);
nor U6757 (N_6757,N_6130,N_6313);
or U6758 (N_6758,N_6332,N_6348);
nor U6759 (N_6759,N_6422,N_6024);
nand U6760 (N_6760,N_6209,N_6325);
nand U6761 (N_6761,N_6462,N_6206);
and U6762 (N_6762,N_6358,N_6430);
nand U6763 (N_6763,N_6304,N_6012);
or U6764 (N_6764,N_6485,N_6424);
or U6765 (N_6765,N_6049,N_6490);
and U6766 (N_6766,N_6241,N_6430);
xor U6767 (N_6767,N_6007,N_6399);
and U6768 (N_6768,N_6392,N_6489);
nand U6769 (N_6769,N_6124,N_6208);
nor U6770 (N_6770,N_6400,N_6063);
and U6771 (N_6771,N_6148,N_6018);
xor U6772 (N_6772,N_6472,N_6443);
nor U6773 (N_6773,N_6114,N_6410);
and U6774 (N_6774,N_6254,N_6397);
nor U6775 (N_6775,N_6481,N_6289);
xor U6776 (N_6776,N_6383,N_6043);
nand U6777 (N_6777,N_6071,N_6188);
and U6778 (N_6778,N_6307,N_6201);
and U6779 (N_6779,N_6193,N_6212);
and U6780 (N_6780,N_6347,N_6288);
or U6781 (N_6781,N_6171,N_6275);
and U6782 (N_6782,N_6000,N_6230);
or U6783 (N_6783,N_6276,N_6131);
or U6784 (N_6784,N_6337,N_6358);
or U6785 (N_6785,N_6007,N_6085);
nand U6786 (N_6786,N_6213,N_6106);
nor U6787 (N_6787,N_6041,N_6254);
nand U6788 (N_6788,N_6181,N_6413);
and U6789 (N_6789,N_6480,N_6290);
nor U6790 (N_6790,N_6098,N_6245);
or U6791 (N_6791,N_6303,N_6421);
or U6792 (N_6792,N_6496,N_6153);
and U6793 (N_6793,N_6314,N_6321);
nand U6794 (N_6794,N_6202,N_6214);
xor U6795 (N_6795,N_6265,N_6446);
nor U6796 (N_6796,N_6284,N_6197);
nand U6797 (N_6797,N_6381,N_6097);
or U6798 (N_6798,N_6076,N_6358);
and U6799 (N_6799,N_6222,N_6269);
or U6800 (N_6800,N_6408,N_6186);
nand U6801 (N_6801,N_6375,N_6407);
nand U6802 (N_6802,N_6282,N_6120);
nor U6803 (N_6803,N_6322,N_6315);
and U6804 (N_6804,N_6427,N_6215);
or U6805 (N_6805,N_6498,N_6108);
or U6806 (N_6806,N_6415,N_6070);
and U6807 (N_6807,N_6299,N_6438);
nor U6808 (N_6808,N_6497,N_6321);
or U6809 (N_6809,N_6116,N_6275);
xor U6810 (N_6810,N_6228,N_6126);
nor U6811 (N_6811,N_6444,N_6239);
nand U6812 (N_6812,N_6115,N_6280);
nand U6813 (N_6813,N_6454,N_6330);
nand U6814 (N_6814,N_6473,N_6472);
nand U6815 (N_6815,N_6344,N_6148);
or U6816 (N_6816,N_6414,N_6388);
or U6817 (N_6817,N_6090,N_6445);
and U6818 (N_6818,N_6301,N_6393);
nor U6819 (N_6819,N_6214,N_6094);
nand U6820 (N_6820,N_6486,N_6348);
nor U6821 (N_6821,N_6153,N_6105);
nor U6822 (N_6822,N_6114,N_6254);
and U6823 (N_6823,N_6210,N_6341);
xnor U6824 (N_6824,N_6128,N_6403);
or U6825 (N_6825,N_6106,N_6434);
nand U6826 (N_6826,N_6141,N_6332);
nor U6827 (N_6827,N_6227,N_6433);
and U6828 (N_6828,N_6073,N_6439);
and U6829 (N_6829,N_6229,N_6209);
nor U6830 (N_6830,N_6205,N_6351);
nand U6831 (N_6831,N_6007,N_6271);
nand U6832 (N_6832,N_6092,N_6341);
or U6833 (N_6833,N_6314,N_6344);
nor U6834 (N_6834,N_6133,N_6064);
nor U6835 (N_6835,N_6383,N_6139);
or U6836 (N_6836,N_6086,N_6087);
nor U6837 (N_6837,N_6226,N_6323);
xnor U6838 (N_6838,N_6468,N_6302);
nor U6839 (N_6839,N_6114,N_6213);
nor U6840 (N_6840,N_6350,N_6206);
and U6841 (N_6841,N_6387,N_6048);
and U6842 (N_6842,N_6338,N_6203);
and U6843 (N_6843,N_6031,N_6082);
nand U6844 (N_6844,N_6244,N_6010);
nor U6845 (N_6845,N_6251,N_6363);
nor U6846 (N_6846,N_6441,N_6142);
nand U6847 (N_6847,N_6403,N_6154);
nand U6848 (N_6848,N_6023,N_6118);
nor U6849 (N_6849,N_6141,N_6169);
nor U6850 (N_6850,N_6292,N_6100);
or U6851 (N_6851,N_6378,N_6423);
nor U6852 (N_6852,N_6419,N_6180);
or U6853 (N_6853,N_6141,N_6426);
nor U6854 (N_6854,N_6492,N_6398);
nand U6855 (N_6855,N_6117,N_6178);
and U6856 (N_6856,N_6299,N_6098);
nand U6857 (N_6857,N_6459,N_6333);
nand U6858 (N_6858,N_6154,N_6120);
or U6859 (N_6859,N_6477,N_6463);
and U6860 (N_6860,N_6321,N_6425);
nor U6861 (N_6861,N_6034,N_6171);
nor U6862 (N_6862,N_6226,N_6202);
nor U6863 (N_6863,N_6184,N_6170);
or U6864 (N_6864,N_6442,N_6199);
nand U6865 (N_6865,N_6182,N_6389);
nand U6866 (N_6866,N_6285,N_6391);
nand U6867 (N_6867,N_6100,N_6096);
and U6868 (N_6868,N_6010,N_6177);
nand U6869 (N_6869,N_6498,N_6295);
nor U6870 (N_6870,N_6065,N_6059);
or U6871 (N_6871,N_6075,N_6096);
nor U6872 (N_6872,N_6370,N_6027);
nor U6873 (N_6873,N_6208,N_6017);
nand U6874 (N_6874,N_6053,N_6383);
and U6875 (N_6875,N_6246,N_6282);
or U6876 (N_6876,N_6388,N_6408);
and U6877 (N_6877,N_6133,N_6456);
nor U6878 (N_6878,N_6474,N_6272);
nand U6879 (N_6879,N_6099,N_6390);
nor U6880 (N_6880,N_6431,N_6469);
nand U6881 (N_6881,N_6221,N_6170);
or U6882 (N_6882,N_6471,N_6406);
nor U6883 (N_6883,N_6335,N_6005);
nor U6884 (N_6884,N_6254,N_6468);
xor U6885 (N_6885,N_6212,N_6130);
nand U6886 (N_6886,N_6291,N_6144);
nor U6887 (N_6887,N_6140,N_6375);
nor U6888 (N_6888,N_6273,N_6471);
nand U6889 (N_6889,N_6194,N_6069);
nand U6890 (N_6890,N_6077,N_6150);
nor U6891 (N_6891,N_6476,N_6075);
or U6892 (N_6892,N_6311,N_6274);
nand U6893 (N_6893,N_6321,N_6171);
and U6894 (N_6894,N_6382,N_6106);
or U6895 (N_6895,N_6256,N_6365);
and U6896 (N_6896,N_6348,N_6255);
and U6897 (N_6897,N_6412,N_6245);
and U6898 (N_6898,N_6228,N_6205);
nor U6899 (N_6899,N_6401,N_6249);
or U6900 (N_6900,N_6120,N_6142);
and U6901 (N_6901,N_6146,N_6463);
xor U6902 (N_6902,N_6197,N_6003);
nand U6903 (N_6903,N_6021,N_6041);
or U6904 (N_6904,N_6201,N_6321);
nor U6905 (N_6905,N_6228,N_6208);
or U6906 (N_6906,N_6262,N_6445);
and U6907 (N_6907,N_6107,N_6379);
or U6908 (N_6908,N_6070,N_6136);
or U6909 (N_6909,N_6186,N_6196);
or U6910 (N_6910,N_6320,N_6085);
nor U6911 (N_6911,N_6416,N_6444);
and U6912 (N_6912,N_6412,N_6410);
and U6913 (N_6913,N_6049,N_6459);
or U6914 (N_6914,N_6007,N_6453);
or U6915 (N_6915,N_6298,N_6143);
and U6916 (N_6916,N_6476,N_6474);
nand U6917 (N_6917,N_6287,N_6314);
nand U6918 (N_6918,N_6413,N_6266);
nand U6919 (N_6919,N_6418,N_6294);
and U6920 (N_6920,N_6132,N_6483);
nand U6921 (N_6921,N_6470,N_6138);
nand U6922 (N_6922,N_6283,N_6052);
nor U6923 (N_6923,N_6166,N_6373);
nand U6924 (N_6924,N_6449,N_6360);
and U6925 (N_6925,N_6486,N_6265);
nor U6926 (N_6926,N_6077,N_6338);
nor U6927 (N_6927,N_6159,N_6382);
nand U6928 (N_6928,N_6458,N_6204);
xor U6929 (N_6929,N_6454,N_6314);
and U6930 (N_6930,N_6469,N_6146);
nor U6931 (N_6931,N_6399,N_6080);
and U6932 (N_6932,N_6181,N_6342);
nor U6933 (N_6933,N_6301,N_6063);
or U6934 (N_6934,N_6112,N_6117);
nand U6935 (N_6935,N_6254,N_6309);
nor U6936 (N_6936,N_6218,N_6319);
or U6937 (N_6937,N_6245,N_6430);
nand U6938 (N_6938,N_6369,N_6016);
or U6939 (N_6939,N_6318,N_6050);
or U6940 (N_6940,N_6016,N_6041);
and U6941 (N_6941,N_6280,N_6173);
nor U6942 (N_6942,N_6159,N_6303);
and U6943 (N_6943,N_6481,N_6189);
and U6944 (N_6944,N_6422,N_6058);
or U6945 (N_6945,N_6159,N_6325);
nand U6946 (N_6946,N_6093,N_6452);
or U6947 (N_6947,N_6326,N_6099);
nand U6948 (N_6948,N_6147,N_6034);
and U6949 (N_6949,N_6240,N_6155);
and U6950 (N_6950,N_6272,N_6111);
and U6951 (N_6951,N_6300,N_6410);
nor U6952 (N_6952,N_6107,N_6374);
or U6953 (N_6953,N_6340,N_6104);
and U6954 (N_6954,N_6298,N_6079);
nor U6955 (N_6955,N_6426,N_6475);
nand U6956 (N_6956,N_6339,N_6027);
nand U6957 (N_6957,N_6475,N_6371);
nand U6958 (N_6958,N_6468,N_6217);
and U6959 (N_6959,N_6063,N_6038);
or U6960 (N_6960,N_6255,N_6005);
nor U6961 (N_6961,N_6099,N_6291);
or U6962 (N_6962,N_6063,N_6290);
and U6963 (N_6963,N_6448,N_6159);
nand U6964 (N_6964,N_6447,N_6091);
and U6965 (N_6965,N_6248,N_6187);
nand U6966 (N_6966,N_6293,N_6359);
or U6967 (N_6967,N_6421,N_6329);
or U6968 (N_6968,N_6429,N_6421);
and U6969 (N_6969,N_6454,N_6274);
nor U6970 (N_6970,N_6169,N_6291);
nor U6971 (N_6971,N_6421,N_6457);
nor U6972 (N_6972,N_6385,N_6497);
and U6973 (N_6973,N_6204,N_6474);
and U6974 (N_6974,N_6469,N_6425);
nand U6975 (N_6975,N_6460,N_6148);
and U6976 (N_6976,N_6322,N_6269);
nor U6977 (N_6977,N_6296,N_6328);
nand U6978 (N_6978,N_6270,N_6126);
nor U6979 (N_6979,N_6058,N_6266);
nor U6980 (N_6980,N_6446,N_6332);
nor U6981 (N_6981,N_6392,N_6222);
and U6982 (N_6982,N_6354,N_6405);
nand U6983 (N_6983,N_6446,N_6337);
nor U6984 (N_6984,N_6096,N_6187);
nor U6985 (N_6985,N_6409,N_6230);
and U6986 (N_6986,N_6069,N_6143);
and U6987 (N_6987,N_6177,N_6093);
nand U6988 (N_6988,N_6451,N_6190);
nand U6989 (N_6989,N_6243,N_6399);
or U6990 (N_6990,N_6472,N_6371);
nand U6991 (N_6991,N_6037,N_6354);
or U6992 (N_6992,N_6442,N_6376);
and U6993 (N_6993,N_6119,N_6065);
and U6994 (N_6994,N_6166,N_6259);
or U6995 (N_6995,N_6485,N_6319);
nor U6996 (N_6996,N_6091,N_6366);
nand U6997 (N_6997,N_6133,N_6034);
nor U6998 (N_6998,N_6450,N_6137);
or U6999 (N_6999,N_6255,N_6408);
or U7000 (N_7000,N_6676,N_6908);
or U7001 (N_7001,N_6708,N_6597);
nand U7002 (N_7002,N_6916,N_6896);
nor U7003 (N_7003,N_6983,N_6873);
or U7004 (N_7004,N_6953,N_6881);
nor U7005 (N_7005,N_6817,N_6756);
nand U7006 (N_7006,N_6914,N_6987);
or U7007 (N_7007,N_6659,N_6872);
nand U7008 (N_7008,N_6792,N_6705);
or U7009 (N_7009,N_6802,N_6982);
nand U7010 (N_7010,N_6605,N_6532);
or U7011 (N_7011,N_6731,N_6910);
nand U7012 (N_7012,N_6939,N_6664);
or U7013 (N_7013,N_6923,N_6500);
nor U7014 (N_7014,N_6846,N_6771);
nand U7015 (N_7015,N_6850,N_6727);
and U7016 (N_7016,N_6685,N_6798);
or U7017 (N_7017,N_6569,N_6822);
and U7018 (N_7018,N_6957,N_6767);
and U7019 (N_7019,N_6578,N_6955);
nor U7020 (N_7020,N_6734,N_6834);
nor U7021 (N_7021,N_6847,N_6996);
and U7022 (N_7022,N_6507,N_6875);
nand U7023 (N_7023,N_6561,N_6815);
or U7024 (N_7024,N_6788,N_6601);
and U7025 (N_7025,N_6512,N_6866);
nand U7026 (N_7026,N_6541,N_6934);
or U7027 (N_7027,N_6775,N_6858);
and U7028 (N_7028,N_6813,N_6820);
nand U7029 (N_7029,N_6511,N_6550);
and U7030 (N_7030,N_6701,N_6535);
nor U7031 (N_7031,N_6743,N_6713);
or U7032 (N_7032,N_6746,N_6593);
and U7033 (N_7033,N_6844,N_6668);
nand U7034 (N_7034,N_6924,N_6869);
nor U7035 (N_7035,N_6629,N_6780);
nor U7036 (N_7036,N_6747,N_6994);
nand U7037 (N_7037,N_6579,N_6964);
nor U7038 (N_7038,N_6645,N_6891);
or U7039 (N_7039,N_6871,N_6922);
nand U7040 (N_7040,N_6962,N_6604);
nor U7041 (N_7041,N_6837,N_6534);
nand U7042 (N_7042,N_6613,N_6735);
nor U7043 (N_7043,N_6989,N_6942);
nand U7044 (N_7044,N_6533,N_6801);
nor U7045 (N_7045,N_6689,N_6918);
nor U7046 (N_7046,N_6588,N_6632);
nor U7047 (N_7047,N_6935,N_6721);
and U7048 (N_7048,N_6856,N_6860);
nand U7049 (N_7049,N_6861,N_6710);
nor U7050 (N_7050,N_6772,N_6599);
nor U7051 (N_7051,N_6811,N_6998);
nand U7052 (N_7052,N_6730,N_6687);
and U7053 (N_7053,N_6696,N_6823);
nand U7054 (N_7054,N_6793,N_6707);
and U7055 (N_7055,N_6821,N_6555);
and U7056 (N_7056,N_6833,N_6724);
nor U7057 (N_7057,N_6651,N_6570);
nor U7058 (N_7058,N_6702,N_6581);
and U7059 (N_7059,N_6819,N_6666);
or U7060 (N_7060,N_6709,N_6516);
or U7061 (N_7061,N_6949,N_6557);
and U7062 (N_7062,N_6531,N_6525);
or U7063 (N_7063,N_6712,N_6648);
nand U7064 (N_7064,N_6976,N_6862);
and U7065 (N_7065,N_6810,N_6562);
nand U7066 (N_7066,N_6538,N_6545);
nor U7067 (N_7067,N_6961,N_6913);
nor U7068 (N_7068,N_6864,N_6673);
nand U7069 (N_7069,N_6971,N_6598);
nand U7070 (N_7070,N_6661,N_6852);
nor U7071 (N_7071,N_6938,N_6754);
and U7072 (N_7072,N_6690,N_6552);
nor U7073 (N_7073,N_6889,N_6768);
xnor U7074 (N_7074,N_6520,N_6654);
nand U7075 (N_7075,N_6585,N_6700);
or U7076 (N_7076,N_6807,N_6510);
xnor U7077 (N_7077,N_6587,N_6635);
or U7078 (N_7078,N_6992,N_6975);
nand U7079 (N_7079,N_6878,N_6519);
or U7080 (N_7080,N_6637,N_6907);
nand U7081 (N_7081,N_6725,N_6655);
nand U7082 (N_7082,N_6703,N_6634);
and U7083 (N_7083,N_6551,N_6619);
nor U7084 (N_7084,N_6733,N_6769);
or U7085 (N_7085,N_6796,N_6610);
xnor U7086 (N_7086,N_6795,N_6740);
or U7087 (N_7087,N_6584,N_6806);
and U7088 (N_7088,N_6715,N_6946);
nand U7089 (N_7089,N_6776,N_6556);
nor U7090 (N_7090,N_6988,N_6506);
nor U7091 (N_7091,N_6867,N_6745);
and U7092 (N_7092,N_6986,N_6773);
or U7093 (N_7093,N_6940,N_6513);
nand U7094 (N_7094,N_6984,N_6699);
and U7095 (N_7095,N_6848,N_6572);
nand U7096 (N_7096,N_6865,N_6919);
and U7097 (N_7097,N_6657,N_6947);
nor U7098 (N_7098,N_6523,N_6517);
nor U7099 (N_7099,N_6602,N_6509);
xor U7100 (N_7100,N_6527,N_6956);
nor U7101 (N_7101,N_6718,N_6717);
and U7102 (N_7102,N_6782,N_6640);
nand U7103 (N_7103,N_6592,N_6893);
xnor U7104 (N_7104,N_6749,N_6722);
nand U7105 (N_7105,N_6894,N_6899);
nand U7106 (N_7106,N_6757,N_6504);
nand U7107 (N_7107,N_6929,N_6609);
xor U7108 (N_7108,N_6620,N_6558);
nor U7109 (N_7109,N_6600,N_6958);
nor U7110 (N_7110,N_6716,N_6933);
and U7111 (N_7111,N_6638,N_6559);
nor U7112 (N_7112,N_6670,N_6571);
and U7113 (N_7113,N_6799,N_6941);
nand U7114 (N_7114,N_6675,N_6627);
nor U7115 (N_7115,N_6880,N_6503);
nor U7116 (N_7116,N_6607,N_6567);
xor U7117 (N_7117,N_6643,N_6658);
nor U7118 (N_7118,N_6783,N_6814);
nor U7119 (N_7119,N_6995,N_6902);
nand U7120 (N_7120,N_6671,N_6892);
and U7121 (N_7121,N_6501,N_6828);
nand U7122 (N_7122,N_6979,N_6662);
or U7123 (N_7123,N_6909,N_6681);
nor U7124 (N_7124,N_6505,N_6750);
nor U7125 (N_7125,N_6800,N_6674);
nor U7126 (N_7126,N_6622,N_6728);
or U7127 (N_7127,N_6583,N_6566);
xor U7128 (N_7128,N_6969,N_6808);
nor U7129 (N_7129,N_6665,N_6830);
or U7130 (N_7130,N_6739,N_6954);
nand U7131 (N_7131,N_6959,N_6835);
or U7132 (N_7132,N_6980,N_6543);
nand U7133 (N_7133,N_6952,N_6568);
or U7134 (N_7134,N_6606,N_6774);
nand U7135 (N_7135,N_6824,N_6649);
or U7136 (N_7136,N_6522,N_6827);
nand U7137 (N_7137,N_6618,N_6762);
and U7138 (N_7138,N_6763,N_6912);
nor U7139 (N_7139,N_6794,N_6879);
nor U7140 (N_7140,N_6832,N_6977);
or U7141 (N_7141,N_6580,N_6732);
or U7142 (N_7142,N_6549,N_6589);
nor U7143 (N_7143,N_6766,N_6921);
nor U7144 (N_7144,N_6777,N_6930);
or U7145 (N_7145,N_6682,N_6943);
nor U7146 (N_7146,N_6925,N_6586);
and U7147 (N_7147,N_6698,N_6626);
and U7148 (N_7148,N_6981,N_6608);
nand U7149 (N_7149,N_6868,N_6797);
nor U7150 (N_7150,N_6960,N_6617);
nor U7151 (N_7151,N_6841,N_6927);
nor U7152 (N_7152,N_6577,N_6787);
nor U7153 (N_7153,N_6818,N_6972);
nor U7154 (N_7154,N_6900,N_6695);
xor U7155 (N_7155,N_6688,N_6529);
nand U7156 (N_7156,N_6677,N_6816);
or U7157 (N_7157,N_6603,N_6853);
and U7158 (N_7158,N_6932,N_6704);
nor U7159 (N_7159,N_6812,N_6784);
nand U7160 (N_7160,N_6755,N_6553);
or U7161 (N_7161,N_6741,N_6697);
nand U7162 (N_7162,N_6778,N_6789);
or U7163 (N_7163,N_6898,N_6886);
nand U7164 (N_7164,N_6874,N_6904);
nand U7165 (N_7165,N_6652,N_6720);
and U7166 (N_7166,N_6653,N_6686);
nor U7167 (N_7167,N_6508,N_6646);
nand U7168 (N_7168,N_6803,N_6680);
and U7169 (N_7169,N_6944,N_6595);
and U7170 (N_7170,N_6905,N_6615);
and U7171 (N_7171,N_6897,N_6758);
and U7172 (N_7172,N_6887,N_6548);
or U7173 (N_7173,N_6694,N_6596);
nor U7174 (N_7174,N_6628,N_6521);
nand U7175 (N_7175,N_6936,N_6781);
or U7176 (N_7176,N_6945,N_6631);
xnor U7177 (N_7177,N_6574,N_6855);
xnor U7178 (N_7178,N_6544,N_6515);
nor U7179 (N_7179,N_6591,N_6966);
nor U7180 (N_7180,N_6711,N_6876);
nand U7181 (N_7181,N_6636,N_6985);
and U7182 (N_7182,N_6642,N_6978);
nand U7183 (N_7183,N_6970,N_6993);
and U7184 (N_7184,N_6920,N_6744);
nor U7185 (N_7185,N_6729,N_6951);
nor U7186 (N_7186,N_6719,N_6616);
or U7187 (N_7187,N_6656,N_6928);
nor U7188 (N_7188,N_6641,N_6890);
and U7189 (N_7189,N_6843,N_6779);
nor U7190 (N_7190,N_6590,N_6693);
and U7191 (N_7191,N_6748,N_6679);
nor U7192 (N_7192,N_6736,N_6851);
nand U7193 (N_7193,N_6594,N_6838);
nand U7194 (N_7194,N_6882,N_6742);
or U7195 (N_7195,N_6915,N_6672);
and U7196 (N_7196,N_6669,N_6564);
or U7197 (N_7197,N_6539,N_6895);
nor U7198 (N_7198,N_6582,N_6528);
nor U7199 (N_7199,N_6963,N_6926);
nand U7200 (N_7200,N_6575,N_6805);
or U7201 (N_7201,N_6565,N_6825);
nor U7202 (N_7202,N_6737,N_6917);
and U7203 (N_7203,N_6804,N_6540);
nor U7204 (N_7204,N_6611,N_6990);
or U7205 (N_7205,N_6831,N_6885);
and U7206 (N_7206,N_6883,N_6790);
or U7207 (N_7207,N_6760,N_6937);
and U7208 (N_7208,N_6621,N_6723);
nor U7209 (N_7209,N_6524,N_6877);
nor U7210 (N_7210,N_6650,N_6931);
and U7211 (N_7211,N_6906,N_6563);
and U7212 (N_7212,N_6859,N_6974);
nor U7213 (N_7213,N_6726,N_6752);
or U7214 (N_7214,N_6842,N_6692);
or U7215 (N_7215,N_6612,N_6968);
and U7216 (N_7216,N_6770,N_6573);
nor U7217 (N_7217,N_6888,N_6826);
nand U7218 (N_7218,N_6546,N_6576);
nand U7219 (N_7219,N_6560,N_6839);
or U7220 (N_7220,N_6870,N_6759);
nor U7221 (N_7221,N_6537,N_6526);
or U7222 (N_7222,N_6765,N_6845);
and U7223 (N_7223,N_6785,N_6836);
or U7224 (N_7224,N_6530,N_6691);
and U7225 (N_7225,N_6863,N_6644);
nand U7226 (N_7226,N_6542,N_6706);
nor U7227 (N_7227,N_6991,N_6663);
nor U7228 (N_7228,N_6684,N_6536);
nor U7229 (N_7229,N_6753,N_6502);
nand U7230 (N_7230,N_6518,N_6547);
nor U7231 (N_7231,N_6809,N_6667);
nand U7232 (N_7232,N_6967,N_6849);
nand U7233 (N_7233,N_6764,N_6623);
nand U7234 (N_7234,N_6554,N_6738);
and U7235 (N_7235,N_6840,N_6614);
xor U7236 (N_7236,N_6630,N_6625);
nand U7237 (N_7237,N_6751,N_6647);
and U7238 (N_7238,N_6854,N_6714);
nor U7239 (N_7239,N_6965,N_6999);
and U7240 (N_7240,N_6911,N_6829);
or U7241 (N_7241,N_6903,N_6514);
or U7242 (N_7242,N_6639,N_6660);
nand U7243 (N_7243,N_6948,N_6761);
or U7244 (N_7244,N_6683,N_6997);
or U7245 (N_7245,N_6791,N_6950);
and U7246 (N_7246,N_6786,N_6857);
or U7247 (N_7247,N_6624,N_6884);
nor U7248 (N_7248,N_6678,N_6633);
nand U7249 (N_7249,N_6973,N_6901);
or U7250 (N_7250,N_6770,N_6907);
and U7251 (N_7251,N_6927,N_6667);
or U7252 (N_7252,N_6650,N_6606);
and U7253 (N_7253,N_6924,N_6621);
xor U7254 (N_7254,N_6648,N_6983);
and U7255 (N_7255,N_6799,N_6503);
or U7256 (N_7256,N_6837,N_6793);
nor U7257 (N_7257,N_6896,N_6628);
or U7258 (N_7258,N_6541,N_6579);
and U7259 (N_7259,N_6636,N_6652);
nand U7260 (N_7260,N_6521,N_6889);
nor U7261 (N_7261,N_6694,N_6715);
nor U7262 (N_7262,N_6817,N_6718);
and U7263 (N_7263,N_6776,N_6908);
nor U7264 (N_7264,N_6577,N_6795);
or U7265 (N_7265,N_6921,N_6912);
or U7266 (N_7266,N_6577,N_6505);
nor U7267 (N_7267,N_6525,N_6556);
nor U7268 (N_7268,N_6575,N_6554);
nand U7269 (N_7269,N_6686,N_6586);
nor U7270 (N_7270,N_6569,N_6683);
or U7271 (N_7271,N_6584,N_6772);
nor U7272 (N_7272,N_6966,N_6765);
and U7273 (N_7273,N_6593,N_6777);
nand U7274 (N_7274,N_6997,N_6726);
nand U7275 (N_7275,N_6708,N_6623);
nand U7276 (N_7276,N_6584,N_6989);
or U7277 (N_7277,N_6932,N_6551);
or U7278 (N_7278,N_6866,N_6774);
or U7279 (N_7279,N_6732,N_6634);
nor U7280 (N_7280,N_6972,N_6648);
and U7281 (N_7281,N_6817,N_6540);
or U7282 (N_7282,N_6933,N_6727);
nor U7283 (N_7283,N_6947,N_6588);
nand U7284 (N_7284,N_6949,N_6816);
or U7285 (N_7285,N_6962,N_6954);
or U7286 (N_7286,N_6727,N_6676);
and U7287 (N_7287,N_6649,N_6832);
or U7288 (N_7288,N_6763,N_6537);
nor U7289 (N_7289,N_6754,N_6521);
or U7290 (N_7290,N_6560,N_6703);
or U7291 (N_7291,N_6736,N_6962);
nand U7292 (N_7292,N_6841,N_6852);
or U7293 (N_7293,N_6560,N_6552);
nand U7294 (N_7294,N_6744,N_6568);
nor U7295 (N_7295,N_6944,N_6816);
and U7296 (N_7296,N_6765,N_6942);
and U7297 (N_7297,N_6740,N_6832);
nor U7298 (N_7298,N_6879,N_6727);
nor U7299 (N_7299,N_6636,N_6676);
or U7300 (N_7300,N_6746,N_6850);
and U7301 (N_7301,N_6999,N_6777);
and U7302 (N_7302,N_6952,N_6989);
nand U7303 (N_7303,N_6704,N_6698);
and U7304 (N_7304,N_6837,N_6815);
or U7305 (N_7305,N_6547,N_6964);
nor U7306 (N_7306,N_6697,N_6813);
or U7307 (N_7307,N_6700,N_6504);
and U7308 (N_7308,N_6634,N_6742);
and U7309 (N_7309,N_6992,N_6657);
nand U7310 (N_7310,N_6790,N_6849);
and U7311 (N_7311,N_6658,N_6639);
nand U7312 (N_7312,N_6575,N_6826);
or U7313 (N_7313,N_6770,N_6858);
nor U7314 (N_7314,N_6509,N_6530);
nand U7315 (N_7315,N_6592,N_6584);
nand U7316 (N_7316,N_6845,N_6955);
or U7317 (N_7317,N_6670,N_6549);
nand U7318 (N_7318,N_6703,N_6773);
xnor U7319 (N_7319,N_6510,N_6783);
nor U7320 (N_7320,N_6887,N_6662);
nand U7321 (N_7321,N_6800,N_6545);
nand U7322 (N_7322,N_6794,N_6558);
nand U7323 (N_7323,N_6828,N_6946);
or U7324 (N_7324,N_6708,N_6749);
and U7325 (N_7325,N_6730,N_6856);
nand U7326 (N_7326,N_6897,N_6841);
and U7327 (N_7327,N_6962,N_6549);
or U7328 (N_7328,N_6742,N_6624);
or U7329 (N_7329,N_6680,N_6812);
nor U7330 (N_7330,N_6828,N_6967);
or U7331 (N_7331,N_6633,N_6909);
nor U7332 (N_7332,N_6612,N_6510);
or U7333 (N_7333,N_6982,N_6729);
nand U7334 (N_7334,N_6802,N_6516);
and U7335 (N_7335,N_6785,N_6884);
nor U7336 (N_7336,N_6711,N_6895);
and U7337 (N_7337,N_6627,N_6576);
xnor U7338 (N_7338,N_6564,N_6932);
and U7339 (N_7339,N_6880,N_6897);
nor U7340 (N_7340,N_6574,N_6711);
nor U7341 (N_7341,N_6947,N_6977);
or U7342 (N_7342,N_6748,N_6784);
nand U7343 (N_7343,N_6610,N_6946);
and U7344 (N_7344,N_6561,N_6510);
or U7345 (N_7345,N_6642,N_6682);
nand U7346 (N_7346,N_6540,N_6918);
and U7347 (N_7347,N_6560,N_6826);
nor U7348 (N_7348,N_6973,N_6746);
or U7349 (N_7349,N_6593,N_6817);
and U7350 (N_7350,N_6732,N_6690);
and U7351 (N_7351,N_6703,N_6570);
nor U7352 (N_7352,N_6779,N_6559);
and U7353 (N_7353,N_6588,N_6854);
or U7354 (N_7354,N_6510,N_6655);
nand U7355 (N_7355,N_6843,N_6956);
or U7356 (N_7356,N_6570,N_6697);
nor U7357 (N_7357,N_6744,N_6820);
or U7358 (N_7358,N_6788,N_6953);
xor U7359 (N_7359,N_6808,N_6736);
nand U7360 (N_7360,N_6701,N_6592);
and U7361 (N_7361,N_6721,N_6574);
nand U7362 (N_7362,N_6795,N_6819);
and U7363 (N_7363,N_6764,N_6655);
or U7364 (N_7364,N_6574,N_6783);
nor U7365 (N_7365,N_6692,N_6955);
nor U7366 (N_7366,N_6699,N_6700);
and U7367 (N_7367,N_6667,N_6938);
and U7368 (N_7368,N_6827,N_6947);
and U7369 (N_7369,N_6504,N_6998);
or U7370 (N_7370,N_6528,N_6945);
nor U7371 (N_7371,N_6830,N_6845);
nor U7372 (N_7372,N_6588,N_6915);
nor U7373 (N_7373,N_6920,N_6741);
nand U7374 (N_7374,N_6525,N_6786);
and U7375 (N_7375,N_6926,N_6571);
nand U7376 (N_7376,N_6609,N_6656);
or U7377 (N_7377,N_6765,N_6601);
or U7378 (N_7378,N_6995,N_6527);
nor U7379 (N_7379,N_6867,N_6863);
nand U7380 (N_7380,N_6738,N_6786);
nand U7381 (N_7381,N_6547,N_6559);
and U7382 (N_7382,N_6969,N_6547);
or U7383 (N_7383,N_6948,N_6711);
and U7384 (N_7384,N_6755,N_6666);
nor U7385 (N_7385,N_6764,N_6586);
nand U7386 (N_7386,N_6768,N_6638);
or U7387 (N_7387,N_6831,N_6606);
nand U7388 (N_7388,N_6825,N_6550);
and U7389 (N_7389,N_6508,N_6835);
and U7390 (N_7390,N_6885,N_6901);
or U7391 (N_7391,N_6665,N_6653);
nand U7392 (N_7392,N_6507,N_6982);
nor U7393 (N_7393,N_6643,N_6921);
and U7394 (N_7394,N_6841,N_6874);
nor U7395 (N_7395,N_6995,N_6500);
nor U7396 (N_7396,N_6944,N_6574);
and U7397 (N_7397,N_6821,N_6928);
xor U7398 (N_7398,N_6738,N_6652);
nor U7399 (N_7399,N_6999,N_6860);
nand U7400 (N_7400,N_6746,N_6922);
or U7401 (N_7401,N_6681,N_6882);
xor U7402 (N_7402,N_6617,N_6709);
nand U7403 (N_7403,N_6825,N_6739);
or U7404 (N_7404,N_6680,N_6703);
nand U7405 (N_7405,N_6825,N_6785);
and U7406 (N_7406,N_6973,N_6753);
and U7407 (N_7407,N_6819,N_6508);
or U7408 (N_7408,N_6638,N_6727);
or U7409 (N_7409,N_6529,N_6987);
and U7410 (N_7410,N_6714,N_6966);
and U7411 (N_7411,N_6691,N_6586);
or U7412 (N_7412,N_6752,N_6894);
or U7413 (N_7413,N_6559,N_6669);
nand U7414 (N_7414,N_6802,N_6964);
and U7415 (N_7415,N_6945,N_6978);
nand U7416 (N_7416,N_6973,N_6593);
and U7417 (N_7417,N_6715,N_6993);
nand U7418 (N_7418,N_6705,N_6858);
nand U7419 (N_7419,N_6640,N_6660);
nand U7420 (N_7420,N_6785,N_6746);
nor U7421 (N_7421,N_6569,N_6550);
xor U7422 (N_7422,N_6587,N_6579);
and U7423 (N_7423,N_6956,N_6977);
nand U7424 (N_7424,N_6517,N_6833);
and U7425 (N_7425,N_6655,N_6643);
nand U7426 (N_7426,N_6923,N_6619);
and U7427 (N_7427,N_6513,N_6615);
and U7428 (N_7428,N_6846,N_6971);
and U7429 (N_7429,N_6799,N_6568);
and U7430 (N_7430,N_6750,N_6952);
nor U7431 (N_7431,N_6814,N_6869);
and U7432 (N_7432,N_6599,N_6560);
or U7433 (N_7433,N_6596,N_6547);
or U7434 (N_7434,N_6870,N_6882);
or U7435 (N_7435,N_6927,N_6902);
and U7436 (N_7436,N_6878,N_6556);
and U7437 (N_7437,N_6763,N_6557);
nor U7438 (N_7438,N_6834,N_6649);
nor U7439 (N_7439,N_6950,N_6646);
nor U7440 (N_7440,N_6613,N_6679);
nand U7441 (N_7441,N_6672,N_6569);
nand U7442 (N_7442,N_6949,N_6714);
nor U7443 (N_7443,N_6704,N_6553);
nor U7444 (N_7444,N_6783,N_6628);
and U7445 (N_7445,N_6625,N_6690);
nor U7446 (N_7446,N_6825,N_6500);
nor U7447 (N_7447,N_6721,N_6934);
and U7448 (N_7448,N_6551,N_6706);
and U7449 (N_7449,N_6818,N_6650);
or U7450 (N_7450,N_6871,N_6879);
and U7451 (N_7451,N_6813,N_6773);
nor U7452 (N_7452,N_6861,N_6907);
nor U7453 (N_7453,N_6722,N_6790);
or U7454 (N_7454,N_6876,N_6752);
and U7455 (N_7455,N_6647,N_6683);
nor U7456 (N_7456,N_6762,N_6946);
nor U7457 (N_7457,N_6619,N_6664);
nand U7458 (N_7458,N_6512,N_6765);
or U7459 (N_7459,N_6614,N_6678);
nand U7460 (N_7460,N_6529,N_6636);
or U7461 (N_7461,N_6572,N_6540);
nand U7462 (N_7462,N_6633,N_6763);
nand U7463 (N_7463,N_6794,N_6753);
nand U7464 (N_7464,N_6949,N_6608);
nand U7465 (N_7465,N_6611,N_6877);
and U7466 (N_7466,N_6519,N_6557);
or U7467 (N_7467,N_6853,N_6842);
and U7468 (N_7468,N_6991,N_6558);
nand U7469 (N_7469,N_6567,N_6796);
or U7470 (N_7470,N_6724,N_6520);
nor U7471 (N_7471,N_6515,N_6955);
nor U7472 (N_7472,N_6738,N_6651);
or U7473 (N_7473,N_6747,N_6518);
nor U7474 (N_7474,N_6877,N_6512);
and U7475 (N_7475,N_6807,N_6823);
and U7476 (N_7476,N_6828,N_6905);
and U7477 (N_7477,N_6606,N_6820);
and U7478 (N_7478,N_6544,N_6854);
nand U7479 (N_7479,N_6848,N_6793);
or U7480 (N_7480,N_6636,N_6605);
nor U7481 (N_7481,N_6557,N_6535);
and U7482 (N_7482,N_6956,N_6737);
or U7483 (N_7483,N_6762,N_6821);
nor U7484 (N_7484,N_6597,N_6967);
nor U7485 (N_7485,N_6624,N_6857);
nand U7486 (N_7486,N_6656,N_6623);
and U7487 (N_7487,N_6898,N_6632);
nor U7488 (N_7488,N_6800,N_6501);
and U7489 (N_7489,N_6529,N_6909);
and U7490 (N_7490,N_6719,N_6933);
nor U7491 (N_7491,N_6961,N_6781);
and U7492 (N_7492,N_6847,N_6703);
nand U7493 (N_7493,N_6834,N_6717);
and U7494 (N_7494,N_6932,N_6647);
nor U7495 (N_7495,N_6701,N_6544);
or U7496 (N_7496,N_6785,N_6998);
nor U7497 (N_7497,N_6745,N_6663);
nor U7498 (N_7498,N_6655,N_6823);
nor U7499 (N_7499,N_6911,N_6971);
and U7500 (N_7500,N_7214,N_7245);
and U7501 (N_7501,N_7140,N_7167);
or U7502 (N_7502,N_7443,N_7078);
and U7503 (N_7503,N_7131,N_7254);
nand U7504 (N_7504,N_7367,N_7386);
or U7505 (N_7505,N_7043,N_7450);
nand U7506 (N_7506,N_7098,N_7217);
and U7507 (N_7507,N_7403,N_7338);
nor U7508 (N_7508,N_7080,N_7392);
or U7509 (N_7509,N_7325,N_7330);
and U7510 (N_7510,N_7289,N_7166);
or U7511 (N_7511,N_7134,N_7455);
and U7512 (N_7512,N_7425,N_7446);
nor U7513 (N_7513,N_7469,N_7086);
or U7514 (N_7514,N_7047,N_7211);
nand U7515 (N_7515,N_7191,N_7288);
and U7516 (N_7516,N_7319,N_7249);
and U7517 (N_7517,N_7116,N_7333);
and U7518 (N_7518,N_7055,N_7454);
and U7519 (N_7519,N_7287,N_7368);
or U7520 (N_7520,N_7421,N_7447);
or U7521 (N_7521,N_7062,N_7173);
or U7522 (N_7522,N_7318,N_7040);
nand U7523 (N_7523,N_7356,N_7073);
nand U7524 (N_7524,N_7076,N_7327);
nor U7525 (N_7525,N_7068,N_7427);
xnor U7526 (N_7526,N_7050,N_7230);
or U7527 (N_7527,N_7185,N_7273);
nor U7528 (N_7528,N_7136,N_7268);
or U7529 (N_7529,N_7188,N_7372);
or U7530 (N_7530,N_7239,N_7498);
and U7531 (N_7531,N_7415,N_7441);
or U7532 (N_7532,N_7381,N_7243);
and U7533 (N_7533,N_7435,N_7194);
and U7534 (N_7534,N_7206,N_7198);
nand U7535 (N_7535,N_7488,N_7432);
and U7536 (N_7536,N_7101,N_7074);
and U7537 (N_7537,N_7046,N_7474);
and U7538 (N_7538,N_7234,N_7100);
nand U7539 (N_7539,N_7088,N_7184);
and U7540 (N_7540,N_7473,N_7277);
nand U7541 (N_7541,N_7144,N_7227);
and U7542 (N_7542,N_7160,N_7499);
nand U7543 (N_7543,N_7495,N_7222);
and U7544 (N_7544,N_7486,N_7020);
and U7545 (N_7545,N_7434,N_7135);
nor U7546 (N_7546,N_7232,N_7099);
or U7547 (N_7547,N_7341,N_7321);
and U7548 (N_7548,N_7155,N_7158);
nor U7549 (N_7549,N_7310,N_7472);
nand U7550 (N_7550,N_7215,N_7260);
and U7551 (N_7551,N_7347,N_7001);
xor U7552 (N_7552,N_7459,N_7458);
nand U7553 (N_7553,N_7487,N_7383);
and U7554 (N_7554,N_7156,N_7219);
or U7555 (N_7555,N_7391,N_7360);
nor U7556 (N_7556,N_7316,N_7393);
nor U7557 (N_7557,N_7023,N_7390);
nor U7558 (N_7558,N_7339,N_7444);
nand U7559 (N_7559,N_7242,N_7352);
xnor U7560 (N_7560,N_7124,N_7409);
or U7561 (N_7561,N_7138,N_7146);
and U7562 (N_7562,N_7478,N_7102);
nor U7563 (N_7563,N_7412,N_7059);
nor U7564 (N_7564,N_7380,N_7344);
nand U7565 (N_7565,N_7428,N_7241);
and U7566 (N_7566,N_7464,N_7233);
and U7567 (N_7567,N_7265,N_7298);
and U7568 (N_7568,N_7027,N_7423);
or U7569 (N_7569,N_7263,N_7125);
and U7570 (N_7570,N_7305,N_7189);
and U7571 (N_7571,N_7448,N_7017);
or U7572 (N_7572,N_7252,N_7422);
nor U7573 (N_7573,N_7104,N_7150);
or U7574 (N_7574,N_7369,N_7121);
or U7575 (N_7575,N_7430,N_7468);
and U7576 (N_7576,N_7250,N_7382);
nor U7577 (N_7577,N_7378,N_7366);
or U7578 (N_7578,N_7183,N_7196);
and U7579 (N_7579,N_7083,N_7168);
nand U7580 (N_7580,N_7304,N_7342);
nand U7581 (N_7581,N_7451,N_7218);
and U7582 (N_7582,N_7373,N_7404);
nand U7583 (N_7583,N_7096,N_7207);
xnor U7584 (N_7584,N_7299,N_7462);
or U7585 (N_7585,N_7240,N_7093);
or U7586 (N_7586,N_7461,N_7034);
or U7587 (N_7587,N_7479,N_7414);
nor U7588 (N_7588,N_7300,N_7110);
nor U7589 (N_7589,N_7351,N_7285);
nor U7590 (N_7590,N_7292,N_7274);
and U7591 (N_7591,N_7114,N_7065);
nand U7592 (N_7592,N_7449,N_7337);
and U7593 (N_7593,N_7037,N_7346);
nand U7594 (N_7594,N_7251,N_7123);
or U7595 (N_7595,N_7008,N_7282);
nand U7596 (N_7596,N_7179,N_7041);
and U7597 (N_7597,N_7259,N_7152);
xnor U7598 (N_7598,N_7332,N_7385);
or U7599 (N_7599,N_7377,N_7416);
nand U7600 (N_7600,N_7224,N_7025);
or U7601 (N_7601,N_7294,N_7089);
nand U7602 (N_7602,N_7496,N_7484);
nand U7603 (N_7603,N_7306,N_7457);
nor U7604 (N_7604,N_7187,N_7405);
and U7605 (N_7605,N_7176,N_7210);
and U7606 (N_7606,N_7220,N_7395);
and U7607 (N_7607,N_7353,N_7445);
or U7608 (N_7608,N_7015,N_7022);
or U7609 (N_7609,N_7387,N_7108);
or U7610 (N_7610,N_7397,N_7112);
nor U7611 (N_7611,N_7328,N_7336);
or U7612 (N_7612,N_7236,N_7293);
xnor U7613 (N_7613,N_7053,N_7313);
nand U7614 (N_7614,N_7141,N_7018);
and U7615 (N_7615,N_7105,N_7154);
nor U7616 (N_7616,N_7480,N_7370);
and U7617 (N_7617,N_7256,N_7401);
nor U7618 (N_7618,N_7231,N_7453);
nor U7619 (N_7619,N_7399,N_7209);
nand U7620 (N_7620,N_7235,N_7129);
nor U7621 (N_7621,N_7054,N_7375);
nor U7622 (N_7622,N_7161,N_7276);
nand U7623 (N_7623,N_7296,N_7190);
or U7624 (N_7624,N_7388,N_7494);
or U7625 (N_7625,N_7085,N_7348);
nor U7626 (N_7626,N_7200,N_7365);
nor U7627 (N_7627,N_7389,N_7255);
nand U7628 (N_7628,N_7270,N_7056);
nand U7629 (N_7629,N_7145,N_7044);
or U7630 (N_7630,N_7402,N_7467);
xor U7631 (N_7631,N_7084,N_7127);
or U7632 (N_7632,N_7005,N_7413);
nand U7633 (N_7633,N_7326,N_7225);
or U7634 (N_7634,N_7315,N_7317);
nand U7635 (N_7635,N_7172,N_7436);
nand U7636 (N_7636,N_7159,N_7475);
xnor U7637 (N_7637,N_7384,N_7364);
or U7638 (N_7638,N_7128,N_7205);
nand U7639 (N_7639,N_7374,N_7257);
nor U7640 (N_7640,N_7039,N_7442);
nand U7641 (N_7641,N_7376,N_7340);
nor U7642 (N_7642,N_7019,N_7262);
and U7643 (N_7643,N_7171,N_7345);
nand U7644 (N_7644,N_7180,N_7379);
and U7645 (N_7645,N_7164,N_7491);
nor U7646 (N_7646,N_7314,N_7106);
nand U7647 (N_7647,N_7320,N_7466);
and U7648 (N_7648,N_7429,N_7431);
nor U7649 (N_7649,N_7186,N_7477);
or U7650 (N_7650,N_7178,N_7117);
nor U7651 (N_7651,N_7290,N_7079);
nand U7652 (N_7652,N_7011,N_7028);
nand U7653 (N_7653,N_7193,N_7440);
nor U7654 (N_7654,N_7077,N_7308);
nand U7655 (N_7655,N_7087,N_7272);
or U7656 (N_7656,N_7036,N_7075);
xor U7657 (N_7657,N_7157,N_7197);
xnor U7658 (N_7658,N_7081,N_7132);
and U7659 (N_7659,N_7139,N_7408);
nand U7660 (N_7660,N_7267,N_7014);
and U7661 (N_7661,N_7358,N_7163);
and U7662 (N_7662,N_7350,N_7226);
nand U7663 (N_7663,N_7174,N_7051);
xor U7664 (N_7664,N_7012,N_7312);
or U7665 (N_7665,N_7029,N_7202);
nand U7666 (N_7666,N_7010,N_7439);
nor U7667 (N_7667,N_7223,N_7357);
or U7668 (N_7668,N_7032,N_7362);
nor U7669 (N_7669,N_7126,N_7109);
and U7670 (N_7670,N_7463,N_7286);
or U7671 (N_7671,N_7063,N_7147);
or U7672 (N_7672,N_7143,N_7323);
nor U7673 (N_7673,N_7301,N_7082);
nand U7674 (N_7674,N_7400,N_7090);
and U7675 (N_7675,N_7111,N_7061);
and U7676 (N_7676,N_7007,N_7302);
nor U7677 (N_7677,N_7275,N_7471);
nor U7678 (N_7678,N_7489,N_7355);
nor U7679 (N_7679,N_7177,N_7066);
and U7680 (N_7680,N_7481,N_7149);
or U7681 (N_7681,N_7057,N_7203);
nand U7682 (N_7682,N_7291,N_7122);
nor U7683 (N_7683,N_7031,N_7004);
nor U7684 (N_7684,N_7070,N_7199);
nor U7685 (N_7685,N_7213,N_7229);
nand U7686 (N_7686,N_7266,N_7006);
nor U7687 (N_7687,N_7192,N_7092);
nand U7688 (N_7688,N_7490,N_7493);
nand U7689 (N_7689,N_7095,N_7411);
nand U7690 (N_7690,N_7151,N_7060);
and U7691 (N_7691,N_7237,N_7309);
nand U7692 (N_7692,N_7281,N_7153);
nand U7693 (N_7693,N_7107,N_7094);
and U7694 (N_7694,N_7212,N_7279);
nand U7695 (N_7695,N_7049,N_7420);
and U7696 (N_7696,N_7331,N_7349);
nor U7697 (N_7697,N_7295,N_7035);
nand U7698 (N_7698,N_7244,N_7119);
nor U7699 (N_7699,N_7284,N_7002);
nor U7700 (N_7700,N_7407,N_7113);
nand U7701 (N_7701,N_7033,N_7115);
and U7702 (N_7702,N_7246,N_7013);
nand U7703 (N_7703,N_7297,N_7137);
nor U7704 (N_7704,N_7433,N_7248);
nor U7705 (N_7705,N_7181,N_7264);
nor U7706 (N_7706,N_7303,N_7394);
nor U7707 (N_7707,N_7465,N_7307);
nand U7708 (N_7708,N_7278,N_7419);
nand U7709 (N_7709,N_7283,N_7361);
nand U7710 (N_7710,N_7343,N_7396);
or U7711 (N_7711,N_7067,N_7359);
and U7712 (N_7712,N_7064,N_7497);
nand U7713 (N_7713,N_7363,N_7120);
nor U7714 (N_7714,N_7335,N_7417);
or U7715 (N_7715,N_7269,N_7485);
xnor U7716 (N_7716,N_7045,N_7170);
nand U7717 (N_7717,N_7118,N_7071);
nor U7718 (N_7718,N_7322,N_7418);
or U7719 (N_7719,N_7334,N_7398);
and U7720 (N_7720,N_7261,N_7311);
and U7721 (N_7721,N_7258,N_7253);
and U7722 (N_7722,N_7072,N_7208);
xor U7723 (N_7723,N_7016,N_7091);
nor U7724 (N_7724,N_7103,N_7042);
and U7725 (N_7725,N_7329,N_7000);
and U7726 (N_7726,N_7476,N_7175);
nand U7727 (N_7727,N_7058,N_7021);
nand U7728 (N_7728,N_7030,N_7182);
and U7729 (N_7729,N_7371,N_7097);
nand U7730 (N_7730,N_7406,N_7201);
nand U7731 (N_7731,N_7026,N_7204);
nand U7732 (N_7732,N_7148,N_7437);
nor U7733 (N_7733,N_7426,N_7228);
nor U7734 (N_7734,N_7354,N_7483);
and U7735 (N_7735,N_7324,N_7162);
nor U7736 (N_7736,N_7424,N_7130);
nand U7737 (N_7737,N_7452,N_7492);
and U7738 (N_7738,N_7169,N_7482);
nor U7739 (N_7739,N_7238,N_7470);
nand U7740 (N_7740,N_7195,N_7410);
nor U7741 (N_7741,N_7271,N_7069);
and U7742 (N_7742,N_7247,N_7165);
nand U7743 (N_7743,N_7038,N_7460);
nor U7744 (N_7744,N_7221,N_7048);
and U7745 (N_7745,N_7133,N_7052);
and U7746 (N_7746,N_7456,N_7003);
nor U7747 (N_7747,N_7009,N_7024);
and U7748 (N_7748,N_7216,N_7280);
or U7749 (N_7749,N_7142,N_7438);
nand U7750 (N_7750,N_7145,N_7260);
and U7751 (N_7751,N_7175,N_7245);
or U7752 (N_7752,N_7200,N_7240);
or U7753 (N_7753,N_7390,N_7483);
nor U7754 (N_7754,N_7174,N_7145);
nand U7755 (N_7755,N_7431,N_7073);
nor U7756 (N_7756,N_7314,N_7216);
or U7757 (N_7757,N_7064,N_7136);
nor U7758 (N_7758,N_7407,N_7339);
nand U7759 (N_7759,N_7198,N_7182);
or U7760 (N_7760,N_7042,N_7437);
or U7761 (N_7761,N_7087,N_7383);
or U7762 (N_7762,N_7206,N_7064);
and U7763 (N_7763,N_7116,N_7447);
and U7764 (N_7764,N_7396,N_7280);
and U7765 (N_7765,N_7040,N_7151);
xor U7766 (N_7766,N_7214,N_7328);
or U7767 (N_7767,N_7083,N_7202);
nor U7768 (N_7768,N_7405,N_7490);
or U7769 (N_7769,N_7029,N_7359);
and U7770 (N_7770,N_7055,N_7146);
nor U7771 (N_7771,N_7073,N_7279);
nor U7772 (N_7772,N_7193,N_7181);
nand U7773 (N_7773,N_7144,N_7017);
nand U7774 (N_7774,N_7198,N_7268);
and U7775 (N_7775,N_7350,N_7426);
nand U7776 (N_7776,N_7132,N_7379);
or U7777 (N_7777,N_7059,N_7137);
or U7778 (N_7778,N_7259,N_7018);
nor U7779 (N_7779,N_7379,N_7213);
and U7780 (N_7780,N_7074,N_7290);
nand U7781 (N_7781,N_7022,N_7078);
nand U7782 (N_7782,N_7388,N_7137);
nor U7783 (N_7783,N_7428,N_7005);
and U7784 (N_7784,N_7076,N_7146);
nand U7785 (N_7785,N_7272,N_7333);
and U7786 (N_7786,N_7176,N_7389);
and U7787 (N_7787,N_7428,N_7205);
nor U7788 (N_7788,N_7048,N_7155);
nor U7789 (N_7789,N_7461,N_7283);
nand U7790 (N_7790,N_7443,N_7199);
nand U7791 (N_7791,N_7375,N_7343);
nand U7792 (N_7792,N_7309,N_7236);
and U7793 (N_7793,N_7220,N_7206);
nand U7794 (N_7794,N_7354,N_7378);
and U7795 (N_7795,N_7336,N_7345);
or U7796 (N_7796,N_7260,N_7376);
nand U7797 (N_7797,N_7206,N_7257);
nor U7798 (N_7798,N_7494,N_7211);
or U7799 (N_7799,N_7279,N_7288);
xor U7800 (N_7800,N_7268,N_7119);
and U7801 (N_7801,N_7058,N_7221);
nand U7802 (N_7802,N_7065,N_7392);
nor U7803 (N_7803,N_7130,N_7289);
nand U7804 (N_7804,N_7437,N_7088);
and U7805 (N_7805,N_7087,N_7232);
or U7806 (N_7806,N_7081,N_7019);
and U7807 (N_7807,N_7493,N_7119);
or U7808 (N_7808,N_7459,N_7249);
and U7809 (N_7809,N_7365,N_7076);
nand U7810 (N_7810,N_7348,N_7478);
nor U7811 (N_7811,N_7438,N_7134);
nand U7812 (N_7812,N_7132,N_7330);
nor U7813 (N_7813,N_7224,N_7197);
nor U7814 (N_7814,N_7472,N_7073);
nand U7815 (N_7815,N_7258,N_7114);
nand U7816 (N_7816,N_7483,N_7240);
or U7817 (N_7817,N_7097,N_7459);
nand U7818 (N_7818,N_7393,N_7239);
and U7819 (N_7819,N_7227,N_7173);
nor U7820 (N_7820,N_7435,N_7392);
and U7821 (N_7821,N_7493,N_7105);
and U7822 (N_7822,N_7239,N_7455);
nand U7823 (N_7823,N_7209,N_7079);
nand U7824 (N_7824,N_7238,N_7365);
nand U7825 (N_7825,N_7263,N_7016);
and U7826 (N_7826,N_7347,N_7353);
and U7827 (N_7827,N_7193,N_7386);
or U7828 (N_7828,N_7262,N_7173);
nor U7829 (N_7829,N_7396,N_7207);
nor U7830 (N_7830,N_7147,N_7202);
nor U7831 (N_7831,N_7486,N_7314);
and U7832 (N_7832,N_7070,N_7148);
and U7833 (N_7833,N_7365,N_7356);
nor U7834 (N_7834,N_7157,N_7382);
nor U7835 (N_7835,N_7339,N_7125);
nor U7836 (N_7836,N_7368,N_7032);
and U7837 (N_7837,N_7456,N_7130);
and U7838 (N_7838,N_7256,N_7459);
nand U7839 (N_7839,N_7442,N_7086);
and U7840 (N_7840,N_7315,N_7000);
nand U7841 (N_7841,N_7127,N_7091);
or U7842 (N_7842,N_7396,N_7179);
nand U7843 (N_7843,N_7461,N_7446);
and U7844 (N_7844,N_7270,N_7207);
nor U7845 (N_7845,N_7350,N_7090);
or U7846 (N_7846,N_7065,N_7211);
nand U7847 (N_7847,N_7281,N_7177);
xnor U7848 (N_7848,N_7026,N_7184);
nand U7849 (N_7849,N_7309,N_7375);
or U7850 (N_7850,N_7218,N_7348);
and U7851 (N_7851,N_7165,N_7019);
or U7852 (N_7852,N_7080,N_7023);
and U7853 (N_7853,N_7274,N_7073);
nor U7854 (N_7854,N_7216,N_7250);
and U7855 (N_7855,N_7337,N_7010);
nand U7856 (N_7856,N_7224,N_7406);
xnor U7857 (N_7857,N_7175,N_7202);
or U7858 (N_7858,N_7346,N_7295);
nor U7859 (N_7859,N_7083,N_7282);
nor U7860 (N_7860,N_7447,N_7207);
or U7861 (N_7861,N_7413,N_7144);
and U7862 (N_7862,N_7263,N_7467);
nor U7863 (N_7863,N_7245,N_7015);
nand U7864 (N_7864,N_7327,N_7386);
or U7865 (N_7865,N_7037,N_7203);
nand U7866 (N_7866,N_7049,N_7326);
nor U7867 (N_7867,N_7230,N_7161);
nand U7868 (N_7868,N_7323,N_7445);
nor U7869 (N_7869,N_7229,N_7221);
or U7870 (N_7870,N_7430,N_7302);
nand U7871 (N_7871,N_7254,N_7026);
nor U7872 (N_7872,N_7479,N_7166);
xor U7873 (N_7873,N_7006,N_7031);
nor U7874 (N_7874,N_7360,N_7207);
or U7875 (N_7875,N_7281,N_7213);
and U7876 (N_7876,N_7060,N_7256);
nand U7877 (N_7877,N_7231,N_7133);
nor U7878 (N_7878,N_7197,N_7269);
nor U7879 (N_7879,N_7164,N_7435);
nand U7880 (N_7880,N_7300,N_7394);
nand U7881 (N_7881,N_7169,N_7175);
nor U7882 (N_7882,N_7282,N_7451);
nor U7883 (N_7883,N_7167,N_7191);
nand U7884 (N_7884,N_7364,N_7183);
or U7885 (N_7885,N_7181,N_7136);
nor U7886 (N_7886,N_7085,N_7247);
and U7887 (N_7887,N_7111,N_7043);
and U7888 (N_7888,N_7047,N_7273);
or U7889 (N_7889,N_7166,N_7322);
nor U7890 (N_7890,N_7142,N_7240);
and U7891 (N_7891,N_7435,N_7360);
nand U7892 (N_7892,N_7498,N_7076);
or U7893 (N_7893,N_7346,N_7012);
nor U7894 (N_7894,N_7194,N_7248);
nor U7895 (N_7895,N_7066,N_7315);
and U7896 (N_7896,N_7408,N_7446);
or U7897 (N_7897,N_7283,N_7435);
and U7898 (N_7898,N_7118,N_7157);
or U7899 (N_7899,N_7307,N_7216);
and U7900 (N_7900,N_7238,N_7369);
or U7901 (N_7901,N_7447,N_7287);
or U7902 (N_7902,N_7242,N_7063);
nor U7903 (N_7903,N_7467,N_7351);
nand U7904 (N_7904,N_7293,N_7038);
and U7905 (N_7905,N_7356,N_7062);
nand U7906 (N_7906,N_7053,N_7409);
and U7907 (N_7907,N_7423,N_7365);
and U7908 (N_7908,N_7048,N_7377);
xor U7909 (N_7909,N_7263,N_7233);
xor U7910 (N_7910,N_7052,N_7498);
nor U7911 (N_7911,N_7491,N_7333);
and U7912 (N_7912,N_7269,N_7058);
or U7913 (N_7913,N_7098,N_7090);
and U7914 (N_7914,N_7065,N_7486);
and U7915 (N_7915,N_7197,N_7027);
nand U7916 (N_7916,N_7229,N_7417);
nand U7917 (N_7917,N_7003,N_7093);
and U7918 (N_7918,N_7159,N_7408);
nor U7919 (N_7919,N_7029,N_7145);
nor U7920 (N_7920,N_7000,N_7336);
or U7921 (N_7921,N_7333,N_7088);
and U7922 (N_7922,N_7231,N_7455);
xor U7923 (N_7923,N_7144,N_7261);
nand U7924 (N_7924,N_7095,N_7363);
nor U7925 (N_7925,N_7324,N_7034);
nand U7926 (N_7926,N_7336,N_7255);
nand U7927 (N_7927,N_7062,N_7357);
nor U7928 (N_7928,N_7396,N_7159);
xnor U7929 (N_7929,N_7365,N_7191);
and U7930 (N_7930,N_7440,N_7035);
and U7931 (N_7931,N_7304,N_7331);
nor U7932 (N_7932,N_7086,N_7488);
nand U7933 (N_7933,N_7295,N_7213);
nor U7934 (N_7934,N_7394,N_7015);
and U7935 (N_7935,N_7302,N_7457);
nand U7936 (N_7936,N_7181,N_7258);
nand U7937 (N_7937,N_7446,N_7160);
nand U7938 (N_7938,N_7116,N_7397);
nor U7939 (N_7939,N_7149,N_7008);
nor U7940 (N_7940,N_7149,N_7188);
nand U7941 (N_7941,N_7127,N_7234);
nor U7942 (N_7942,N_7002,N_7194);
and U7943 (N_7943,N_7217,N_7184);
nand U7944 (N_7944,N_7007,N_7345);
and U7945 (N_7945,N_7282,N_7377);
or U7946 (N_7946,N_7485,N_7117);
nor U7947 (N_7947,N_7077,N_7039);
nand U7948 (N_7948,N_7063,N_7240);
nand U7949 (N_7949,N_7276,N_7449);
nor U7950 (N_7950,N_7484,N_7416);
nor U7951 (N_7951,N_7112,N_7460);
nand U7952 (N_7952,N_7435,N_7156);
and U7953 (N_7953,N_7195,N_7138);
and U7954 (N_7954,N_7202,N_7484);
nand U7955 (N_7955,N_7185,N_7236);
and U7956 (N_7956,N_7402,N_7389);
nand U7957 (N_7957,N_7493,N_7200);
or U7958 (N_7958,N_7281,N_7161);
and U7959 (N_7959,N_7001,N_7336);
or U7960 (N_7960,N_7250,N_7274);
nor U7961 (N_7961,N_7185,N_7154);
nand U7962 (N_7962,N_7214,N_7009);
nor U7963 (N_7963,N_7392,N_7422);
and U7964 (N_7964,N_7432,N_7024);
nor U7965 (N_7965,N_7222,N_7423);
or U7966 (N_7966,N_7221,N_7434);
nand U7967 (N_7967,N_7185,N_7250);
nor U7968 (N_7968,N_7349,N_7147);
and U7969 (N_7969,N_7159,N_7479);
and U7970 (N_7970,N_7380,N_7452);
or U7971 (N_7971,N_7024,N_7263);
or U7972 (N_7972,N_7150,N_7419);
nor U7973 (N_7973,N_7174,N_7034);
nor U7974 (N_7974,N_7376,N_7009);
xnor U7975 (N_7975,N_7142,N_7051);
nor U7976 (N_7976,N_7360,N_7127);
nor U7977 (N_7977,N_7060,N_7176);
nor U7978 (N_7978,N_7153,N_7173);
or U7979 (N_7979,N_7357,N_7191);
or U7980 (N_7980,N_7366,N_7471);
or U7981 (N_7981,N_7205,N_7146);
nor U7982 (N_7982,N_7326,N_7218);
and U7983 (N_7983,N_7362,N_7262);
and U7984 (N_7984,N_7050,N_7060);
or U7985 (N_7985,N_7361,N_7001);
and U7986 (N_7986,N_7070,N_7197);
nor U7987 (N_7987,N_7074,N_7053);
nor U7988 (N_7988,N_7419,N_7079);
and U7989 (N_7989,N_7085,N_7324);
nor U7990 (N_7990,N_7209,N_7216);
nand U7991 (N_7991,N_7171,N_7388);
nand U7992 (N_7992,N_7331,N_7341);
nor U7993 (N_7993,N_7089,N_7469);
or U7994 (N_7994,N_7294,N_7040);
nor U7995 (N_7995,N_7016,N_7456);
or U7996 (N_7996,N_7350,N_7292);
and U7997 (N_7997,N_7422,N_7006);
or U7998 (N_7998,N_7242,N_7325);
nand U7999 (N_7999,N_7237,N_7010);
and U8000 (N_8000,N_7735,N_7693);
nor U8001 (N_8001,N_7800,N_7560);
nor U8002 (N_8002,N_7563,N_7908);
nand U8003 (N_8003,N_7681,N_7902);
or U8004 (N_8004,N_7596,N_7981);
and U8005 (N_8005,N_7538,N_7533);
nand U8006 (N_8006,N_7948,N_7620);
and U8007 (N_8007,N_7973,N_7879);
and U8008 (N_8008,N_7933,N_7992);
nand U8009 (N_8009,N_7710,N_7860);
nor U8010 (N_8010,N_7656,N_7896);
and U8011 (N_8011,N_7674,N_7816);
nor U8012 (N_8012,N_7988,N_7873);
nor U8013 (N_8013,N_7904,N_7773);
nand U8014 (N_8014,N_7820,N_7787);
nand U8015 (N_8015,N_7959,N_7892);
nand U8016 (N_8016,N_7612,N_7502);
xnor U8017 (N_8017,N_7545,N_7601);
nor U8018 (N_8018,N_7870,N_7853);
and U8019 (N_8019,N_7962,N_7554);
and U8020 (N_8020,N_7876,N_7742);
nand U8021 (N_8021,N_7914,N_7971);
nor U8022 (N_8022,N_7659,N_7878);
nand U8023 (N_8023,N_7778,N_7667);
nand U8024 (N_8024,N_7907,N_7516);
or U8025 (N_8025,N_7635,N_7969);
nand U8026 (N_8026,N_7552,N_7996);
nand U8027 (N_8027,N_7805,N_7759);
nand U8028 (N_8028,N_7950,N_7544);
nor U8029 (N_8029,N_7925,N_7994);
and U8030 (N_8030,N_7526,N_7866);
and U8031 (N_8031,N_7966,N_7883);
and U8032 (N_8032,N_7676,N_7776);
nor U8033 (N_8033,N_7529,N_7758);
or U8034 (N_8034,N_7649,N_7802);
nand U8035 (N_8035,N_7891,N_7855);
nor U8036 (N_8036,N_7786,N_7598);
nand U8037 (N_8037,N_7650,N_7827);
or U8038 (N_8038,N_7595,N_7726);
nor U8039 (N_8039,N_7846,N_7520);
nand U8040 (N_8040,N_7568,N_7509);
nor U8041 (N_8041,N_7547,N_7647);
and U8042 (N_8042,N_7572,N_7641);
or U8043 (N_8043,N_7909,N_7843);
nor U8044 (N_8044,N_7872,N_7818);
nand U8045 (N_8045,N_7690,N_7968);
or U8046 (N_8046,N_7721,N_7922);
or U8047 (N_8047,N_7637,N_7817);
xnor U8048 (N_8048,N_7849,N_7588);
nand U8049 (N_8049,N_7730,N_7836);
xor U8050 (N_8050,N_7956,N_7862);
xor U8051 (N_8051,N_7986,N_7884);
or U8052 (N_8052,N_7675,N_7734);
and U8053 (N_8053,N_7915,N_7643);
nor U8054 (N_8054,N_7731,N_7688);
and U8055 (N_8055,N_7889,N_7733);
and U8056 (N_8056,N_7718,N_7506);
nor U8057 (N_8057,N_7508,N_7597);
nor U8058 (N_8058,N_7703,N_7753);
and U8059 (N_8059,N_7871,N_7531);
xnor U8060 (N_8060,N_7662,N_7697);
nand U8061 (N_8061,N_7760,N_7723);
and U8062 (N_8062,N_7581,N_7685);
nand U8063 (N_8063,N_7768,N_7946);
nor U8064 (N_8064,N_7522,N_7897);
or U8065 (N_8065,N_7608,N_7527);
nor U8066 (N_8066,N_7928,N_7737);
nand U8067 (N_8067,N_7864,N_7744);
or U8068 (N_8068,N_7810,N_7574);
nor U8069 (N_8069,N_7642,N_7717);
nand U8070 (N_8070,N_7664,N_7792);
and U8071 (N_8071,N_7652,N_7648);
nor U8072 (N_8072,N_7706,N_7829);
or U8073 (N_8073,N_7622,N_7705);
nor U8074 (N_8074,N_7707,N_7566);
or U8075 (N_8075,N_7793,N_7765);
and U8076 (N_8076,N_7540,N_7606);
and U8077 (N_8077,N_7580,N_7607);
nand U8078 (N_8078,N_7628,N_7974);
or U8079 (N_8079,N_7539,N_7809);
nand U8080 (N_8080,N_7811,N_7854);
xnor U8081 (N_8081,N_7761,N_7739);
nor U8082 (N_8082,N_7720,N_7813);
and U8083 (N_8083,N_7774,N_7747);
xnor U8084 (N_8084,N_7752,N_7562);
nand U8085 (N_8085,N_7625,N_7558);
xnor U8086 (N_8086,N_7541,N_7646);
nor U8087 (N_8087,N_7746,N_7632);
and U8088 (N_8088,N_7513,N_7828);
and U8089 (N_8089,N_7847,N_7672);
or U8090 (N_8090,N_7604,N_7535);
and U8091 (N_8091,N_7963,N_7900);
nand U8092 (N_8092,N_7748,N_7947);
or U8093 (N_8093,N_7848,N_7831);
and U8094 (N_8094,N_7594,N_7781);
nand U8095 (N_8095,N_7824,N_7934);
or U8096 (N_8096,N_7964,N_7939);
nand U8097 (N_8097,N_7658,N_7957);
or U8098 (N_8098,N_7832,N_7624);
nand U8099 (N_8099,N_7584,N_7524);
nor U8100 (N_8100,N_7655,N_7867);
nand U8101 (N_8101,N_7954,N_7755);
or U8102 (N_8102,N_7953,N_7923);
and U8103 (N_8103,N_7905,N_7521);
xnor U8104 (N_8104,N_7851,N_7979);
nand U8105 (N_8105,N_7769,N_7729);
nor U8106 (N_8106,N_7791,N_7633);
nor U8107 (N_8107,N_7906,N_7546);
nand U8108 (N_8108,N_7550,N_7770);
and U8109 (N_8109,N_7927,N_7715);
or U8110 (N_8110,N_7615,N_7743);
nor U8111 (N_8111,N_7796,N_7868);
or U8112 (N_8112,N_7570,N_7921);
xnor U8113 (N_8113,N_7799,N_7943);
or U8114 (N_8114,N_7949,N_7998);
nand U8115 (N_8115,N_7630,N_7689);
or U8116 (N_8116,N_7888,N_7789);
nor U8117 (N_8117,N_7670,N_7602);
nand U8118 (N_8118,N_7865,N_7727);
nor U8119 (N_8119,N_7579,N_7911);
or U8120 (N_8120,N_7750,N_7638);
and U8121 (N_8121,N_7525,N_7702);
nand U8122 (N_8122,N_7712,N_7698);
or U8123 (N_8123,N_7826,N_7795);
nand U8124 (N_8124,N_7627,N_7859);
and U8125 (N_8125,N_7543,N_7593);
and U8126 (N_8126,N_7610,N_7919);
or U8127 (N_8127,N_7852,N_7980);
nor U8128 (N_8128,N_7613,N_7977);
nand U8129 (N_8129,N_7775,N_7751);
nand U8130 (N_8130,N_7634,N_7970);
or U8131 (N_8131,N_7600,N_7975);
and U8132 (N_8132,N_7993,N_7619);
nor U8133 (N_8133,N_7893,N_7640);
and U8134 (N_8134,N_7504,N_7930);
and U8135 (N_8135,N_7571,N_7519);
or U8136 (N_8136,N_7987,N_7589);
nor U8137 (N_8137,N_7567,N_7823);
nand U8138 (N_8138,N_7825,N_7585);
and U8139 (N_8139,N_7976,N_7569);
or U8140 (N_8140,N_7515,N_7808);
or U8141 (N_8141,N_7575,N_7917);
and U8142 (N_8142,N_7740,N_7532);
nor U8143 (N_8143,N_7679,N_7621);
and U8144 (N_8144,N_7582,N_7666);
and U8145 (N_8145,N_7645,N_7784);
nor U8146 (N_8146,N_7899,N_7565);
or U8147 (N_8147,N_7590,N_7777);
nor U8148 (N_8148,N_7901,N_7938);
or U8149 (N_8149,N_7537,N_7653);
nand U8150 (N_8150,N_7920,N_7629);
nand U8151 (N_8151,N_7686,N_7944);
and U8152 (N_8152,N_7834,N_7680);
and U8153 (N_8153,N_7692,N_7991);
nand U8154 (N_8154,N_7678,N_7910);
and U8155 (N_8155,N_7814,N_7704);
nand U8156 (N_8156,N_7912,N_7591);
nor U8157 (N_8157,N_7644,N_7534);
or U8158 (N_8158,N_7983,N_7687);
or U8159 (N_8159,N_7990,N_7833);
nand U8160 (N_8160,N_7728,N_7882);
or U8161 (N_8161,N_7556,N_7790);
nand U8162 (N_8162,N_7766,N_7738);
nor U8163 (N_8163,N_7941,N_7623);
and U8164 (N_8164,N_7945,N_7995);
nor U8165 (N_8165,N_7691,N_7609);
or U8166 (N_8166,N_7542,N_7782);
nand U8167 (N_8167,N_7783,N_7505);
and U8168 (N_8168,N_7756,N_7835);
and U8169 (N_8169,N_7788,N_7564);
nor U8170 (N_8170,N_7815,N_7618);
nand U8171 (N_8171,N_7603,N_7955);
nor U8172 (N_8172,N_7812,N_7931);
nand U8173 (N_8173,N_7952,N_7741);
nand U8174 (N_8174,N_7695,N_7951);
nor U8175 (N_8175,N_7654,N_7576);
and U8176 (N_8176,N_7785,N_7772);
or U8177 (N_8177,N_7821,N_7507);
and U8178 (N_8178,N_7699,N_7555);
or U8179 (N_8179,N_7913,N_7780);
nor U8180 (N_8180,N_7757,N_7985);
and U8181 (N_8181,N_7557,N_7840);
or U8182 (N_8182,N_7561,N_7961);
nand U8183 (N_8183,N_7500,N_7663);
or U8184 (N_8184,N_7617,N_7665);
and U8185 (N_8185,N_7551,N_7965);
nand U8186 (N_8186,N_7982,N_7709);
nand U8187 (N_8187,N_7501,N_7577);
nor U8188 (N_8188,N_7794,N_7745);
or U8189 (N_8189,N_7850,N_7586);
and U8190 (N_8190,N_7837,N_7636);
nor U8191 (N_8191,N_7510,N_7762);
nor U8192 (N_8192,N_7935,N_7578);
and U8193 (N_8193,N_7881,N_7696);
nor U8194 (N_8194,N_7651,N_7940);
nand U8195 (N_8195,N_7845,N_7708);
or U8196 (N_8196,N_7536,N_7682);
and U8197 (N_8197,N_7725,N_7803);
and U8198 (N_8198,N_7503,N_7918);
or U8199 (N_8199,N_7839,N_7895);
nor U8200 (N_8200,N_7523,N_7880);
or U8201 (N_8201,N_7858,N_7989);
nor U8202 (N_8202,N_7614,N_7926);
nand U8203 (N_8203,N_7886,N_7916);
nor U8204 (N_8204,N_7749,N_7631);
nand U8205 (N_8205,N_7877,N_7937);
and U8206 (N_8206,N_7771,N_7830);
nor U8207 (N_8207,N_7801,N_7549);
or U8208 (N_8208,N_7657,N_7804);
and U8209 (N_8209,N_7700,N_7898);
nand U8210 (N_8210,N_7514,N_7713);
or U8211 (N_8211,N_7517,N_7716);
and U8212 (N_8212,N_7626,N_7719);
or U8213 (N_8213,N_7863,N_7844);
nand U8214 (N_8214,N_7605,N_7779);
and U8215 (N_8215,N_7997,N_7885);
nor U8216 (N_8216,N_7819,N_7714);
nor U8217 (N_8217,N_7861,N_7677);
nand U8218 (N_8218,N_7763,N_7967);
or U8219 (N_8219,N_7694,N_7512);
nand U8220 (N_8220,N_7932,N_7684);
nand U8221 (N_8221,N_7924,N_7936);
nor U8222 (N_8222,N_7806,N_7972);
or U8223 (N_8223,N_7999,N_7559);
or U8224 (N_8224,N_7583,N_7856);
nor U8225 (N_8225,N_7869,N_7822);
nor U8226 (N_8226,N_7671,N_7838);
or U8227 (N_8227,N_7736,N_7875);
nand U8228 (N_8228,N_7669,N_7530);
nor U8229 (N_8229,N_7668,N_7661);
and U8230 (N_8230,N_7890,N_7528);
or U8231 (N_8231,N_7599,N_7857);
nand U8232 (N_8232,N_7978,N_7660);
or U8233 (N_8233,N_7611,N_7767);
or U8234 (N_8234,N_7683,N_7797);
nor U8235 (N_8235,N_7894,N_7842);
or U8236 (N_8236,N_7722,N_7732);
or U8237 (N_8237,N_7553,N_7887);
nand U8238 (N_8238,N_7841,N_7548);
nand U8239 (N_8239,N_7616,N_7701);
or U8240 (N_8240,N_7807,N_7673);
and U8241 (N_8241,N_7724,N_7874);
or U8242 (N_8242,N_7798,N_7764);
or U8243 (N_8243,N_7754,N_7518);
and U8244 (N_8244,N_7592,N_7639);
or U8245 (N_8245,N_7711,N_7984);
or U8246 (N_8246,N_7587,N_7942);
nand U8247 (N_8247,N_7960,N_7511);
nor U8248 (N_8248,N_7573,N_7929);
nand U8249 (N_8249,N_7958,N_7903);
or U8250 (N_8250,N_7712,N_7629);
nor U8251 (N_8251,N_7957,N_7843);
and U8252 (N_8252,N_7656,N_7729);
nor U8253 (N_8253,N_7889,N_7912);
nand U8254 (N_8254,N_7927,N_7977);
and U8255 (N_8255,N_7538,N_7544);
nand U8256 (N_8256,N_7889,N_7719);
or U8257 (N_8257,N_7968,N_7595);
nand U8258 (N_8258,N_7896,N_7863);
nor U8259 (N_8259,N_7573,N_7778);
or U8260 (N_8260,N_7853,N_7652);
xnor U8261 (N_8261,N_7794,N_7687);
nand U8262 (N_8262,N_7522,N_7590);
or U8263 (N_8263,N_7551,N_7692);
nand U8264 (N_8264,N_7766,N_7934);
nor U8265 (N_8265,N_7697,N_7803);
nand U8266 (N_8266,N_7602,N_7660);
nand U8267 (N_8267,N_7666,N_7500);
nand U8268 (N_8268,N_7521,N_7652);
nand U8269 (N_8269,N_7861,N_7685);
nand U8270 (N_8270,N_7801,N_7800);
nor U8271 (N_8271,N_7552,N_7595);
xor U8272 (N_8272,N_7821,N_7820);
and U8273 (N_8273,N_7968,N_7800);
nand U8274 (N_8274,N_7759,N_7695);
nor U8275 (N_8275,N_7757,N_7760);
and U8276 (N_8276,N_7671,N_7647);
nand U8277 (N_8277,N_7804,N_7582);
or U8278 (N_8278,N_7654,N_7627);
xor U8279 (N_8279,N_7532,N_7938);
nand U8280 (N_8280,N_7982,N_7614);
xnor U8281 (N_8281,N_7612,N_7694);
and U8282 (N_8282,N_7616,N_7596);
nor U8283 (N_8283,N_7592,N_7574);
nand U8284 (N_8284,N_7901,N_7549);
or U8285 (N_8285,N_7630,N_7777);
and U8286 (N_8286,N_7801,N_7794);
nor U8287 (N_8287,N_7508,N_7773);
nand U8288 (N_8288,N_7776,N_7521);
nor U8289 (N_8289,N_7832,N_7596);
nand U8290 (N_8290,N_7882,N_7863);
and U8291 (N_8291,N_7617,N_7989);
or U8292 (N_8292,N_7993,N_7802);
or U8293 (N_8293,N_7937,N_7611);
and U8294 (N_8294,N_7902,N_7660);
and U8295 (N_8295,N_7920,N_7550);
nand U8296 (N_8296,N_7964,N_7723);
nor U8297 (N_8297,N_7911,N_7644);
and U8298 (N_8298,N_7774,N_7729);
nand U8299 (N_8299,N_7985,N_7834);
nor U8300 (N_8300,N_7631,N_7521);
or U8301 (N_8301,N_7934,N_7731);
nand U8302 (N_8302,N_7505,N_7601);
nand U8303 (N_8303,N_7950,N_7780);
nand U8304 (N_8304,N_7879,N_7530);
nor U8305 (N_8305,N_7695,N_7691);
xnor U8306 (N_8306,N_7923,N_7637);
nand U8307 (N_8307,N_7989,N_7820);
and U8308 (N_8308,N_7801,N_7707);
xnor U8309 (N_8309,N_7699,N_7892);
nand U8310 (N_8310,N_7904,N_7582);
or U8311 (N_8311,N_7992,N_7919);
or U8312 (N_8312,N_7715,N_7740);
nand U8313 (N_8313,N_7755,N_7559);
or U8314 (N_8314,N_7719,N_7591);
or U8315 (N_8315,N_7962,N_7891);
and U8316 (N_8316,N_7601,N_7633);
nand U8317 (N_8317,N_7983,N_7744);
nor U8318 (N_8318,N_7634,N_7655);
nor U8319 (N_8319,N_7574,N_7747);
nor U8320 (N_8320,N_7933,N_7881);
or U8321 (N_8321,N_7559,N_7869);
nand U8322 (N_8322,N_7656,N_7861);
or U8323 (N_8323,N_7978,N_7921);
nor U8324 (N_8324,N_7844,N_7520);
and U8325 (N_8325,N_7797,N_7534);
or U8326 (N_8326,N_7767,N_7534);
nor U8327 (N_8327,N_7882,N_7983);
and U8328 (N_8328,N_7914,N_7534);
nand U8329 (N_8329,N_7881,N_7692);
and U8330 (N_8330,N_7842,N_7973);
or U8331 (N_8331,N_7905,N_7955);
and U8332 (N_8332,N_7706,N_7739);
and U8333 (N_8333,N_7742,N_7508);
nor U8334 (N_8334,N_7987,N_7774);
and U8335 (N_8335,N_7509,N_7891);
nand U8336 (N_8336,N_7633,N_7518);
nor U8337 (N_8337,N_7849,N_7570);
nand U8338 (N_8338,N_7722,N_7533);
nor U8339 (N_8339,N_7657,N_7625);
and U8340 (N_8340,N_7670,N_7699);
or U8341 (N_8341,N_7759,N_7751);
nor U8342 (N_8342,N_7833,N_7982);
and U8343 (N_8343,N_7818,N_7896);
and U8344 (N_8344,N_7659,N_7795);
nand U8345 (N_8345,N_7721,N_7630);
nand U8346 (N_8346,N_7515,N_7771);
nand U8347 (N_8347,N_7919,N_7675);
nand U8348 (N_8348,N_7621,N_7885);
and U8349 (N_8349,N_7919,N_7757);
nor U8350 (N_8350,N_7882,N_7877);
or U8351 (N_8351,N_7504,N_7835);
nand U8352 (N_8352,N_7752,N_7576);
and U8353 (N_8353,N_7697,N_7717);
nor U8354 (N_8354,N_7635,N_7627);
or U8355 (N_8355,N_7574,N_7889);
and U8356 (N_8356,N_7928,N_7875);
or U8357 (N_8357,N_7848,N_7631);
and U8358 (N_8358,N_7520,N_7513);
or U8359 (N_8359,N_7931,N_7792);
and U8360 (N_8360,N_7599,N_7922);
nand U8361 (N_8361,N_7703,N_7986);
nand U8362 (N_8362,N_7944,N_7518);
nand U8363 (N_8363,N_7860,N_7933);
nand U8364 (N_8364,N_7894,N_7600);
nand U8365 (N_8365,N_7925,N_7820);
and U8366 (N_8366,N_7959,N_7980);
or U8367 (N_8367,N_7857,N_7554);
and U8368 (N_8368,N_7743,N_7751);
nand U8369 (N_8369,N_7504,N_7641);
or U8370 (N_8370,N_7831,N_7641);
or U8371 (N_8371,N_7782,N_7547);
or U8372 (N_8372,N_7759,N_7575);
xnor U8373 (N_8373,N_7860,N_7764);
nor U8374 (N_8374,N_7902,N_7609);
nand U8375 (N_8375,N_7757,N_7740);
nor U8376 (N_8376,N_7604,N_7796);
nor U8377 (N_8377,N_7967,N_7544);
and U8378 (N_8378,N_7567,N_7783);
nor U8379 (N_8379,N_7719,N_7598);
nor U8380 (N_8380,N_7954,N_7935);
or U8381 (N_8381,N_7702,N_7913);
nand U8382 (N_8382,N_7591,N_7564);
nand U8383 (N_8383,N_7935,N_7570);
or U8384 (N_8384,N_7534,N_7615);
nor U8385 (N_8385,N_7560,N_7690);
or U8386 (N_8386,N_7576,N_7545);
and U8387 (N_8387,N_7941,N_7525);
and U8388 (N_8388,N_7658,N_7980);
or U8389 (N_8389,N_7841,N_7740);
nand U8390 (N_8390,N_7868,N_7905);
nor U8391 (N_8391,N_7990,N_7827);
nor U8392 (N_8392,N_7639,N_7885);
nand U8393 (N_8393,N_7895,N_7632);
nor U8394 (N_8394,N_7882,N_7516);
nor U8395 (N_8395,N_7840,N_7731);
and U8396 (N_8396,N_7567,N_7975);
or U8397 (N_8397,N_7817,N_7955);
and U8398 (N_8398,N_7999,N_7614);
nor U8399 (N_8399,N_7563,N_7582);
and U8400 (N_8400,N_7906,N_7514);
xnor U8401 (N_8401,N_7932,N_7759);
nand U8402 (N_8402,N_7586,N_7972);
nand U8403 (N_8403,N_7755,N_7706);
and U8404 (N_8404,N_7559,N_7872);
or U8405 (N_8405,N_7804,N_7525);
nor U8406 (N_8406,N_7594,N_7628);
and U8407 (N_8407,N_7556,N_7749);
nor U8408 (N_8408,N_7520,N_7821);
nor U8409 (N_8409,N_7737,N_7857);
nand U8410 (N_8410,N_7725,N_7736);
and U8411 (N_8411,N_7827,N_7751);
or U8412 (N_8412,N_7633,N_7712);
and U8413 (N_8413,N_7672,N_7709);
nor U8414 (N_8414,N_7585,N_7784);
and U8415 (N_8415,N_7978,N_7552);
nand U8416 (N_8416,N_7699,N_7894);
nor U8417 (N_8417,N_7584,N_7972);
or U8418 (N_8418,N_7711,N_7769);
nor U8419 (N_8419,N_7847,N_7999);
xor U8420 (N_8420,N_7915,N_7664);
nand U8421 (N_8421,N_7861,N_7739);
or U8422 (N_8422,N_7870,N_7527);
nor U8423 (N_8423,N_7810,N_7546);
nand U8424 (N_8424,N_7999,N_7654);
and U8425 (N_8425,N_7651,N_7615);
nand U8426 (N_8426,N_7920,N_7600);
or U8427 (N_8427,N_7717,N_7700);
and U8428 (N_8428,N_7747,N_7674);
or U8429 (N_8429,N_7574,N_7880);
nand U8430 (N_8430,N_7930,N_7911);
and U8431 (N_8431,N_7971,N_7691);
and U8432 (N_8432,N_7543,N_7566);
nor U8433 (N_8433,N_7534,N_7724);
and U8434 (N_8434,N_7602,N_7570);
and U8435 (N_8435,N_7757,N_7743);
and U8436 (N_8436,N_7582,N_7784);
or U8437 (N_8437,N_7966,N_7710);
nand U8438 (N_8438,N_7946,N_7726);
and U8439 (N_8439,N_7645,N_7728);
or U8440 (N_8440,N_7822,N_7955);
nand U8441 (N_8441,N_7520,N_7644);
nand U8442 (N_8442,N_7975,N_7662);
nand U8443 (N_8443,N_7810,N_7746);
or U8444 (N_8444,N_7769,N_7557);
nor U8445 (N_8445,N_7675,N_7849);
xor U8446 (N_8446,N_7737,N_7564);
and U8447 (N_8447,N_7583,N_7512);
or U8448 (N_8448,N_7977,N_7691);
and U8449 (N_8449,N_7572,N_7871);
nand U8450 (N_8450,N_7559,N_7949);
nand U8451 (N_8451,N_7588,N_7548);
or U8452 (N_8452,N_7673,N_7961);
and U8453 (N_8453,N_7650,N_7671);
nor U8454 (N_8454,N_7821,N_7956);
or U8455 (N_8455,N_7533,N_7694);
nor U8456 (N_8456,N_7742,N_7931);
and U8457 (N_8457,N_7579,N_7659);
nand U8458 (N_8458,N_7571,N_7665);
or U8459 (N_8459,N_7536,N_7881);
or U8460 (N_8460,N_7512,N_7849);
nor U8461 (N_8461,N_7922,N_7501);
or U8462 (N_8462,N_7568,N_7870);
nand U8463 (N_8463,N_7622,N_7568);
nand U8464 (N_8464,N_7807,N_7983);
nor U8465 (N_8465,N_7579,N_7523);
nor U8466 (N_8466,N_7589,N_7706);
nor U8467 (N_8467,N_7806,N_7648);
nand U8468 (N_8468,N_7632,N_7822);
nor U8469 (N_8469,N_7775,N_7789);
or U8470 (N_8470,N_7655,N_7938);
and U8471 (N_8471,N_7606,N_7631);
and U8472 (N_8472,N_7532,N_7537);
nor U8473 (N_8473,N_7721,N_7954);
and U8474 (N_8474,N_7582,N_7980);
nor U8475 (N_8475,N_7774,N_7633);
and U8476 (N_8476,N_7799,N_7793);
nand U8477 (N_8477,N_7884,N_7524);
xnor U8478 (N_8478,N_7551,N_7632);
or U8479 (N_8479,N_7766,N_7588);
or U8480 (N_8480,N_7872,N_7538);
nor U8481 (N_8481,N_7765,N_7569);
or U8482 (N_8482,N_7735,N_7924);
and U8483 (N_8483,N_7703,N_7576);
nand U8484 (N_8484,N_7860,N_7879);
and U8485 (N_8485,N_7750,N_7838);
and U8486 (N_8486,N_7994,N_7748);
nor U8487 (N_8487,N_7982,N_7969);
and U8488 (N_8488,N_7725,N_7603);
nor U8489 (N_8489,N_7717,N_7569);
or U8490 (N_8490,N_7534,N_7994);
nor U8491 (N_8491,N_7982,N_7673);
nor U8492 (N_8492,N_7538,N_7589);
and U8493 (N_8493,N_7534,N_7952);
nor U8494 (N_8494,N_7710,N_7524);
nor U8495 (N_8495,N_7679,N_7964);
nor U8496 (N_8496,N_7621,N_7668);
nand U8497 (N_8497,N_7926,N_7869);
xnor U8498 (N_8498,N_7795,N_7828);
and U8499 (N_8499,N_7682,N_7519);
and U8500 (N_8500,N_8356,N_8350);
nor U8501 (N_8501,N_8334,N_8216);
or U8502 (N_8502,N_8025,N_8084);
or U8503 (N_8503,N_8442,N_8094);
or U8504 (N_8504,N_8336,N_8403);
nand U8505 (N_8505,N_8453,N_8152);
or U8506 (N_8506,N_8103,N_8440);
and U8507 (N_8507,N_8110,N_8002);
nor U8508 (N_8508,N_8281,N_8024);
and U8509 (N_8509,N_8470,N_8142);
and U8510 (N_8510,N_8046,N_8223);
nand U8511 (N_8511,N_8112,N_8164);
xor U8512 (N_8512,N_8466,N_8222);
nor U8513 (N_8513,N_8310,N_8132);
xnor U8514 (N_8514,N_8478,N_8118);
nor U8515 (N_8515,N_8316,N_8225);
nand U8516 (N_8516,N_8198,N_8185);
nand U8517 (N_8517,N_8295,N_8059);
or U8518 (N_8518,N_8416,N_8385);
and U8519 (N_8519,N_8378,N_8375);
nand U8520 (N_8520,N_8069,N_8459);
nand U8521 (N_8521,N_8269,N_8499);
and U8522 (N_8522,N_8192,N_8364);
nor U8523 (N_8523,N_8101,N_8017);
nor U8524 (N_8524,N_8394,N_8031);
or U8525 (N_8525,N_8467,N_8100);
and U8526 (N_8526,N_8287,N_8087);
or U8527 (N_8527,N_8245,N_8181);
and U8528 (N_8528,N_8167,N_8159);
nor U8529 (N_8529,N_8048,N_8476);
or U8530 (N_8530,N_8251,N_8109);
or U8531 (N_8531,N_8398,N_8257);
nand U8532 (N_8532,N_8395,N_8073);
and U8533 (N_8533,N_8401,N_8066);
and U8534 (N_8534,N_8033,N_8119);
nor U8535 (N_8535,N_8408,N_8137);
or U8536 (N_8536,N_8209,N_8487);
nor U8537 (N_8537,N_8201,N_8270);
and U8538 (N_8538,N_8340,N_8229);
nor U8539 (N_8539,N_8303,N_8197);
nor U8540 (N_8540,N_8352,N_8188);
and U8541 (N_8541,N_8157,N_8376);
and U8542 (N_8542,N_8099,N_8441);
or U8543 (N_8543,N_8232,N_8362);
or U8544 (N_8544,N_8126,N_8173);
nand U8545 (N_8545,N_8077,N_8381);
nor U8546 (N_8546,N_8194,N_8455);
xnor U8547 (N_8547,N_8256,N_8200);
and U8548 (N_8548,N_8346,N_8241);
or U8549 (N_8549,N_8212,N_8307);
nor U8550 (N_8550,N_8431,N_8484);
and U8551 (N_8551,N_8124,N_8210);
xnor U8552 (N_8552,N_8373,N_8231);
and U8553 (N_8553,N_8050,N_8293);
or U8554 (N_8554,N_8289,N_8178);
or U8555 (N_8555,N_8391,N_8387);
nand U8556 (N_8556,N_8120,N_8389);
nor U8557 (N_8557,N_8088,N_8432);
or U8558 (N_8558,N_8106,N_8266);
or U8559 (N_8559,N_8288,N_8371);
or U8560 (N_8560,N_8186,N_8405);
or U8561 (N_8561,N_8146,N_8353);
or U8562 (N_8562,N_8445,N_8193);
nor U8563 (N_8563,N_8382,N_8436);
and U8564 (N_8564,N_8218,N_8425);
and U8565 (N_8565,N_8187,N_8037);
nor U8566 (N_8566,N_8083,N_8298);
and U8567 (N_8567,N_8238,N_8207);
nand U8568 (N_8568,N_8317,N_8246);
nor U8569 (N_8569,N_8323,N_8093);
or U8570 (N_8570,N_8003,N_8426);
or U8571 (N_8571,N_8052,N_8355);
nand U8572 (N_8572,N_8195,N_8275);
xnor U8573 (N_8573,N_8244,N_8030);
nand U8574 (N_8574,N_8013,N_8019);
nand U8575 (N_8575,N_8020,N_8368);
or U8576 (N_8576,N_8308,N_8253);
nor U8577 (N_8577,N_8023,N_8343);
and U8578 (N_8578,N_8461,N_8473);
nand U8579 (N_8579,N_8324,N_8064);
nor U8580 (N_8580,N_8444,N_8300);
or U8581 (N_8581,N_8189,N_8175);
and U8582 (N_8582,N_8053,N_8452);
nor U8583 (N_8583,N_8070,N_8339);
nand U8584 (N_8584,N_8045,N_8264);
nor U8585 (N_8585,N_8117,N_8361);
and U8586 (N_8586,N_8249,N_8004);
and U8587 (N_8587,N_8057,N_8213);
or U8588 (N_8588,N_8147,N_8498);
nor U8589 (N_8589,N_8479,N_8162);
nand U8590 (N_8590,N_8265,N_8370);
nand U8591 (N_8591,N_8133,N_8468);
and U8592 (N_8592,N_8263,N_8042);
nand U8593 (N_8593,N_8018,N_8301);
nand U8594 (N_8594,N_8434,N_8477);
nand U8595 (N_8595,N_8414,N_8273);
and U8596 (N_8596,N_8016,N_8296);
or U8597 (N_8597,N_8495,N_8486);
nand U8598 (N_8598,N_8297,N_8302);
and U8599 (N_8599,N_8060,N_8366);
nor U8600 (N_8600,N_8451,N_8335);
nand U8601 (N_8601,N_8319,N_8151);
or U8602 (N_8602,N_8490,N_8227);
xor U8603 (N_8603,N_8292,N_8421);
or U8604 (N_8604,N_8135,N_8111);
or U8605 (N_8605,N_8294,N_8404);
nand U8606 (N_8606,N_8127,N_8344);
nor U8607 (N_8607,N_8221,N_8092);
nor U8608 (N_8608,N_8014,N_8333);
xor U8609 (N_8609,N_8482,N_8261);
nand U8610 (N_8610,N_8234,N_8420);
nand U8611 (N_8611,N_8199,N_8305);
or U8612 (N_8612,N_8114,N_8250);
nor U8613 (N_8613,N_8328,N_8131);
nor U8614 (N_8614,N_8446,N_8347);
or U8615 (N_8615,N_8011,N_8454);
and U8616 (N_8616,N_8150,N_8078);
nor U8617 (N_8617,N_8074,N_8423);
and U8618 (N_8618,N_8471,N_8034);
and U8619 (N_8619,N_8215,N_8149);
and U8620 (N_8620,N_8182,N_8260);
and U8621 (N_8621,N_8214,N_8304);
nand U8622 (N_8622,N_8367,N_8429);
nand U8623 (N_8623,N_8415,N_8230);
nor U8624 (N_8624,N_8392,N_8001);
nor U8625 (N_8625,N_8242,N_8326);
nor U8626 (N_8626,N_8176,N_8158);
nand U8627 (N_8627,N_8399,N_8321);
nand U8628 (N_8628,N_8049,N_8035);
or U8629 (N_8629,N_8277,N_8309);
nor U8630 (N_8630,N_8386,N_8240);
or U8631 (N_8631,N_8354,N_8433);
or U8632 (N_8632,N_8130,N_8104);
nor U8633 (N_8633,N_8254,N_8475);
or U8634 (N_8634,N_8397,N_8450);
or U8635 (N_8635,N_8140,N_8105);
nor U8636 (N_8636,N_8255,N_8460);
nand U8637 (N_8637,N_8372,N_8233);
or U8638 (N_8638,N_8123,N_8204);
nand U8639 (N_8639,N_8054,N_8449);
and U8640 (N_8640,N_8276,N_8143);
or U8641 (N_8641,N_8329,N_8079);
and U8642 (N_8642,N_8072,N_8107);
and U8643 (N_8643,N_8125,N_8009);
nand U8644 (N_8644,N_8464,N_8272);
and U8645 (N_8645,N_8091,N_8267);
nor U8646 (N_8646,N_8055,N_8306);
and U8647 (N_8647,N_8437,N_8174);
or U8648 (N_8648,N_8172,N_8396);
or U8649 (N_8649,N_8236,N_8365);
and U8650 (N_8650,N_8315,N_8012);
or U8651 (N_8651,N_8235,N_8492);
and U8652 (N_8652,N_8076,N_8338);
nand U8653 (N_8653,N_8156,N_8122);
nand U8654 (N_8654,N_8312,N_8062);
and U8655 (N_8655,N_8044,N_8283);
nor U8656 (N_8656,N_8342,N_8191);
nor U8657 (N_8657,N_8349,N_8322);
nand U8658 (N_8658,N_8252,N_8015);
nand U8659 (N_8659,N_8005,N_8211);
nor U8660 (N_8660,N_8248,N_8458);
nor U8661 (N_8661,N_8485,N_8051);
nor U8662 (N_8662,N_8121,N_8168);
and U8663 (N_8663,N_8141,N_8331);
nor U8664 (N_8664,N_8280,N_8138);
or U8665 (N_8665,N_8068,N_8374);
or U8666 (N_8666,N_8043,N_8357);
or U8667 (N_8667,N_8029,N_8489);
or U8668 (N_8668,N_8418,N_8438);
nor U8669 (N_8669,N_8026,N_8056);
or U8670 (N_8670,N_8496,N_8379);
nor U8671 (N_8671,N_8180,N_8417);
and U8672 (N_8672,N_8184,N_8285);
and U8673 (N_8673,N_8424,N_8190);
xnor U8674 (N_8674,N_8032,N_8359);
xor U8675 (N_8675,N_8330,N_8228);
or U8676 (N_8676,N_8428,N_8393);
and U8677 (N_8677,N_8239,N_8000);
or U8678 (N_8678,N_8098,N_8465);
and U8679 (N_8679,N_8113,N_8208);
and U8680 (N_8680,N_8063,N_8337);
xor U8681 (N_8681,N_8153,N_8040);
nand U8682 (N_8682,N_8067,N_8047);
and U8683 (N_8683,N_8481,N_8435);
and U8684 (N_8684,N_8413,N_8412);
xor U8685 (N_8685,N_8075,N_8202);
nand U8686 (N_8686,N_8369,N_8430);
and U8687 (N_8687,N_8291,N_8036);
xnor U8688 (N_8688,N_8217,N_8080);
nor U8689 (N_8689,N_8144,N_8129);
nor U8690 (N_8690,N_8170,N_8377);
nand U8691 (N_8691,N_8472,N_8097);
or U8692 (N_8692,N_8116,N_8085);
nand U8693 (N_8693,N_8325,N_8061);
nand U8694 (N_8694,N_8203,N_8447);
nor U8695 (N_8695,N_8341,N_8409);
or U8696 (N_8696,N_8383,N_8493);
or U8697 (N_8697,N_8038,N_8345);
nand U8698 (N_8698,N_8448,N_8071);
and U8699 (N_8699,N_8406,N_8021);
nor U8700 (N_8700,N_8163,N_8271);
and U8701 (N_8701,N_8081,N_8096);
nor U8702 (N_8702,N_8407,N_8226);
nand U8703 (N_8703,N_8388,N_8314);
and U8704 (N_8704,N_8134,N_8411);
nand U8705 (N_8705,N_8320,N_8279);
or U8706 (N_8706,N_8196,N_8443);
and U8707 (N_8707,N_8166,N_8183);
nor U8708 (N_8708,N_8237,N_8205);
or U8709 (N_8709,N_8041,N_8318);
nor U8710 (N_8710,N_8278,N_8311);
nor U8711 (N_8711,N_8384,N_8402);
or U8712 (N_8712,N_8010,N_8474);
nand U8713 (N_8713,N_8427,N_8258);
and U8714 (N_8714,N_8390,N_8058);
and U8715 (N_8715,N_8262,N_8115);
xor U8716 (N_8716,N_8286,N_8259);
nand U8717 (N_8717,N_8220,N_8462);
nand U8718 (N_8718,N_8155,N_8165);
or U8719 (N_8719,N_8177,N_8169);
nand U8720 (N_8720,N_8102,N_8494);
and U8721 (N_8721,N_8219,N_8136);
and U8722 (N_8722,N_8171,N_8419);
nor U8723 (N_8723,N_8360,N_8422);
nor U8724 (N_8724,N_8488,N_8206);
nand U8725 (N_8725,N_8491,N_8410);
nor U8726 (N_8726,N_8327,N_8299);
or U8727 (N_8727,N_8089,N_8154);
nor U8728 (N_8728,N_8348,N_8006);
and U8729 (N_8729,N_8332,N_8351);
nor U8730 (N_8730,N_8247,N_8086);
nand U8731 (N_8731,N_8139,N_8497);
nor U8732 (N_8732,N_8463,N_8457);
or U8733 (N_8733,N_8469,N_8284);
nand U8734 (N_8734,N_8008,N_8082);
xor U8735 (N_8735,N_8380,N_8095);
or U8736 (N_8736,N_8022,N_8313);
or U8737 (N_8737,N_8090,N_8456);
nand U8738 (N_8738,N_8145,N_8480);
nand U8739 (N_8739,N_8108,N_8027);
or U8740 (N_8740,N_8028,N_8358);
xnor U8741 (N_8741,N_8282,N_8148);
and U8742 (N_8742,N_8268,N_8065);
or U8743 (N_8743,N_8363,N_8224);
nor U8744 (N_8744,N_8179,N_8439);
and U8745 (N_8745,N_8400,N_8039);
and U8746 (N_8746,N_8161,N_8483);
and U8747 (N_8747,N_8243,N_8290);
and U8748 (N_8748,N_8007,N_8274);
and U8749 (N_8749,N_8160,N_8128);
and U8750 (N_8750,N_8362,N_8066);
nor U8751 (N_8751,N_8398,N_8076);
or U8752 (N_8752,N_8136,N_8070);
xnor U8753 (N_8753,N_8423,N_8198);
nor U8754 (N_8754,N_8258,N_8186);
or U8755 (N_8755,N_8055,N_8043);
nor U8756 (N_8756,N_8363,N_8378);
and U8757 (N_8757,N_8296,N_8409);
or U8758 (N_8758,N_8211,N_8159);
and U8759 (N_8759,N_8093,N_8225);
nand U8760 (N_8760,N_8076,N_8309);
and U8761 (N_8761,N_8074,N_8453);
nand U8762 (N_8762,N_8070,N_8277);
and U8763 (N_8763,N_8278,N_8138);
nor U8764 (N_8764,N_8215,N_8020);
nand U8765 (N_8765,N_8324,N_8153);
or U8766 (N_8766,N_8052,N_8107);
or U8767 (N_8767,N_8171,N_8100);
and U8768 (N_8768,N_8220,N_8260);
or U8769 (N_8769,N_8126,N_8384);
nor U8770 (N_8770,N_8368,N_8428);
nand U8771 (N_8771,N_8042,N_8344);
or U8772 (N_8772,N_8217,N_8049);
nand U8773 (N_8773,N_8496,N_8334);
nor U8774 (N_8774,N_8416,N_8057);
nor U8775 (N_8775,N_8414,N_8496);
nor U8776 (N_8776,N_8231,N_8236);
nand U8777 (N_8777,N_8258,N_8241);
and U8778 (N_8778,N_8064,N_8119);
nand U8779 (N_8779,N_8016,N_8114);
and U8780 (N_8780,N_8260,N_8315);
or U8781 (N_8781,N_8432,N_8054);
or U8782 (N_8782,N_8233,N_8350);
nor U8783 (N_8783,N_8405,N_8027);
nor U8784 (N_8784,N_8279,N_8218);
and U8785 (N_8785,N_8032,N_8121);
nand U8786 (N_8786,N_8069,N_8300);
or U8787 (N_8787,N_8090,N_8230);
xnor U8788 (N_8788,N_8440,N_8457);
nand U8789 (N_8789,N_8067,N_8450);
or U8790 (N_8790,N_8410,N_8463);
nand U8791 (N_8791,N_8087,N_8257);
and U8792 (N_8792,N_8021,N_8227);
nor U8793 (N_8793,N_8249,N_8244);
nand U8794 (N_8794,N_8125,N_8024);
nor U8795 (N_8795,N_8098,N_8290);
nor U8796 (N_8796,N_8372,N_8049);
nand U8797 (N_8797,N_8153,N_8106);
and U8798 (N_8798,N_8179,N_8057);
nand U8799 (N_8799,N_8121,N_8147);
nor U8800 (N_8800,N_8426,N_8266);
and U8801 (N_8801,N_8222,N_8057);
nand U8802 (N_8802,N_8402,N_8438);
nor U8803 (N_8803,N_8256,N_8323);
or U8804 (N_8804,N_8283,N_8191);
or U8805 (N_8805,N_8347,N_8313);
nand U8806 (N_8806,N_8018,N_8337);
or U8807 (N_8807,N_8007,N_8152);
or U8808 (N_8808,N_8012,N_8232);
nand U8809 (N_8809,N_8212,N_8001);
or U8810 (N_8810,N_8249,N_8116);
or U8811 (N_8811,N_8010,N_8244);
nor U8812 (N_8812,N_8245,N_8427);
or U8813 (N_8813,N_8448,N_8123);
and U8814 (N_8814,N_8457,N_8114);
nor U8815 (N_8815,N_8077,N_8257);
or U8816 (N_8816,N_8182,N_8318);
xor U8817 (N_8817,N_8030,N_8221);
nor U8818 (N_8818,N_8034,N_8433);
nand U8819 (N_8819,N_8167,N_8324);
or U8820 (N_8820,N_8471,N_8387);
nand U8821 (N_8821,N_8437,N_8301);
nor U8822 (N_8822,N_8011,N_8029);
and U8823 (N_8823,N_8226,N_8221);
and U8824 (N_8824,N_8184,N_8104);
nand U8825 (N_8825,N_8287,N_8140);
and U8826 (N_8826,N_8391,N_8120);
nor U8827 (N_8827,N_8076,N_8468);
and U8828 (N_8828,N_8056,N_8111);
and U8829 (N_8829,N_8375,N_8413);
or U8830 (N_8830,N_8173,N_8099);
and U8831 (N_8831,N_8026,N_8420);
or U8832 (N_8832,N_8441,N_8292);
or U8833 (N_8833,N_8254,N_8079);
nor U8834 (N_8834,N_8046,N_8032);
or U8835 (N_8835,N_8116,N_8038);
nand U8836 (N_8836,N_8185,N_8242);
nand U8837 (N_8837,N_8210,N_8102);
or U8838 (N_8838,N_8198,N_8456);
nand U8839 (N_8839,N_8013,N_8467);
and U8840 (N_8840,N_8329,N_8421);
and U8841 (N_8841,N_8213,N_8028);
nand U8842 (N_8842,N_8136,N_8104);
nor U8843 (N_8843,N_8399,N_8132);
or U8844 (N_8844,N_8491,N_8053);
nor U8845 (N_8845,N_8465,N_8059);
nor U8846 (N_8846,N_8299,N_8454);
and U8847 (N_8847,N_8273,N_8095);
and U8848 (N_8848,N_8124,N_8118);
or U8849 (N_8849,N_8080,N_8152);
nand U8850 (N_8850,N_8324,N_8217);
nor U8851 (N_8851,N_8437,N_8015);
nand U8852 (N_8852,N_8178,N_8484);
or U8853 (N_8853,N_8324,N_8433);
nor U8854 (N_8854,N_8236,N_8319);
nor U8855 (N_8855,N_8152,N_8343);
or U8856 (N_8856,N_8141,N_8387);
and U8857 (N_8857,N_8230,N_8082);
and U8858 (N_8858,N_8371,N_8112);
or U8859 (N_8859,N_8470,N_8216);
and U8860 (N_8860,N_8322,N_8012);
or U8861 (N_8861,N_8459,N_8180);
nor U8862 (N_8862,N_8426,N_8230);
and U8863 (N_8863,N_8351,N_8124);
nor U8864 (N_8864,N_8168,N_8359);
nand U8865 (N_8865,N_8207,N_8182);
or U8866 (N_8866,N_8406,N_8128);
or U8867 (N_8867,N_8172,N_8400);
or U8868 (N_8868,N_8019,N_8381);
nor U8869 (N_8869,N_8353,N_8157);
nand U8870 (N_8870,N_8100,N_8226);
nor U8871 (N_8871,N_8142,N_8258);
xor U8872 (N_8872,N_8250,N_8482);
nor U8873 (N_8873,N_8432,N_8329);
xnor U8874 (N_8874,N_8196,N_8175);
xor U8875 (N_8875,N_8127,N_8075);
or U8876 (N_8876,N_8403,N_8158);
and U8877 (N_8877,N_8388,N_8484);
nor U8878 (N_8878,N_8155,N_8237);
nand U8879 (N_8879,N_8188,N_8063);
nor U8880 (N_8880,N_8323,N_8437);
nor U8881 (N_8881,N_8262,N_8436);
and U8882 (N_8882,N_8424,N_8453);
nor U8883 (N_8883,N_8325,N_8031);
and U8884 (N_8884,N_8483,N_8259);
nand U8885 (N_8885,N_8386,N_8196);
or U8886 (N_8886,N_8480,N_8494);
or U8887 (N_8887,N_8171,N_8157);
or U8888 (N_8888,N_8406,N_8414);
xnor U8889 (N_8889,N_8494,N_8269);
xor U8890 (N_8890,N_8246,N_8041);
and U8891 (N_8891,N_8000,N_8012);
and U8892 (N_8892,N_8479,N_8093);
and U8893 (N_8893,N_8260,N_8125);
nand U8894 (N_8894,N_8141,N_8240);
nand U8895 (N_8895,N_8275,N_8303);
and U8896 (N_8896,N_8063,N_8393);
nand U8897 (N_8897,N_8163,N_8377);
xnor U8898 (N_8898,N_8156,N_8084);
nand U8899 (N_8899,N_8225,N_8427);
and U8900 (N_8900,N_8482,N_8105);
nand U8901 (N_8901,N_8401,N_8336);
nand U8902 (N_8902,N_8388,N_8027);
or U8903 (N_8903,N_8167,N_8229);
or U8904 (N_8904,N_8482,N_8030);
nand U8905 (N_8905,N_8117,N_8183);
nand U8906 (N_8906,N_8214,N_8294);
and U8907 (N_8907,N_8427,N_8018);
nor U8908 (N_8908,N_8230,N_8201);
nor U8909 (N_8909,N_8224,N_8046);
nand U8910 (N_8910,N_8215,N_8010);
xnor U8911 (N_8911,N_8475,N_8151);
or U8912 (N_8912,N_8380,N_8075);
nand U8913 (N_8913,N_8257,N_8210);
nor U8914 (N_8914,N_8297,N_8224);
nand U8915 (N_8915,N_8241,N_8483);
or U8916 (N_8916,N_8426,N_8459);
or U8917 (N_8917,N_8158,N_8102);
nor U8918 (N_8918,N_8392,N_8434);
or U8919 (N_8919,N_8422,N_8381);
nand U8920 (N_8920,N_8008,N_8076);
or U8921 (N_8921,N_8008,N_8285);
nor U8922 (N_8922,N_8261,N_8203);
nand U8923 (N_8923,N_8413,N_8449);
and U8924 (N_8924,N_8302,N_8039);
nor U8925 (N_8925,N_8422,N_8456);
or U8926 (N_8926,N_8454,N_8419);
and U8927 (N_8927,N_8459,N_8050);
and U8928 (N_8928,N_8090,N_8020);
nand U8929 (N_8929,N_8296,N_8311);
nor U8930 (N_8930,N_8178,N_8111);
or U8931 (N_8931,N_8184,N_8156);
nand U8932 (N_8932,N_8331,N_8432);
and U8933 (N_8933,N_8242,N_8443);
nand U8934 (N_8934,N_8040,N_8449);
and U8935 (N_8935,N_8480,N_8117);
and U8936 (N_8936,N_8147,N_8140);
or U8937 (N_8937,N_8259,N_8085);
and U8938 (N_8938,N_8122,N_8037);
or U8939 (N_8939,N_8231,N_8397);
xnor U8940 (N_8940,N_8014,N_8267);
xor U8941 (N_8941,N_8062,N_8258);
and U8942 (N_8942,N_8275,N_8320);
and U8943 (N_8943,N_8435,N_8045);
nor U8944 (N_8944,N_8290,N_8491);
nor U8945 (N_8945,N_8478,N_8313);
and U8946 (N_8946,N_8109,N_8466);
and U8947 (N_8947,N_8387,N_8286);
nor U8948 (N_8948,N_8486,N_8196);
nor U8949 (N_8949,N_8034,N_8105);
or U8950 (N_8950,N_8050,N_8123);
nor U8951 (N_8951,N_8363,N_8393);
and U8952 (N_8952,N_8015,N_8034);
or U8953 (N_8953,N_8220,N_8059);
nor U8954 (N_8954,N_8412,N_8235);
or U8955 (N_8955,N_8479,N_8019);
nor U8956 (N_8956,N_8411,N_8289);
nand U8957 (N_8957,N_8381,N_8288);
or U8958 (N_8958,N_8356,N_8263);
or U8959 (N_8959,N_8356,N_8218);
nor U8960 (N_8960,N_8032,N_8444);
nand U8961 (N_8961,N_8023,N_8190);
or U8962 (N_8962,N_8442,N_8179);
nand U8963 (N_8963,N_8336,N_8183);
nand U8964 (N_8964,N_8118,N_8078);
nand U8965 (N_8965,N_8115,N_8020);
or U8966 (N_8966,N_8311,N_8158);
and U8967 (N_8967,N_8216,N_8362);
or U8968 (N_8968,N_8483,N_8067);
nand U8969 (N_8969,N_8168,N_8025);
nor U8970 (N_8970,N_8041,N_8475);
or U8971 (N_8971,N_8165,N_8229);
or U8972 (N_8972,N_8173,N_8466);
or U8973 (N_8973,N_8213,N_8040);
and U8974 (N_8974,N_8375,N_8298);
nor U8975 (N_8975,N_8080,N_8223);
or U8976 (N_8976,N_8042,N_8334);
or U8977 (N_8977,N_8057,N_8313);
nor U8978 (N_8978,N_8408,N_8060);
or U8979 (N_8979,N_8205,N_8375);
nor U8980 (N_8980,N_8436,N_8168);
nor U8981 (N_8981,N_8082,N_8033);
or U8982 (N_8982,N_8190,N_8382);
or U8983 (N_8983,N_8168,N_8407);
and U8984 (N_8984,N_8072,N_8424);
nand U8985 (N_8985,N_8042,N_8046);
and U8986 (N_8986,N_8439,N_8373);
nor U8987 (N_8987,N_8366,N_8037);
nand U8988 (N_8988,N_8251,N_8379);
and U8989 (N_8989,N_8191,N_8079);
and U8990 (N_8990,N_8157,N_8122);
nor U8991 (N_8991,N_8007,N_8097);
nor U8992 (N_8992,N_8102,N_8352);
nor U8993 (N_8993,N_8151,N_8084);
or U8994 (N_8994,N_8003,N_8407);
nor U8995 (N_8995,N_8077,N_8289);
nand U8996 (N_8996,N_8330,N_8123);
and U8997 (N_8997,N_8066,N_8021);
and U8998 (N_8998,N_8226,N_8271);
nand U8999 (N_8999,N_8258,N_8179);
and U9000 (N_9000,N_8945,N_8851);
and U9001 (N_9001,N_8603,N_8991);
nand U9002 (N_9002,N_8859,N_8784);
nand U9003 (N_9003,N_8728,N_8576);
nor U9004 (N_9004,N_8725,N_8843);
and U9005 (N_9005,N_8904,N_8636);
or U9006 (N_9006,N_8755,N_8794);
nor U9007 (N_9007,N_8540,N_8955);
nor U9008 (N_9008,N_8870,N_8522);
and U9009 (N_9009,N_8631,N_8644);
or U9010 (N_9010,N_8674,N_8586);
or U9011 (N_9011,N_8591,N_8681);
nand U9012 (N_9012,N_8960,N_8504);
nor U9013 (N_9013,N_8726,N_8930);
or U9014 (N_9014,N_8561,N_8800);
and U9015 (N_9015,N_8969,N_8617);
nor U9016 (N_9016,N_8640,N_8592);
and U9017 (N_9017,N_8750,N_8787);
nand U9018 (N_9018,N_8700,N_8763);
or U9019 (N_9019,N_8811,N_8925);
or U9020 (N_9020,N_8663,N_8935);
and U9021 (N_9021,N_8970,N_8938);
nor U9022 (N_9022,N_8505,N_8828);
or U9023 (N_9023,N_8780,N_8822);
nand U9024 (N_9024,N_8704,N_8824);
and U9025 (N_9025,N_8807,N_8774);
nor U9026 (N_9026,N_8581,N_8745);
nor U9027 (N_9027,N_8911,N_8873);
or U9028 (N_9028,N_8776,N_8886);
or U9029 (N_9029,N_8585,N_8931);
nand U9030 (N_9030,N_8547,N_8670);
or U9031 (N_9031,N_8952,N_8629);
xnor U9032 (N_9032,N_8769,N_8791);
and U9033 (N_9033,N_8940,N_8778);
nand U9034 (N_9034,N_8786,N_8574);
and U9035 (N_9035,N_8679,N_8537);
and U9036 (N_9036,N_8860,N_8983);
xnor U9037 (N_9037,N_8968,N_8772);
and U9038 (N_9038,N_8577,N_8804);
and U9039 (N_9039,N_8819,N_8775);
or U9040 (N_9040,N_8703,N_8543);
nor U9041 (N_9041,N_8916,N_8521);
or U9042 (N_9042,N_8688,N_8953);
nand U9043 (N_9043,N_8947,N_8805);
nor U9044 (N_9044,N_8874,N_8924);
and U9045 (N_9045,N_8509,N_8734);
nor U9046 (N_9046,N_8920,N_8706);
and U9047 (N_9047,N_8746,N_8835);
or U9048 (N_9048,N_8914,N_8880);
or U9049 (N_9049,N_8587,N_8643);
nand U9050 (N_9050,N_8579,N_8906);
and U9051 (N_9051,N_8927,N_8690);
nor U9052 (N_9052,N_8651,N_8545);
nand U9053 (N_9053,N_8825,N_8714);
nor U9054 (N_9054,N_8936,N_8994);
and U9055 (N_9055,N_8678,N_8753);
or U9056 (N_9056,N_8502,N_8623);
or U9057 (N_9057,N_8608,N_8512);
or U9058 (N_9058,N_8826,N_8619);
nand U9059 (N_9059,N_8610,N_8546);
or U9060 (N_9060,N_8913,N_8907);
nor U9061 (N_9061,N_8864,N_8900);
nor U9062 (N_9062,N_8564,N_8721);
xnor U9063 (N_9063,N_8736,N_8558);
and U9064 (N_9064,N_8588,N_8757);
or U9065 (N_9065,N_8515,N_8532);
and U9066 (N_9066,N_8611,N_8812);
or U9067 (N_9067,N_8854,N_8666);
nand U9068 (N_9068,N_8883,N_8777);
or U9069 (N_9069,N_8555,N_8878);
nor U9070 (N_9070,N_8998,N_8985);
nor U9071 (N_9071,N_8871,N_8575);
and U9072 (N_9072,N_8553,N_8858);
or U9073 (N_9073,N_8554,N_8877);
or U9074 (N_9074,N_8751,N_8869);
nand U9075 (N_9075,N_8524,N_8604);
and U9076 (N_9076,N_8642,N_8535);
nand U9077 (N_9077,N_8709,N_8648);
or U9078 (N_9078,N_8992,N_8536);
or U9079 (N_9079,N_8672,N_8715);
nor U9080 (N_9080,N_8823,N_8645);
nand U9081 (N_9081,N_8990,N_8798);
nand U9082 (N_9082,N_8731,N_8989);
or U9083 (N_9083,N_8818,N_8961);
nor U9084 (N_9084,N_8519,N_8712);
or U9085 (N_9085,N_8950,N_8887);
nand U9086 (N_9086,N_8565,N_8977);
nor U9087 (N_9087,N_8956,N_8973);
nor U9088 (N_9088,N_8821,N_8905);
nor U9089 (N_9089,N_8866,N_8694);
nand U9090 (N_9090,N_8695,N_8979);
nor U9091 (N_9091,N_8687,N_8910);
nor U9092 (N_9092,N_8659,N_8626);
nor U9093 (N_9093,N_8785,N_8958);
nand U9094 (N_9094,N_8607,N_8813);
nand U9095 (N_9095,N_8538,N_8976);
xnor U9096 (N_9096,N_8669,N_8738);
nor U9097 (N_9097,N_8705,N_8868);
or U9098 (N_9098,N_8901,N_8997);
or U9099 (N_9099,N_8594,N_8937);
nand U9100 (N_9100,N_8526,N_8595);
nor U9101 (N_9101,N_8556,N_8981);
or U9102 (N_9102,N_8891,N_8966);
nor U9103 (N_9103,N_8572,N_8987);
nor U9104 (N_9104,N_8514,N_8507);
nor U9105 (N_9105,N_8779,N_8896);
nor U9106 (N_9106,N_8550,N_8657);
and U9107 (N_9107,N_8609,N_8820);
xor U9108 (N_9108,N_8732,N_8530);
nor U9109 (N_9109,N_8963,N_8692);
nand U9110 (N_9110,N_8582,N_8801);
and U9111 (N_9111,N_8542,N_8809);
nor U9112 (N_9112,N_8735,N_8838);
and U9113 (N_9113,N_8962,N_8501);
and U9114 (N_9114,N_8840,N_8766);
or U9115 (N_9115,N_8844,N_8718);
and U9116 (N_9116,N_8861,N_8600);
xor U9117 (N_9117,N_8918,N_8999);
or U9118 (N_9118,N_8523,N_8827);
nor U9119 (N_9119,N_8944,N_8872);
or U9120 (N_9120,N_8803,N_8957);
and U9121 (N_9121,N_8783,N_8656);
nand U9122 (N_9122,N_8889,N_8684);
nand U9123 (N_9123,N_8764,N_8909);
nand U9124 (N_9124,N_8544,N_8899);
or U9125 (N_9125,N_8597,N_8921);
or U9126 (N_9126,N_8857,N_8830);
or U9127 (N_9127,N_8885,N_8510);
nor U9128 (N_9128,N_8618,N_8503);
or U9129 (N_9129,N_8759,N_8567);
and U9130 (N_9130,N_8964,N_8863);
and U9131 (N_9131,N_8730,N_8749);
and U9132 (N_9132,N_8702,N_8641);
nand U9133 (N_9133,N_8653,N_8634);
nand U9134 (N_9134,N_8762,N_8954);
or U9135 (N_9135,N_8673,N_8848);
nor U9136 (N_9136,N_8949,N_8984);
nor U9137 (N_9137,N_8768,N_8747);
or U9138 (N_9138,N_8792,N_8517);
nand U9139 (N_9139,N_8833,N_8894);
nor U9140 (N_9140,N_8928,N_8948);
or U9141 (N_9141,N_8884,N_8566);
and U9142 (N_9142,N_8606,N_8799);
and U9143 (N_9143,N_8852,N_8511);
nand U9144 (N_9144,N_8520,N_8590);
and U9145 (N_9145,N_8630,N_8685);
nand U9146 (N_9146,N_8570,N_8668);
or U9147 (N_9147,N_8754,N_8902);
or U9148 (N_9148,N_8919,N_8500);
and U9149 (N_9149,N_8855,N_8845);
and U9150 (N_9150,N_8797,N_8717);
nand U9151 (N_9151,N_8978,N_8516);
or U9152 (N_9152,N_8563,N_8710);
nand U9153 (N_9153,N_8518,N_8729);
and U9154 (N_9154,N_8806,N_8525);
nand U9155 (N_9155,N_8951,N_8995);
or U9156 (N_9156,N_8727,N_8881);
and U9157 (N_9157,N_8737,N_8980);
and U9158 (N_9158,N_8676,N_8917);
or U9159 (N_9159,N_8601,N_8767);
nor U9160 (N_9160,N_8667,N_8761);
and U9161 (N_9161,N_8665,N_8599);
nand U9162 (N_9162,N_8568,N_8584);
nor U9163 (N_9163,N_8614,N_8817);
and U9164 (N_9164,N_8639,N_8625);
nand U9165 (N_9165,N_8982,N_8627);
or U9166 (N_9166,N_8815,N_8770);
nor U9167 (N_9167,N_8596,N_8789);
and U9168 (N_9168,N_8739,N_8865);
xor U9169 (N_9169,N_8646,N_8557);
or U9170 (N_9170,N_8686,N_8895);
or U9171 (N_9171,N_8708,N_8740);
nand U9172 (N_9172,N_8898,N_8699);
nor U9173 (N_9173,N_8650,N_8612);
or U9174 (N_9174,N_8660,N_8971);
nor U9175 (N_9175,N_8652,N_8580);
nand U9176 (N_9176,N_8808,N_8689);
or U9177 (N_9177,N_8897,N_8834);
nor U9178 (N_9178,N_8814,N_8862);
and U9179 (N_9179,N_8633,N_8593);
or U9180 (N_9180,N_8573,N_8842);
nor U9181 (N_9181,N_8701,N_8635);
and U9182 (N_9182,N_8893,N_8661);
and U9183 (N_9183,N_8693,N_8733);
or U9184 (N_9184,N_8831,N_8765);
nor U9185 (N_9185,N_8959,N_8856);
or U9186 (N_9186,N_8677,N_8771);
nand U9187 (N_9187,N_8758,N_8988);
nand U9188 (N_9188,N_8836,N_8796);
or U9189 (N_9189,N_8975,N_8781);
nand U9190 (N_9190,N_8680,N_8993);
or U9191 (N_9191,N_8867,N_8846);
and U9192 (N_9192,N_8624,N_8720);
nand U9193 (N_9193,N_8598,N_8841);
nand U9194 (N_9194,N_8926,N_8662);
nor U9195 (N_9195,N_8915,N_8589);
nand U9196 (N_9196,N_8748,N_8691);
xnor U9197 (N_9197,N_8923,N_8847);
nor U9198 (N_9198,N_8571,N_8903);
nor U9199 (N_9199,N_8551,N_8912);
nand U9200 (N_9200,N_8892,N_8756);
and U9201 (N_9201,N_8647,N_8802);
nor U9202 (N_9202,N_8527,N_8698);
or U9203 (N_9203,N_8882,N_8637);
nor U9204 (N_9204,N_8943,N_8743);
and U9205 (N_9205,N_8853,N_8569);
nor U9206 (N_9206,N_8996,N_8810);
or U9207 (N_9207,N_8932,N_8888);
nand U9208 (N_9208,N_8790,N_8533);
nand U9209 (N_9209,N_8529,N_8837);
or U9210 (N_9210,N_8760,N_8559);
nor U9211 (N_9211,N_8506,N_8539);
and U9212 (N_9212,N_8513,N_8583);
nor U9213 (N_9213,N_8658,N_8632);
nor U9214 (N_9214,N_8628,N_8741);
or U9215 (N_9215,N_8528,N_8934);
nor U9216 (N_9216,N_8605,N_8615);
and U9217 (N_9217,N_8638,N_8816);
and U9218 (N_9218,N_8649,N_8908);
nand U9219 (N_9219,N_8829,N_8752);
or U9220 (N_9220,N_8922,N_8620);
nor U9221 (N_9221,N_8716,N_8675);
and U9222 (N_9222,N_8773,N_8664);
or U9223 (N_9223,N_8541,N_8724);
nor U9224 (N_9224,N_8719,N_8967);
or U9225 (N_9225,N_8683,N_8879);
nand U9226 (N_9226,N_8946,N_8578);
nor U9227 (N_9227,N_8613,N_8793);
and U9228 (N_9228,N_8876,N_8744);
nor U9229 (N_9229,N_8549,N_8616);
or U9230 (N_9230,N_8548,N_8711);
nor U9231 (N_9231,N_8713,N_8875);
nand U9232 (N_9232,N_8508,N_8602);
nand U9233 (N_9233,N_8534,N_8742);
and U9234 (N_9234,N_8890,N_8965);
and U9235 (N_9235,N_8696,N_8655);
or U9236 (N_9236,N_8531,N_8562);
nand U9237 (N_9237,N_8941,N_8654);
or U9238 (N_9238,N_8795,N_8560);
nor U9239 (N_9239,N_8682,N_8707);
nor U9240 (N_9240,N_8986,N_8722);
nor U9241 (N_9241,N_8839,N_8622);
nor U9242 (N_9242,N_8939,N_8849);
or U9243 (N_9243,N_8929,N_8621);
or U9244 (N_9244,N_8972,N_8782);
and U9245 (N_9245,N_8697,N_8671);
or U9246 (N_9246,N_8552,N_8974);
and U9247 (N_9247,N_8942,N_8723);
xor U9248 (N_9248,N_8788,N_8850);
nand U9249 (N_9249,N_8832,N_8933);
or U9250 (N_9250,N_8960,N_8907);
and U9251 (N_9251,N_8645,N_8607);
and U9252 (N_9252,N_8917,N_8914);
nand U9253 (N_9253,N_8689,N_8868);
nor U9254 (N_9254,N_8660,N_8601);
nor U9255 (N_9255,N_8877,N_8544);
nand U9256 (N_9256,N_8747,N_8602);
nand U9257 (N_9257,N_8875,N_8785);
nor U9258 (N_9258,N_8530,N_8507);
nor U9259 (N_9259,N_8695,N_8633);
nor U9260 (N_9260,N_8563,N_8692);
xnor U9261 (N_9261,N_8581,N_8645);
and U9262 (N_9262,N_8972,N_8643);
xor U9263 (N_9263,N_8663,N_8553);
nor U9264 (N_9264,N_8921,N_8685);
and U9265 (N_9265,N_8759,N_8717);
and U9266 (N_9266,N_8566,N_8694);
nor U9267 (N_9267,N_8761,N_8830);
or U9268 (N_9268,N_8525,N_8715);
or U9269 (N_9269,N_8872,N_8798);
or U9270 (N_9270,N_8910,N_8660);
or U9271 (N_9271,N_8942,N_8608);
or U9272 (N_9272,N_8609,N_8607);
and U9273 (N_9273,N_8923,N_8764);
or U9274 (N_9274,N_8541,N_8925);
and U9275 (N_9275,N_8538,N_8744);
xnor U9276 (N_9276,N_8924,N_8529);
and U9277 (N_9277,N_8954,N_8553);
and U9278 (N_9278,N_8719,N_8860);
or U9279 (N_9279,N_8544,N_8979);
nor U9280 (N_9280,N_8803,N_8950);
or U9281 (N_9281,N_8869,N_8976);
nor U9282 (N_9282,N_8660,N_8906);
nor U9283 (N_9283,N_8786,N_8595);
nand U9284 (N_9284,N_8511,N_8948);
or U9285 (N_9285,N_8957,N_8635);
nand U9286 (N_9286,N_8880,N_8655);
nor U9287 (N_9287,N_8737,N_8550);
and U9288 (N_9288,N_8656,N_8565);
nand U9289 (N_9289,N_8846,N_8914);
nor U9290 (N_9290,N_8514,N_8937);
or U9291 (N_9291,N_8915,N_8797);
or U9292 (N_9292,N_8948,N_8823);
nand U9293 (N_9293,N_8818,N_8604);
or U9294 (N_9294,N_8520,N_8513);
and U9295 (N_9295,N_8911,N_8845);
and U9296 (N_9296,N_8757,N_8566);
or U9297 (N_9297,N_8907,N_8956);
or U9298 (N_9298,N_8854,N_8684);
nor U9299 (N_9299,N_8618,N_8777);
xor U9300 (N_9300,N_8598,N_8752);
nor U9301 (N_9301,N_8610,N_8690);
and U9302 (N_9302,N_8904,N_8941);
or U9303 (N_9303,N_8525,N_8539);
nand U9304 (N_9304,N_8640,N_8655);
xor U9305 (N_9305,N_8769,N_8944);
nor U9306 (N_9306,N_8990,N_8788);
or U9307 (N_9307,N_8885,N_8749);
or U9308 (N_9308,N_8888,N_8662);
and U9309 (N_9309,N_8825,N_8804);
nor U9310 (N_9310,N_8564,N_8894);
or U9311 (N_9311,N_8838,N_8679);
nand U9312 (N_9312,N_8782,N_8921);
and U9313 (N_9313,N_8946,N_8900);
nor U9314 (N_9314,N_8949,N_8580);
nand U9315 (N_9315,N_8885,N_8609);
or U9316 (N_9316,N_8551,N_8638);
nor U9317 (N_9317,N_8642,N_8523);
or U9318 (N_9318,N_8663,N_8898);
xor U9319 (N_9319,N_8588,N_8929);
or U9320 (N_9320,N_8795,N_8570);
or U9321 (N_9321,N_8777,N_8539);
nor U9322 (N_9322,N_8752,N_8677);
nand U9323 (N_9323,N_8690,N_8721);
and U9324 (N_9324,N_8659,N_8990);
and U9325 (N_9325,N_8987,N_8997);
or U9326 (N_9326,N_8689,N_8845);
nor U9327 (N_9327,N_8508,N_8708);
nor U9328 (N_9328,N_8839,N_8851);
or U9329 (N_9329,N_8623,N_8711);
or U9330 (N_9330,N_8554,N_8917);
and U9331 (N_9331,N_8599,N_8928);
nor U9332 (N_9332,N_8780,N_8655);
and U9333 (N_9333,N_8812,N_8647);
nor U9334 (N_9334,N_8937,N_8949);
nand U9335 (N_9335,N_8792,N_8689);
nand U9336 (N_9336,N_8614,N_8505);
nor U9337 (N_9337,N_8675,N_8610);
and U9338 (N_9338,N_8648,N_8953);
xnor U9339 (N_9339,N_8918,N_8506);
nor U9340 (N_9340,N_8517,N_8570);
nor U9341 (N_9341,N_8548,N_8648);
nand U9342 (N_9342,N_8721,N_8604);
xnor U9343 (N_9343,N_8809,N_8807);
or U9344 (N_9344,N_8570,N_8854);
nor U9345 (N_9345,N_8886,N_8950);
and U9346 (N_9346,N_8752,N_8777);
and U9347 (N_9347,N_8880,N_8572);
or U9348 (N_9348,N_8761,N_8629);
nor U9349 (N_9349,N_8661,N_8837);
nor U9350 (N_9350,N_8927,N_8602);
or U9351 (N_9351,N_8588,N_8516);
nor U9352 (N_9352,N_8754,N_8511);
and U9353 (N_9353,N_8993,N_8544);
and U9354 (N_9354,N_8531,N_8876);
nand U9355 (N_9355,N_8671,N_8863);
or U9356 (N_9356,N_8823,N_8628);
and U9357 (N_9357,N_8785,N_8796);
nor U9358 (N_9358,N_8835,N_8611);
or U9359 (N_9359,N_8636,N_8848);
nand U9360 (N_9360,N_8626,N_8796);
or U9361 (N_9361,N_8582,N_8788);
nor U9362 (N_9362,N_8812,N_8631);
or U9363 (N_9363,N_8836,N_8788);
xnor U9364 (N_9364,N_8781,N_8934);
or U9365 (N_9365,N_8511,N_8848);
or U9366 (N_9366,N_8588,N_8699);
and U9367 (N_9367,N_8657,N_8690);
and U9368 (N_9368,N_8739,N_8759);
nor U9369 (N_9369,N_8843,N_8572);
nand U9370 (N_9370,N_8728,N_8582);
or U9371 (N_9371,N_8870,N_8540);
nand U9372 (N_9372,N_8806,N_8642);
and U9373 (N_9373,N_8923,N_8623);
or U9374 (N_9374,N_8967,N_8873);
and U9375 (N_9375,N_8861,N_8561);
nor U9376 (N_9376,N_8882,N_8604);
nor U9377 (N_9377,N_8641,N_8850);
nor U9378 (N_9378,N_8831,N_8758);
nor U9379 (N_9379,N_8570,N_8552);
nor U9380 (N_9380,N_8963,N_8921);
nand U9381 (N_9381,N_8671,N_8865);
or U9382 (N_9382,N_8832,N_8798);
nor U9383 (N_9383,N_8626,N_8886);
nor U9384 (N_9384,N_8575,N_8965);
or U9385 (N_9385,N_8601,N_8874);
nand U9386 (N_9386,N_8561,N_8633);
and U9387 (N_9387,N_8575,N_8989);
nand U9388 (N_9388,N_8827,N_8994);
or U9389 (N_9389,N_8513,N_8601);
and U9390 (N_9390,N_8593,N_8695);
and U9391 (N_9391,N_8612,N_8867);
nor U9392 (N_9392,N_8565,N_8723);
xnor U9393 (N_9393,N_8727,N_8570);
nand U9394 (N_9394,N_8660,N_8934);
nand U9395 (N_9395,N_8637,N_8869);
nand U9396 (N_9396,N_8747,N_8785);
and U9397 (N_9397,N_8789,N_8979);
and U9398 (N_9398,N_8874,N_8751);
or U9399 (N_9399,N_8617,N_8865);
and U9400 (N_9400,N_8908,N_8971);
nor U9401 (N_9401,N_8722,N_8736);
nor U9402 (N_9402,N_8874,N_8861);
or U9403 (N_9403,N_8532,N_8907);
nand U9404 (N_9404,N_8810,N_8823);
and U9405 (N_9405,N_8805,N_8686);
and U9406 (N_9406,N_8994,N_8675);
nand U9407 (N_9407,N_8921,N_8879);
or U9408 (N_9408,N_8637,N_8871);
or U9409 (N_9409,N_8702,N_8535);
and U9410 (N_9410,N_8991,N_8590);
nor U9411 (N_9411,N_8613,N_8741);
nor U9412 (N_9412,N_8580,N_8827);
xor U9413 (N_9413,N_8879,N_8933);
nand U9414 (N_9414,N_8968,N_8583);
nor U9415 (N_9415,N_8755,N_8608);
xnor U9416 (N_9416,N_8673,N_8744);
and U9417 (N_9417,N_8594,N_8639);
xnor U9418 (N_9418,N_8871,N_8728);
nor U9419 (N_9419,N_8600,N_8844);
or U9420 (N_9420,N_8905,N_8912);
nand U9421 (N_9421,N_8641,N_8839);
nor U9422 (N_9422,N_8899,N_8916);
or U9423 (N_9423,N_8650,N_8510);
nor U9424 (N_9424,N_8643,N_8515);
and U9425 (N_9425,N_8707,N_8830);
or U9426 (N_9426,N_8701,N_8996);
or U9427 (N_9427,N_8523,N_8992);
or U9428 (N_9428,N_8929,N_8805);
nor U9429 (N_9429,N_8642,N_8983);
nand U9430 (N_9430,N_8917,N_8559);
nor U9431 (N_9431,N_8535,N_8579);
and U9432 (N_9432,N_8798,N_8543);
nand U9433 (N_9433,N_8665,N_8524);
xor U9434 (N_9434,N_8904,N_8773);
and U9435 (N_9435,N_8931,N_8945);
and U9436 (N_9436,N_8801,N_8664);
nand U9437 (N_9437,N_8697,N_8717);
nor U9438 (N_9438,N_8979,N_8905);
nor U9439 (N_9439,N_8902,N_8776);
xnor U9440 (N_9440,N_8537,N_8682);
nor U9441 (N_9441,N_8810,N_8891);
or U9442 (N_9442,N_8669,N_8613);
and U9443 (N_9443,N_8998,N_8911);
nand U9444 (N_9444,N_8622,N_8659);
and U9445 (N_9445,N_8584,N_8829);
and U9446 (N_9446,N_8864,N_8685);
and U9447 (N_9447,N_8760,N_8932);
or U9448 (N_9448,N_8601,N_8894);
or U9449 (N_9449,N_8716,N_8620);
and U9450 (N_9450,N_8938,N_8989);
and U9451 (N_9451,N_8830,N_8848);
nand U9452 (N_9452,N_8529,N_8967);
nand U9453 (N_9453,N_8754,N_8708);
nor U9454 (N_9454,N_8657,N_8796);
or U9455 (N_9455,N_8589,N_8803);
nand U9456 (N_9456,N_8789,N_8838);
nand U9457 (N_9457,N_8882,N_8731);
and U9458 (N_9458,N_8541,N_8972);
and U9459 (N_9459,N_8661,N_8529);
and U9460 (N_9460,N_8576,N_8952);
or U9461 (N_9461,N_8795,N_8661);
and U9462 (N_9462,N_8828,N_8830);
nand U9463 (N_9463,N_8964,N_8665);
or U9464 (N_9464,N_8727,N_8718);
nand U9465 (N_9465,N_8686,N_8919);
or U9466 (N_9466,N_8597,N_8653);
nand U9467 (N_9467,N_8563,N_8967);
nand U9468 (N_9468,N_8505,N_8837);
nand U9469 (N_9469,N_8517,N_8637);
nor U9470 (N_9470,N_8873,N_8826);
or U9471 (N_9471,N_8929,N_8589);
nand U9472 (N_9472,N_8886,N_8599);
nor U9473 (N_9473,N_8799,N_8970);
and U9474 (N_9474,N_8720,N_8887);
nor U9475 (N_9475,N_8737,N_8680);
nor U9476 (N_9476,N_8994,N_8579);
and U9477 (N_9477,N_8553,N_8926);
nor U9478 (N_9478,N_8687,N_8901);
nor U9479 (N_9479,N_8718,N_8679);
nand U9480 (N_9480,N_8773,N_8970);
nand U9481 (N_9481,N_8677,N_8687);
nand U9482 (N_9482,N_8676,N_8963);
or U9483 (N_9483,N_8881,N_8731);
or U9484 (N_9484,N_8966,N_8515);
nor U9485 (N_9485,N_8637,N_8898);
nand U9486 (N_9486,N_8734,N_8883);
nor U9487 (N_9487,N_8736,N_8929);
nor U9488 (N_9488,N_8962,N_8780);
nand U9489 (N_9489,N_8629,N_8968);
and U9490 (N_9490,N_8560,N_8826);
and U9491 (N_9491,N_8903,N_8950);
or U9492 (N_9492,N_8703,N_8771);
nor U9493 (N_9493,N_8825,N_8865);
nor U9494 (N_9494,N_8671,N_8837);
nor U9495 (N_9495,N_8821,N_8621);
and U9496 (N_9496,N_8919,N_8955);
and U9497 (N_9497,N_8814,N_8891);
nand U9498 (N_9498,N_8942,N_8929);
and U9499 (N_9499,N_8500,N_8641);
or U9500 (N_9500,N_9428,N_9367);
or U9501 (N_9501,N_9199,N_9131);
or U9502 (N_9502,N_9204,N_9089);
and U9503 (N_9503,N_9295,N_9290);
and U9504 (N_9504,N_9383,N_9285);
nor U9505 (N_9505,N_9117,N_9123);
or U9506 (N_9506,N_9375,N_9087);
or U9507 (N_9507,N_9387,N_9161);
and U9508 (N_9508,N_9398,N_9318);
nor U9509 (N_9509,N_9358,N_9075);
and U9510 (N_9510,N_9036,N_9132);
and U9511 (N_9511,N_9254,N_9452);
nor U9512 (N_9512,N_9491,N_9060);
and U9513 (N_9513,N_9122,N_9044);
nand U9514 (N_9514,N_9463,N_9342);
nor U9515 (N_9515,N_9340,N_9183);
nand U9516 (N_9516,N_9413,N_9421);
or U9517 (N_9517,N_9308,N_9113);
or U9518 (N_9518,N_9346,N_9135);
and U9519 (N_9519,N_9269,N_9162);
or U9520 (N_9520,N_9159,N_9454);
and U9521 (N_9521,N_9414,N_9102);
or U9522 (N_9522,N_9443,N_9478);
and U9523 (N_9523,N_9418,N_9294);
and U9524 (N_9524,N_9012,N_9480);
nand U9525 (N_9525,N_9195,N_9144);
or U9526 (N_9526,N_9000,N_9083);
nand U9527 (N_9527,N_9069,N_9292);
nor U9528 (N_9528,N_9265,N_9333);
and U9529 (N_9529,N_9149,N_9481);
or U9530 (N_9530,N_9499,N_9279);
nor U9531 (N_9531,N_9050,N_9289);
or U9532 (N_9532,N_9167,N_9234);
nor U9533 (N_9533,N_9406,N_9474);
nand U9534 (N_9534,N_9098,N_9311);
nand U9535 (N_9535,N_9194,N_9011);
nor U9536 (N_9536,N_9412,N_9403);
nand U9537 (N_9537,N_9091,N_9457);
xor U9538 (N_9538,N_9205,N_9051);
and U9539 (N_9539,N_9399,N_9324);
nand U9540 (N_9540,N_9298,N_9227);
nor U9541 (N_9541,N_9465,N_9444);
nor U9542 (N_9542,N_9001,N_9497);
nor U9543 (N_9543,N_9389,N_9170);
or U9544 (N_9544,N_9219,N_9355);
or U9545 (N_9545,N_9467,N_9202);
nor U9546 (N_9546,N_9006,N_9140);
and U9547 (N_9547,N_9109,N_9025);
and U9548 (N_9548,N_9392,N_9074);
or U9549 (N_9549,N_9068,N_9238);
nor U9550 (N_9550,N_9479,N_9411);
and U9551 (N_9551,N_9276,N_9158);
or U9552 (N_9552,N_9339,N_9314);
nor U9553 (N_9553,N_9095,N_9024);
or U9554 (N_9554,N_9013,N_9459);
nor U9555 (N_9555,N_9281,N_9280);
or U9556 (N_9556,N_9005,N_9246);
or U9557 (N_9557,N_9105,N_9248);
or U9558 (N_9558,N_9448,N_9084);
or U9559 (N_9559,N_9156,N_9350);
nand U9560 (N_9560,N_9488,N_9129);
or U9561 (N_9561,N_9142,N_9472);
and U9562 (N_9562,N_9049,N_9407);
or U9563 (N_9563,N_9125,N_9464);
and U9564 (N_9564,N_9435,N_9243);
nand U9565 (N_9565,N_9192,N_9316);
nand U9566 (N_9566,N_9237,N_9450);
and U9567 (N_9567,N_9460,N_9483);
nor U9568 (N_9568,N_9033,N_9317);
and U9569 (N_9569,N_9458,N_9208);
or U9570 (N_9570,N_9286,N_9059);
nor U9571 (N_9571,N_9228,N_9048);
nand U9572 (N_9572,N_9273,N_9240);
xor U9573 (N_9573,N_9203,N_9076);
or U9574 (N_9574,N_9482,N_9309);
or U9575 (N_9575,N_9128,N_9388);
xnor U9576 (N_9576,N_9189,N_9152);
or U9577 (N_9577,N_9410,N_9141);
or U9578 (N_9578,N_9155,N_9232);
and U9579 (N_9579,N_9364,N_9072);
nor U9580 (N_9580,N_9390,N_9267);
nand U9581 (N_9581,N_9046,N_9114);
or U9582 (N_9582,N_9035,N_9283);
nor U9583 (N_9583,N_9221,N_9090);
nor U9584 (N_9584,N_9485,N_9224);
or U9585 (N_9585,N_9016,N_9165);
nand U9586 (N_9586,N_9430,N_9334);
nand U9587 (N_9587,N_9453,N_9190);
or U9588 (N_9588,N_9034,N_9198);
nor U9589 (N_9589,N_9368,N_9081);
or U9590 (N_9590,N_9395,N_9101);
nor U9591 (N_9591,N_9301,N_9381);
nand U9592 (N_9592,N_9391,N_9096);
nor U9593 (N_9593,N_9266,N_9326);
or U9594 (N_9594,N_9030,N_9052);
nor U9595 (N_9595,N_9337,N_9042);
nand U9596 (N_9596,N_9146,N_9218);
nor U9597 (N_9597,N_9233,N_9402);
nor U9598 (N_9598,N_9422,N_9196);
nand U9599 (N_9599,N_9160,N_9213);
and U9600 (N_9600,N_9370,N_9211);
or U9601 (N_9601,N_9121,N_9477);
or U9602 (N_9602,N_9262,N_9099);
nand U9603 (N_9603,N_9201,N_9085);
nand U9604 (N_9604,N_9111,N_9078);
or U9605 (N_9605,N_9116,N_9047);
nand U9606 (N_9606,N_9376,N_9029);
or U9607 (N_9607,N_9304,N_9476);
or U9608 (N_9608,N_9360,N_9139);
or U9609 (N_9609,N_9222,N_9447);
nor U9610 (N_9610,N_9057,N_9297);
nor U9611 (N_9611,N_9186,N_9063);
nor U9612 (N_9612,N_9118,N_9372);
nand U9613 (N_9613,N_9495,N_9425);
nand U9614 (N_9614,N_9181,N_9185);
and U9615 (N_9615,N_9349,N_9451);
nand U9616 (N_9616,N_9404,N_9150);
and U9617 (N_9617,N_9020,N_9242);
and U9618 (N_9618,N_9385,N_9409);
nand U9619 (N_9619,N_9007,N_9126);
xnor U9620 (N_9620,N_9200,N_9369);
and U9621 (N_9621,N_9217,N_9168);
and U9622 (N_9622,N_9303,N_9380);
and U9623 (N_9623,N_9462,N_9055);
nand U9624 (N_9624,N_9359,N_9426);
nor U9625 (N_9625,N_9470,N_9362);
nor U9626 (N_9626,N_9032,N_9147);
and U9627 (N_9627,N_9115,N_9230);
and U9628 (N_9628,N_9361,N_9241);
nand U9629 (N_9629,N_9256,N_9154);
and U9630 (N_9630,N_9252,N_9037);
and U9631 (N_9631,N_9107,N_9377);
or U9632 (N_9632,N_9302,N_9438);
nand U9633 (N_9633,N_9093,N_9344);
and U9634 (N_9634,N_9420,N_9176);
nor U9635 (N_9635,N_9193,N_9282);
and U9636 (N_9636,N_9374,N_9382);
or U9637 (N_9637,N_9226,N_9145);
or U9638 (N_9638,N_9363,N_9475);
nand U9639 (N_9639,N_9010,N_9215);
nand U9640 (N_9640,N_9274,N_9394);
nor U9641 (N_9641,N_9306,N_9133);
nor U9642 (N_9642,N_9332,N_9264);
or U9643 (N_9643,N_9124,N_9424);
nor U9644 (N_9644,N_9088,N_9053);
and U9645 (N_9645,N_9319,N_9251);
nand U9646 (N_9646,N_9436,N_9094);
and U9647 (N_9647,N_9287,N_9003);
or U9648 (N_9648,N_9261,N_9174);
nand U9649 (N_9649,N_9148,N_9489);
nand U9650 (N_9650,N_9079,N_9338);
nand U9651 (N_9651,N_9157,N_9207);
nor U9652 (N_9652,N_9209,N_9429);
nor U9653 (N_9653,N_9027,N_9106);
or U9654 (N_9654,N_9250,N_9330);
or U9655 (N_9655,N_9313,N_9347);
nor U9656 (N_9656,N_9405,N_9427);
and U9657 (N_9657,N_9056,N_9073);
nor U9658 (N_9658,N_9416,N_9239);
nor U9659 (N_9659,N_9197,N_9379);
and U9660 (N_9660,N_9112,N_9041);
nor U9661 (N_9661,N_9366,N_9268);
xnor U9662 (N_9662,N_9004,N_9080);
nor U9663 (N_9663,N_9278,N_9293);
or U9664 (N_9664,N_9373,N_9164);
nand U9665 (N_9665,N_9229,N_9247);
or U9666 (N_9666,N_9082,N_9271);
nor U9667 (N_9667,N_9067,N_9323);
nand U9668 (N_9668,N_9259,N_9014);
or U9669 (N_9669,N_9419,N_9245);
nand U9670 (N_9670,N_9178,N_9216);
or U9671 (N_9671,N_9335,N_9321);
nor U9672 (N_9672,N_9408,N_9345);
or U9673 (N_9673,N_9300,N_9498);
nor U9674 (N_9674,N_9225,N_9393);
and U9675 (N_9675,N_9028,N_9432);
or U9676 (N_9676,N_9172,N_9466);
nor U9677 (N_9677,N_9396,N_9356);
or U9678 (N_9678,N_9487,N_9138);
nand U9679 (N_9679,N_9108,N_9103);
nand U9680 (N_9680,N_9312,N_9026);
nand U9681 (N_9681,N_9015,N_9320);
nor U9682 (N_9682,N_9253,N_9184);
or U9683 (N_9683,N_9299,N_9493);
nor U9684 (N_9684,N_9441,N_9401);
or U9685 (N_9685,N_9275,N_9214);
and U9686 (N_9686,N_9433,N_9163);
nor U9687 (N_9687,N_9327,N_9328);
or U9688 (N_9688,N_9352,N_9065);
or U9689 (N_9689,N_9040,N_9449);
nand U9690 (N_9690,N_9070,N_9066);
and U9691 (N_9691,N_9166,N_9354);
or U9692 (N_9692,N_9191,N_9104);
or U9693 (N_9693,N_9315,N_9439);
and U9694 (N_9694,N_9351,N_9494);
nor U9695 (N_9695,N_9455,N_9022);
or U9696 (N_9696,N_9179,N_9336);
nand U9697 (N_9697,N_9062,N_9446);
nor U9698 (N_9698,N_9456,N_9322);
nand U9699 (N_9699,N_9143,N_9177);
nand U9700 (N_9700,N_9009,N_9086);
nand U9701 (N_9701,N_9008,N_9038);
xnor U9702 (N_9702,N_9021,N_9423);
nand U9703 (N_9703,N_9169,N_9110);
nand U9704 (N_9704,N_9490,N_9097);
nor U9705 (N_9705,N_9305,N_9236);
nor U9706 (N_9706,N_9325,N_9263);
or U9707 (N_9707,N_9017,N_9031);
and U9708 (N_9708,N_9341,N_9175);
and U9709 (N_9709,N_9365,N_9058);
nand U9710 (N_9710,N_9137,N_9249);
or U9711 (N_9711,N_9136,N_9244);
nand U9712 (N_9712,N_9277,N_9417);
or U9713 (N_9713,N_9077,N_9255);
nand U9714 (N_9714,N_9484,N_9023);
or U9715 (N_9715,N_9331,N_9486);
nor U9716 (N_9716,N_9296,N_9210);
or U9717 (N_9717,N_9496,N_9182);
or U9718 (N_9718,N_9187,N_9437);
or U9719 (N_9719,N_9386,N_9348);
or U9720 (N_9720,N_9288,N_9343);
nor U9721 (N_9721,N_9206,N_9492);
nor U9722 (N_9722,N_9134,N_9153);
nor U9723 (N_9723,N_9002,N_9468);
nor U9724 (N_9724,N_9054,N_9039);
nor U9725 (N_9725,N_9119,N_9235);
nor U9726 (N_9726,N_9284,N_9442);
or U9727 (N_9727,N_9173,N_9272);
nor U9728 (N_9728,N_9018,N_9120);
nand U9729 (N_9729,N_9257,N_9220);
and U9730 (N_9730,N_9415,N_9469);
nand U9731 (N_9731,N_9473,N_9357);
or U9732 (N_9732,N_9384,N_9400);
nand U9733 (N_9733,N_9019,N_9434);
nor U9734 (N_9734,N_9307,N_9371);
nand U9735 (N_9735,N_9397,N_9378);
and U9736 (N_9736,N_9045,N_9127);
and U9737 (N_9737,N_9231,N_9310);
or U9738 (N_9738,N_9188,N_9260);
or U9739 (N_9739,N_9431,N_9471);
or U9740 (N_9740,N_9180,N_9171);
and U9741 (N_9741,N_9130,N_9043);
nand U9742 (N_9742,N_9270,N_9329);
or U9743 (N_9743,N_9064,N_9461);
nor U9744 (N_9744,N_9061,N_9445);
or U9745 (N_9745,N_9092,N_9071);
nand U9746 (N_9746,N_9100,N_9258);
or U9747 (N_9747,N_9440,N_9291);
nor U9748 (N_9748,N_9223,N_9151);
nor U9749 (N_9749,N_9212,N_9353);
and U9750 (N_9750,N_9492,N_9258);
nand U9751 (N_9751,N_9437,N_9490);
nand U9752 (N_9752,N_9169,N_9279);
and U9753 (N_9753,N_9252,N_9485);
nor U9754 (N_9754,N_9215,N_9363);
nand U9755 (N_9755,N_9316,N_9011);
and U9756 (N_9756,N_9223,N_9414);
nand U9757 (N_9757,N_9047,N_9006);
nor U9758 (N_9758,N_9155,N_9018);
nor U9759 (N_9759,N_9440,N_9039);
and U9760 (N_9760,N_9402,N_9261);
nor U9761 (N_9761,N_9215,N_9311);
or U9762 (N_9762,N_9366,N_9474);
or U9763 (N_9763,N_9435,N_9249);
and U9764 (N_9764,N_9352,N_9228);
nor U9765 (N_9765,N_9167,N_9215);
nand U9766 (N_9766,N_9496,N_9294);
nor U9767 (N_9767,N_9052,N_9453);
or U9768 (N_9768,N_9339,N_9416);
or U9769 (N_9769,N_9332,N_9042);
xnor U9770 (N_9770,N_9215,N_9371);
nor U9771 (N_9771,N_9354,N_9033);
xnor U9772 (N_9772,N_9484,N_9432);
xnor U9773 (N_9773,N_9041,N_9021);
and U9774 (N_9774,N_9099,N_9019);
nand U9775 (N_9775,N_9363,N_9109);
nand U9776 (N_9776,N_9024,N_9166);
nor U9777 (N_9777,N_9377,N_9233);
nand U9778 (N_9778,N_9479,N_9433);
nand U9779 (N_9779,N_9266,N_9436);
and U9780 (N_9780,N_9408,N_9144);
xnor U9781 (N_9781,N_9020,N_9207);
nand U9782 (N_9782,N_9330,N_9123);
nand U9783 (N_9783,N_9134,N_9326);
nor U9784 (N_9784,N_9459,N_9425);
nor U9785 (N_9785,N_9100,N_9307);
nor U9786 (N_9786,N_9261,N_9267);
or U9787 (N_9787,N_9060,N_9288);
nor U9788 (N_9788,N_9144,N_9233);
or U9789 (N_9789,N_9405,N_9446);
or U9790 (N_9790,N_9014,N_9132);
nor U9791 (N_9791,N_9468,N_9347);
or U9792 (N_9792,N_9018,N_9083);
nor U9793 (N_9793,N_9021,N_9213);
nand U9794 (N_9794,N_9376,N_9178);
and U9795 (N_9795,N_9147,N_9062);
and U9796 (N_9796,N_9360,N_9156);
nand U9797 (N_9797,N_9390,N_9352);
nor U9798 (N_9798,N_9479,N_9052);
nor U9799 (N_9799,N_9166,N_9026);
nand U9800 (N_9800,N_9109,N_9018);
or U9801 (N_9801,N_9099,N_9413);
or U9802 (N_9802,N_9373,N_9121);
and U9803 (N_9803,N_9141,N_9083);
or U9804 (N_9804,N_9360,N_9296);
nand U9805 (N_9805,N_9406,N_9323);
and U9806 (N_9806,N_9274,N_9034);
nor U9807 (N_9807,N_9129,N_9481);
or U9808 (N_9808,N_9004,N_9360);
and U9809 (N_9809,N_9289,N_9391);
nand U9810 (N_9810,N_9148,N_9116);
and U9811 (N_9811,N_9440,N_9390);
and U9812 (N_9812,N_9355,N_9134);
nor U9813 (N_9813,N_9204,N_9085);
nand U9814 (N_9814,N_9259,N_9159);
nand U9815 (N_9815,N_9371,N_9350);
nand U9816 (N_9816,N_9318,N_9083);
and U9817 (N_9817,N_9348,N_9336);
nand U9818 (N_9818,N_9206,N_9328);
nand U9819 (N_9819,N_9174,N_9052);
and U9820 (N_9820,N_9281,N_9477);
nand U9821 (N_9821,N_9260,N_9075);
nand U9822 (N_9822,N_9108,N_9149);
or U9823 (N_9823,N_9256,N_9049);
nand U9824 (N_9824,N_9315,N_9348);
nand U9825 (N_9825,N_9158,N_9013);
or U9826 (N_9826,N_9137,N_9332);
nor U9827 (N_9827,N_9499,N_9204);
or U9828 (N_9828,N_9283,N_9173);
or U9829 (N_9829,N_9259,N_9114);
and U9830 (N_9830,N_9385,N_9366);
and U9831 (N_9831,N_9288,N_9148);
xnor U9832 (N_9832,N_9141,N_9132);
nor U9833 (N_9833,N_9227,N_9063);
nor U9834 (N_9834,N_9319,N_9392);
nor U9835 (N_9835,N_9312,N_9307);
nor U9836 (N_9836,N_9238,N_9113);
nand U9837 (N_9837,N_9328,N_9373);
or U9838 (N_9838,N_9323,N_9074);
nor U9839 (N_9839,N_9437,N_9470);
nand U9840 (N_9840,N_9146,N_9184);
nand U9841 (N_9841,N_9103,N_9400);
nor U9842 (N_9842,N_9181,N_9069);
nand U9843 (N_9843,N_9019,N_9237);
or U9844 (N_9844,N_9013,N_9116);
and U9845 (N_9845,N_9196,N_9075);
and U9846 (N_9846,N_9118,N_9371);
nor U9847 (N_9847,N_9106,N_9093);
nor U9848 (N_9848,N_9288,N_9336);
and U9849 (N_9849,N_9250,N_9149);
or U9850 (N_9850,N_9491,N_9125);
xnor U9851 (N_9851,N_9317,N_9328);
and U9852 (N_9852,N_9140,N_9371);
nand U9853 (N_9853,N_9343,N_9282);
nand U9854 (N_9854,N_9445,N_9451);
and U9855 (N_9855,N_9019,N_9316);
nand U9856 (N_9856,N_9084,N_9153);
nand U9857 (N_9857,N_9358,N_9292);
and U9858 (N_9858,N_9143,N_9362);
nand U9859 (N_9859,N_9456,N_9072);
and U9860 (N_9860,N_9493,N_9385);
nor U9861 (N_9861,N_9009,N_9282);
nand U9862 (N_9862,N_9341,N_9296);
nand U9863 (N_9863,N_9082,N_9179);
nand U9864 (N_9864,N_9303,N_9377);
xnor U9865 (N_9865,N_9279,N_9284);
nand U9866 (N_9866,N_9229,N_9429);
or U9867 (N_9867,N_9207,N_9139);
and U9868 (N_9868,N_9416,N_9319);
nor U9869 (N_9869,N_9330,N_9203);
nor U9870 (N_9870,N_9082,N_9367);
or U9871 (N_9871,N_9313,N_9408);
nor U9872 (N_9872,N_9473,N_9122);
or U9873 (N_9873,N_9126,N_9467);
and U9874 (N_9874,N_9369,N_9280);
nor U9875 (N_9875,N_9387,N_9284);
and U9876 (N_9876,N_9466,N_9240);
nor U9877 (N_9877,N_9292,N_9351);
nor U9878 (N_9878,N_9055,N_9476);
nor U9879 (N_9879,N_9288,N_9185);
nand U9880 (N_9880,N_9078,N_9172);
and U9881 (N_9881,N_9042,N_9476);
nand U9882 (N_9882,N_9111,N_9258);
nor U9883 (N_9883,N_9027,N_9446);
nor U9884 (N_9884,N_9148,N_9189);
or U9885 (N_9885,N_9324,N_9188);
nor U9886 (N_9886,N_9117,N_9280);
nand U9887 (N_9887,N_9256,N_9157);
and U9888 (N_9888,N_9149,N_9122);
nor U9889 (N_9889,N_9383,N_9251);
nor U9890 (N_9890,N_9243,N_9290);
and U9891 (N_9891,N_9006,N_9180);
nand U9892 (N_9892,N_9065,N_9191);
or U9893 (N_9893,N_9033,N_9413);
or U9894 (N_9894,N_9036,N_9125);
and U9895 (N_9895,N_9285,N_9455);
and U9896 (N_9896,N_9244,N_9270);
and U9897 (N_9897,N_9359,N_9391);
or U9898 (N_9898,N_9033,N_9041);
and U9899 (N_9899,N_9299,N_9484);
or U9900 (N_9900,N_9311,N_9252);
and U9901 (N_9901,N_9173,N_9361);
or U9902 (N_9902,N_9351,N_9162);
and U9903 (N_9903,N_9112,N_9059);
or U9904 (N_9904,N_9224,N_9486);
and U9905 (N_9905,N_9224,N_9491);
or U9906 (N_9906,N_9312,N_9108);
or U9907 (N_9907,N_9123,N_9030);
nor U9908 (N_9908,N_9435,N_9295);
nand U9909 (N_9909,N_9296,N_9170);
nor U9910 (N_9910,N_9138,N_9159);
nor U9911 (N_9911,N_9375,N_9011);
nor U9912 (N_9912,N_9105,N_9251);
nand U9913 (N_9913,N_9045,N_9115);
nand U9914 (N_9914,N_9267,N_9344);
or U9915 (N_9915,N_9223,N_9362);
nor U9916 (N_9916,N_9434,N_9137);
nor U9917 (N_9917,N_9299,N_9324);
and U9918 (N_9918,N_9262,N_9361);
or U9919 (N_9919,N_9027,N_9196);
nor U9920 (N_9920,N_9285,N_9111);
nor U9921 (N_9921,N_9137,N_9170);
and U9922 (N_9922,N_9225,N_9423);
and U9923 (N_9923,N_9128,N_9048);
nand U9924 (N_9924,N_9401,N_9066);
and U9925 (N_9925,N_9225,N_9131);
nor U9926 (N_9926,N_9384,N_9248);
or U9927 (N_9927,N_9173,N_9135);
or U9928 (N_9928,N_9122,N_9204);
and U9929 (N_9929,N_9296,N_9444);
and U9930 (N_9930,N_9101,N_9462);
or U9931 (N_9931,N_9364,N_9012);
nand U9932 (N_9932,N_9077,N_9119);
nor U9933 (N_9933,N_9010,N_9287);
nand U9934 (N_9934,N_9088,N_9426);
nor U9935 (N_9935,N_9110,N_9229);
nor U9936 (N_9936,N_9176,N_9367);
and U9937 (N_9937,N_9496,N_9369);
nor U9938 (N_9938,N_9314,N_9205);
and U9939 (N_9939,N_9174,N_9049);
nor U9940 (N_9940,N_9280,N_9488);
nor U9941 (N_9941,N_9128,N_9040);
or U9942 (N_9942,N_9048,N_9365);
or U9943 (N_9943,N_9070,N_9113);
nand U9944 (N_9944,N_9225,N_9023);
nand U9945 (N_9945,N_9220,N_9493);
nand U9946 (N_9946,N_9163,N_9259);
nand U9947 (N_9947,N_9035,N_9098);
nor U9948 (N_9948,N_9087,N_9418);
or U9949 (N_9949,N_9345,N_9207);
and U9950 (N_9950,N_9474,N_9480);
nand U9951 (N_9951,N_9145,N_9156);
and U9952 (N_9952,N_9156,N_9257);
or U9953 (N_9953,N_9457,N_9352);
nand U9954 (N_9954,N_9364,N_9425);
and U9955 (N_9955,N_9461,N_9411);
or U9956 (N_9956,N_9198,N_9022);
and U9957 (N_9957,N_9206,N_9129);
nand U9958 (N_9958,N_9190,N_9015);
nand U9959 (N_9959,N_9326,N_9035);
nand U9960 (N_9960,N_9120,N_9084);
or U9961 (N_9961,N_9240,N_9123);
and U9962 (N_9962,N_9203,N_9217);
and U9963 (N_9963,N_9463,N_9303);
and U9964 (N_9964,N_9457,N_9225);
or U9965 (N_9965,N_9023,N_9093);
and U9966 (N_9966,N_9350,N_9209);
or U9967 (N_9967,N_9499,N_9027);
and U9968 (N_9968,N_9362,N_9309);
nand U9969 (N_9969,N_9275,N_9203);
or U9970 (N_9970,N_9212,N_9397);
or U9971 (N_9971,N_9306,N_9414);
nor U9972 (N_9972,N_9361,N_9240);
nor U9973 (N_9973,N_9437,N_9145);
and U9974 (N_9974,N_9278,N_9455);
nor U9975 (N_9975,N_9359,N_9067);
nor U9976 (N_9976,N_9360,N_9214);
and U9977 (N_9977,N_9195,N_9400);
nor U9978 (N_9978,N_9469,N_9113);
and U9979 (N_9979,N_9191,N_9255);
nand U9980 (N_9980,N_9337,N_9393);
and U9981 (N_9981,N_9094,N_9204);
or U9982 (N_9982,N_9126,N_9253);
or U9983 (N_9983,N_9293,N_9171);
and U9984 (N_9984,N_9246,N_9482);
or U9985 (N_9985,N_9297,N_9347);
nand U9986 (N_9986,N_9380,N_9018);
and U9987 (N_9987,N_9482,N_9121);
or U9988 (N_9988,N_9371,N_9163);
and U9989 (N_9989,N_9008,N_9002);
or U9990 (N_9990,N_9289,N_9029);
nor U9991 (N_9991,N_9407,N_9493);
or U9992 (N_9992,N_9478,N_9366);
nor U9993 (N_9993,N_9433,N_9346);
nand U9994 (N_9994,N_9106,N_9028);
nor U9995 (N_9995,N_9143,N_9233);
and U9996 (N_9996,N_9025,N_9337);
nand U9997 (N_9997,N_9443,N_9232);
and U9998 (N_9998,N_9389,N_9122);
nor U9999 (N_9999,N_9352,N_9179);
nand U10000 (N_10000,N_9951,N_9572);
and U10001 (N_10001,N_9931,N_9971);
or U10002 (N_10002,N_9631,N_9768);
and U10003 (N_10003,N_9911,N_9502);
and U10004 (N_10004,N_9942,N_9763);
or U10005 (N_10005,N_9505,N_9541);
nor U10006 (N_10006,N_9937,N_9816);
or U10007 (N_10007,N_9757,N_9566);
nand U10008 (N_10008,N_9758,N_9944);
and U10009 (N_10009,N_9679,N_9531);
nand U10010 (N_10010,N_9526,N_9953);
nand U10011 (N_10011,N_9610,N_9893);
and U10012 (N_10012,N_9929,N_9964);
nand U10013 (N_10013,N_9614,N_9875);
nand U10014 (N_10014,N_9690,N_9878);
and U10015 (N_10015,N_9984,N_9595);
nor U10016 (N_10016,N_9829,N_9688);
nor U10017 (N_10017,N_9990,N_9556);
or U10018 (N_10018,N_9969,N_9537);
or U10019 (N_10019,N_9930,N_9504);
or U10020 (N_10020,N_9926,N_9613);
or U10021 (N_10021,N_9745,N_9698);
or U10022 (N_10022,N_9542,N_9821);
xnor U10023 (N_10023,N_9822,N_9905);
nor U10024 (N_10024,N_9854,N_9594);
nand U10025 (N_10025,N_9810,N_9887);
and U10026 (N_10026,N_9622,N_9922);
nor U10027 (N_10027,N_9928,N_9647);
and U10028 (N_10028,N_9949,N_9507);
nand U10029 (N_10029,N_9718,N_9766);
or U10030 (N_10030,N_9644,N_9805);
or U10031 (N_10031,N_9597,N_9569);
or U10032 (N_10032,N_9714,N_9914);
nand U10033 (N_10033,N_9722,N_9789);
and U10034 (N_10034,N_9880,N_9624);
and U10035 (N_10035,N_9909,N_9847);
and U10036 (N_10036,N_9617,N_9574);
and U10037 (N_10037,N_9856,N_9790);
nand U10038 (N_10038,N_9673,N_9589);
or U10039 (N_10039,N_9948,N_9976);
and U10040 (N_10040,N_9642,N_9511);
and U10041 (N_10041,N_9888,N_9695);
nor U10042 (N_10042,N_9962,N_9648);
nor U10043 (N_10043,N_9588,N_9960);
or U10044 (N_10044,N_9662,N_9533);
nand U10045 (N_10045,N_9573,N_9672);
nand U10046 (N_10046,N_9958,N_9705);
and U10047 (N_10047,N_9635,N_9515);
or U10048 (N_10048,N_9711,N_9826);
nor U10049 (N_10049,N_9563,N_9774);
nor U10050 (N_10050,N_9756,N_9978);
or U10051 (N_10051,N_9609,N_9568);
xnor U10052 (N_10052,N_9667,N_9837);
and U10053 (N_10053,N_9501,N_9550);
or U10054 (N_10054,N_9967,N_9830);
or U10055 (N_10055,N_9834,N_9866);
and U10056 (N_10056,N_9643,N_9625);
nor U10057 (N_10057,N_9612,N_9770);
nor U10058 (N_10058,N_9818,N_9655);
and U10059 (N_10059,N_9611,N_9882);
or U10060 (N_10060,N_9862,N_9513);
nand U10061 (N_10061,N_9633,N_9986);
nor U10062 (N_10062,N_9927,N_9831);
nand U10063 (N_10063,N_9736,N_9925);
nor U10064 (N_10064,N_9506,N_9733);
and U10065 (N_10065,N_9970,N_9699);
or U10066 (N_10066,N_9913,N_9720);
and U10067 (N_10067,N_9751,N_9988);
nor U10068 (N_10068,N_9889,N_9605);
nand U10069 (N_10069,N_9656,N_9580);
nand U10070 (N_10070,N_9686,N_9972);
or U10071 (N_10071,N_9744,N_9777);
or U10072 (N_10072,N_9823,N_9529);
nand U10073 (N_10073,N_9665,N_9702);
and U10074 (N_10074,N_9739,N_9780);
nand U10075 (N_10075,N_9668,N_9606);
nor U10076 (N_10076,N_9833,N_9982);
and U10077 (N_10077,N_9973,N_9754);
and U10078 (N_10078,N_9527,N_9747);
or U10079 (N_10079,N_9968,N_9996);
and U10080 (N_10080,N_9868,N_9576);
nor U10081 (N_10081,N_9603,N_9808);
or U10082 (N_10082,N_9799,N_9782);
or U10083 (N_10083,N_9728,N_9985);
nor U10084 (N_10084,N_9998,N_9784);
nand U10085 (N_10085,N_9678,N_9932);
nor U10086 (N_10086,N_9734,N_9980);
nand U10087 (N_10087,N_9650,N_9508);
nor U10088 (N_10088,N_9737,N_9957);
and U10089 (N_10089,N_9836,N_9634);
nor U10090 (N_10090,N_9850,N_9883);
nand U10091 (N_10091,N_9864,N_9807);
nand U10092 (N_10092,N_9917,N_9682);
nand U10093 (N_10093,N_9583,N_9760);
and U10094 (N_10094,N_9947,N_9955);
or U10095 (N_10095,N_9706,N_9767);
xor U10096 (N_10096,N_9865,N_9729);
nor U10097 (N_10097,N_9628,N_9881);
nand U10098 (N_10098,N_9709,N_9540);
nor U10099 (N_10099,N_9886,N_9804);
nand U10100 (N_10100,N_9708,N_9559);
and U10101 (N_10101,N_9906,N_9590);
or U10102 (N_10102,N_9997,N_9827);
nand U10103 (N_10103,N_9994,N_9658);
or U10104 (N_10104,N_9901,N_9908);
nand U10105 (N_10105,N_9910,N_9983);
or U10106 (N_10106,N_9748,N_9840);
nand U10107 (N_10107,N_9602,N_9579);
nand U10108 (N_10108,N_9921,N_9661);
and U10109 (N_10109,N_9918,N_9731);
and U10110 (N_10110,N_9548,N_9727);
nor U10111 (N_10111,N_9759,N_9891);
nand U10112 (N_10112,N_9564,N_9813);
nand U10113 (N_10113,N_9554,N_9623);
nor U10114 (N_10114,N_9752,N_9920);
and U10115 (N_10115,N_9743,N_9538);
and U10116 (N_10116,N_9860,N_9870);
nand U10117 (N_10117,N_9794,N_9512);
or U10118 (N_10118,N_9943,N_9730);
or U10119 (N_10119,N_9534,N_9791);
nor U10120 (N_10120,N_9692,N_9697);
or U10121 (N_10121,N_9773,N_9859);
xnor U10122 (N_10122,N_9669,N_9523);
and U10123 (N_10123,N_9663,N_9638);
nor U10124 (N_10124,N_9771,N_9520);
or U10125 (N_10125,N_9849,N_9577);
nor U10126 (N_10126,N_9786,N_9549);
or U10127 (N_10127,N_9629,N_9912);
or U10128 (N_10128,N_9660,N_9919);
nand U10129 (N_10129,N_9500,N_9735);
nand U10130 (N_10130,N_9558,N_9867);
or U10131 (N_10131,N_9701,N_9959);
xnor U10132 (N_10132,N_9599,N_9879);
nand U10133 (N_10133,N_9936,N_9788);
xor U10134 (N_10134,N_9700,N_9664);
and U10135 (N_10135,N_9578,N_9899);
nand U10136 (N_10136,N_9800,N_9845);
nand U10137 (N_10137,N_9832,N_9570);
nand U10138 (N_10138,N_9896,N_9704);
and U10139 (N_10139,N_9809,N_9979);
nand U10140 (N_10140,N_9607,N_9742);
nand U10141 (N_10141,N_9503,N_9726);
or U10142 (N_10142,N_9544,N_9975);
or U10143 (N_10143,N_9966,N_9584);
nor U10144 (N_10144,N_9924,N_9934);
nand U10145 (N_10145,N_9820,N_9645);
or U10146 (N_10146,N_9546,N_9775);
and U10147 (N_10147,N_9941,N_9749);
or U10148 (N_10148,N_9684,N_9898);
nor U10149 (N_10149,N_9819,N_9871);
nor U10150 (N_10150,N_9670,N_9939);
nand U10151 (N_10151,N_9761,N_9565);
nor U10152 (N_10152,N_9999,N_9853);
nand U10153 (N_10153,N_9619,N_9516);
nand U10154 (N_10154,N_9715,N_9659);
and U10155 (N_10155,N_9600,N_9872);
and U10156 (N_10156,N_9876,N_9591);
and U10157 (N_10157,N_9769,N_9646);
and U10158 (N_10158,N_9765,N_9935);
nand U10159 (N_10159,N_9651,N_9802);
or U10160 (N_10160,N_9993,N_9553);
nor U10161 (N_10161,N_9618,N_9779);
nor U10162 (N_10162,N_9904,N_9547);
or U10163 (N_10163,N_9676,N_9518);
or U10164 (N_10164,N_9992,N_9521);
xor U10165 (N_10165,N_9693,N_9626);
nand U10166 (N_10166,N_9861,N_9963);
and U10167 (N_10167,N_9776,N_9652);
nor U10168 (N_10168,N_9680,N_9723);
and U10169 (N_10169,N_9815,N_9630);
and U10170 (N_10170,N_9848,N_9687);
and U10171 (N_10171,N_9787,N_9894);
and U10172 (N_10172,N_9961,N_9778);
nor U10173 (N_10173,N_9838,N_9923);
and U10174 (N_10174,N_9863,N_9907);
and U10175 (N_10175,N_9689,N_9694);
nand U10176 (N_10176,N_9677,N_9890);
and U10177 (N_10177,N_9916,N_9965);
and U10178 (N_10178,N_9915,N_9873);
and U10179 (N_10179,N_9892,N_9811);
nor U10180 (N_10180,N_9545,N_9795);
or U10181 (N_10181,N_9675,N_9674);
and U10182 (N_10182,N_9987,N_9510);
and U10183 (N_10183,N_9741,N_9536);
nor U10184 (N_10184,N_9524,N_9842);
nand U10185 (N_10185,N_9707,N_9902);
and U10186 (N_10186,N_9637,N_9897);
nor U10187 (N_10187,N_9683,N_9828);
nor U10188 (N_10188,N_9575,N_9552);
nor U10189 (N_10189,N_9785,N_9596);
nor U10190 (N_10190,N_9940,N_9641);
or U10191 (N_10191,N_9514,N_9846);
and U10192 (N_10192,N_9657,N_9781);
xor U10193 (N_10193,N_9627,N_9817);
nor U10194 (N_10194,N_9592,N_9582);
nor U10195 (N_10195,N_9843,N_9814);
nand U10196 (N_10196,N_9855,N_9806);
or U10197 (N_10197,N_9793,N_9710);
and U10198 (N_10198,N_9740,N_9945);
nand U10199 (N_10199,N_9933,N_9654);
nand U10200 (N_10200,N_9801,N_9532);
nand U10201 (N_10201,N_9604,N_9798);
and U10202 (N_10202,N_9825,N_9716);
nand U10203 (N_10203,N_9750,N_9525);
nor U10204 (N_10204,N_9571,N_9858);
xnor U10205 (N_10205,N_9632,N_9703);
or U10206 (N_10206,N_9835,N_9903);
or U10207 (N_10207,N_9666,N_9755);
nor U10208 (N_10208,N_9974,N_9621);
nor U10209 (N_10209,N_9713,N_9803);
nor U10210 (N_10210,N_9608,N_9691);
and U10211 (N_10211,N_9989,N_9995);
or U10212 (N_10212,N_9952,N_9732);
nand U10213 (N_10213,N_9685,N_9885);
or U10214 (N_10214,N_9696,N_9567);
and U10215 (N_10215,N_9681,N_9796);
and U10216 (N_10216,N_9649,N_9519);
and U10217 (N_10217,N_9551,N_9581);
and U10218 (N_10218,N_9852,N_9844);
or U10219 (N_10219,N_9585,N_9509);
nand U10220 (N_10220,N_9764,N_9772);
nand U10221 (N_10221,N_9762,N_9517);
or U10222 (N_10222,N_9620,N_9528);
and U10223 (N_10223,N_9938,N_9555);
nand U10224 (N_10224,N_9981,N_9535);
nor U10225 (N_10225,N_9562,N_9869);
and U10226 (N_10226,N_9719,N_9560);
xnor U10227 (N_10227,N_9851,N_9616);
or U10228 (N_10228,N_9950,N_9615);
nand U10229 (N_10229,N_9530,N_9839);
or U10230 (N_10230,N_9753,N_9812);
nor U10231 (N_10231,N_9783,N_9598);
xnor U10232 (N_10232,N_9954,N_9522);
nor U10233 (N_10233,N_9671,N_9601);
nand U10234 (N_10234,N_9946,N_9653);
nand U10235 (N_10235,N_9561,N_9895);
and U10236 (N_10236,N_9874,N_9586);
nand U10237 (N_10237,N_9725,N_9539);
nor U10238 (N_10238,N_9721,N_9877);
or U10239 (N_10239,N_9956,N_9991);
or U10240 (N_10240,N_9557,N_9841);
nor U10241 (N_10241,N_9977,N_9797);
nor U10242 (N_10242,N_9543,N_9640);
nand U10243 (N_10243,N_9738,N_9746);
or U10244 (N_10244,N_9792,N_9593);
nor U10245 (N_10245,N_9724,N_9587);
nor U10246 (N_10246,N_9636,N_9824);
nor U10247 (N_10247,N_9717,N_9712);
and U10248 (N_10248,N_9900,N_9639);
nor U10249 (N_10249,N_9857,N_9884);
or U10250 (N_10250,N_9649,N_9645);
nand U10251 (N_10251,N_9530,N_9949);
and U10252 (N_10252,N_9635,N_9977);
nand U10253 (N_10253,N_9795,N_9735);
and U10254 (N_10254,N_9531,N_9981);
or U10255 (N_10255,N_9698,N_9563);
nor U10256 (N_10256,N_9698,N_9839);
xnor U10257 (N_10257,N_9863,N_9616);
and U10258 (N_10258,N_9704,N_9520);
and U10259 (N_10259,N_9793,N_9792);
and U10260 (N_10260,N_9553,N_9507);
or U10261 (N_10261,N_9819,N_9993);
or U10262 (N_10262,N_9553,N_9564);
nor U10263 (N_10263,N_9855,N_9893);
and U10264 (N_10264,N_9977,N_9647);
or U10265 (N_10265,N_9539,N_9782);
xnor U10266 (N_10266,N_9933,N_9601);
nor U10267 (N_10267,N_9674,N_9695);
or U10268 (N_10268,N_9640,N_9635);
or U10269 (N_10269,N_9963,N_9742);
or U10270 (N_10270,N_9740,N_9532);
or U10271 (N_10271,N_9527,N_9703);
or U10272 (N_10272,N_9580,N_9920);
nand U10273 (N_10273,N_9762,N_9814);
or U10274 (N_10274,N_9867,N_9525);
or U10275 (N_10275,N_9828,N_9858);
or U10276 (N_10276,N_9773,N_9523);
nand U10277 (N_10277,N_9833,N_9795);
or U10278 (N_10278,N_9678,N_9973);
nor U10279 (N_10279,N_9507,N_9558);
and U10280 (N_10280,N_9582,N_9833);
nor U10281 (N_10281,N_9949,N_9782);
and U10282 (N_10282,N_9608,N_9589);
nor U10283 (N_10283,N_9631,N_9821);
xor U10284 (N_10284,N_9958,N_9838);
or U10285 (N_10285,N_9893,N_9939);
or U10286 (N_10286,N_9557,N_9678);
xor U10287 (N_10287,N_9552,N_9634);
or U10288 (N_10288,N_9754,N_9549);
or U10289 (N_10289,N_9678,N_9525);
nand U10290 (N_10290,N_9548,N_9705);
nand U10291 (N_10291,N_9942,N_9619);
nor U10292 (N_10292,N_9543,N_9632);
or U10293 (N_10293,N_9806,N_9647);
nand U10294 (N_10294,N_9943,N_9602);
and U10295 (N_10295,N_9512,N_9528);
nand U10296 (N_10296,N_9656,N_9977);
and U10297 (N_10297,N_9860,N_9934);
and U10298 (N_10298,N_9925,N_9602);
or U10299 (N_10299,N_9969,N_9750);
and U10300 (N_10300,N_9580,N_9555);
nor U10301 (N_10301,N_9599,N_9707);
nor U10302 (N_10302,N_9748,N_9533);
nor U10303 (N_10303,N_9652,N_9592);
and U10304 (N_10304,N_9535,N_9879);
and U10305 (N_10305,N_9682,N_9816);
xnor U10306 (N_10306,N_9919,N_9986);
and U10307 (N_10307,N_9797,N_9641);
nor U10308 (N_10308,N_9814,N_9604);
nand U10309 (N_10309,N_9678,N_9584);
or U10310 (N_10310,N_9712,N_9805);
nor U10311 (N_10311,N_9912,N_9811);
nand U10312 (N_10312,N_9728,N_9993);
nor U10313 (N_10313,N_9665,N_9923);
and U10314 (N_10314,N_9703,N_9532);
nor U10315 (N_10315,N_9938,N_9728);
nand U10316 (N_10316,N_9773,N_9837);
and U10317 (N_10317,N_9561,N_9736);
or U10318 (N_10318,N_9967,N_9818);
nand U10319 (N_10319,N_9753,N_9695);
or U10320 (N_10320,N_9586,N_9730);
or U10321 (N_10321,N_9653,N_9924);
nor U10322 (N_10322,N_9675,N_9667);
and U10323 (N_10323,N_9556,N_9861);
nor U10324 (N_10324,N_9848,N_9898);
nor U10325 (N_10325,N_9949,N_9739);
or U10326 (N_10326,N_9579,N_9724);
and U10327 (N_10327,N_9891,N_9722);
and U10328 (N_10328,N_9663,N_9974);
nor U10329 (N_10329,N_9781,N_9593);
xnor U10330 (N_10330,N_9890,N_9672);
nand U10331 (N_10331,N_9892,N_9775);
nand U10332 (N_10332,N_9659,N_9661);
nand U10333 (N_10333,N_9665,N_9567);
nor U10334 (N_10334,N_9745,N_9619);
or U10335 (N_10335,N_9777,N_9506);
and U10336 (N_10336,N_9836,N_9600);
or U10337 (N_10337,N_9942,N_9887);
and U10338 (N_10338,N_9624,N_9824);
or U10339 (N_10339,N_9853,N_9789);
and U10340 (N_10340,N_9579,N_9781);
nand U10341 (N_10341,N_9501,N_9786);
nand U10342 (N_10342,N_9802,N_9541);
and U10343 (N_10343,N_9557,N_9769);
nand U10344 (N_10344,N_9787,N_9542);
and U10345 (N_10345,N_9744,N_9674);
xor U10346 (N_10346,N_9741,N_9624);
nand U10347 (N_10347,N_9722,N_9552);
nand U10348 (N_10348,N_9618,N_9754);
nor U10349 (N_10349,N_9666,N_9928);
or U10350 (N_10350,N_9918,N_9657);
and U10351 (N_10351,N_9548,N_9930);
or U10352 (N_10352,N_9565,N_9823);
or U10353 (N_10353,N_9779,N_9823);
nand U10354 (N_10354,N_9581,N_9638);
nor U10355 (N_10355,N_9887,N_9969);
or U10356 (N_10356,N_9992,N_9750);
and U10357 (N_10357,N_9981,N_9904);
nor U10358 (N_10358,N_9862,N_9848);
or U10359 (N_10359,N_9574,N_9861);
and U10360 (N_10360,N_9713,N_9840);
nor U10361 (N_10361,N_9602,N_9580);
and U10362 (N_10362,N_9665,N_9691);
and U10363 (N_10363,N_9743,N_9537);
and U10364 (N_10364,N_9855,N_9844);
nor U10365 (N_10365,N_9958,N_9537);
and U10366 (N_10366,N_9739,N_9732);
nor U10367 (N_10367,N_9629,N_9978);
and U10368 (N_10368,N_9617,N_9560);
nor U10369 (N_10369,N_9949,N_9778);
or U10370 (N_10370,N_9567,N_9566);
or U10371 (N_10371,N_9863,N_9608);
and U10372 (N_10372,N_9519,N_9775);
and U10373 (N_10373,N_9811,N_9966);
nor U10374 (N_10374,N_9793,N_9517);
nor U10375 (N_10375,N_9864,N_9949);
and U10376 (N_10376,N_9736,N_9792);
nor U10377 (N_10377,N_9552,N_9969);
nor U10378 (N_10378,N_9668,N_9821);
or U10379 (N_10379,N_9802,N_9963);
and U10380 (N_10380,N_9675,N_9552);
nand U10381 (N_10381,N_9673,N_9573);
nand U10382 (N_10382,N_9568,N_9957);
nand U10383 (N_10383,N_9743,N_9753);
xnor U10384 (N_10384,N_9818,N_9963);
nand U10385 (N_10385,N_9885,N_9726);
or U10386 (N_10386,N_9881,N_9592);
and U10387 (N_10387,N_9829,N_9504);
nor U10388 (N_10388,N_9548,N_9604);
nor U10389 (N_10389,N_9559,N_9779);
nand U10390 (N_10390,N_9965,N_9702);
and U10391 (N_10391,N_9871,N_9550);
or U10392 (N_10392,N_9708,N_9902);
or U10393 (N_10393,N_9925,N_9812);
nand U10394 (N_10394,N_9985,N_9950);
nor U10395 (N_10395,N_9565,N_9864);
or U10396 (N_10396,N_9834,N_9774);
or U10397 (N_10397,N_9912,N_9982);
nor U10398 (N_10398,N_9634,N_9900);
nor U10399 (N_10399,N_9796,N_9803);
nand U10400 (N_10400,N_9818,N_9607);
nor U10401 (N_10401,N_9533,N_9727);
and U10402 (N_10402,N_9967,N_9748);
nor U10403 (N_10403,N_9523,N_9508);
or U10404 (N_10404,N_9967,N_9803);
or U10405 (N_10405,N_9882,N_9573);
and U10406 (N_10406,N_9708,N_9738);
or U10407 (N_10407,N_9918,N_9733);
and U10408 (N_10408,N_9581,N_9636);
nand U10409 (N_10409,N_9905,N_9580);
xor U10410 (N_10410,N_9614,N_9725);
and U10411 (N_10411,N_9997,N_9666);
xor U10412 (N_10412,N_9853,N_9602);
and U10413 (N_10413,N_9575,N_9728);
nand U10414 (N_10414,N_9584,N_9608);
and U10415 (N_10415,N_9931,N_9944);
or U10416 (N_10416,N_9701,N_9832);
or U10417 (N_10417,N_9704,N_9808);
nor U10418 (N_10418,N_9879,N_9576);
nor U10419 (N_10419,N_9977,N_9946);
nor U10420 (N_10420,N_9589,N_9683);
or U10421 (N_10421,N_9722,N_9555);
and U10422 (N_10422,N_9703,N_9879);
nand U10423 (N_10423,N_9955,N_9746);
or U10424 (N_10424,N_9750,N_9626);
nand U10425 (N_10425,N_9535,N_9544);
nor U10426 (N_10426,N_9974,N_9803);
nor U10427 (N_10427,N_9962,N_9526);
or U10428 (N_10428,N_9717,N_9549);
and U10429 (N_10429,N_9608,N_9732);
nor U10430 (N_10430,N_9600,N_9800);
nand U10431 (N_10431,N_9884,N_9625);
and U10432 (N_10432,N_9531,N_9777);
or U10433 (N_10433,N_9643,N_9692);
nand U10434 (N_10434,N_9743,N_9918);
or U10435 (N_10435,N_9661,N_9998);
nand U10436 (N_10436,N_9641,N_9647);
nor U10437 (N_10437,N_9982,N_9918);
nor U10438 (N_10438,N_9534,N_9571);
nand U10439 (N_10439,N_9908,N_9857);
nor U10440 (N_10440,N_9683,N_9923);
nor U10441 (N_10441,N_9591,N_9921);
or U10442 (N_10442,N_9584,N_9580);
and U10443 (N_10443,N_9536,N_9933);
nor U10444 (N_10444,N_9655,N_9743);
and U10445 (N_10445,N_9858,N_9517);
and U10446 (N_10446,N_9834,N_9668);
nor U10447 (N_10447,N_9810,N_9635);
nand U10448 (N_10448,N_9540,N_9851);
nand U10449 (N_10449,N_9969,N_9764);
nor U10450 (N_10450,N_9622,N_9501);
nor U10451 (N_10451,N_9631,N_9502);
and U10452 (N_10452,N_9518,N_9630);
nand U10453 (N_10453,N_9594,N_9917);
and U10454 (N_10454,N_9734,N_9852);
and U10455 (N_10455,N_9597,N_9841);
and U10456 (N_10456,N_9583,N_9667);
nand U10457 (N_10457,N_9705,N_9670);
nor U10458 (N_10458,N_9883,N_9786);
nor U10459 (N_10459,N_9794,N_9519);
and U10460 (N_10460,N_9809,N_9852);
and U10461 (N_10461,N_9601,N_9727);
nand U10462 (N_10462,N_9965,N_9535);
nor U10463 (N_10463,N_9748,N_9929);
nand U10464 (N_10464,N_9934,N_9905);
and U10465 (N_10465,N_9931,N_9925);
nor U10466 (N_10466,N_9859,N_9669);
or U10467 (N_10467,N_9639,N_9693);
nand U10468 (N_10468,N_9790,N_9968);
nand U10469 (N_10469,N_9554,N_9540);
nor U10470 (N_10470,N_9567,N_9562);
or U10471 (N_10471,N_9994,N_9892);
and U10472 (N_10472,N_9770,N_9734);
and U10473 (N_10473,N_9613,N_9790);
or U10474 (N_10474,N_9561,N_9525);
and U10475 (N_10475,N_9856,N_9797);
or U10476 (N_10476,N_9954,N_9899);
and U10477 (N_10477,N_9802,N_9746);
and U10478 (N_10478,N_9537,N_9962);
and U10479 (N_10479,N_9512,N_9822);
nor U10480 (N_10480,N_9878,N_9990);
nor U10481 (N_10481,N_9636,N_9509);
and U10482 (N_10482,N_9928,N_9599);
or U10483 (N_10483,N_9807,N_9908);
nor U10484 (N_10484,N_9922,N_9939);
nor U10485 (N_10485,N_9736,N_9697);
nor U10486 (N_10486,N_9964,N_9588);
and U10487 (N_10487,N_9541,N_9791);
or U10488 (N_10488,N_9939,N_9867);
or U10489 (N_10489,N_9634,N_9992);
and U10490 (N_10490,N_9910,N_9881);
nand U10491 (N_10491,N_9826,N_9681);
nor U10492 (N_10492,N_9871,N_9539);
or U10493 (N_10493,N_9916,N_9942);
nand U10494 (N_10494,N_9748,N_9724);
nor U10495 (N_10495,N_9586,N_9566);
nand U10496 (N_10496,N_9562,N_9652);
and U10497 (N_10497,N_9659,N_9534);
and U10498 (N_10498,N_9751,N_9602);
nor U10499 (N_10499,N_9763,N_9693);
nor U10500 (N_10500,N_10101,N_10108);
and U10501 (N_10501,N_10320,N_10382);
nand U10502 (N_10502,N_10274,N_10360);
nand U10503 (N_10503,N_10296,N_10275);
and U10504 (N_10504,N_10017,N_10450);
nor U10505 (N_10505,N_10457,N_10227);
or U10506 (N_10506,N_10151,N_10342);
and U10507 (N_10507,N_10386,N_10220);
or U10508 (N_10508,N_10150,N_10468);
and U10509 (N_10509,N_10381,N_10188);
or U10510 (N_10510,N_10399,N_10126);
nand U10511 (N_10511,N_10347,N_10025);
and U10512 (N_10512,N_10070,N_10125);
nand U10513 (N_10513,N_10333,N_10395);
nand U10514 (N_10514,N_10096,N_10475);
nor U10515 (N_10515,N_10470,N_10169);
nand U10516 (N_10516,N_10272,N_10459);
or U10517 (N_10517,N_10303,N_10435);
or U10518 (N_10518,N_10001,N_10461);
nand U10519 (N_10519,N_10196,N_10172);
nor U10520 (N_10520,N_10261,N_10400);
nand U10521 (N_10521,N_10350,N_10094);
and U10522 (N_10522,N_10484,N_10144);
nand U10523 (N_10523,N_10233,N_10408);
or U10524 (N_10524,N_10106,N_10492);
nor U10525 (N_10525,N_10203,N_10329);
and U10526 (N_10526,N_10281,N_10288);
or U10527 (N_10527,N_10002,N_10341);
nor U10528 (N_10528,N_10077,N_10011);
nor U10529 (N_10529,N_10121,N_10195);
nor U10530 (N_10530,N_10419,N_10112);
or U10531 (N_10531,N_10302,N_10117);
nor U10532 (N_10532,N_10184,N_10310);
nor U10533 (N_10533,N_10279,N_10245);
nor U10534 (N_10534,N_10149,N_10388);
xor U10535 (N_10535,N_10438,N_10051);
nand U10536 (N_10536,N_10278,N_10130);
nand U10537 (N_10537,N_10217,N_10481);
or U10538 (N_10538,N_10029,N_10028);
or U10539 (N_10539,N_10050,N_10043);
nor U10540 (N_10540,N_10476,N_10344);
nand U10541 (N_10541,N_10204,N_10058);
or U10542 (N_10542,N_10016,N_10346);
and U10543 (N_10543,N_10014,N_10053);
and U10544 (N_10544,N_10390,N_10452);
xnor U10545 (N_10545,N_10006,N_10467);
or U10546 (N_10546,N_10335,N_10059);
and U10547 (N_10547,N_10009,N_10191);
and U10548 (N_10548,N_10349,N_10216);
or U10549 (N_10549,N_10116,N_10298);
or U10550 (N_10550,N_10198,N_10123);
nand U10551 (N_10551,N_10215,N_10308);
and U10552 (N_10552,N_10205,N_10165);
and U10553 (N_10553,N_10113,N_10371);
or U10554 (N_10554,N_10404,N_10389);
and U10555 (N_10555,N_10361,N_10460);
xor U10556 (N_10556,N_10328,N_10482);
and U10557 (N_10557,N_10474,N_10441);
nand U10558 (N_10558,N_10238,N_10168);
and U10559 (N_10559,N_10148,N_10127);
xor U10560 (N_10560,N_10192,N_10005);
nand U10561 (N_10561,N_10301,N_10283);
nand U10562 (N_10562,N_10102,N_10264);
nand U10563 (N_10563,N_10250,N_10396);
nor U10564 (N_10564,N_10115,N_10407);
nor U10565 (N_10565,N_10498,N_10224);
and U10566 (N_10566,N_10472,N_10182);
or U10567 (N_10567,N_10236,N_10253);
or U10568 (N_10568,N_10026,N_10131);
nand U10569 (N_10569,N_10416,N_10294);
or U10570 (N_10570,N_10495,N_10060);
nand U10571 (N_10571,N_10242,N_10097);
nand U10572 (N_10572,N_10075,N_10318);
or U10573 (N_10573,N_10260,N_10269);
nor U10574 (N_10574,N_10199,N_10212);
nor U10575 (N_10575,N_10262,N_10120);
or U10576 (N_10576,N_10339,N_10083);
and U10577 (N_10577,N_10426,N_10249);
nand U10578 (N_10578,N_10417,N_10081);
nor U10579 (N_10579,N_10047,N_10137);
or U10580 (N_10580,N_10394,N_10436);
and U10581 (N_10581,N_10041,N_10076);
and U10582 (N_10582,N_10143,N_10122);
nand U10583 (N_10583,N_10379,N_10183);
and U10584 (N_10584,N_10422,N_10478);
nand U10585 (N_10585,N_10378,N_10248);
or U10586 (N_10586,N_10138,N_10145);
nand U10587 (N_10587,N_10013,N_10035);
and U10588 (N_10588,N_10255,N_10045);
xor U10589 (N_10589,N_10099,N_10104);
nor U10590 (N_10590,N_10370,N_10038);
nand U10591 (N_10591,N_10052,N_10219);
nor U10592 (N_10592,N_10202,N_10268);
nand U10593 (N_10593,N_10048,N_10454);
and U10594 (N_10594,N_10114,N_10331);
nand U10595 (N_10595,N_10312,N_10374);
or U10596 (N_10596,N_10237,N_10166);
and U10597 (N_10597,N_10488,N_10140);
or U10598 (N_10598,N_10392,N_10164);
nand U10599 (N_10599,N_10092,N_10209);
and U10600 (N_10600,N_10133,N_10355);
nand U10601 (N_10601,N_10037,N_10000);
or U10602 (N_10602,N_10107,N_10230);
nand U10603 (N_10603,N_10086,N_10152);
nor U10604 (N_10604,N_10229,N_10483);
nor U10605 (N_10605,N_10193,N_10464);
nand U10606 (N_10606,N_10291,N_10336);
xnor U10607 (N_10607,N_10421,N_10240);
nor U10608 (N_10608,N_10020,N_10067);
or U10609 (N_10609,N_10247,N_10410);
or U10610 (N_10610,N_10056,N_10080);
or U10611 (N_10611,N_10073,N_10187);
xnor U10612 (N_10612,N_10443,N_10289);
or U10613 (N_10613,N_10429,N_10027);
or U10614 (N_10614,N_10155,N_10411);
nor U10615 (N_10615,N_10449,N_10089);
and U10616 (N_10616,N_10218,N_10437);
or U10617 (N_10617,N_10458,N_10087);
or U10618 (N_10618,N_10161,N_10095);
and U10619 (N_10619,N_10175,N_10031);
or U10620 (N_10620,N_10316,N_10466);
or U10621 (N_10621,N_10100,N_10063);
or U10622 (N_10622,N_10489,N_10069);
nor U10623 (N_10623,N_10469,N_10362);
nor U10624 (N_10624,N_10030,N_10351);
nand U10625 (N_10625,N_10345,N_10284);
and U10626 (N_10626,N_10295,N_10257);
nor U10627 (N_10627,N_10424,N_10018);
nor U10628 (N_10628,N_10010,N_10032);
nand U10629 (N_10629,N_10430,N_10314);
nor U10630 (N_10630,N_10496,N_10366);
xor U10631 (N_10631,N_10185,N_10354);
and U10632 (N_10632,N_10231,N_10153);
and U10633 (N_10633,N_10397,N_10334);
xor U10634 (N_10634,N_10118,N_10444);
xor U10635 (N_10635,N_10486,N_10179);
or U10636 (N_10636,N_10071,N_10139);
or U10637 (N_10637,N_10226,N_10447);
xor U10638 (N_10638,N_10085,N_10084);
nor U10639 (N_10639,N_10451,N_10007);
nor U10640 (N_10640,N_10340,N_10364);
and U10641 (N_10641,N_10015,N_10129);
nand U10642 (N_10642,N_10046,N_10243);
and U10643 (N_10643,N_10485,N_10348);
nor U10644 (N_10644,N_10338,N_10082);
and U10645 (N_10645,N_10276,N_10207);
nor U10646 (N_10646,N_10033,N_10305);
nand U10647 (N_10647,N_10190,N_10431);
and U10648 (N_10648,N_10146,N_10124);
nor U10649 (N_10649,N_10251,N_10103);
nand U10650 (N_10650,N_10163,N_10271);
nand U10651 (N_10651,N_10049,N_10414);
and U10652 (N_10652,N_10270,N_10311);
nor U10653 (N_10653,N_10074,N_10324);
and U10654 (N_10654,N_10369,N_10241);
nand U10655 (N_10655,N_10256,N_10440);
or U10656 (N_10656,N_10228,N_10293);
nand U10657 (N_10657,N_10021,N_10066);
nand U10658 (N_10658,N_10427,N_10405);
nand U10659 (N_10659,N_10330,N_10003);
nand U10660 (N_10660,N_10036,N_10235);
or U10661 (N_10661,N_10157,N_10480);
or U10662 (N_10662,N_10189,N_10307);
nand U10663 (N_10663,N_10497,N_10353);
or U10664 (N_10664,N_10008,N_10042);
and U10665 (N_10665,N_10208,N_10455);
and U10666 (N_10666,N_10194,N_10322);
and U10667 (N_10667,N_10055,N_10313);
and U10668 (N_10668,N_10068,N_10323);
and U10669 (N_10669,N_10326,N_10280);
nand U10670 (N_10670,N_10343,N_10211);
nor U10671 (N_10671,N_10376,N_10337);
xor U10672 (N_10672,N_10057,N_10359);
nor U10673 (N_10673,N_10439,N_10453);
nand U10674 (N_10674,N_10093,N_10160);
nor U10675 (N_10675,N_10132,N_10304);
and U10676 (N_10676,N_10383,N_10490);
nand U10677 (N_10677,N_10158,N_10176);
or U10678 (N_10678,N_10022,N_10465);
nand U10679 (N_10679,N_10266,N_10325);
or U10680 (N_10680,N_10171,N_10356);
nand U10681 (N_10681,N_10141,N_10040);
nand U10682 (N_10682,N_10154,N_10418);
nand U10683 (N_10683,N_10200,N_10456);
nand U10684 (N_10684,N_10254,N_10134);
nand U10685 (N_10685,N_10128,N_10368);
and U10686 (N_10686,N_10263,N_10462);
and U10687 (N_10687,N_10119,N_10287);
xnor U10688 (N_10688,N_10292,N_10088);
and U10689 (N_10689,N_10415,N_10434);
nor U10690 (N_10690,N_10135,N_10181);
nand U10691 (N_10691,N_10012,N_10223);
and U10692 (N_10692,N_10147,N_10413);
nand U10693 (N_10693,N_10259,N_10306);
nor U10694 (N_10694,N_10023,N_10373);
nor U10695 (N_10695,N_10109,N_10065);
and U10696 (N_10696,N_10448,N_10406);
or U10697 (N_10697,N_10197,N_10039);
nor U10698 (N_10698,N_10210,N_10428);
nor U10699 (N_10699,N_10024,N_10299);
or U10700 (N_10700,N_10079,N_10380);
or U10701 (N_10701,N_10290,N_10387);
nor U10702 (N_10702,N_10432,N_10425);
nand U10703 (N_10703,N_10479,N_10258);
nor U10704 (N_10704,N_10321,N_10174);
nand U10705 (N_10705,N_10232,N_10319);
nand U10706 (N_10706,N_10159,N_10471);
nand U10707 (N_10707,N_10473,N_10167);
and U10708 (N_10708,N_10178,N_10463);
nor U10709 (N_10709,N_10170,N_10352);
nand U10710 (N_10710,N_10078,N_10365);
and U10711 (N_10711,N_10401,N_10244);
and U10712 (N_10712,N_10064,N_10442);
and U10713 (N_10713,N_10213,N_10225);
xnor U10714 (N_10714,N_10239,N_10412);
nand U10715 (N_10715,N_10409,N_10034);
or U10716 (N_10716,N_10494,N_10357);
and U10717 (N_10717,N_10162,N_10173);
nor U10718 (N_10718,N_10423,N_10267);
or U10719 (N_10719,N_10019,N_10300);
nor U10720 (N_10720,N_10391,N_10487);
or U10721 (N_10721,N_10206,N_10252);
nor U10722 (N_10722,N_10377,N_10372);
or U10723 (N_10723,N_10110,N_10214);
or U10724 (N_10724,N_10277,N_10234);
nor U10725 (N_10725,N_10393,N_10477);
or U10726 (N_10726,N_10054,N_10156);
nor U10727 (N_10727,N_10286,N_10285);
and U10728 (N_10728,N_10222,N_10327);
nand U10729 (N_10729,N_10375,N_10420);
or U10730 (N_10730,N_10363,N_10446);
or U10731 (N_10731,N_10265,N_10072);
nand U10732 (N_10732,N_10367,N_10062);
or U10733 (N_10733,N_10180,N_10402);
nand U10734 (N_10734,N_10221,N_10493);
and U10735 (N_10735,N_10385,N_10090);
nor U10736 (N_10736,N_10142,N_10246);
and U10737 (N_10737,N_10186,N_10445);
nor U10738 (N_10738,N_10105,N_10398);
or U10739 (N_10739,N_10111,N_10282);
and U10740 (N_10740,N_10433,N_10309);
xor U10741 (N_10741,N_10403,N_10004);
nand U10742 (N_10742,N_10061,N_10091);
and U10743 (N_10743,N_10098,N_10297);
nor U10744 (N_10744,N_10201,N_10315);
nor U10745 (N_10745,N_10491,N_10499);
nor U10746 (N_10746,N_10384,N_10136);
and U10747 (N_10747,N_10358,N_10332);
nor U10748 (N_10748,N_10273,N_10177);
nor U10749 (N_10749,N_10044,N_10317);
or U10750 (N_10750,N_10215,N_10106);
nor U10751 (N_10751,N_10429,N_10088);
and U10752 (N_10752,N_10313,N_10196);
nor U10753 (N_10753,N_10192,N_10120);
nand U10754 (N_10754,N_10466,N_10358);
nor U10755 (N_10755,N_10186,N_10054);
nand U10756 (N_10756,N_10491,N_10060);
and U10757 (N_10757,N_10170,N_10052);
and U10758 (N_10758,N_10063,N_10273);
and U10759 (N_10759,N_10074,N_10441);
nor U10760 (N_10760,N_10433,N_10138);
or U10761 (N_10761,N_10389,N_10250);
and U10762 (N_10762,N_10017,N_10171);
and U10763 (N_10763,N_10419,N_10149);
nand U10764 (N_10764,N_10449,N_10494);
and U10765 (N_10765,N_10333,N_10052);
nand U10766 (N_10766,N_10120,N_10410);
nand U10767 (N_10767,N_10309,N_10036);
and U10768 (N_10768,N_10090,N_10449);
nor U10769 (N_10769,N_10228,N_10215);
or U10770 (N_10770,N_10035,N_10348);
and U10771 (N_10771,N_10050,N_10190);
nor U10772 (N_10772,N_10227,N_10316);
xor U10773 (N_10773,N_10010,N_10215);
nand U10774 (N_10774,N_10097,N_10168);
nor U10775 (N_10775,N_10315,N_10183);
nand U10776 (N_10776,N_10214,N_10207);
nor U10777 (N_10777,N_10405,N_10384);
xor U10778 (N_10778,N_10248,N_10359);
nor U10779 (N_10779,N_10300,N_10087);
and U10780 (N_10780,N_10342,N_10048);
nand U10781 (N_10781,N_10116,N_10312);
or U10782 (N_10782,N_10177,N_10480);
or U10783 (N_10783,N_10122,N_10079);
and U10784 (N_10784,N_10326,N_10357);
or U10785 (N_10785,N_10179,N_10283);
nor U10786 (N_10786,N_10371,N_10490);
and U10787 (N_10787,N_10048,N_10246);
or U10788 (N_10788,N_10331,N_10110);
nand U10789 (N_10789,N_10013,N_10164);
nor U10790 (N_10790,N_10395,N_10030);
or U10791 (N_10791,N_10254,N_10384);
or U10792 (N_10792,N_10419,N_10353);
nand U10793 (N_10793,N_10457,N_10336);
nor U10794 (N_10794,N_10080,N_10427);
and U10795 (N_10795,N_10361,N_10152);
and U10796 (N_10796,N_10459,N_10407);
or U10797 (N_10797,N_10149,N_10405);
xnor U10798 (N_10798,N_10358,N_10225);
and U10799 (N_10799,N_10394,N_10164);
nor U10800 (N_10800,N_10411,N_10096);
xor U10801 (N_10801,N_10409,N_10411);
nand U10802 (N_10802,N_10346,N_10277);
nand U10803 (N_10803,N_10142,N_10092);
or U10804 (N_10804,N_10044,N_10123);
and U10805 (N_10805,N_10270,N_10222);
nor U10806 (N_10806,N_10095,N_10423);
or U10807 (N_10807,N_10494,N_10066);
and U10808 (N_10808,N_10164,N_10111);
nand U10809 (N_10809,N_10177,N_10170);
nor U10810 (N_10810,N_10308,N_10443);
and U10811 (N_10811,N_10186,N_10288);
nand U10812 (N_10812,N_10313,N_10229);
and U10813 (N_10813,N_10205,N_10351);
nor U10814 (N_10814,N_10014,N_10143);
or U10815 (N_10815,N_10110,N_10064);
or U10816 (N_10816,N_10169,N_10413);
or U10817 (N_10817,N_10386,N_10191);
or U10818 (N_10818,N_10021,N_10476);
nand U10819 (N_10819,N_10258,N_10034);
nand U10820 (N_10820,N_10090,N_10082);
or U10821 (N_10821,N_10350,N_10433);
or U10822 (N_10822,N_10200,N_10092);
or U10823 (N_10823,N_10006,N_10327);
or U10824 (N_10824,N_10486,N_10395);
or U10825 (N_10825,N_10336,N_10447);
and U10826 (N_10826,N_10495,N_10259);
and U10827 (N_10827,N_10042,N_10401);
nand U10828 (N_10828,N_10110,N_10206);
and U10829 (N_10829,N_10478,N_10369);
nor U10830 (N_10830,N_10015,N_10108);
nor U10831 (N_10831,N_10150,N_10046);
or U10832 (N_10832,N_10104,N_10253);
or U10833 (N_10833,N_10253,N_10380);
or U10834 (N_10834,N_10255,N_10100);
nand U10835 (N_10835,N_10376,N_10189);
nor U10836 (N_10836,N_10236,N_10054);
nand U10837 (N_10837,N_10015,N_10433);
nand U10838 (N_10838,N_10143,N_10313);
nor U10839 (N_10839,N_10072,N_10007);
or U10840 (N_10840,N_10220,N_10258);
nor U10841 (N_10841,N_10273,N_10048);
or U10842 (N_10842,N_10021,N_10254);
nor U10843 (N_10843,N_10435,N_10021);
and U10844 (N_10844,N_10078,N_10037);
or U10845 (N_10845,N_10182,N_10372);
nand U10846 (N_10846,N_10296,N_10434);
nand U10847 (N_10847,N_10019,N_10284);
nand U10848 (N_10848,N_10412,N_10068);
and U10849 (N_10849,N_10178,N_10088);
nor U10850 (N_10850,N_10225,N_10041);
and U10851 (N_10851,N_10138,N_10300);
or U10852 (N_10852,N_10105,N_10234);
and U10853 (N_10853,N_10322,N_10440);
and U10854 (N_10854,N_10004,N_10014);
or U10855 (N_10855,N_10400,N_10438);
nand U10856 (N_10856,N_10134,N_10393);
and U10857 (N_10857,N_10102,N_10042);
nand U10858 (N_10858,N_10318,N_10230);
nor U10859 (N_10859,N_10293,N_10449);
nand U10860 (N_10860,N_10002,N_10322);
or U10861 (N_10861,N_10330,N_10168);
nand U10862 (N_10862,N_10186,N_10350);
nor U10863 (N_10863,N_10265,N_10407);
and U10864 (N_10864,N_10224,N_10307);
and U10865 (N_10865,N_10349,N_10324);
nand U10866 (N_10866,N_10166,N_10167);
or U10867 (N_10867,N_10392,N_10049);
and U10868 (N_10868,N_10244,N_10420);
nor U10869 (N_10869,N_10291,N_10419);
nand U10870 (N_10870,N_10420,N_10409);
or U10871 (N_10871,N_10293,N_10292);
nor U10872 (N_10872,N_10082,N_10178);
nor U10873 (N_10873,N_10029,N_10206);
and U10874 (N_10874,N_10162,N_10286);
nand U10875 (N_10875,N_10090,N_10119);
nand U10876 (N_10876,N_10100,N_10404);
nand U10877 (N_10877,N_10193,N_10142);
and U10878 (N_10878,N_10229,N_10212);
nand U10879 (N_10879,N_10498,N_10232);
or U10880 (N_10880,N_10386,N_10496);
nor U10881 (N_10881,N_10494,N_10097);
nor U10882 (N_10882,N_10358,N_10080);
nor U10883 (N_10883,N_10274,N_10318);
and U10884 (N_10884,N_10273,N_10054);
nor U10885 (N_10885,N_10057,N_10177);
and U10886 (N_10886,N_10132,N_10341);
or U10887 (N_10887,N_10243,N_10210);
nor U10888 (N_10888,N_10007,N_10425);
and U10889 (N_10889,N_10081,N_10352);
and U10890 (N_10890,N_10222,N_10091);
and U10891 (N_10891,N_10093,N_10237);
or U10892 (N_10892,N_10376,N_10330);
or U10893 (N_10893,N_10219,N_10479);
or U10894 (N_10894,N_10073,N_10207);
nor U10895 (N_10895,N_10156,N_10256);
nand U10896 (N_10896,N_10195,N_10047);
and U10897 (N_10897,N_10069,N_10106);
xnor U10898 (N_10898,N_10107,N_10495);
or U10899 (N_10899,N_10160,N_10021);
nand U10900 (N_10900,N_10308,N_10234);
or U10901 (N_10901,N_10335,N_10442);
and U10902 (N_10902,N_10080,N_10127);
and U10903 (N_10903,N_10191,N_10018);
nand U10904 (N_10904,N_10181,N_10323);
nand U10905 (N_10905,N_10360,N_10079);
nor U10906 (N_10906,N_10249,N_10453);
or U10907 (N_10907,N_10315,N_10343);
or U10908 (N_10908,N_10318,N_10103);
nand U10909 (N_10909,N_10475,N_10266);
or U10910 (N_10910,N_10081,N_10338);
nand U10911 (N_10911,N_10072,N_10159);
and U10912 (N_10912,N_10145,N_10237);
nand U10913 (N_10913,N_10387,N_10147);
nor U10914 (N_10914,N_10061,N_10498);
nor U10915 (N_10915,N_10097,N_10203);
nand U10916 (N_10916,N_10212,N_10006);
nand U10917 (N_10917,N_10212,N_10140);
or U10918 (N_10918,N_10490,N_10014);
or U10919 (N_10919,N_10020,N_10057);
or U10920 (N_10920,N_10346,N_10137);
nor U10921 (N_10921,N_10276,N_10268);
nand U10922 (N_10922,N_10012,N_10268);
and U10923 (N_10923,N_10142,N_10397);
nor U10924 (N_10924,N_10433,N_10394);
nor U10925 (N_10925,N_10057,N_10056);
or U10926 (N_10926,N_10145,N_10124);
or U10927 (N_10927,N_10267,N_10459);
nand U10928 (N_10928,N_10347,N_10454);
nand U10929 (N_10929,N_10084,N_10280);
nand U10930 (N_10930,N_10284,N_10221);
nand U10931 (N_10931,N_10054,N_10376);
and U10932 (N_10932,N_10063,N_10133);
nand U10933 (N_10933,N_10355,N_10286);
and U10934 (N_10934,N_10311,N_10472);
nand U10935 (N_10935,N_10246,N_10457);
and U10936 (N_10936,N_10062,N_10043);
nand U10937 (N_10937,N_10299,N_10395);
or U10938 (N_10938,N_10146,N_10375);
or U10939 (N_10939,N_10448,N_10394);
and U10940 (N_10940,N_10263,N_10168);
and U10941 (N_10941,N_10077,N_10472);
nand U10942 (N_10942,N_10406,N_10269);
and U10943 (N_10943,N_10433,N_10379);
nor U10944 (N_10944,N_10241,N_10448);
nor U10945 (N_10945,N_10277,N_10006);
nand U10946 (N_10946,N_10284,N_10247);
and U10947 (N_10947,N_10322,N_10476);
and U10948 (N_10948,N_10179,N_10245);
nand U10949 (N_10949,N_10243,N_10309);
xor U10950 (N_10950,N_10458,N_10079);
or U10951 (N_10951,N_10034,N_10287);
and U10952 (N_10952,N_10220,N_10070);
and U10953 (N_10953,N_10259,N_10261);
nor U10954 (N_10954,N_10460,N_10481);
or U10955 (N_10955,N_10215,N_10499);
nor U10956 (N_10956,N_10018,N_10415);
or U10957 (N_10957,N_10157,N_10484);
and U10958 (N_10958,N_10373,N_10001);
nand U10959 (N_10959,N_10189,N_10285);
nor U10960 (N_10960,N_10378,N_10214);
nand U10961 (N_10961,N_10443,N_10232);
or U10962 (N_10962,N_10110,N_10440);
nand U10963 (N_10963,N_10061,N_10423);
nor U10964 (N_10964,N_10176,N_10086);
and U10965 (N_10965,N_10192,N_10022);
and U10966 (N_10966,N_10382,N_10055);
or U10967 (N_10967,N_10494,N_10041);
or U10968 (N_10968,N_10115,N_10331);
nand U10969 (N_10969,N_10267,N_10307);
nor U10970 (N_10970,N_10295,N_10141);
nor U10971 (N_10971,N_10383,N_10161);
or U10972 (N_10972,N_10272,N_10435);
nor U10973 (N_10973,N_10202,N_10127);
and U10974 (N_10974,N_10187,N_10118);
or U10975 (N_10975,N_10184,N_10123);
and U10976 (N_10976,N_10403,N_10461);
nand U10977 (N_10977,N_10058,N_10082);
nand U10978 (N_10978,N_10002,N_10264);
and U10979 (N_10979,N_10260,N_10163);
or U10980 (N_10980,N_10325,N_10297);
nor U10981 (N_10981,N_10470,N_10251);
nor U10982 (N_10982,N_10140,N_10388);
and U10983 (N_10983,N_10256,N_10068);
nand U10984 (N_10984,N_10333,N_10355);
or U10985 (N_10985,N_10103,N_10082);
nand U10986 (N_10986,N_10074,N_10488);
nor U10987 (N_10987,N_10137,N_10332);
and U10988 (N_10988,N_10367,N_10419);
and U10989 (N_10989,N_10010,N_10080);
nand U10990 (N_10990,N_10454,N_10187);
nor U10991 (N_10991,N_10201,N_10388);
and U10992 (N_10992,N_10417,N_10496);
nand U10993 (N_10993,N_10290,N_10275);
or U10994 (N_10994,N_10095,N_10192);
and U10995 (N_10995,N_10396,N_10426);
nor U10996 (N_10996,N_10465,N_10304);
and U10997 (N_10997,N_10143,N_10362);
xor U10998 (N_10998,N_10381,N_10060);
or U10999 (N_10999,N_10439,N_10342);
and U11000 (N_11000,N_10633,N_10988);
nand U11001 (N_11001,N_10514,N_10709);
nor U11002 (N_11002,N_10939,N_10547);
nand U11003 (N_11003,N_10665,N_10906);
nand U11004 (N_11004,N_10756,N_10559);
nand U11005 (N_11005,N_10673,N_10824);
nor U11006 (N_11006,N_10802,N_10664);
or U11007 (N_11007,N_10975,N_10923);
nor U11008 (N_11008,N_10517,N_10875);
nand U11009 (N_11009,N_10831,N_10896);
nand U11010 (N_11010,N_10555,N_10880);
nand U11011 (N_11011,N_10606,N_10783);
nand U11012 (N_11012,N_10786,N_10674);
nand U11013 (N_11013,N_10767,N_10803);
nand U11014 (N_11014,N_10602,N_10582);
and U11015 (N_11015,N_10693,N_10640);
nor U11016 (N_11016,N_10937,N_10926);
or U11017 (N_11017,N_10535,N_10741);
and U11018 (N_11018,N_10849,N_10727);
or U11019 (N_11019,N_10779,N_10776);
and U11020 (N_11020,N_10591,N_10903);
and U11021 (N_11021,N_10945,N_10502);
nor U11022 (N_11022,N_10688,N_10782);
or U11023 (N_11023,N_10639,N_10840);
nor U11024 (N_11024,N_10877,N_10548);
or U11025 (N_11025,N_10611,N_10984);
nand U11026 (N_11026,N_10768,N_10683);
nand U11027 (N_11027,N_10809,N_10750);
nor U11028 (N_11028,N_10503,N_10949);
or U11029 (N_11029,N_10520,N_10560);
or U11030 (N_11030,N_10960,N_10533);
or U11031 (N_11031,N_10852,N_10554);
nor U11032 (N_11032,N_10881,N_10909);
nor U11033 (N_11033,N_10543,N_10738);
nor U11034 (N_11034,N_10842,N_10597);
or U11035 (N_11035,N_10653,N_10626);
and U11036 (N_11036,N_10759,N_10793);
nand U11037 (N_11037,N_10947,N_10836);
or U11038 (N_11038,N_10961,N_10980);
nand U11039 (N_11039,N_10792,N_10825);
and U11040 (N_11040,N_10858,N_10883);
nor U11041 (N_11041,N_10837,N_10821);
nor U11042 (N_11042,N_10922,N_10609);
and U11043 (N_11043,N_10715,N_10734);
or U11044 (N_11044,N_10652,N_10585);
nand U11045 (N_11045,N_10718,N_10890);
or U11046 (N_11046,N_10619,N_10780);
nand U11047 (N_11047,N_10931,N_10695);
and U11048 (N_11048,N_10642,N_10868);
or U11049 (N_11049,N_10904,N_10967);
nor U11050 (N_11050,N_10704,N_10889);
nor U11051 (N_11051,N_10789,N_10726);
nor U11052 (N_11052,N_10509,N_10919);
nand U11053 (N_11053,N_10616,N_10818);
or U11054 (N_11054,N_10798,N_10747);
nor U11055 (N_11055,N_10743,N_10932);
and U11056 (N_11056,N_10971,N_10927);
and U11057 (N_11057,N_10970,N_10964);
nand U11058 (N_11058,N_10902,N_10826);
or U11059 (N_11059,N_10636,N_10784);
nor U11060 (N_11060,N_10617,N_10615);
or U11061 (N_11061,N_10605,N_10807);
or U11062 (N_11062,N_10815,N_10518);
and U11063 (N_11063,N_10530,N_10590);
and U11064 (N_11064,N_10536,N_10879);
nand U11065 (N_11065,N_10834,N_10714);
nand U11066 (N_11066,N_10552,N_10913);
nor U11067 (N_11067,N_10671,N_10812);
nand U11068 (N_11068,N_10746,N_10978);
and U11069 (N_11069,N_10878,N_10655);
nor U11070 (N_11070,N_10788,N_10706);
nor U11071 (N_11071,N_10504,N_10568);
nor U11072 (N_11072,N_10928,N_10887);
nor U11073 (N_11073,N_10647,N_10992);
or U11074 (N_11074,N_10716,N_10696);
nor U11075 (N_11075,N_10675,N_10733);
nand U11076 (N_11076,N_10659,N_10774);
nand U11077 (N_11077,N_10566,N_10833);
or U11078 (N_11078,N_10730,N_10843);
nor U11079 (N_11079,N_10524,N_10965);
nor U11080 (N_11080,N_10613,N_10565);
nand U11081 (N_11081,N_10894,N_10791);
xnor U11082 (N_11082,N_10999,N_10805);
nor U11083 (N_11083,N_10711,N_10884);
and U11084 (N_11084,N_10827,N_10736);
nor U11085 (N_11085,N_10943,N_10893);
nor U11086 (N_11086,N_10863,N_10583);
or U11087 (N_11087,N_10771,N_10562);
or U11088 (N_11088,N_10513,N_10853);
nand U11089 (N_11089,N_10628,N_10669);
or U11090 (N_11090,N_10822,N_10512);
nand U11091 (N_11091,N_10963,N_10646);
xor U11092 (N_11092,N_10627,N_10526);
xnor U11093 (N_11093,N_10620,N_10869);
nor U11094 (N_11094,N_10731,N_10740);
and U11095 (N_11095,N_10685,N_10510);
nand U11096 (N_11096,N_10871,N_10629);
nor U11097 (N_11097,N_10592,N_10921);
or U11098 (N_11098,N_10918,N_10643);
or U11099 (N_11099,N_10765,N_10761);
nand U11100 (N_11100,N_10755,N_10800);
or U11101 (N_11101,N_10787,N_10811);
nor U11102 (N_11102,N_10556,N_10850);
nand U11103 (N_11103,N_10691,N_10569);
and U11104 (N_11104,N_10682,N_10694);
and U11105 (N_11105,N_10933,N_10969);
and U11106 (N_11106,N_10816,N_10703);
nand U11107 (N_11107,N_10546,N_10575);
or U11108 (N_11108,N_10985,N_10845);
nor U11109 (N_11109,N_10766,N_10678);
or U11110 (N_11110,N_10580,N_10550);
xor U11111 (N_11111,N_10672,N_10966);
nor U11112 (N_11112,N_10942,N_10534);
nor U11113 (N_11113,N_10676,N_10995);
nand U11114 (N_11114,N_10707,N_10697);
nand U11115 (N_11115,N_10680,N_10956);
and U11116 (N_11116,N_10832,N_10855);
nand U11117 (N_11117,N_10873,N_10705);
nor U11118 (N_11118,N_10870,N_10677);
nand U11119 (N_11119,N_10660,N_10857);
nor U11120 (N_11120,N_10977,N_10814);
nand U11121 (N_11121,N_10915,N_10544);
nor U11122 (N_11122,N_10573,N_10618);
and U11123 (N_11123,N_10872,N_10522);
nor U11124 (N_11124,N_10912,N_10631);
or U11125 (N_11125,N_10772,N_10981);
nand U11126 (N_11126,N_10581,N_10936);
and U11127 (N_11127,N_10684,N_10935);
nor U11128 (N_11128,N_10621,N_10925);
or U11129 (N_11129,N_10770,N_10957);
nor U11130 (N_11130,N_10892,N_10905);
nor U11131 (N_11131,N_10844,N_10940);
nor U11132 (N_11132,N_10701,N_10724);
nand U11133 (N_11133,N_10846,N_10690);
xnor U11134 (N_11134,N_10588,N_10866);
nor U11135 (N_11135,N_10570,N_10594);
and U11136 (N_11136,N_10601,N_10589);
nand U11137 (N_11137,N_10593,N_10819);
or U11138 (N_11138,N_10641,N_10763);
and U11139 (N_11139,N_10865,N_10542);
or U11140 (N_11140,N_10523,N_10700);
nand U11141 (N_11141,N_10951,N_10861);
nand U11142 (N_11142,N_10571,N_10668);
nor U11143 (N_11143,N_10994,N_10507);
or U11144 (N_11144,N_10917,N_10976);
or U11145 (N_11145,N_10598,N_10799);
nor U11146 (N_11146,N_10501,N_10658);
nand U11147 (N_11147,N_10910,N_10895);
xnor U11148 (N_11148,N_10528,N_10525);
xor U11149 (N_11149,N_10998,N_10929);
and U11150 (N_11150,N_10962,N_10508);
and U11151 (N_11151,N_10720,N_10721);
or U11152 (N_11152,N_10993,N_10948);
nor U11153 (N_11153,N_10713,N_10996);
or U11154 (N_11154,N_10670,N_10661);
or U11155 (N_11155,N_10952,N_10710);
or U11156 (N_11156,N_10778,N_10614);
nor U11157 (N_11157,N_10924,N_10564);
nand U11158 (N_11158,N_10773,N_10649);
nor U11159 (N_11159,N_10644,N_10603);
and U11160 (N_11160,N_10986,N_10859);
nor U11161 (N_11161,N_10775,N_10801);
and U11162 (N_11162,N_10916,N_10539);
and U11163 (N_11163,N_10867,N_10891);
nand U11164 (N_11164,N_10579,N_10898);
nor U11165 (N_11165,N_10930,N_10541);
nand U11166 (N_11166,N_10578,N_10717);
or U11167 (N_11167,N_10900,N_10654);
and U11168 (N_11168,N_10864,N_10797);
nor U11169 (N_11169,N_10595,N_10735);
nor U11170 (N_11170,N_10862,N_10612);
xor U11171 (N_11171,N_10681,N_10607);
nand U11172 (N_11172,N_10886,N_10972);
or U11173 (N_11173,N_10702,N_10838);
and U11174 (N_11174,N_10604,N_10723);
nor U11175 (N_11175,N_10830,N_10848);
or U11176 (N_11176,N_10532,N_10897);
nand U11177 (N_11177,N_10656,N_10666);
nand U11178 (N_11178,N_10551,N_10820);
nor U11179 (N_11179,N_10973,N_10645);
or U11180 (N_11180,N_10739,N_10529);
and U11181 (N_11181,N_10692,N_10899);
or U11182 (N_11182,N_10549,N_10794);
or U11183 (N_11183,N_10637,N_10987);
nor U11184 (N_11184,N_10608,N_10856);
or U11185 (N_11185,N_10625,N_10990);
and U11186 (N_11186,N_10781,N_10982);
and U11187 (N_11187,N_10650,N_10835);
nor U11188 (N_11188,N_10908,N_10806);
nand U11189 (N_11189,N_10531,N_10979);
and U11190 (N_11190,N_10938,N_10795);
and U11191 (N_11191,N_10829,N_10689);
and U11192 (N_11192,N_10920,N_10584);
nand U11193 (N_11193,N_10632,N_10847);
nand U11194 (N_11194,N_10828,N_10860);
and U11195 (N_11195,N_10997,N_10553);
or U11196 (N_11196,N_10959,N_10744);
nand U11197 (N_11197,N_10785,N_10732);
or U11198 (N_11198,N_10648,N_10708);
nor U11199 (N_11199,N_10914,N_10762);
and U11200 (N_11200,N_10558,N_10989);
nor U11201 (N_11201,N_10624,N_10599);
and U11202 (N_11202,N_10941,N_10561);
or U11203 (N_11203,N_10634,N_10841);
xor U11204 (N_11204,N_10752,N_10769);
or U11205 (N_11205,N_10719,N_10729);
nor U11206 (N_11206,N_10622,N_10753);
or U11207 (N_11207,N_10823,N_10687);
nor U11208 (N_11208,N_10817,N_10728);
or U11209 (N_11209,N_10586,N_10725);
nor U11210 (N_11210,N_10574,N_10662);
nand U11211 (N_11211,N_10538,N_10983);
or U11212 (N_11212,N_10698,N_10950);
nand U11213 (N_11213,N_10748,N_10667);
and U11214 (N_11214,N_10777,N_10623);
or U11215 (N_11215,N_10519,N_10511);
nand U11216 (N_11216,N_10790,N_10888);
nand U11217 (N_11217,N_10737,N_10630);
and U11218 (N_11218,N_10567,N_10934);
nand U11219 (N_11219,N_10563,N_10635);
or U11220 (N_11220,N_10610,N_10953);
nand U11221 (N_11221,N_10946,N_10749);
nor U11222 (N_11222,N_10958,N_10954);
nand U11223 (N_11223,N_10663,N_10577);
nor U11224 (N_11224,N_10882,N_10540);
nand U11225 (N_11225,N_10907,N_10796);
nor U11226 (N_11226,N_10712,N_10751);
nand U11227 (N_11227,N_10991,N_10760);
nand U11228 (N_11228,N_10506,N_10587);
or U11229 (N_11229,N_10516,N_10657);
nand U11230 (N_11230,N_10521,N_10974);
or U11231 (N_11231,N_10885,N_10876);
and U11232 (N_11232,N_10505,N_10851);
or U11233 (N_11233,N_10742,N_10600);
and U11234 (N_11234,N_10810,N_10968);
nand U11235 (N_11235,N_10537,N_10839);
nor U11236 (N_11236,N_10596,N_10754);
or U11237 (N_11237,N_10679,N_10874);
or U11238 (N_11238,N_10808,N_10557);
or U11239 (N_11239,N_10651,N_10638);
nor U11240 (N_11240,N_10901,N_10515);
nand U11241 (N_11241,N_10944,N_10955);
nand U11242 (N_11242,N_10745,N_10527);
nor U11243 (N_11243,N_10764,N_10911);
nand U11244 (N_11244,N_10576,N_10500);
nand U11245 (N_11245,N_10758,N_10686);
or U11246 (N_11246,N_10722,N_10757);
and U11247 (N_11247,N_10804,N_10545);
nor U11248 (N_11248,N_10699,N_10572);
nand U11249 (N_11249,N_10854,N_10813);
nor U11250 (N_11250,N_10770,N_10776);
nand U11251 (N_11251,N_10696,N_10704);
or U11252 (N_11252,N_10927,N_10957);
or U11253 (N_11253,N_10695,N_10794);
or U11254 (N_11254,N_10680,N_10734);
or U11255 (N_11255,N_10835,N_10719);
and U11256 (N_11256,N_10822,N_10505);
and U11257 (N_11257,N_10903,N_10588);
nand U11258 (N_11258,N_10911,N_10527);
or U11259 (N_11259,N_10515,N_10764);
nand U11260 (N_11260,N_10717,N_10783);
and U11261 (N_11261,N_10866,N_10917);
xor U11262 (N_11262,N_10994,N_10575);
nor U11263 (N_11263,N_10872,N_10859);
xnor U11264 (N_11264,N_10728,N_10888);
nand U11265 (N_11265,N_10949,N_10780);
and U11266 (N_11266,N_10789,N_10698);
nor U11267 (N_11267,N_10665,N_10754);
and U11268 (N_11268,N_10943,N_10561);
and U11269 (N_11269,N_10811,N_10887);
or U11270 (N_11270,N_10642,N_10736);
nand U11271 (N_11271,N_10631,N_10781);
and U11272 (N_11272,N_10871,N_10897);
and U11273 (N_11273,N_10693,N_10975);
or U11274 (N_11274,N_10528,N_10910);
or U11275 (N_11275,N_10858,N_10714);
nor U11276 (N_11276,N_10691,N_10560);
nand U11277 (N_11277,N_10836,N_10691);
and U11278 (N_11278,N_10576,N_10928);
nor U11279 (N_11279,N_10705,N_10837);
nor U11280 (N_11280,N_10938,N_10930);
and U11281 (N_11281,N_10954,N_10530);
and U11282 (N_11282,N_10872,N_10575);
nor U11283 (N_11283,N_10940,N_10744);
or U11284 (N_11284,N_10759,N_10792);
xor U11285 (N_11285,N_10662,N_10948);
and U11286 (N_11286,N_10960,N_10952);
and U11287 (N_11287,N_10847,N_10844);
and U11288 (N_11288,N_10994,N_10624);
and U11289 (N_11289,N_10926,N_10609);
and U11290 (N_11290,N_10970,N_10551);
and U11291 (N_11291,N_10560,N_10693);
and U11292 (N_11292,N_10819,N_10935);
nand U11293 (N_11293,N_10960,N_10780);
xor U11294 (N_11294,N_10879,N_10807);
nand U11295 (N_11295,N_10926,N_10694);
nand U11296 (N_11296,N_10719,N_10601);
nand U11297 (N_11297,N_10840,N_10996);
or U11298 (N_11298,N_10878,N_10949);
or U11299 (N_11299,N_10895,N_10810);
or U11300 (N_11300,N_10799,N_10989);
nor U11301 (N_11301,N_10559,N_10700);
and U11302 (N_11302,N_10738,N_10841);
nand U11303 (N_11303,N_10641,N_10706);
nand U11304 (N_11304,N_10502,N_10786);
nor U11305 (N_11305,N_10619,N_10787);
and U11306 (N_11306,N_10536,N_10694);
nor U11307 (N_11307,N_10505,N_10654);
or U11308 (N_11308,N_10599,N_10984);
nor U11309 (N_11309,N_10678,N_10634);
xnor U11310 (N_11310,N_10630,N_10802);
nand U11311 (N_11311,N_10507,N_10591);
nand U11312 (N_11312,N_10684,N_10529);
nand U11313 (N_11313,N_10680,N_10907);
and U11314 (N_11314,N_10827,N_10795);
and U11315 (N_11315,N_10976,N_10592);
nand U11316 (N_11316,N_10611,N_10607);
or U11317 (N_11317,N_10755,N_10846);
nand U11318 (N_11318,N_10903,N_10924);
nand U11319 (N_11319,N_10598,N_10795);
and U11320 (N_11320,N_10615,N_10805);
nand U11321 (N_11321,N_10637,N_10729);
nand U11322 (N_11322,N_10507,N_10631);
or U11323 (N_11323,N_10701,N_10515);
and U11324 (N_11324,N_10655,N_10824);
nand U11325 (N_11325,N_10830,N_10536);
nand U11326 (N_11326,N_10562,N_10598);
nor U11327 (N_11327,N_10584,N_10879);
nor U11328 (N_11328,N_10997,N_10656);
or U11329 (N_11329,N_10697,N_10747);
and U11330 (N_11330,N_10671,N_10866);
nand U11331 (N_11331,N_10672,N_10814);
nor U11332 (N_11332,N_10848,N_10838);
nand U11333 (N_11333,N_10588,N_10548);
nor U11334 (N_11334,N_10740,N_10558);
nand U11335 (N_11335,N_10772,N_10544);
nor U11336 (N_11336,N_10700,N_10724);
nor U11337 (N_11337,N_10875,N_10955);
or U11338 (N_11338,N_10783,N_10604);
and U11339 (N_11339,N_10915,N_10966);
and U11340 (N_11340,N_10776,N_10640);
nand U11341 (N_11341,N_10554,N_10538);
nor U11342 (N_11342,N_10526,N_10572);
nor U11343 (N_11343,N_10809,N_10709);
nand U11344 (N_11344,N_10652,N_10909);
and U11345 (N_11345,N_10946,N_10778);
nand U11346 (N_11346,N_10659,N_10723);
nor U11347 (N_11347,N_10665,N_10570);
and U11348 (N_11348,N_10693,N_10916);
xnor U11349 (N_11349,N_10561,N_10501);
nor U11350 (N_11350,N_10945,N_10737);
and U11351 (N_11351,N_10767,N_10808);
or U11352 (N_11352,N_10664,N_10624);
and U11353 (N_11353,N_10608,N_10914);
and U11354 (N_11354,N_10931,N_10563);
nor U11355 (N_11355,N_10732,N_10883);
nand U11356 (N_11356,N_10937,N_10998);
nand U11357 (N_11357,N_10574,N_10501);
nand U11358 (N_11358,N_10655,N_10906);
and U11359 (N_11359,N_10883,N_10957);
and U11360 (N_11360,N_10944,N_10937);
or U11361 (N_11361,N_10812,N_10876);
or U11362 (N_11362,N_10881,N_10938);
or U11363 (N_11363,N_10538,N_10911);
or U11364 (N_11364,N_10535,N_10774);
or U11365 (N_11365,N_10532,N_10992);
nor U11366 (N_11366,N_10908,N_10847);
nand U11367 (N_11367,N_10519,N_10753);
nor U11368 (N_11368,N_10700,N_10766);
and U11369 (N_11369,N_10741,N_10937);
nand U11370 (N_11370,N_10966,N_10563);
or U11371 (N_11371,N_10990,N_10610);
nand U11372 (N_11372,N_10821,N_10944);
or U11373 (N_11373,N_10877,N_10658);
and U11374 (N_11374,N_10563,N_10699);
and U11375 (N_11375,N_10541,N_10716);
and U11376 (N_11376,N_10508,N_10993);
nand U11377 (N_11377,N_10996,N_10933);
nand U11378 (N_11378,N_10964,N_10829);
and U11379 (N_11379,N_10796,N_10827);
nor U11380 (N_11380,N_10739,N_10518);
nand U11381 (N_11381,N_10806,N_10509);
or U11382 (N_11382,N_10945,N_10941);
nor U11383 (N_11383,N_10959,N_10954);
and U11384 (N_11384,N_10668,N_10817);
xor U11385 (N_11385,N_10820,N_10947);
nand U11386 (N_11386,N_10703,N_10968);
and U11387 (N_11387,N_10586,N_10548);
nor U11388 (N_11388,N_10803,N_10853);
and U11389 (N_11389,N_10617,N_10797);
nand U11390 (N_11390,N_10639,N_10663);
and U11391 (N_11391,N_10555,N_10669);
and U11392 (N_11392,N_10623,N_10587);
and U11393 (N_11393,N_10844,N_10956);
and U11394 (N_11394,N_10829,N_10515);
and U11395 (N_11395,N_10658,N_10920);
nand U11396 (N_11396,N_10775,N_10693);
or U11397 (N_11397,N_10548,N_10981);
nand U11398 (N_11398,N_10645,N_10633);
nand U11399 (N_11399,N_10529,N_10544);
nor U11400 (N_11400,N_10613,N_10642);
or U11401 (N_11401,N_10554,N_10726);
nand U11402 (N_11402,N_10815,N_10654);
nor U11403 (N_11403,N_10831,N_10792);
nor U11404 (N_11404,N_10745,N_10622);
nand U11405 (N_11405,N_10620,N_10914);
and U11406 (N_11406,N_10898,N_10667);
and U11407 (N_11407,N_10621,N_10909);
xnor U11408 (N_11408,N_10727,N_10609);
and U11409 (N_11409,N_10907,N_10533);
nor U11410 (N_11410,N_10592,N_10948);
or U11411 (N_11411,N_10834,N_10664);
or U11412 (N_11412,N_10675,N_10801);
or U11413 (N_11413,N_10847,N_10651);
nand U11414 (N_11414,N_10755,N_10892);
or U11415 (N_11415,N_10819,N_10848);
or U11416 (N_11416,N_10699,N_10956);
and U11417 (N_11417,N_10986,N_10572);
or U11418 (N_11418,N_10661,N_10751);
and U11419 (N_11419,N_10777,N_10744);
nor U11420 (N_11420,N_10892,N_10686);
nor U11421 (N_11421,N_10897,N_10668);
nor U11422 (N_11422,N_10553,N_10959);
nand U11423 (N_11423,N_10779,N_10532);
nor U11424 (N_11424,N_10850,N_10992);
nand U11425 (N_11425,N_10750,N_10967);
or U11426 (N_11426,N_10745,N_10676);
and U11427 (N_11427,N_10965,N_10533);
or U11428 (N_11428,N_10802,N_10548);
or U11429 (N_11429,N_10787,N_10962);
nand U11430 (N_11430,N_10586,N_10520);
nand U11431 (N_11431,N_10795,N_10908);
nand U11432 (N_11432,N_10749,N_10827);
or U11433 (N_11433,N_10717,N_10943);
or U11434 (N_11434,N_10682,N_10622);
and U11435 (N_11435,N_10912,N_10801);
or U11436 (N_11436,N_10524,N_10736);
and U11437 (N_11437,N_10856,N_10878);
nand U11438 (N_11438,N_10574,N_10603);
or U11439 (N_11439,N_10631,N_10536);
or U11440 (N_11440,N_10995,N_10610);
xor U11441 (N_11441,N_10794,N_10752);
and U11442 (N_11442,N_10840,N_10930);
nand U11443 (N_11443,N_10559,N_10644);
nand U11444 (N_11444,N_10824,N_10752);
nand U11445 (N_11445,N_10609,N_10643);
nor U11446 (N_11446,N_10576,N_10814);
or U11447 (N_11447,N_10686,N_10516);
and U11448 (N_11448,N_10993,N_10906);
and U11449 (N_11449,N_10590,N_10716);
nor U11450 (N_11450,N_10667,N_10752);
and U11451 (N_11451,N_10979,N_10713);
or U11452 (N_11452,N_10607,N_10898);
nand U11453 (N_11453,N_10994,N_10587);
and U11454 (N_11454,N_10538,N_10734);
nor U11455 (N_11455,N_10535,N_10711);
nand U11456 (N_11456,N_10854,N_10527);
or U11457 (N_11457,N_10929,N_10503);
nor U11458 (N_11458,N_10937,N_10943);
nor U11459 (N_11459,N_10863,N_10870);
nand U11460 (N_11460,N_10677,N_10795);
nand U11461 (N_11461,N_10792,N_10571);
nand U11462 (N_11462,N_10871,N_10734);
or U11463 (N_11463,N_10678,N_10890);
or U11464 (N_11464,N_10683,N_10766);
nand U11465 (N_11465,N_10702,N_10856);
nor U11466 (N_11466,N_10854,N_10715);
and U11467 (N_11467,N_10650,N_10984);
nand U11468 (N_11468,N_10748,N_10726);
or U11469 (N_11469,N_10810,N_10881);
and U11470 (N_11470,N_10602,N_10883);
or U11471 (N_11471,N_10990,N_10519);
and U11472 (N_11472,N_10645,N_10989);
nor U11473 (N_11473,N_10951,N_10556);
nor U11474 (N_11474,N_10931,N_10705);
and U11475 (N_11475,N_10819,N_10908);
nor U11476 (N_11476,N_10689,N_10996);
or U11477 (N_11477,N_10603,N_10512);
or U11478 (N_11478,N_10808,N_10674);
and U11479 (N_11479,N_10615,N_10804);
and U11480 (N_11480,N_10768,N_10902);
nor U11481 (N_11481,N_10764,N_10695);
xor U11482 (N_11482,N_10708,N_10908);
nor U11483 (N_11483,N_10958,N_10760);
nor U11484 (N_11484,N_10675,N_10604);
nand U11485 (N_11485,N_10666,N_10831);
xnor U11486 (N_11486,N_10631,N_10524);
or U11487 (N_11487,N_10698,N_10578);
nor U11488 (N_11488,N_10683,N_10881);
and U11489 (N_11489,N_10951,N_10692);
nand U11490 (N_11490,N_10687,N_10942);
nor U11491 (N_11491,N_10504,N_10724);
or U11492 (N_11492,N_10573,N_10622);
nor U11493 (N_11493,N_10652,N_10957);
nor U11494 (N_11494,N_10791,N_10992);
and U11495 (N_11495,N_10781,N_10844);
and U11496 (N_11496,N_10805,N_10575);
nor U11497 (N_11497,N_10697,N_10970);
nand U11498 (N_11498,N_10535,N_10987);
or U11499 (N_11499,N_10539,N_10966);
or U11500 (N_11500,N_11107,N_11137);
nand U11501 (N_11501,N_11344,N_11213);
or U11502 (N_11502,N_11279,N_11007);
and U11503 (N_11503,N_11413,N_11112);
or U11504 (N_11504,N_11399,N_11443);
or U11505 (N_11505,N_11187,N_11299);
nand U11506 (N_11506,N_11428,N_11166);
or U11507 (N_11507,N_11458,N_11357);
nand U11508 (N_11508,N_11421,N_11289);
nand U11509 (N_11509,N_11330,N_11026);
and U11510 (N_11510,N_11309,N_11093);
or U11511 (N_11511,N_11387,N_11483);
nor U11512 (N_11512,N_11047,N_11308);
nor U11513 (N_11513,N_11391,N_11262);
nand U11514 (N_11514,N_11392,N_11478);
or U11515 (N_11515,N_11046,N_11084);
and U11516 (N_11516,N_11304,N_11296);
or U11517 (N_11517,N_11172,N_11141);
or U11518 (N_11518,N_11003,N_11264);
nand U11519 (N_11519,N_11381,N_11200);
or U11520 (N_11520,N_11398,N_11063);
nand U11521 (N_11521,N_11044,N_11177);
xnor U11522 (N_11522,N_11179,N_11411);
nor U11523 (N_11523,N_11097,N_11088);
and U11524 (N_11524,N_11286,N_11184);
nand U11525 (N_11525,N_11131,N_11369);
nor U11526 (N_11526,N_11250,N_11336);
nand U11527 (N_11527,N_11120,N_11065);
and U11528 (N_11528,N_11104,N_11416);
nand U11529 (N_11529,N_11293,N_11454);
and U11530 (N_11530,N_11247,N_11307);
or U11531 (N_11531,N_11339,N_11487);
and U11532 (N_11532,N_11069,N_11477);
and U11533 (N_11533,N_11362,N_11110);
and U11534 (N_11534,N_11465,N_11189);
or U11535 (N_11535,N_11237,N_11356);
and U11536 (N_11536,N_11175,N_11291);
and U11537 (N_11537,N_11027,N_11319);
nand U11538 (N_11538,N_11019,N_11022);
nand U11539 (N_11539,N_11354,N_11129);
nor U11540 (N_11540,N_11052,N_11225);
and U11541 (N_11541,N_11002,N_11275);
and U11542 (N_11542,N_11091,N_11498);
nor U11543 (N_11543,N_11193,N_11371);
or U11544 (N_11544,N_11313,N_11431);
or U11545 (N_11545,N_11417,N_11033);
nand U11546 (N_11546,N_11375,N_11230);
nor U11547 (N_11547,N_11457,N_11248);
or U11548 (N_11548,N_11318,N_11292);
nor U11549 (N_11549,N_11464,N_11456);
or U11550 (N_11550,N_11281,N_11241);
nand U11551 (N_11551,N_11195,N_11364);
and U11552 (N_11552,N_11390,N_11143);
or U11553 (N_11553,N_11485,N_11316);
or U11554 (N_11554,N_11385,N_11178);
nand U11555 (N_11555,N_11395,N_11058);
nor U11556 (N_11556,N_11072,N_11315);
or U11557 (N_11557,N_11270,N_11089);
nor U11558 (N_11558,N_11102,N_11242);
or U11559 (N_11559,N_11243,N_11150);
nand U11560 (N_11560,N_11186,N_11015);
and U11561 (N_11561,N_11448,N_11438);
nor U11562 (N_11562,N_11071,N_11301);
nor U11563 (N_11563,N_11410,N_11139);
xnor U11564 (N_11564,N_11461,N_11087);
nand U11565 (N_11565,N_11174,N_11473);
or U11566 (N_11566,N_11401,N_11359);
nor U11567 (N_11567,N_11469,N_11476);
nor U11568 (N_11568,N_11310,N_11300);
or U11569 (N_11569,N_11155,N_11470);
or U11570 (N_11570,N_11060,N_11151);
and U11571 (N_11571,N_11018,N_11235);
or U11572 (N_11572,N_11266,N_11408);
and U11573 (N_11573,N_11445,N_11441);
or U11574 (N_11574,N_11467,N_11386);
nor U11575 (N_11575,N_11199,N_11430);
or U11576 (N_11576,N_11118,N_11349);
xnor U11577 (N_11577,N_11372,N_11073);
nand U11578 (N_11578,N_11043,N_11092);
nand U11579 (N_11579,N_11489,N_11348);
or U11580 (N_11580,N_11331,N_11329);
nand U11581 (N_11581,N_11338,N_11149);
nor U11582 (N_11582,N_11163,N_11185);
nor U11583 (N_11583,N_11366,N_11215);
or U11584 (N_11584,N_11459,N_11358);
or U11585 (N_11585,N_11032,N_11351);
nor U11586 (N_11586,N_11271,N_11034);
xor U11587 (N_11587,N_11312,N_11379);
or U11588 (N_11588,N_11254,N_11100);
or U11589 (N_11589,N_11037,N_11446);
and U11590 (N_11590,N_11497,N_11420);
or U11591 (N_11591,N_11136,N_11482);
or U11592 (N_11592,N_11332,N_11085);
and U11593 (N_11593,N_11378,N_11158);
nor U11594 (N_11594,N_11340,N_11059);
nand U11595 (N_11595,N_11249,N_11406);
nand U11596 (N_11596,N_11165,N_11140);
or U11597 (N_11597,N_11014,N_11011);
nand U11598 (N_11598,N_11402,N_11363);
nor U11599 (N_11599,N_11083,N_11463);
nor U11600 (N_11600,N_11409,N_11077);
nor U11601 (N_11601,N_11006,N_11125);
nor U11602 (N_11602,N_11181,N_11353);
nand U11603 (N_11603,N_11272,N_11370);
nor U11604 (N_11604,N_11196,N_11075);
nand U11605 (N_11605,N_11162,N_11216);
nand U11606 (N_11606,N_11295,N_11218);
or U11607 (N_11607,N_11440,N_11276);
or U11608 (N_11608,N_11012,N_11415);
nand U11609 (N_11609,N_11324,N_11285);
nand U11610 (N_11610,N_11206,N_11377);
nor U11611 (N_11611,N_11156,N_11444);
nor U11612 (N_11612,N_11115,N_11452);
and U11613 (N_11613,N_11474,N_11236);
nor U11614 (N_11614,N_11244,N_11197);
or U11615 (N_11615,N_11122,N_11154);
and U11616 (N_11616,N_11374,N_11278);
and U11617 (N_11617,N_11439,N_11035);
nor U11618 (N_11618,N_11050,N_11062);
nand U11619 (N_11619,N_11350,N_11038);
nor U11620 (N_11620,N_11499,N_11161);
xnor U11621 (N_11621,N_11297,N_11096);
and U11622 (N_11622,N_11397,N_11145);
nand U11623 (N_11623,N_11255,N_11273);
and U11624 (N_11624,N_11393,N_11423);
and U11625 (N_11625,N_11265,N_11368);
nor U11626 (N_11626,N_11067,N_11116);
and U11627 (N_11627,N_11159,N_11451);
xnor U11628 (N_11628,N_11016,N_11442);
nor U11629 (N_11629,N_11494,N_11082);
and U11630 (N_11630,N_11433,N_11090);
nor U11631 (N_11631,N_11167,N_11039);
xor U11632 (N_11632,N_11475,N_11490);
or U11633 (N_11633,N_11404,N_11495);
nand U11634 (N_11634,N_11394,N_11260);
or U11635 (N_11635,N_11234,N_11064);
nand U11636 (N_11636,N_11238,N_11045);
xnor U11637 (N_11637,N_11280,N_11124);
or U11638 (N_11638,N_11383,N_11269);
nor U11639 (N_11639,N_11209,N_11079);
or U11640 (N_11640,N_11169,N_11203);
nor U11641 (N_11641,N_11211,N_11396);
nand U11642 (N_11642,N_11101,N_11054);
or U11643 (N_11643,N_11025,N_11194);
nand U11644 (N_11644,N_11068,N_11078);
nand U11645 (N_11645,N_11214,N_11041);
nor U11646 (N_11646,N_11466,N_11480);
nor U11647 (N_11647,N_11347,N_11335);
or U11648 (N_11648,N_11412,N_11282);
nor U11649 (N_11649,N_11182,N_11231);
and U11650 (N_11650,N_11076,N_11245);
nor U11651 (N_11651,N_11384,N_11133);
or U11652 (N_11652,N_11382,N_11001);
and U11653 (N_11653,N_11201,N_11171);
nor U11654 (N_11654,N_11367,N_11388);
xnor U11655 (N_11655,N_11017,N_11496);
or U11656 (N_11656,N_11227,N_11147);
nor U11657 (N_11657,N_11294,N_11325);
and U11658 (N_11658,N_11121,N_11258);
and U11659 (N_11659,N_11128,N_11337);
or U11660 (N_11660,N_11000,N_11488);
nand U11661 (N_11661,N_11481,N_11029);
nand U11662 (N_11662,N_11191,N_11414);
or U11663 (N_11663,N_11328,N_11432);
nand U11664 (N_11664,N_11020,N_11326);
nand U11665 (N_11665,N_11455,N_11119);
nand U11666 (N_11666,N_11010,N_11468);
nand U11667 (N_11667,N_11219,N_11228);
nor U11668 (N_11668,N_11263,N_11239);
or U11669 (N_11669,N_11148,N_11051);
nor U11670 (N_11670,N_11352,N_11327);
nand U11671 (N_11671,N_11126,N_11251);
and U11672 (N_11672,N_11341,N_11220);
or U11673 (N_11673,N_11111,N_11009);
nor U11674 (N_11674,N_11261,N_11424);
nor U11675 (N_11675,N_11055,N_11426);
or U11676 (N_11676,N_11256,N_11491);
or U11677 (N_11677,N_11080,N_11212);
nor U11678 (N_11678,N_11049,N_11074);
nand U11679 (N_11679,N_11346,N_11005);
nand U11680 (N_11680,N_11407,N_11302);
nand U11681 (N_11681,N_11138,N_11323);
nor U11682 (N_11682,N_11204,N_11283);
or U11683 (N_11683,N_11134,N_11036);
nor U11684 (N_11684,N_11434,N_11048);
or U11685 (N_11685,N_11170,N_11284);
and U11686 (N_11686,N_11061,N_11405);
nand U11687 (N_11687,N_11376,N_11042);
or U11688 (N_11688,N_11109,N_11168);
nor U11689 (N_11689,N_11180,N_11450);
nand U11690 (N_11690,N_11117,N_11253);
nor U11691 (N_11691,N_11274,N_11355);
or U11692 (N_11692,N_11246,N_11257);
or U11693 (N_11693,N_11004,N_11361);
or U11694 (N_11694,N_11240,N_11202);
nor U11695 (N_11695,N_11290,N_11208);
and U11696 (N_11696,N_11157,N_11221);
nor U11697 (N_11697,N_11132,N_11190);
nor U11698 (N_11698,N_11188,N_11380);
nor U11699 (N_11699,N_11070,N_11210);
nand U11700 (N_11700,N_11106,N_11030);
nand U11701 (N_11701,N_11094,N_11287);
nand U11702 (N_11702,N_11427,N_11343);
nand U11703 (N_11703,N_11217,N_11031);
nand U11704 (N_11704,N_11471,N_11298);
or U11705 (N_11705,N_11311,N_11453);
and U11706 (N_11706,N_11127,N_11153);
nand U11707 (N_11707,N_11460,N_11142);
and U11708 (N_11708,N_11233,N_11226);
and U11709 (N_11709,N_11277,N_11114);
nor U11710 (N_11710,N_11146,N_11268);
and U11711 (N_11711,N_11322,N_11024);
or U11712 (N_11712,N_11086,N_11152);
nor U11713 (N_11713,N_11056,N_11081);
and U11714 (N_11714,N_11223,N_11314);
or U11715 (N_11715,N_11207,N_11333);
nor U11716 (N_11716,N_11192,N_11449);
nand U11717 (N_11717,N_11403,N_11436);
nor U11718 (N_11718,N_11342,N_11160);
or U11719 (N_11719,N_11013,N_11040);
nor U11720 (N_11720,N_11422,N_11303);
and U11721 (N_11721,N_11021,N_11144);
nand U11722 (N_11722,N_11135,N_11224);
and U11723 (N_11723,N_11267,N_11437);
nor U11724 (N_11724,N_11472,N_11176);
or U11725 (N_11725,N_11320,N_11103);
nor U11726 (N_11726,N_11229,N_11492);
nor U11727 (N_11727,N_11105,N_11205);
and U11728 (N_11728,N_11057,N_11173);
or U11729 (N_11729,N_11066,N_11373);
nor U11730 (N_11730,N_11345,N_11429);
nor U11731 (N_11731,N_11360,N_11232);
nand U11732 (N_11732,N_11317,N_11486);
nand U11733 (N_11733,N_11435,N_11198);
and U11734 (N_11734,N_11108,N_11493);
nand U11735 (N_11735,N_11130,N_11095);
and U11736 (N_11736,N_11321,N_11418);
nand U11737 (N_11737,N_11164,N_11425);
and U11738 (N_11738,N_11306,N_11222);
and U11739 (N_11739,N_11462,N_11113);
and U11740 (N_11740,N_11123,N_11183);
nor U11741 (N_11741,N_11252,N_11028);
and U11742 (N_11742,N_11099,N_11023);
nor U11743 (N_11743,N_11479,N_11098);
and U11744 (N_11744,N_11259,N_11447);
or U11745 (N_11745,N_11008,N_11419);
nor U11746 (N_11746,N_11288,N_11305);
or U11747 (N_11747,N_11400,N_11053);
or U11748 (N_11748,N_11484,N_11365);
or U11749 (N_11749,N_11389,N_11334);
and U11750 (N_11750,N_11482,N_11181);
nand U11751 (N_11751,N_11384,N_11383);
and U11752 (N_11752,N_11209,N_11226);
and U11753 (N_11753,N_11086,N_11137);
or U11754 (N_11754,N_11025,N_11397);
nor U11755 (N_11755,N_11174,N_11322);
or U11756 (N_11756,N_11353,N_11270);
xnor U11757 (N_11757,N_11239,N_11165);
nor U11758 (N_11758,N_11204,N_11417);
nand U11759 (N_11759,N_11241,N_11178);
nor U11760 (N_11760,N_11312,N_11094);
or U11761 (N_11761,N_11125,N_11146);
or U11762 (N_11762,N_11218,N_11298);
or U11763 (N_11763,N_11168,N_11475);
and U11764 (N_11764,N_11102,N_11353);
or U11765 (N_11765,N_11210,N_11363);
nor U11766 (N_11766,N_11050,N_11457);
and U11767 (N_11767,N_11320,N_11128);
or U11768 (N_11768,N_11391,N_11256);
and U11769 (N_11769,N_11178,N_11080);
nand U11770 (N_11770,N_11424,N_11462);
nor U11771 (N_11771,N_11227,N_11414);
or U11772 (N_11772,N_11479,N_11367);
or U11773 (N_11773,N_11206,N_11179);
or U11774 (N_11774,N_11165,N_11164);
nor U11775 (N_11775,N_11149,N_11326);
nand U11776 (N_11776,N_11268,N_11261);
and U11777 (N_11777,N_11277,N_11329);
nand U11778 (N_11778,N_11438,N_11142);
nor U11779 (N_11779,N_11239,N_11081);
nor U11780 (N_11780,N_11137,N_11293);
nor U11781 (N_11781,N_11177,N_11255);
nand U11782 (N_11782,N_11304,N_11244);
and U11783 (N_11783,N_11460,N_11411);
and U11784 (N_11784,N_11381,N_11217);
and U11785 (N_11785,N_11029,N_11334);
and U11786 (N_11786,N_11335,N_11060);
or U11787 (N_11787,N_11080,N_11072);
and U11788 (N_11788,N_11294,N_11164);
nand U11789 (N_11789,N_11433,N_11270);
nand U11790 (N_11790,N_11116,N_11267);
nand U11791 (N_11791,N_11006,N_11168);
nor U11792 (N_11792,N_11150,N_11137);
and U11793 (N_11793,N_11056,N_11355);
or U11794 (N_11794,N_11153,N_11118);
or U11795 (N_11795,N_11050,N_11279);
nand U11796 (N_11796,N_11110,N_11218);
or U11797 (N_11797,N_11259,N_11181);
and U11798 (N_11798,N_11183,N_11442);
nand U11799 (N_11799,N_11195,N_11391);
or U11800 (N_11800,N_11316,N_11489);
or U11801 (N_11801,N_11186,N_11357);
nor U11802 (N_11802,N_11214,N_11371);
nand U11803 (N_11803,N_11041,N_11378);
and U11804 (N_11804,N_11250,N_11405);
nor U11805 (N_11805,N_11367,N_11222);
xor U11806 (N_11806,N_11418,N_11101);
nor U11807 (N_11807,N_11164,N_11138);
nand U11808 (N_11808,N_11167,N_11417);
xnor U11809 (N_11809,N_11465,N_11384);
or U11810 (N_11810,N_11443,N_11272);
and U11811 (N_11811,N_11361,N_11373);
nand U11812 (N_11812,N_11334,N_11330);
nor U11813 (N_11813,N_11096,N_11270);
or U11814 (N_11814,N_11095,N_11316);
nor U11815 (N_11815,N_11065,N_11263);
or U11816 (N_11816,N_11310,N_11255);
and U11817 (N_11817,N_11397,N_11061);
nand U11818 (N_11818,N_11116,N_11041);
or U11819 (N_11819,N_11021,N_11201);
nand U11820 (N_11820,N_11492,N_11447);
or U11821 (N_11821,N_11492,N_11317);
nor U11822 (N_11822,N_11211,N_11271);
nor U11823 (N_11823,N_11435,N_11444);
nand U11824 (N_11824,N_11015,N_11233);
nor U11825 (N_11825,N_11443,N_11244);
nand U11826 (N_11826,N_11396,N_11121);
and U11827 (N_11827,N_11382,N_11358);
xor U11828 (N_11828,N_11392,N_11408);
nor U11829 (N_11829,N_11485,N_11014);
or U11830 (N_11830,N_11137,N_11149);
nand U11831 (N_11831,N_11003,N_11249);
nand U11832 (N_11832,N_11337,N_11127);
nor U11833 (N_11833,N_11422,N_11190);
or U11834 (N_11834,N_11384,N_11412);
and U11835 (N_11835,N_11315,N_11095);
or U11836 (N_11836,N_11324,N_11089);
xor U11837 (N_11837,N_11120,N_11165);
nand U11838 (N_11838,N_11353,N_11070);
and U11839 (N_11839,N_11009,N_11110);
or U11840 (N_11840,N_11460,N_11465);
or U11841 (N_11841,N_11499,N_11125);
or U11842 (N_11842,N_11074,N_11354);
or U11843 (N_11843,N_11157,N_11135);
or U11844 (N_11844,N_11186,N_11065);
nand U11845 (N_11845,N_11420,N_11192);
nand U11846 (N_11846,N_11478,N_11114);
nand U11847 (N_11847,N_11066,N_11269);
nor U11848 (N_11848,N_11438,N_11474);
or U11849 (N_11849,N_11441,N_11418);
nor U11850 (N_11850,N_11064,N_11146);
nand U11851 (N_11851,N_11141,N_11458);
nor U11852 (N_11852,N_11295,N_11007);
and U11853 (N_11853,N_11034,N_11257);
or U11854 (N_11854,N_11058,N_11292);
nor U11855 (N_11855,N_11386,N_11177);
and U11856 (N_11856,N_11255,N_11477);
and U11857 (N_11857,N_11143,N_11309);
nand U11858 (N_11858,N_11474,N_11362);
nand U11859 (N_11859,N_11126,N_11229);
and U11860 (N_11860,N_11086,N_11136);
nor U11861 (N_11861,N_11081,N_11474);
or U11862 (N_11862,N_11167,N_11199);
nor U11863 (N_11863,N_11339,N_11408);
and U11864 (N_11864,N_11486,N_11306);
or U11865 (N_11865,N_11240,N_11142);
nor U11866 (N_11866,N_11409,N_11246);
or U11867 (N_11867,N_11336,N_11341);
or U11868 (N_11868,N_11013,N_11478);
nand U11869 (N_11869,N_11021,N_11429);
or U11870 (N_11870,N_11099,N_11141);
nor U11871 (N_11871,N_11272,N_11364);
and U11872 (N_11872,N_11200,N_11117);
or U11873 (N_11873,N_11082,N_11475);
and U11874 (N_11874,N_11215,N_11086);
and U11875 (N_11875,N_11226,N_11326);
or U11876 (N_11876,N_11192,N_11108);
nand U11877 (N_11877,N_11164,N_11304);
or U11878 (N_11878,N_11230,N_11151);
or U11879 (N_11879,N_11435,N_11335);
nand U11880 (N_11880,N_11422,N_11222);
nand U11881 (N_11881,N_11364,N_11468);
or U11882 (N_11882,N_11458,N_11173);
nand U11883 (N_11883,N_11067,N_11283);
nand U11884 (N_11884,N_11197,N_11271);
xnor U11885 (N_11885,N_11008,N_11172);
nor U11886 (N_11886,N_11323,N_11213);
or U11887 (N_11887,N_11371,N_11433);
nand U11888 (N_11888,N_11108,N_11152);
or U11889 (N_11889,N_11068,N_11248);
or U11890 (N_11890,N_11348,N_11053);
nand U11891 (N_11891,N_11003,N_11102);
and U11892 (N_11892,N_11096,N_11202);
or U11893 (N_11893,N_11351,N_11136);
nor U11894 (N_11894,N_11400,N_11224);
nand U11895 (N_11895,N_11086,N_11369);
nand U11896 (N_11896,N_11213,N_11225);
and U11897 (N_11897,N_11378,N_11296);
nand U11898 (N_11898,N_11234,N_11205);
and U11899 (N_11899,N_11192,N_11066);
nand U11900 (N_11900,N_11215,N_11240);
nand U11901 (N_11901,N_11370,N_11049);
nor U11902 (N_11902,N_11053,N_11393);
nand U11903 (N_11903,N_11332,N_11440);
nor U11904 (N_11904,N_11394,N_11060);
nor U11905 (N_11905,N_11007,N_11287);
and U11906 (N_11906,N_11041,N_11374);
or U11907 (N_11907,N_11254,N_11248);
or U11908 (N_11908,N_11325,N_11343);
and U11909 (N_11909,N_11129,N_11175);
nor U11910 (N_11910,N_11233,N_11201);
nand U11911 (N_11911,N_11443,N_11254);
nand U11912 (N_11912,N_11226,N_11023);
and U11913 (N_11913,N_11261,N_11203);
and U11914 (N_11914,N_11420,N_11348);
or U11915 (N_11915,N_11321,N_11434);
nor U11916 (N_11916,N_11094,N_11480);
nor U11917 (N_11917,N_11470,N_11086);
or U11918 (N_11918,N_11186,N_11173);
nand U11919 (N_11919,N_11439,N_11327);
or U11920 (N_11920,N_11174,N_11209);
and U11921 (N_11921,N_11276,N_11481);
nor U11922 (N_11922,N_11288,N_11021);
nand U11923 (N_11923,N_11334,N_11016);
and U11924 (N_11924,N_11062,N_11162);
nor U11925 (N_11925,N_11417,N_11252);
nor U11926 (N_11926,N_11463,N_11246);
nor U11927 (N_11927,N_11284,N_11304);
nand U11928 (N_11928,N_11427,N_11138);
nand U11929 (N_11929,N_11274,N_11024);
and U11930 (N_11930,N_11202,N_11161);
nand U11931 (N_11931,N_11489,N_11218);
nand U11932 (N_11932,N_11051,N_11421);
nand U11933 (N_11933,N_11064,N_11363);
nor U11934 (N_11934,N_11465,N_11318);
nand U11935 (N_11935,N_11175,N_11446);
or U11936 (N_11936,N_11016,N_11343);
or U11937 (N_11937,N_11297,N_11293);
and U11938 (N_11938,N_11111,N_11240);
nor U11939 (N_11939,N_11458,N_11013);
and U11940 (N_11940,N_11457,N_11089);
nand U11941 (N_11941,N_11447,N_11385);
or U11942 (N_11942,N_11311,N_11283);
nor U11943 (N_11943,N_11452,N_11012);
and U11944 (N_11944,N_11039,N_11302);
nand U11945 (N_11945,N_11196,N_11285);
nand U11946 (N_11946,N_11456,N_11258);
nand U11947 (N_11947,N_11421,N_11317);
nor U11948 (N_11948,N_11227,N_11318);
and U11949 (N_11949,N_11205,N_11300);
nor U11950 (N_11950,N_11366,N_11054);
nand U11951 (N_11951,N_11109,N_11062);
and U11952 (N_11952,N_11177,N_11144);
or U11953 (N_11953,N_11141,N_11246);
and U11954 (N_11954,N_11262,N_11234);
xor U11955 (N_11955,N_11015,N_11202);
nand U11956 (N_11956,N_11378,N_11077);
and U11957 (N_11957,N_11464,N_11183);
or U11958 (N_11958,N_11455,N_11214);
and U11959 (N_11959,N_11458,N_11387);
or U11960 (N_11960,N_11053,N_11492);
nand U11961 (N_11961,N_11045,N_11142);
nor U11962 (N_11962,N_11389,N_11222);
nor U11963 (N_11963,N_11028,N_11133);
nand U11964 (N_11964,N_11215,N_11376);
nor U11965 (N_11965,N_11243,N_11030);
nand U11966 (N_11966,N_11236,N_11260);
or U11967 (N_11967,N_11226,N_11143);
nand U11968 (N_11968,N_11299,N_11038);
xor U11969 (N_11969,N_11235,N_11267);
or U11970 (N_11970,N_11444,N_11359);
or U11971 (N_11971,N_11159,N_11210);
and U11972 (N_11972,N_11053,N_11213);
or U11973 (N_11973,N_11324,N_11360);
nor U11974 (N_11974,N_11027,N_11248);
nor U11975 (N_11975,N_11212,N_11244);
and U11976 (N_11976,N_11091,N_11097);
and U11977 (N_11977,N_11087,N_11141);
or U11978 (N_11978,N_11425,N_11133);
or U11979 (N_11979,N_11392,N_11202);
or U11980 (N_11980,N_11401,N_11151);
or U11981 (N_11981,N_11359,N_11078);
and U11982 (N_11982,N_11498,N_11235);
xnor U11983 (N_11983,N_11029,N_11343);
nand U11984 (N_11984,N_11158,N_11280);
and U11985 (N_11985,N_11393,N_11205);
or U11986 (N_11986,N_11382,N_11410);
nand U11987 (N_11987,N_11162,N_11237);
and U11988 (N_11988,N_11264,N_11093);
nand U11989 (N_11989,N_11443,N_11078);
nand U11990 (N_11990,N_11073,N_11227);
and U11991 (N_11991,N_11412,N_11226);
and U11992 (N_11992,N_11096,N_11319);
nand U11993 (N_11993,N_11449,N_11484);
nor U11994 (N_11994,N_11467,N_11146);
nor U11995 (N_11995,N_11129,N_11374);
nand U11996 (N_11996,N_11093,N_11424);
nand U11997 (N_11997,N_11067,N_11458);
nand U11998 (N_11998,N_11357,N_11172);
nand U11999 (N_11999,N_11277,N_11490);
nand U12000 (N_12000,N_11790,N_11646);
xor U12001 (N_12001,N_11758,N_11562);
nand U12002 (N_12002,N_11647,N_11601);
nor U12003 (N_12003,N_11753,N_11616);
and U12004 (N_12004,N_11577,N_11864);
nor U12005 (N_12005,N_11913,N_11984);
and U12006 (N_12006,N_11779,N_11809);
and U12007 (N_12007,N_11846,N_11935);
and U12008 (N_12008,N_11835,N_11681);
xnor U12009 (N_12009,N_11757,N_11624);
nand U12010 (N_12010,N_11697,N_11664);
and U12011 (N_12011,N_11806,N_11620);
nor U12012 (N_12012,N_11986,N_11659);
and U12013 (N_12013,N_11805,N_11511);
or U12014 (N_12014,N_11612,N_11791);
and U12015 (N_12015,N_11800,N_11759);
or U12016 (N_12016,N_11535,N_11936);
and U12017 (N_12017,N_11585,N_11726);
and U12018 (N_12018,N_11582,N_11884);
or U12019 (N_12019,N_11554,N_11702);
and U12020 (N_12020,N_11823,N_11506);
nand U12021 (N_12021,N_11748,N_11827);
and U12022 (N_12022,N_11849,N_11880);
or U12023 (N_12023,N_11614,N_11816);
xnor U12024 (N_12024,N_11636,N_11843);
nor U12025 (N_12025,N_11866,N_11642);
xor U12026 (N_12026,N_11902,N_11547);
nor U12027 (N_12027,N_11596,N_11609);
nor U12028 (N_12028,N_11696,N_11847);
and U12029 (N_12029,N_11715,N_11894);
and U12030 (N_12030,N_11645,N_11522);
or U12031 (N_12031,N_11574,N_11896);
nand U12032 (N_12032,N_11649,N_11873);
and U12033 (N_12033,N_11676,N_11889);
and U12034 (N_12034,N_11524,N_11818);
and U12035 (N_12035,N_11989,N_11760);
and U12036 (N_12036,N_11743,N_11716);
and U12037 (N_12037,N_11611,N_11797);
or U12038 (N_12038,N_11631,N_11950);
and U12039 (N_12039,N_11739,N_11794);
nor U12040 (N_12040,N_11576,N_11970);
nor U12041 (N_12041,N_11639,N_11878);
or U12042 (N_12042,N_11851,N_11803);
nor U12043 (N_12043,N_11982,N_11543);
and U12044 (N_12044,N_11888,N_11708);
or U12045 (N_12045,N_11922,N_11865);
nand U12046 (N_12046,N_11597,N_11802);
nand U12047 (N_12047,N_11555,N_11980);
nand U12048 (N_12048,N_11774,N_11660);
nand U12049 (N_12049,N_11625,N_11912);
nor U12050 (N_12050,N_11523,N_11682);
or U12051 (N_12051,N_11749,N_11537);
and U12052 (N_12052,N_11714,N_11583);
nor U12053 (N_12053,N_11668,N_11921);
or U12054 (N_12054,N_11500,N_11837);
and U12055 (N_12055,N_11530,N_11958);
nor U12056 (N_12056,N_11915,N_11767);
nand U12057 (N_12057,N_11569,N_11613);
or U12058 (N_12058,N_11956,N_11819);
or U12059 (N_12059,N_11557,N_11877);
nand U12060 (N_12060,N_11890,N_11538);
or U12061 (N_12061,N_11804,N_11992);
nand U12062 (N_12062,N_11776,N_11814);
nor U12063 (N_12063,N_11505,N_11868);
xor U12064 (N_12064,N_11870,N_11990);
nand U12065 (N_12065,N_11504,N_11656);
or U12066 (N_12066,N_11947,N_11940);
nor U12067 (N_12067,N_11644,N_11633);
nand U12068 (N_12068,N_11897,N_11648);
and U12069 (N_12069,N_11684,N_11693);
nand U12070 (N_12070,N_11752,N_11669);
nor U12071 (N_12071,N_11605,N_11775);
and U12072 (N_12072,N_11621,N_11512);
or U12073 (N_12073,N_11626,N_11699);
or U12074 (N_12074,N_11813,N_11534);
nor U12075 (N_12075,N_11590,N_11763);
or U12076 (N_12076,N_11799,N_11903);
or U12077 (N_12077,N_11661,N_11706);
and U12078 (N_12078,N_11928,N_11932);
nand U12079 (N_12079,N_11727,N_11824);
nor U12080 (N_12080,N_11677,N_11939);
xnor U12081 (N_12081,N_11501,N_11793);
nand U12082 (N_12082,N_11899,N_11937);
nand U12083 (N_12083,N_11925,N_11919);
or U12084 (N_12084,N_11549,N_11988);
nand U12085 (N_12085,N_11658,N_11617);
or U12086 (N_12086,N_11862,N_11623);
nand U12087 (N_12087,N_11721,N_11967);
and U12088 (N_12088,N_11858,N_11671);
or U12089 (N_12089,N_11550,N_11879);
or U12090 (N_12090,N_11917,N_11575);
and U12091 (N_12091,N_11996,N_11971);
and U12092 (N_12092,N_11729,N_11540);
and U12093 (N_12093,N_11783,N_11964);
or U12094 (N_12094,N_11876,N_11717);
and U12095 (N_12095,N_11856,N_11694);
or U12096 (N_12096,N_11586,N_11825);
nor U12097 (N_12097,N_11587,N_11869);
or U12098 (N_12098,N_11909,N_11568);
nand U12099 (N_12099,N_11834,N_11503);
nor U12100 (N_12100,N_11777,N_11755);
and U12101 (N_12101,N_11675,N_11691);
nor U12102 (N_12102,N_11854,N_11926);
and U12103 (N_12103,N_11598,N_11718);
nand U12104 (N_12104,N_11859,N_11638);
nor U12105 (N_12105,N_11732,N_11904);
and U12106 (N_12106,N_11728,N_11987);
and U12107 (N_12107,N_11667,N_11544);
nand U12108 (N_12108,N_11910,N_11704);
nor U12109 (N_12109,N_11978,N_11931);
nand U12110 (N_12110,N_11997,N_11891);
nor U12111 (N_12111,N_11999,N_11578);
nand U12112 (N_12112,N_11957,N_11746);
or U12113 (N_12113,N_11563,N_11772);
nor U12114 (N_12114,N_11705,N_11829);
or U12115 (N_12115,N_11769,N_11845);
and U12116 (N_12116,N_11558,N_11968);
or U12117 (N_12117,N_11740,N_11579);
nand U12118 (N_12118,N_11528,N_11942);
nand U12119 (N_12119,N_11887,N_11632);
or U12120 (N_12120,N_11828,N_11710);
and U12121 (N_12121,N_11863,N_11961);
nor U12122 (N_12122,N_11559,N_11949);
and U12123 (N_12123,N_11874,N_11798);
nor U12124 (N_12124,N_11853,N_11965);
nor U12125 (N_12125,N_11692,N_11654);
or U12126 (N_12126,N_11548,N_11741);
nand U12127 (N_12127,N_11857,N_11689);
nand U12128 (N_12128,N_11698,N_11588);
xor U12129 (N_12129,N_11627,N_11551);
xnor U12130 (N_12130,N_11966,N_11589);
or U12131 (N_12131,N_11720,N_11652);
and U12132 (N_12132,N_11572,N_11541);
and U12133 (N_12133,N_11519,N_11820);
nand U12134 (N_12134,N_11521,N_11566);
and U12135 (N_12135,N_11738,N_11893);
nor U12136 (N_12136,N_11665,N_11606);
nand U12137 (N_12137,N_11977,N_11930);
or U12138 (N_12138,N_11860,N_11607);
xor U12139 (N_12139,N_11836,N_11680);
or U12140 (N_12140,N_11513,N_11539);
or U12141 (N_12141,N_11510,N_11918);
nor U12142 (N_12142,N_11810,N_11945);
or U12143 (N_12143,N_11686,N_11604);
nor U12144 (N_12144,N_11831,N_11952);
nand U12145 (N_12145,N_11591,N_11507);
nand U12146 (N_12146,N_11593,N_11920);
nand U12147 (N_12147,N_11975,N_11595);
or U12148 (N_12148,N_11842,N_11885);
and U12149 (N_12149,N_11784,N_11653);
nand U12150 (N_12150,N_11754,N_11666);
and U12151 (N_12151,N_11969,N_11788);
and U12152 (N_12152,N_11599,N_11985);
nor U12153 (N_12153,N_11929,N_11946);
or U12154 (N_12154,N_11592,N_11542);
and U12155 (N_12155,N_11608,N_11619);
nand U12156 (N_12156,N_11905,N_11695);
or U12157 (N_12157,N_11815,N_11995);
nor U12158 (N_12158,N_11580,N_11672);
or U12159 (N_12159,N_11841,N_11976);
nand U12160 (N_12160,N_11941,N_11955);
or U12161 (N_12161,N_11944,N_11745);
nor U12162 (N_12162,N_11839,N_11737);
and U12163 (N_12163,N_11933,N_11657);
or U12164 (N_12164,N_11571,N_11622);
nor U12165 (N_12165,N_11525,N_11822);
and U12166 (N_12166,N_11734,N_11807);
or U12167 (N_12167,N_11640,N_11795);
and U12168 (N_12168,N_11679,N_11785);
and U12169 (N_12169,N_11520,N_11981);
nor U12170 (N_12170,N_11786,N_11993);
nor U12171 (N_12171,N_11735,N_11650);
and U12172 (N_12172,N_11764,N_11526);
nor U12173 (N_12173,N_11855,N_11983);
nor U12174 (N_12174,N_11951,N_11736);
nor U12175 (N_12175,N_11532,N_11934);
or U12176 (N_12176,N_11778,N_11960);
nand U12177 (N_12177,N_11709,N_11895);
or U12178 (N_12178,N_11908,N_11529);
nand U12179 (N_12179,N_11773,N_11723);
or U12180 (N_12180,N_11954,N_11923);
and U12181 (N_12181,N_11712,N_11871);
nor U12182 (N_12182,N_11561,N_11581);
nor U12183 (N_12183,N_11643,N_11898);
nor U12184 (N_12184,N_11801,N_11906);
or U12185 (N_12185,N_11911,N_11655);
nor U12186 (N_12186,N_11938,N_11508);
nor U12187 (N_12187,N_11610,N_11766);
nand U12188 (N_12188,N_11635,N_11750);
nand U12189 (N_12189,N_11509,N_11924);
nor U12190 (N_12190,N_11570,N_11628);
nor U12191 (N_12191,N_11796,N_11687);
xnor U12192 (N_12192,N_11678,N_11603);
and U12193 (N_12193,N_11780,N_11546);
or U12194 (N_12194,N_11707,N_11916);
and U12195 (N_12195,N_11670,N_11567);
and U12196 (N_12196,N_11812,N_11700);
nor U12197 (N_12197,N_11531,N_11744);
and U12198 (N_12198,N_11556,N_11517);
nor U12199 (N_12199,N_11527,N_11761);
and U12200 (N_12200,N_11892,N_11875);
xnor U12201 (N_12201,N_11782,N_11713);
and U12202 (N_12202,N_11900,N_11787);
nor U12203 (N_12203,N_11789,N_11770);
nand U12204 (N_12204,N_11882,N_11553);
nor U12205 (N_12205,N_11768,N_11830);
nor U12206 (N_12206,N_11808,N_11881);
and U12207 (N_12207,N_11685,N_11848);
nand U12208 (N_12208,N_11914,N_11711);
and U12209 (N_12209,N_11536,N_11565);
and U12210 (N_12210,N_11771,N_11733);
or U12211 (N_12211,N_11742,N_11637);
nor U12212 (N_12212,N_11762,N_11533);
nor U12213 (N_12213,N_11959,N_11615);
nor U12214 (N_12214,N_11991,N_11518);
nor U12215 (N_12215,N_11634,N_11972);
nor U12216 (N_12216,N_11701,N_11979);
and U12217 (N_12217,N_11886,N_11618);
nand U12218 (N_12218,N_11630,N_11674);
or U12219 (N_12219,N_11751,N_11974);
and U12220 (N_12220,N_11560,N_11833);
nand U12221 (N_12221,N_11826,N_11725);
and U12222 (N_12222,N_11821,N_11883);
nand U12223 (N_12223,N_11514,N_11564);
and U12224 (N_12224,N_11584,N_11963);
nor U12225 (N_12225,N_11731,N_11724);
nor U12226 (N_12226,N_11852,N_11690);
and U12227 (N_12227,N_11927,N_11722);
or U12228 (N_12228,N_11948,N_11844);
and U12229 (N_12229,N_11545,N_11662);
and U12230 (N_12230,N_11641,N_11756);
nand U12231 (N_12231,N_11673,N_11953);
nor U12232 (N_12232,N_11502,N_11907);
and U12233 (N_12233,N_11998,N_11872);
nand U12234 (N_12234,N_11663,N_11850);
or U12235 (N_12235,N_11683,N_11747);
or U12236 (N_12236,N_11688,N_11861);
nor U12237 (N_12237,N_11792,N_11867);
and U12238 (N_12238,N_11962,N_11552);
nor U12239 (N_12239,N_11943,N_11973);
and U12240 (N_12240,N_11651,N_11703);
nor U12241 (N_12241,N_11994,N_11840);
nand U12242 (N_12242,N_11730,N_11817);
nand U12243 (N_12243,N_11781,N_11594);
nor U12244 (N_12244,N_11832,N_11515);
nand U12245 (N_12245,N_11838,N_11516);
or U12246 (N_12246,N_11811,N_11901);
and U12247 (N_12247,N_11719,N_11765);
and U12248 (N_12248,N_11629,N_11602);
or U12249 (N_12249,N_11573,N_11600);
and U12250 (N_12250,N_11585,N_11595);
or U12251 (N_12251,N_11555,N_11714);
and U12252 (N_12252,N_11745,N_11661);
nand U12253 (N_12253,N_11884,N_11629);
or U12254 (N_12254,N_11638,N_11948);
nor U12255 (N_12255,N_11569,N_11846);
nor U12256 (N_12256,N_11813,N_11803);
nor U12257 (N_12257,N_11642,N_11992);
nand U12258 (N_12258,N_11847,N_11852);
nand U12259 (N_12259,N_11853,N_11922);
and U12260 (N_12260,N_11833,N_11538);
and U12261 (N_12261,N_11753,N_11812);
and U12262 (N_12262,N_11998,N_11659);
nand U12263 (N_12263,N_11551,N_11809);
and U12264 (N_12264,N_11765,N_11999);
and U12265 (N_12265,N_11587,N_11594);
nor U12266 (N_12266,N_11588,N_11548);
or U12267 (N_12267,N_11621,N_11862);
and U12268 (N_12268,N_11923,N_11693);
nand U12269 (N_12269,N_11655,N_11865);
nand U12270 (N_12270,N_11610,N_11763);
and U12271 (N_12271,N_11776,N_11793);
nand U12272 (N_12272,N_11522,N_11640);
nor U12273 (N_12273,N_11886,N_11616);
nor U12274 (N_12274,N_11888,N_11595);
and U12275 (N_12275,N_11902,N_11502);
nor U12276 (N_12276,N_11852,N_11572);
xor U12277 (N_12277,N_11881,N_11507);
nand U12278 (N_12278,N_11986,N_11972);
or U12279 (N_12279,N_11922,N_11591);
nand U12280 (N_12280,N_11542,N_11851);
and U12281 (N_12281,N_11942,N_11860);
nor U12282 (N_12282,N_11920,N_11778);
xor U12283 (N_12283,N_11589,N_11832);
and U12284 (N_12284,N_11749,N_11555);
or U12285 (N_12285,N_11919,N_11932);
nor U12286 (N_12286,N_11992,N_11816);
nor U12287 (N_12287,N_11612,N_11590);
and U12288 (N_12288,N_11917,N_11588);
nor U12289 (N_12289,N_11519,N_11978);
or U12290 (N_12290,N_11520,N_11843);
nand U12291 (N_12291,N_11948,N_11726);
nor U12292 (N_12292,N_11977,N_11883);
or U12293 (N_12293,N_11616,N_11897);
and U12294 (N_12294,N_11576,N_11823);
or U12295 (N_12295,N_11866,N_11613);
and U12296 (N_12296,N_11574,N_11932);
nor U12297 (N_12297,N_11677,N_11654);
nor U12298 (N_12298,N_11748,N_11991);
or U12299 (N_12299,N_11659,N_11897);
or U12300 (N_12300,N_11948,N_11755);
nor U12301 (N_12301,N_11870,N_11939);
nor U12302 (N_12302,N_11937,N_11903);
nand U12303 (N_12303,N_11533,N_11860);
nand U12304 (N_12304,N_11566,N_11748);
nand U12305 (N_12305,N_11933,N_11754);
nor U12306 (N_12306,N_11653,N_11697);
or U12307 (N_12307,N_11908,N_11619);
nand U12308 (N_12308,N_11849,N_11920);
and U12309 (N_12309,N_11932,N_11580);
nor U12310 (N_12310,N_11888,N_11503);
or U12311 (N_12311,N_11544,N_11832);
or U12312 (N_12312,N_11591,N_11698);
nand U12313 (N_12313,N_11505,N_11832);
nand U12314 (N_12314,N_11845,N_11976);
nor U12315 (N_12315,N_11940,N_11633);
nor U12316 (N_12316,N_11639,N_11713);
nor U12317 (N_12317,N_11532,N_11644);
or U12318 (N_12318,N_11623,N_11935);
nand U12319 (N_12319,N_11691,N_11711);
nor U12320 (N_12320,N_11780,N_11678);
or U12321 (N_12321,N_11692,N_11777);
and U12322 (N_12322,N_11550,N_11761);
xnor U12323 (N_12323,N_11844,N_11925);
nor U12324 (N_12324,N_11772,N_11942);
or U12325 (N_12325,N_11674,N_11629);
nand U12326 (N_12326,N_11983,N_11748);
and U12327 (N_12327,N_11893,N_11562);
or U12328 (N_12328,N_11849,N_11540);
nor U12329 (N_12329,N_11730,N_11791);
nor U12330 (N_12330,N_11968,N_11872);
or U12331 (N_12331,N_11730,N_11965);
nand U12332 (N_12332,N_11921,N_11604);
or U12333 (N_12333,N_11909,N_11816);
or U12334 (N_12334,N_11727,N_11605);
and U12335 (N_12335,N_11759,N_11683);
and U12336 (N_12336,N_11762,N_11778);
nor U12337 (N_12337,N_11873,N_11652);
nand U12338 (N_12338,N_11830,N_11978);
and U12339 (N_12339,N_11994,N_11672);
nand U12340 (N_12340,N_11819,N_11908);
or U12341 (N_12341,N_11655,N_11666);
nand U12342 (N_12342,N_11912,N_11934);
or U12343 (N_12343,N_11849,N_11782);
nor U12344 (N_12344,N_11858,N_11510);
nand U12345 (N_12345,N_11939,N_11923);
nor U12346 (N_12346,N_11771,N_11820);
and U12347 (N_12347,N_11660,N_11958);
or U12348 (N_12348,N_11901,N_11730);
nor U12349 (N_12349,N_11546,N_11525);
or U12350 (N_12350,N_11703,N_11877);
nand U12351 (N_12351,N_11816,N_11759);
and U12352 (N_12352,N_11979,N_11980);
nor U12353 (N_12353,N_11613,N_11576);
nand U12354 (N_12354,N_11857,N_11631);
and U12355 (N_12355,N_11820,N_11527);
nand U12356 (N_12356,N_11571,N_11775);
or U12357 (N_12357,N_11924,N_11538);
nor U12358 (N_12358,N_11797,N_11731);
nor U12359 (N_12359,N_11656,N_11810);
or U12360 (N_12360,N_11576,N_11711);
and U12361 (N_12361,N_11705,N_11973);
nor U12362 (N_12362,N_11622,N_11827);
nand U12363 (N_12363,N_11976,N_11851);
nand U12364 (N_12364,N_11799,N_11884);
nor U12365 (N_12365,N_11698,N_11810);
nor U12366 (N_12366,N_11504,N_11586);
nor U12367 (N_12367,N_11702,N_11765);
or U12368 (N_12368,N_11647,N_11713);
and U12369 (N_12369,N_11616,N_11630);
and U12370 (N_12370,N_11807,N_11518);
or U12371 (N_12371,N_11567,N_11673);
nor U12372 (N_12372,N_11700,N_11847);
nand U12373 (N_12373,N_11931,N_11966);
nand U12374 (N_12374,N_11621,N_11813);
and U12375 (N_12375,N_11751,N_11571);
and U12376 (N_12376,N_11916,N_11807);
nor U12377 (N_12377,N_11812,N_11664);
nor U12378 (N_12378,N_11700,N_11569);
nor U12379 (N_12379,N_11883,N_11731);
or U12380 (N_12380,N_11658,N_11887);
nor U12381 (N_12381,N_11529,N_11537);
nor U12382 (N_12382,N_11537,N_11868);
or U12383 (N_12383,N_11830,N_11886);
nor U12384 (N_12384,N_11583,N_11890);
nor U12385 (N_12385,N_11529,N_11829);
xnor U12386 (N_12386,N_11950,N_11782);
or U12387 (N_12387,N_11624,N_11867);
nand U12388 (N_12388,N_11772,N_11870);
nand U12389 (N_12389,N_11859,N_11815);
nand U12390 (N_12390,N_11643,N_11819);
nor U12391 (N_12391,N_11912,N_11684);
nand U12392 (N_12392,N_11631,N_11603);
nand U12393 (N_12393,N_11532,N_11618);
nand U12394 (N_12394,N_11627,N_11936);
xor U12395 (N_12395,N_11601,N_11664);
nand U12396 (N_12396,N_11714,N_11658);
xnor U12397 (N_12397,N_11593,N_11879);
nand U12398 (N_12398,N_11854,N_11797);
nand U12399 (N_12399,N_11557,N_11688);
nand U12400 (N_12400,N_11847,N_11837);
nor U12401 (N_12401,N_11704,N_11803);
or U12402 (N_12402,N_11839,N_11713);
or U12403 (N_12403,N_11964,N_11822);
and U12404 (N_12404,N_11539,N_11720);
nor U12405 (N_12405,N_11993,N_11605);
nand U12406 (N_12406,N_11585,N_11822);
or U12407 (N_12407,N_11536,N_11611);
and U12408 (N_12408,N_11796,N_11650);
nor U12409 (N_12409,N_11961,N_11927);
nand U12410 (N_12410,N_11531,N_11513);
and U12411 (N_12411,N_11524,N_11692);
nor U12412 (N_12412,N_11545,N_11621);
or U12413 (N_12413,N_11669,N_11634);
nor U12414 (N_12414,N_11543,N_11671);
nand U12415 (N_12415,N_11995,N_11521);
or U12416 (N_12416,N_11731,N_11604);
or U12417 (N_12417,N_11962,N_11816);
nor U12418 (N_12418,N_11793,N_11881);
nor U12419 (N_12419,N_11672,N_11756);
nor U12420 (N_12420,N_11624,N_11613);
and U12421 (N_12421,N_11952,N_11872);
nor U12422 (N_12422,N_11640,N_11683);
or U12423 (N_12423,N_11840,N_11905);
nand U12424 (N_12424,N_11990,N_11864);
nand U12425 (N_12425,N_11767,N_11793);
nand U12426 (N_12426,N_11922,N_11891);
or U12427 (N_12427,N_11525,N_11596);
nor U12428 (N_12428,N_11737,N_11822);
nand U12429 (N_12429,N_11980,N_11933);
or U12430 (N_12430,N_11587,N_11640);
and U12431 (N_12431,N_11574,N_11693);
nand U12432 (N_12432,N_11954,N_11943);
nor U12433 (N_12433,N_11803,N_11878);
nand U12434 (N_12434,N_11558,N_11977);
nand U12435 (N_12435,N_11953,N_11995);
nand U12436 (N_12436,N_11534,N_11876);
or U12437 (N_12437,N_11818,N_11584);
nand U12438 (N_12438,N_11996,N_11952);
nand U12439 (N_12439,N_11899,N_11614);
nor U12440 (N_12440,N_11987,N_11634);
nor U12441 (N_12441,N_11617,N_11882);
xnor U12442 (N_12442,N_11696,N_11931);
and U12443 (N_12443,N_11916,N_11960);
nor U12444 (N_12444,N_11541,N_11855);
nor U12445 (N_12445,N_11506,N_11718);
and U12446 (N_12446,N_11569,N_11994);
or U12447 (N_12447,N_11917,N_11909);
or U12448 (N_12448,N_11979,N_11840);
nand U12449 (N_12449,N_11513,N_11814);
or U12450 (N_12450,N_11598,N_11646);
nor U12451 (N_12451,N_11663,N_11915);
nor U12452 (N_12452,N_11525,N_11980);
and U12453 (N_12453,N_11531,N_11950);
or U12454 (N_12454,N_11920,N_11812);
and U12455 (N_12455,N_11776,N_11584);
nor U12456 (N_12456,N_11881,N_11694);
nand U12457 (N_12457,N_11690,N_11828);
nand U12458 (N_12458,N_11696,N_11766);
or U12459 (N_12459,N_11511,N_11868);
nand U12460 (N_12460,N_11782,N_11721);
nor U12461 (N_12461,N_11953,N_11878);
nor U12462 (N_12462,N_11652,N_11904);
nand U12463 (N_12463,N_11926,N_11748);
nand U12464 (N_12464,N_11577,N_11824);
or U12465 (N_12465,N_11788,N_11909);
and U12466 (N_12466,N_11868,N_11614);
nand U12467 (N_12467,N_11695,N_11953);
nor U12468 (N_12468,N_11809,N_11916);
and U12469 (N_12469,N_11780,N_11592);
xor U12470 (N_12470,N_11835,N_11684);
and U12471 (N_12471,N_11587,N_11589);
nand U12472 (N_12472,N_11938,N_11633);
or U12473 (N_12473,N_11895,N_11797);
nand U12474 (N_12474,N_11932,N_11732);
and U12475 (N_12475,N_11970,N_11811);
xnor U12476 (N_12476,N_11608,N_11938);
and U12477 (N_12477,N_11711,N_11906);
or U12478 (N_12478,N_11933,N_11592);
or U12479 (N_12479,N_11607,N_11877);
or U12480 (N_12480,N_11625,N_11658);
nand U12481 (N_12481,N_11927,N_11858);
nand U12482 (N_12482,N_11701,N_11792);
nor U12483 (N_12483,N_11649,N_11506);
nor U12484 (N_12484,N_11724,N_11823);
nor U12485 (N_12485,N_11701,N_11798);
nand U12486 (N_12486,N_11839,N_11812);
nand U12487 (N_12487,N_11820,N_11635);
and U12488 (N_12488,N_11930,N_11621);
nand U12489 (N_12489,N_11711,N_11572);
or U12490 (N_12490,N_11917,N_11854);
nor U12491 (N_12491,N_11895,N_11523);
xor U12492 (N_12492,N_11840,N_11546);
nor U12493 (N_12493,N_11553,N_11821);
and U12494 (N_12494,N_11934,N_11555);
and U12495 (N_12495,N_11504,N_11655);
or U12496 (N_12496,N_11992,N_11942);
nand U12497 (N_12497,N_11630,N_11676);
nand U12498 (N_12498,N_11914,N_11819);
nand U12499 (N_12499,N_11806,N_11778);
nand U12500 (N_12500,N_12491,N_12039);
or U12501 (N_12501,N_12482,N_12191);
nor U12502 (N_12502,N_12384,N_12286);
and U12503 (N_12503,N_12228,N_12147);
and U12504 (N_12504,N_12262,N_12208);
xor U12505 (N_12505,N_12156,N_12352);
and U12506 (N_12506,N_12238,N_12211);
and U12507 (N_12507,N_12284,N_12389);
nand U12508 (N_12508,N_12251,N_12323);
or U12509 (N_12509,N_12429,N_12124);
or U12510 (N_12510,N_12485,N_12223);
or U12511 (N_12511,N_12473,N_12250);
or U12512 (N_12512,N_12050,N_12186);
nand U12513 (N_12513,N_12302,N_12413);
nor U12514 (N_12514,N_12259,N_12014);
and U12515 (N_12515,N_12012,N_12112);
nor U12516 (N_12516,N_12455,N_12493);
and U12517 (N_12517,N_12280,N_12283);
or U12518 (N_12518,N_12111,N_12037);
and U12519 (N_12519,N_12380,N_12201);
or U12520 (N_12520,N_12232,N_12486);
and U12521 (N_12521,N_12433,N_12324);
nand U12522 (N_12522,N_12479,N_12080);
xor U12523 (N_12523,N_12436,N_12071);
and U12524 (N_12524,N_12133,N_12487);
and U12525 (N_12525,N_12265,N_12119);
nor U12526 (N_12526,N_12178,N_12464);
nand U12527 (N_12527,N_12372,N_12184);
or U12528 (N_12528,N_12008,N_12297);
nand U12529 (N_12529,N_12396,N_12020);
or U12530 (N_12530,N_12195,N_12469);
nor U12531 (N_12531,N_12356,N_12047);
nand U12532 (N_12532,N_12225,N_12398);
nor U12533 (N_12533,N_12375,N_12086);
and U12534 (N_12534,N_12214,N_12160);
nor U12535 (N_12535,N_12062,N_12472);
or U12536 (N_12536,N_12296,N_12377);
nor U12537 (N_12537,N_12040,N_12237);
and U12538 (N_12538,N_12365,N_12104);
and U12539 (N_12539,N_12064,N_12350);
xnor U12540 (N_12540,N_12338,N_12094);
nor U12541 (N_12541,N_12371,N_12194);
nor U12542 (N_12542,N_12461,N_12107);
or U12543 (N_12543,N_12084,N_12068);
nor U12544 (N_12544,N_12139,N_12411);
and U12545 (N_12545,N_12041,N_12340);
or U12546 (N_12546,N_12495,N_12034);
nor U12547 (N_12547,N_12131,N_12373);
or U12548 (N_12548,N_12336,N_12056);
and U12549 (N_12549,N_12305,N_12307);
nand U12550 (N_12550,N_12113,N_12101);
nor U12551 (N_12551,N_12349,N_12256);
and U12552 (N_12552,N_12418,N_12183);
and U12553 (N_12553,N_12480,N_12221);
nor U12554 (N_12554,N_12368,N_12278);
nor U12555 (N_12555,N_12177,N_12029);
nor U12556 (N_12556,N_12312,N_12125);
and U12557 (N_12557,N_12002,N_12153);
nor U12558 (N_12558,N_12016,N_12386);
and U12559 (N_12559,N_12341,N_12154);
or U12560 (N_12560,N_12437,N_12328);
nand U12561 (N_12561,N_12116,N_12475);
nand U12562 (N_12562,N_12360,N_12110);
and U12563 (N_12563,N_12400,N_12130);
or U12564 (N_12564,N_12248,N_12488);
nor U12565 (N_12565,N_12310,N_12209);
or U12566 (N_12566,N_12009,N_12026);
and U12567 (N_12567,N_12106,N_12048);
nand U12568 (N_12568,N_12388,N_12244);
and U12569 (N_12569,N_12440,N_12145);
nand U12570 (N_12570,N_12367,N_12152);
or U12571 (N_12571,N_12192,N_12355);
and U12572 (N_12572,N_12470,N_12369);
xor U12573 (N_12573,N_12281,N_12406);
and U12574 (N_12574,N_12415,N_12474);
nand U12575 (N_12575,N_12067,N_12462);
nor U12576 (N_12576,N_12300,N_12035);
or U12577 (N_12577,N_12490,N_12379);
nor U12578 (N_12578,N_12290,N_12199);
nand U12579 (N_12579,N_12254,N_12174);
and U12580 (N_12580,N_12291,N_12212);
and U12581 (N_12581,N_12424,N_12091);
and U12582 (N_12582,N_12230,N_12046);
and U12583 (N_12583,N_12391,N_12031);
xor U12584 (N_12584,N_12070,N_12481);
nor U12585 (N_12585,N_12011,N_12477);
or U12586 (N_12586,N_12332,N_12466);
nor U12587 (N_12587,N_12025,N_12401);
or U12588 (N_12588,N_12090,N_12024);
nand U12589 (N_12589,N_12102,N_12122);
or U12590 (N_12590,N_12412,N_12061);
nand U12591 (N_12591,N_12150,N_12497);
nand U12592 (N_12592,N_12361,N_12081);
and U12593 (N_12593,N_12088,N_12492);
and U12594 (N_12594,N_12202,N_12337);
nand U12595 (N_12595,N_12326,N_12357);
nand U12596 (N_12596,N_12393,N_12456);
nand U12597 (N_12597,N_12231,N_12077);
and U12598 (N_12598,N_12489,N_12144);
and U12599 (N_12599,N_12022,N_12451);
xor U12600 (N_12600,N_12051,N_12318);
nand U12601 (N_12601,N_12193,N_12459);
nor U12602 (N_12602,N_12141,N_12364);
or U12603 (N_12603,N_12348,N_12120);
nor U12604 (N_12604,N_12273,N_12353);
nor U12605 (N_12605,N_12172,N_12285);
nand U12606 (N_12606,N_12204,N_12158);
nor U12607 (N_12607,N_12423,N_12115);
or U12608 (N_12608,N_12381,N_12319);
nor U12609 (N_12609,N_12460,N_12288);
nand U12610 (N_12610,N_12496,N_12042);
and U12611 (N_12611,N_12339,N_12181);
nand U12612 (N_12612,N_12015,N_12374);
or U12613 (N_12613,N_12126,N_12498);
and U12614 (N_12614,N_12478,N_12171);
and U12615 (N_12615,N_12260,N_12180);
and U12616 (N_12616,N_12007,N_12074);
and U12617 (N_12617,N_12200,N_12175);
nand U12618 (N_12618,N_12151,N_12216);
or U12619 (N_12619,N_12394,N_12438);
nor U12620 (N_12620,N_12358,N_12004);
nor U12621 (N_12621,N_12279,N_12027);
and U12622 (N_12622,N_12434,N_12155);
nor U12623 (N_12623,N_12162,N_12363);
nor U12624 (N_12624,N_12142,N_12347);
nand U12625 (N_12625,N_12370,N_12079);
or U12626 (N_12626,N_12096,N_12114);
or U12627 (N_12627,N_12419,N_12241);
nand U12628 (N_12628,N_12019,N_12330);
nor U12629 (N_12629,N_12089,N_12117);
nand U12630 (N_12630,N_12063,N_12137);
nand U12631 (N_12631,N_12315,N_12446);
or U12632 (N_12632,N_12058,N_12021);
nand U12633 (N_12633,N_12435,N_12399);
or U12634 (N_12634,N_12476,N_12448);
or U12635 (N_12635,N_12207,N_12320);
or U12636 (N_12636,N_12210,N_12416);
nor U12637 (N_12637,N_12409,N_12093);
or U12638 (N_12638,N_12390,N_12030);
and U12639 (N_12639,N_12168,N_12043);
nand U12640 (N_12640,N_12407,N_12165);
xor U12641 (N_12641,N_12362,N_12057);
nand U12642 (N_12642,N_12161,N_12342);
nand U12643 (N_12643,N_12309,N_12032);
xor U12644 (N_12644,N_12299,N_12135);
nand U12645 (N_12645,N_12454,N_12376);
nand U12646 (N_12646,N_12306,N_12322);
nand U12647 (N_12647,N_12366,N_12001);
and U12648 (N_12648,N_12308,N_12494);
or U12649 (N_12649,N_12421,N_12234);
nor U12650 (N_12650,N_12313,N_12245);
and U12651 (N_12651,N_12382,N_12257);
nand U12652 (N_12652,N_12410,N_12123);
and U12653 (N_12653,N_12268,N_12303);
nor U12654 (N_12654,N_12065,N_12447);
nor U12655 (N_12655,N_12233,N_12452);
and U12656 (N_12656,N_12203,N_12134);
nor U12657 (N_12657,N_12346,N_12182);
and U12658 (N_12658,N_12264,N_12054);
or U12659 (N_12659,N_12321,N_12427);
nor U12660 (N_12660,N_12439,N_12270);
or U12661 (N_12661,N_12017,N_12138);
and U12662 (N_12662,N_12185,N_12467);
and U12663 (N_12663,N_12457,N_12404);
xnor U12664 (N_12664,N_12100,N_12463);
nor U12665 (N_12665,N_12010,N_12468);
nor U12666 (N_12666,N_12003,N_12235);
or U12667 (N_12667,N_12060,N_12149);
or U12668 (N_12668,N_12219,N_12227);
nand U12669 (N_12669,N_12426,N_12450);
nor U12670 (N_12670,N_12073,N_12325);
xnor U12671 (N_12671,N_12222,N_12044);
and U12672 (N_12672,N_12217,N_12164);
nand U12673 (N_12673,N_12099,N_12197);
nand U12674 (N_12674,N_12092,N_12213);
or U12675 (N_12675,N_12229,N_12255);
nand U12676 (N_12676,N_12188,N_12000);
nand U12677 (N_12677,N_12189,N_12148);
or U12678 (N_12678,N_12392,N_12301);
nor U12679 (N_12679,N_12395,N_12275);
nor U12680 (N_12680,N_12387,N_12432);
nor U12681 (N_12681,N_12287,N_12095);
nor U12682 (N_12682,N_12103,N_12179);
nand U12683 (N_12683,N_12484,N_12397);
or U12684 (N_12684,N_12176,N_12163);
or U12685 (N_12685,N_12499,N_12140);
and U12686 (N_12686,N_12239,N_12276);
nand U12687 (N_12687,N_12267,N_12205);
and U12688 (N_12688,N_12072,N_12127);
or U12689 (N_12689,N_12403,N_12220);
nand U12690 (N_12690,N_12458,N_12344);
or U12691 (N_12691,N_12097,N_12075);
nor U12692 (N_12692,N_12453,N_12243);
nand U12693 (N_12693,N_12258,N_12261);
nor U12694 (N_12694,N_12274,N_12298);
nand U12695 (N_12695,N_12483,N_12085);
xor U12696 (N_12696,N_12083,N_12129);
and U12697 (N_12697,N_12218,N_12441);
nor U12698 (N_12698,N_12249,N_12187);
or U12699 (N_12699,N_12335,N_12331);
nand U12700 (N_12700,N_12078,N_12069);
nand U12701 (N_12701,N_12028,N_12005);
nor U12702 (N_12702,N_12018,N_12334);
xnor U12703 (N_12703,N_12170,N_12121);
nand U12704 (N_12704,N_12049,N_12240);
nand U12705 (N_12705,N_12289,N_12428);
nand U12706 (N_12706,N_12157,N_12343);
nor U12707 (N_12707,N_12449,N_12082);
xor U12708 (N_12708,N_12442,N_12402);
nand U12709 (N_12709,N_12294,N_12173);
nand U12710 (N_12710,N_12118,N_12226);
nor U12711 (N_12711,N_12053,N_12045);
nor U12712 (N_12712,N_12277,N_12143);
nand U12713 (N_12713,N_12059,N_12408);
or U12714 (N_12714,N_12445,N_12354);
nand U12715 (N_12715,N_12351,N_12292);
or U12716 (N_12716,N_12417,N_12242);
nand U12717 (N_12717,N_12444,N_12036);
nor U12718 (N_12718,N_12405,N_12304);
nand U12719 (N_12719,N_12420,N_12167);
nand U12720 (N_12720,N_12169,N_12317);
and U12721 (N_12721,N_12443,N_12345);
nor U12722 (N_12722,N_12266,N_12431);
nand U12723 (N_12723,N_12033,N_12314);
nand U12724 (N_12724,N_12269,N_12146);
nand U12725 (N_12725,N_12293,N_12066);
nor U12726 (N_12726,N_12196,N_12087);
and U12727 (N_12727,N_12378,N_12108);
nor U12728 (N_12728,N_12359,N_12023);
or U12729 (N_12729,N_12166,N_12206);
nand U12730 (N_12730,N_12271,N_12159);
nand U12731 (N_12731,N_12006,N_12215);
xor U12732 (N_12732,N_12327,N_12414);
nand U12733 (N_12733,N_12422,N_12471);
and U12734 (N_12734,N_12295,N_12425);
or U12735 (N_12735,N_12136,N_12055);
nor U12736 (N_12736,N_12109,N_12190);
or U12737 (N_12737,N_12311,N_12098);
or U12738 (N_12738,N_12263,N_12465);
nor U12739 (N_12739,N_12253,N_12385);
or U12740 (N_12740,N_12013,N_12198);
nor U12741 (N_12741,N_12224,N_12038);
nor U12742 (N_12742,N_12132,N_12128);
nor U12743 (N_12743,N_12076,N_12236);
nor U12744 (N_12744,N_12252,N_12430);
or U12745 (N_12745,N_12247,N_12272);
and U12746 (N_12746,N_12383,N_12333);
or U12747 (N_12747,N_12246,N_12105);
nor U12748 (N_12748,N_12282,N_12329);
nor U12749 (N_12749,N_12052,N_12316);
nand U12750 (N_12750,N_12278,N_12331);
and U12751 (N_12751,N_12415,N_12003);
nand U12752 (N_12752,N_12333,N_12414);
and U12753 (N_12753,N_12197,N_12067);
nor U12754 (N_12754,N_12315,N_12267);
or U12755 (N_12755,N_12003,N_12457);
or U12756 (N_12756,N_12125,N_12349);
nand U12757 (N_12757,N_12436,N_12433);
or U12758 (N_12758,N_12467,N_12099);
and U12759 (N_12759,N_12346,N_12099);
and U12760 (N_12760,N_12194,N_12139);
and U12761 (N_12761,N_12299,N_12333);
or U12762 (N_12762,N_12175,N_12061);
and U12763 (N_12763,N_12029,N_12266);
nor U12764 (N_12764,N_12336,N_12113);
nand U12765 (N_12765,N_12190,N_12483);
nor U12766 (N_12766,N_12247,N_12293);
and U12767 (N_12767,N_12487,N_12456);
and U12768 (N_12768,N_12040,N_12429);
nor U12769 (N_12769,N_12452,N_12484);
or U12770 (N_12770,N_12463,N_12257);
nand U12771 (N_12771,N_12441,N_12358);
or U12772 (N_12772,N_12083,N_12047);
nor U12773 (N_12773,N_12463,N_12365);
nand U12774 (N_12774,N_12447,N_12318);
and U12775 (N_12775,N_12126,N_12246);
nand U12776 (N_12776,N_12279,N_12223);
nor U12777 (N_12777,N_12256,N_12137);
nor U12778 (N_12778,N_12219,N_12202);
and U12779 (N_12779,N_12391,N_12290);
nor U12780 (N_12780,N_12306,N_12134);
nor U12781 (N_12781,N_12137,N_12453);
or U12782 (N_12782,N_12276,N_12255);
or U12783 (N_12783,N_12028,N_12303);
nor U12784 (N_12784,N_12322,N_12351);
nor U12785 (N_12785,N_12419,N_12074);
or U12786 (N_12786,N_12377,N_12215);
or U12787 (N_12787,N_12298,N_12016);
nand U12788 (N_12788,N_12358,N_12046);
or U12789 (N_12789,N_12307,N_12257);
or U12790 (N_12790,N_12105,N_12164);
and U12791 (N_12791,N_12496,N_12404);
nor U12792 (N_12792,N_12484,N_12329);
nand U12793 (N_12793,N_12079,N_12244);
xnor U12794 (N_12794,N_12127,N_12083);
nand U12795 (N_12795,N_12473,N_12380);
or U12796 (N_12796,N_12421,N_12038);
or U12797 (N_12797,N_12183,N_12403);
nor U12798 (N_12798,N_12273,N_12453);
nand U12799 (N_12799,N_12240,N_12430);
and U12800 (N_12800,N_12390,N_12398);
nor U12801 (N_12801,N_12384,N_12200);
xor U12802 (N_12802,N_12359,N_12091);
and U12803 (N_12803,N_12464,N_12109);
nor U12804 (N_12804,N_12193,N_12264);
xnor U12805 (N_12805,N_12244,N_12304);
and U12806 (N_12806,N_12273,N_12361);
and U12807 (N_12807,N_12152,N_12343);
nand U12808 (N_12808,N_12142,N_12041);
nand U12809 (N_12809,N_12492,N_12438);
nor U12810 (N_12810,N_12200,N_12443);
xor U12811 (N_12811,N_12365,N_12431);
and U12812 (N_12812,N_12317,N_12162);
nand U12813 (N_12813,N_12140,N_12284);
and U12814 (N_12814,N_12286,N_12267);
nand U12815 (N_12815,N_12257,N_12252);
and U12816 (N_12816,N_12241,N_12033);
or U12817 (N_12817,N_12198,N_12194);
nand U12818 (N_12818,N_12485,N_12405);
nand U12819 (N_12819,N_12371,N_12206);
or U12820 (N_12820,N_12237,N_12178);
or U12821 (N_12821,N_12022,N_12476);
nor U12822 (N_12822,N_12493,N_12276);
xor U12823 (N_12823,N_12245,N_12217);
nand U12824 (N_12824,N_12335,N_12339);
and U12825 (N_12825,N_12274,N_12341);
nand U12826 (N_12826,N_12141,N_12016);
nand U12827 (N_12827,N_12470,N_12273);
and U12828 (N_12828,N_12345,N_12373);
nand U12829 (N_12829,N_12190,N_12147);
nor U12830 (N_12830,N_12342,N_12176);
and U12831 (N_12831,N_12085,N_12425);
nand U12832 (N_12832,N_12455,N_12074);
and U12833 (N_12833,N_12391,N_12493);
or U12834 (N_12834,N_12177,N_12248);
nand U12835 (N_12835,N_12340,N_12263);
nor U12836 (N_12836,N_12417,N_12279);
or U12837 (N_12837,N_12483,N_12207);
nor U12838 (N_12838,N_12197,N_12354);
nor U12839 (N_12839,N_12049,N_12213);
nand U12840 (N_12840,N_12366,N_12053);
nor U12841 (N_12841,N_12358,N_12388);
and U12842 (N_12842,N_12137,N_12242);
or U12843 (N_12843,N_12464,N_12214);
and U12844 (N_12844,N_12105,N_12365);
nand U12845 (N_12845,N_12301,N_12042);
and U12846 (N_12846,N_12185,N_12054);
or U12847 (N_12847,N_12120,N_12139);
and U12848 (N_12848,N_12286,N_12241);
and U12849 (N_12849,N_12279,N_12216);
and U12850 (N_12850,N_12486,N_12495);
and U12851 (N_12851,N_12455,N_12458);
nor U12852 (N_12852,N_12393,N_12345);
nand U12853 (N_12853,N_12078,N_12012);
or U12854 (N_12854,N_12056,N_12431);
nor U12855 (N_12855,N_12190,N_12382);
and U12856 (N_12856,N_12090,N_12110);
nor U12857 (N_12857,N_12426,N_12243);
and U12858 (N_12858,N_12369,N_12121);
nand U12859 (N_12859,N_12185,N_12023);
nor U12860 (N_12860,N_12301,N_12193);
nand U12861 (N_12861,N_12332,N_12235);
and U12862 (N_12862,N_12354,N_12303);
and U12863 (N_12863,N_12148,N_12488);
nor U12864 (N_12864,N_12464,N_12085);
or U12865 (N_12865,N_12295,N_12332);
nand U12866 (N_12866,N_12327,N_12099);
nand U12867 (N_12867,N_12300,N_12419);
nor U12868 (N_12868,N_12310,N_12125);
nand U12869 (N_12869,N_12011,N_12235);
or U12870 (N_12870,N_12156,N_12356);
and U12871 (N_12871,N_12304,N_12443);
or U12872 (N_12872,N_12478,N_12324);
or U12873 (N_12873,N_12038,N_12067);
or U12874 (N_12874,N_12364,N_12269);
nand U12875 (N_12875,N_12330,N_12386);
nor U12876 (N_12876,N_12361,N_12244);
and U12877 (N_12877,N_12273,N_12213);
or U12878 (N_12878,N_12302,N_12066);
and U12879 (N_12879,N_12386,N_12085);
nand U12880 (N_12880,N_12299,N_12124);
and U12881 (N_12881,N_12210,N_12269);
and U12882 (N_12882,N_12287,N_12182);
or U12883 (N_12883,N_12127,N_12288);
and U12884 (N_12884,N_12427,N_12205);
and U12885 (N_12885,N_12476,N_12063);
nand U12886 (N_12886,N_12330,N_12122);
nand U12887 (N_12887,N_12394,N_12122);
nand U12888 (N_12888,N_12291,N_12241);
nand U12889 (N_12889,N_12269,N_12101);
nand U12890 (N_12890,N_12464,N_12401);
or U12891 (N_12891,N_12111,N_12287);
or U12892 (N_12892,N_12233,N_12312);
or U12893 (N_12893,N_12198,N_12250);
and U12894 (N_12894,N_12459,N_12047);
or U12895 (N_12895,N_12244,N_12185);
nor U12896 (N_12896,N_12327,N_12483);
or U12897 (N_12897,N_12166,N_12163);
nor U12898 (N_12898,N_12312,N_12234);
xnor U12899 (N_12899,N_12162,N_12335);
and U12900 (N_12900,N_12404,N_12297);
nor U12901 (N_12901,N_12300,N_12234);
and U12902 (N_12902,N_12201,N_12434);
or U12903 (N_12903,N_12065,N_12101);
or U12904 (N_12904,N_12144,N_12338);
xnor U12905 (N_12905,N_12168,N_12123);
and U12906 (N_12906,N_12125,N_12249);
nand U12907 (N_12907,N_12213,N_12088);
nand U12908 (N_12908,N_12393,N_12136);
and U12909 (N_12909,N_12493,N_12129);
and U12910 (N_12910,N_12013,N_12491);
or U12911 (N_12911,N_12271,N_12256);
and U12912 (N_12912,N_12021,N_12492);
and U12913 (N_12913,N_12496,N_12214);
or U12914 (N_12914,N_12067,N_12106);
nand U12915 (N_12915,N_12074,N_12048);
or U12916 (N_12916,N_12239,N_12363);
xor U12917 (N_12917,N_12371,N_12081);
nor U12918 (N_12918,N_12420,N_12158);
or U12919 (N_12919,N_12483,N_12290);
or U12920 (N_12920,N_12217,N_12094);
and U12921 (N_12921,N_12323,N_12056);
nor U12922 (N_12922,N_12173,N_12119);
nor U12923 (N_12923,N_12417,N_12175);
nor U12924 (N_12924,N_12234,N_12432);
or U12925 (N_12925,N_12400,N_12010);
and U12926 (N_12926,N_12424,N_12143);
nor U12927 (N_12927,N_12070,N_12199);
and U12928 (N_12928,N_12382,N_12211);
nor U12929 (N_12929,N_12139,N_12437);
nand U12930 (N_12930,N_12009,N_12470);
nor U12931 (N_12931,N_12242,N_12346);
nand U12932 (N_12932,N_12497,N_12322);
nor U12933 (N_12933,N_12449,N_12056);
or U12934 (N_12934,N_12237,N_12111);
or U12935 (N_12935,N_12397,N_12291);
xnor U12936 (N_12936,N_12456,N_12413);
xnor U12937 (N_12937,N_12171,N_12301);
nand U12938 (N_12938,N_12001,N_12487);
and U12939 (N_12939,N_12223,N_12439);
or U12940 (N_12940,N_12260,N_12089);
and U12941 (N_12941,N_12292,N_12469);
nand U12942 (N_12942,N_12373,N_12258);
nor U12943 (N_12943,N_12164,N_12331);
nand U12944 (N_12944,N_12063,N_12462);
and U12945 (N_12945,N_12080,N_12359);
or U12946 (N_12946,N_12007,N_12008);
or U12947 (N_12947,N_12432,N_12331);
nor U12948 (N_12948,N_12252,N_12230);
xor U12949 (N_12949,N_12309,N_12449);
nand U12950 (N_12950,N_12498,N_12201);
and U12951 (N_12951,N_12222,N_12405);
and U12952 (N_12952,N_12338,N_12288);
and U12953 (N_12953,N_12162,N_12043);
or U12954 (N_12954,N_12168,N_12074);
nand U12955 (N_12955,N_12410,N_12289);
nand U12956 (N_12956,N_12097,N_12217);
nand U12957 (N_12957,N_12203,N_12455);
nor U12958 (N_12958,N_12050,N_12370);
nand U12959 (N_12959,N_12316,N_12167);
nand U12960 (N_12960,N_12276,N_12302);
nor U12961 (N_12961,N_12397,N_12062);
and U12962 (N_12962,N_12213,N_12225);
and U12963 (N_12963,N_12112,N_12162);
nor U12964 (N_12964,N_12474,N_12448);
or U12965 (N_12965,N_12138,N_12452);
nor U12966 (N_12966,N_12328,N_12331);
and U12967 (N_12967,N_12206,N_12139);
or U12968 (N_12968,N_12260,N_12436);
or U12969 (N_12969,N_12375,N_12420);
and U12970 (N_12970,N_12471,N_12076);
and U12971 (N_12971,N_12151,N_12342);
nand U12972 (N_12972,N_12201,N_12310);
nand U12973 (N_12973,N_12485,N_12003);
and U12974 (N_12974,N_12039,N_12496);
nor U12975 (N_12975,N_12103,N_12098);
and U12976 (N_12976,N_12116,N_12269);
nor U12977 (N_12977,N_12243,N_12221);
nand U12978 (N_12978,N_12083,N_12357);
nand U12979 (N_12979,N_12039,N_12327);
and U12980 (N_12980,N_12192,N_12178);
or U12981 (N_12981,N_12414,N_12466);
xnor U12982 (N_12982,N_12266,N_12175);
nor U12983 (N_12983,N_12071,N_12229);
and U12984 (N_12984,N_12474,N_12027);
and U12985 (N_12985,N_12351,N_12491);
and U12986 (N_12986,N_12265,N_12068);
or U12987 (N_12987,N_12447,N_12255);
and U12988 (N_12988,N_12055,N_12261);
or U12989 (N_12989,N_12136,N_12040);
or U12990 (N_12990,N_12158,N_12150);
nor U12991 (N_12991,N_12092,N_12083);
or U12992 (N_12992,N_12372,N_12058);
nand U12993 (N_12993,N_12487,N_12097);
and U12994 (N_12994,N_12489,N_12365);
and U12995 (N_12995,N_12478,N_12334);
nor U12996 (N_12996,N_12055,N_12457);
xor U12997 (N_12997,N_12283,N_12304);
and U12998 (N_12998,N_12406,N_12044);
nor U12999 (N_12999,N_12483,N_12015);
and U13000 (N_13000,N_12503,N_12734);
nand U13001 (N_13001,N_12682,N_12733);
nor U13002 (N_13002,N_12901,N_12980);
nand U13003 (N_13003,N_12654,N_12889);
nor U13004 (N_13004,N_12912,N_12863);
nand U13005 (N_13005,N_12514,N_12783);
and U13006 (N_13006,N_12862,N_12669);
and U13007 (N_13007,N_12976,N_12743);
or U13008 (N_13008,N_12906,N_12642);
nand U13009 (N_13009,N_12721,N_12577);
nor U13010 (N_13010,N_12678,N_12681);
and U13011 (N_13011,N_12575,N_12967);
and U13012 (N_13012,N_12811,N_12596);
nor U13013 (N_13013,N_12739,N_12786);
or U13014 (N_13014,N_12991,N_12799);
or U13015 (N_13015,N_12515,N_12546);
or U13016 (N_13016,N_12689,N_12968);
nand U13017 (N_13017,N_12572,N_12939);
nand U13018 (N_13018,N_12926,N_12886);
nor U13019 (N_13019,N_12717,N_12639);
xnor U13020 (N_13020,N_12970,N_12581);
nor U13021 (N_13021,N_12608,N_12938);
or U13022 (N_13022,N_12684,N_12606);
nand U13023 (N_13023,N_12561,N_12955);
xor U13024 (N_13024,N_12807,N_12512);
or U13025 (N_13025,N_12957,N_12533);
xnor U13026 (N_13026,N_12550,N_12853);
and U13027 (N_13027,N_12997,N_12604);
nand U13028 (N_13028,N_12999,N_12752);
nand U13029 (N_13029,N_12929,N_12992);
xor U13030 (N_13030,N_12755,N_12990);
nand U13031 (N_13031,N_12709,N_12907);
nor U13032 (N_13032,N_12539,N_12788);
nor U13033 (N_13033,N_12825,N_12890);
xor U13034 (N_13034,N_12954,N_12824);
nand U13035 (N_13035,N_12756,N_12768);
or U13036 (N_13036,N_12645,N_12818);
or U13037 (N_13037,N_12802,N_12795);
or U13038 (N_13038,N_12838,N_12896);
nor U13039 (N_13039,N_12944,N_12918);
and U13040 (N_13040,N_12854,N_12844);
or U13041 (N_13041,N_12961,N_12949);
nor U13042 (N_13042,N_12979,N_12930);
nor U13043 (N_13043,N_12840,N_12599);
nor U13044 (N_13044,N_12615,N_12568);
nor U13045 (N_13045,N_12507,N_12866);
nand U13046 (N_13046,N_12777,N_12774);
or U13047 (N_13047,N_12859,N_12611);
nand U13048 (N_13048,N_12922,N_12917);
and U13049 (N_13049,N_12765,N_12660);
or U13050 (N_13050,N_12775,N_12751);
nand U13051 (N_13051,N_12879,N_12500);
or U13052 (N_13052,N_12989,N_12827);
and U13053 (N_13053,N_12839,N_12972);
nor U13054 (N_13054,N_12624,N_12842);
and U13055 (N_13055,N_12952,N_12760);
and U13056 (N_13056,N_12740,N_12644);
xnor U13057 (N_13057,N_12510,N_12711);
and U13058 (N_13058,N_12509,N_12594);
xnor U13059 (N_13059,N_12796,N_12536);
nor U13060 (N_13060,N_12753,N_12958);
nand U13061 (N_13061,N_12580,N_12610);
and U13062 (N_13062,N_12663,N_12826);
nand U13063 (N_13063,N_12529,N_12694);
nor U13064 (N_13064,N_12987,N_12877);
and U13065 (N_13065,N_12903,N_12787);
nand U13066 (N_13066,N_12659,N_12592);
nor U13067 (N_13067,N_12962,N_12705);
nor U13068 (N_13068,N_12505,N_12723);
nor U13069 (N_13069,N_12937,N_12549);
nand U13070 (N_13070,N_12563,N_12932);
nor U13071 (N_13071,N_12870,N_12857);
nor U13072 (N_13072,N_12523,N_12762);
nand U13073 (N_13073,N_12649,N_12819);
nand U13074 (N_13074,N_12770,N_12766);
nand U13075 (N_13075,N_12746,N_12915);
or U13076 (N_13076,N_12526,N_12865);
nand U13077 (N_13077,N_12916,N_12813);
and U13078 (N_13078,N_12833,N_12931);
and U13079 (N_13079,N_12612,N_12789);
nor U13080 (N_13080,N_12562,N_12714);
and U13081 (N_13081,N_12548,N_12666);
or U13082 (N_13082,N_12727,N_12693);
and U13083 (N_13083,N_12782,N_12994);
nand U13084 (N_13084,N_12506,N_12908);
nor U13085 (N_13085,N_12969,N_12983);
nand U13086 (N_13086,N_12633,N_12758);
nor U13087 (N_13087,N_12974,N_12793);
nand U13088 (N_13088,N_12810,N_12590);
or U13089 (N_13089,N_12812,N_12898);
nand U13090 (N_13090,N_12528,N_12587);
nand U13091 (N_13091,N_12545,N_12704);
nor U13092 (N_13092,N_12888,N_12892);
nor U13093 (N_13093,N_12626,N_12518);
or U13094 (N_13094,N_12557,N_12643);
nand U13095 (N_13095,N_12532,N_12894);
or U13096 (N_13096,N_12607,N_12832);
and U13097 (N_13097,N_12715,N_12982);
nor U13098 (N_13098,N_12609,N_12924);
nor U13099 (N_13099,N_12502,N_12530);
and U13100 (N_13100,N_12686,N_12692);
nor U13101 (N_13101,N_12848,N_12623);
nor U13102 (N_13102,N_12656,N_12946);
and U13103 (N_13103,N_12593,N_12700);
nand U13104 (N_13104,N_12736,N_12747);
nor U13105 (N_13105,N_12618,N_12657);
nand U13106 (N_13106,N_12614,N_12801);
nand U13107 (N_13107,N_12951,N_12790);
nor U13108 (N_13108,N_12570,N_12638);
nor U13109 (N_13109,N_12792,N_12525);
nand U13110 (N_13110,N_12621,N_12835);
and U13111 (N_13111,N_12841,N_12828);
and U13112 (N_13112,N_12672,N_12584);
nor U13113 (N_13113,N_12662,N_12820);
nor U13114 (N_13114,N_12710,N_12628);
nor U13115 (N_13115,N_12742,N_12858);
xnor U13116 (N_13116,N_12869,N_12749);
nor U13117 (N_13117,N_12874,N_12647);
nor U13118 (N_13118,N_12978,N_12551);
and U13119 (N_13119,N_12808,N_12920);
nand U13120 (N_13120,N_12941,N_12757);
nand U13121 (N_13121,N_12847,N_12670);
or U13122 (N_13122,N_12578,N_12966);
or U13123 (N_13123,N_12933,N_12867);
nand U13124 (N_13124,N_12893,N_12535);
nand U13125 (N_13125,N_12873,N_12861);
or U13126 (N_13126,N_12583,N_12542);
nand U13127 (N_13127,N_12527,N_12846);
nor U13128 (N_13128,N_12959,N_12940);
or U13129 (N_13129,N_12695,N_12794);
or U13130 (N_13130,N_12636,N_12560);
nand U13131 (N_13131,N_12652,N_12665);
nor U13132 (N_13132,N_12914,N_12803);
and U13133 (N_13133,N_12555,N_12698);
nand U13134 (N_13134,N_12516,N_12911);
and U13135 (N_13135,N_12702,N_12771);
nand U13136 (N_13136,N_12701,N_12860);
nor U13137 (N_13137,N_12830,N_12683);
or U13138 (N_13138,N_12823,N_12664);
and U13139 (N_13139,N_12817,N_12910);
and U13140 (N_13140,N_12691,N_12696);
nor U13141 (N_13141,N_12759,N_12960);
nor U13142 (N_13142,N_12754,N_12541);
xor U13143 (N_13143,N_12646,N_12620);
nand U13144 (N_13144,N_12619,N_12556);
or U13145 (N_13145,N_12852,N_12804);
nand U13146 (N_13146,N_12741,N_12780);
and U13147 (N_13147,N_12935,N_12745);
or U13148 (N_13148,N_12945,N_12781);
nor U13149 (N_13149,N_12868,N_12772);
or U13150 (N_13150,N_12653,N_12637);
nor U13151 (N_13151,N_12569,N_12554);
and U13152 (N_13152,N_12631,N_12885);
nor U13153 (N_13153,N_12534,N_12688);
nand U13154 (N_13154,N_12522,N_12806);
nand U13155 (N_13155,N_12719,N_12553);
and U13156 (N_13156,N_12845,N_12680);
or U13157 (N_13157,N_12778,N_12899);
nor U13158 (N_13158,N_12591,N_12928);
nor U13159 (N_13159,N_12750,N_12995);
nand U13160 (N_13160,N_12735,N_12690);
and U13161 (N_13161,N_12558,N_12779);
nand U13162 (N_13162,N_12730,N_12891);
or U13163 (N_13163,N_12658,N_12773);
nor U13164 (N_13164,N_12737,N_12586);
and U13165 (N_13165,N_12634,N_12965);
and U13166 (N_13166,N_12708,N_12785);
nor U13167 (N_13167,N_12707,N_12998);
nor U13168 (N_13168,N_12720,N_12630);
and U13169 (N_13169,N_12687,N_12520);
nand U13170 (N_13170,N_12981,N_12504);
nand U13171 (N_13171,N_12876,N_12576);
or U13172 (N_13172,N_12511,N_12724);
nand U13173 (N_13173,N_12871,N_12597);
xnor U13174 (N_13174,N_12769,N_12531);
nor U13175 (N_13175,N_12884,N_12718);
and U13176 (N_13176,N_12573,N_12988);
and U13177 (N_13177,N_12763,N_12963);
nand U13178 (N_13178,N_12685,N_12947);
nand U13179 (N_13179,N_12934,N_12517);
or U13180 (N_13180,N_12800,N_12521);
and U13181 (N_13181,N_12677,N_12601);
and U13182 (N_13182,N_12950,N_12831);
or U13183 (N_13183,N_12872,N_12864);
and U13184 (N_13184,N_12722,N_12559);
or U13185 (N_13185,N_12895,N_12815);
nor U13186 (N_13186,N_12851,N_12501);
nor U13187 (N_13187,N_12699,N_12613);
and U13188 (N_13188,N_12882,N_12519);
nor U13189 (N_13189,N_12798,N_12964);
nor U13190 (N_13190,N_12834,N_12728);
or U13191 (N_13191,N_12679,N_12821);
nand U13192 (N_13192,N_12706,N_12641);
and U13193 (N_13193,N_12887,N_12971);
nand U13194 (N_13194,N_12668,N_12675);
nor U13195 (N_13195,N_12880,N_12881);
xor U13196 (N_13196,N_12676,N_12977);
and U13197 (N_13197,N_12805,N_12674);
nand U13198 (N_13198,N_12565,N_12716);
nand U13199 (N_13199,N_12598,N_12936);
and U13200 (N_13200,N_12673,N_12849);
nor U13201 (N_13201,N_12927,N_12843);
nand U13202 (N_13202,N_12567,N_12797);
and U13203 (N_13203,N_12629,N_12875);
and U13204 (N_13204,N_12632,N_12897);
and U13205 (N_13205,N_12791,N_12524);
and U13206 (N_13206,N_12809,N_12761);
nor U13207 (N_13207,N_12725,N_12574);
nor U13208 (N_13208,N_12953,N_12996);
nand U13209 (N_13209,N_12640,N_12776);
or U13210 (N_13210,N_12732,N_12712);
nor U13211 (N_13211,N_12921,N_12850);
nor U13212 (N_13212,N_12731,N_12588);
nor U13213 (N_13213,N_12571,N_12605);
and U13214 (N_13214,N_12985,N_12595);
nand U13215 (N_13215,N_12973,N_12902);
nor U13216 (N_13216,N_12617,N_12589);
or U13217 (N_13217,N_12814,N_12540);
or U13218 (N_13218,N_12919,N_12671);
nor U13219 (N_13219,N_12942,N_12622);
or U13220 (N_13220,N_12508,N_12855);
nand U13221 (N_13221,N_12837,N_12905);
or U13222 (N_13222,N_12543,N_12651);
nand U13223 (N_13223,N_12956,N_12748);
nor U13224 (N_13224,N_12713,N_12585);
nand U13225 (N_13225,N_12744,N_12764);
nor U13226 (N_13226,N_12661,N_12547);
and U13227 (N_13227,N_12697,N_12625);
and U13228 (N_13228,N_12729,N_12909);
nor U13229 (N_13229,N_12726,N_12767);
and U13230 (N_13230,N_12784,N_12738);
and U13231 (N_13231,N_12822,N_12602);
or U13232 (N_13232,N_12900,N_12635);
or U13233 (N_13233,N_12913,N_12600);
and U13234 (N_13234,N_12650,N_12943);
or U13235 (N_13235,N_12538,N_12986);
nor U13236 (N_13236,N_12904,N_12836);
nor U13237 (N_13237,N_12648,N_12582);
xor U13238 (N_13238,N_12984,N_12703);
or U13239 (N_13239,N_12655,N_12948);
xnor U13240 (N_13240,N_12856,N_12975);
and U13241 (N_13241,N_12513,N_12616);
nand U13242 (N_13242,N_12564,N_12816);
or U13243 (N_13243,N_12667,N_12923);
and U13244 (N_13244,N_12883,N_12829);
and U13245 (N_13245,N_12627,N_12925);
xnor U13246 (N_13246,N_12878,N_12566);
and U13247 (N_13247,N_12552,N_12544);
and U13248 (N_13248,N_12993,N_12603);
or U13249 (N_13249,N_12579,N_12537);
nand U13250 (N_13250,N_12922,N_12753);
and U13251 (N_13251,N_12681,N_12632);
nor U13252 (N_13252,N_12939,N_12966);
nor U13253 (N_13253,N_12922,N_12513);
nand U13254 (N_13254,N_12902,N_12554);
and U13255 (N_13255,N_12780,N_12774);
or U13256 (N_13256,N_12737,N_12992);
or U13257 (N_13257,N_12649,N_12616);
or U13258 (N_13258,N_12975,N_12966);
nor U13259 (N_13259,N_12761,N_12909);
nor U13260 (N_13260,N_12620,N_12811);
or U13261 (N_13261,N_12750,N_12968);
nor U13262 (N_13262,N_12818,N_12506);
and U13263 (N_13263,N_12546,N_12782);
nand U13264 (N_13264,N_12663,N_12637);
nor U13265 (N_13265,N_12615,N_12897);
and U13266 (N_13266,N_12618,N_12974);
or U13267 (N_13267,N_12750,N_12797);
and U13268 (N_13268,N_12532,N_12813);
and U13269 (N_13269,N_12578,N_12637);
nor U13270 (N_13270,N_12545,N_12858);
nor U13271 (N_13271,N_12690,N_12764);
and U13272 (N_13272,N_12700,N_12531);
nor U13273 (N_13273,N_12846,N_12711);
nor U13274 (N_13274,N_12912,N_12870);
or U13275 (N_13275,N_12883,N_12923);
nor U13276 (N_13276,N_12946,N_12927);
nor U13277 (N_13277,N_12711,N_12853);
nand U13278 (N_13278,N_12945,N_12641);
nand U13279 (N_13279,N_12702,N_12919);
nor U13280 (N_13280,N_12680,N_12826);
nand U13281 (N_13281,N_12857,N_12699);
xnor U13282 (N_13282,N_12777,N_12780);
nor U13283 (N_13283,N_12716,N_12879);
nand U13284 (N_13284,N_12562,N_12827);
nand U13285 (N_13285,N_12944,N_12788);
or U13286 (N_13286,N_12544,N_12569);
nand U13287 (N_13287,N_12989,N_12885);
nor U13288 (N_13288,N_12669,N_12713);
nor U13289 (N_13289,N_12728,N_12749);
nand U13290 (N_13290,N_12744,N_12755);
or U13291 (N_13291,N_12794,N_12564);
nand U13292 (N_13292,N_12551,N_12614);
nor U13293 (N_13293,N_12588,N_12892);
and U13294 (N_13294,N_12601,N_12800);
nand U13295 (N_13295,N_12501,N_12893);
and U13296 (N_13296,N_12690,N_12625);
xnor U13297 (N_13297,N_12685,N_12776);
and U13298 (N_13298,N_12767,N_12967);
nor U13299 (N_13299,N_12817,N_12975);
and U13300 (N_13300,N_12926,N_12796);
nand U13301 (N_13301,N_12690,N_12602);
nor U13302 (N_13302,N_12580,N_12627);
nand U13303 (N_13303,N_12706,N_12914);
or U13304 (N_13304,N_12747,N_12944);
or U13305 (N_13305,N_12948,N_12715);
nand U13306 (N_13306,N_12912,N_12596);
nand U13307 (N_13307,N_12735,N_12996);
nor U13308 (N_13308,N_12929,N_12896);
or U13309 (N_13309,N_12932,N_12623);
nand U13310 (N_13310,N_12870,N_12791);
nand U13311 (N_13311,N_12656,N_12851);
nor U13312 (N_13312,N_12539,N_12617);
nand U13313 (N_13313,N_12701,N_12512);
nor U13314 (N_13314,N_12707,N_12654);
and U13315 (N_13315,N_12796,N_12945);
or U13316 (N_13316,N_12520,N_12997);
or U13317 (N_13317,N_12622,N_12594);
nand U13318 (N_13318,N_12809,N_12953);
and U13319 (N_13319,N_12556,N_12509);
nand U13320 (N_13320,N_12688,N_12549);
nand U13321 (N_13321,N_12663,N_12973);
and U13322 (N_13322,N_12727,N_12825);
and U13323 (N_13323,N_12694,N_12540);
or U13324 (N_13324,N_12841,N_12766);
and U13325 (N_13325,N_12702,N_12965);
and U13326 (N_13326,N_12999,N_12710);
and U13327 (N_13327,N_12501,N_12582);
and U13328 (N_13328,N_12611,N_12744);
and U13329 (N_13329,N_12642,N_12825);
and U13330 (N_13330,N_12677,N_12935);
xnor U13331 (N_13331,N_12589,N_12537);
or U13332 (N_13332,N_12650,N_12994);
nand U13333 (N_13333,N_12796,N_12500);
or U13334 (N_13334,N_12876,N_12731);
nor U13335 (N_13335,N_12510,N_12969);
nand U13336 (N_13336,N_12661,N_12837);
and U13337 (N_13337,N_12755,N_12842);
and U13338 (N_13338,N_12922,N_12911);
and U13339 (N_13339,N_12536,N_12648);
nand U13340 (N_13340,N_12862,N_12791);
or U13341 (N_13341,N_12705,N_12900);
or U13342 (N_13342,N_12748,N_12750);
nand U13343 (N_13343,N_12968,N_12603);
or U13344 (N_13344,N_12952,N_12814);
nand U13345 (N_13345,N_12983,N_12879);
nand U13346 (N_13346,N_12683,N_12764);
or U13347 (N_13347,N_12939,N_12796);
nor U13348 (N_13348,N_12928,N_12691);
or U13349 (N_13349,N_12955,N_12536);
or U13350 (N_13350,N_12969,N_12768);
and U13351 (N_13351,N_12628,N_12918);
nand U13352 (N_13352,N_12827,N_12742);
nand U13353 (N_13353,N_12558,N_12881);
xor U13354 (N_13354,N_12767,N_12916);
nor U13355 (N_13355,N_12685,N_12546);
and U13356 (N_13356,N_12692,N_12653);
nor U13357 (N_13357,N_12541,N_12695);
or U13358 (N_13358,N_12719,N_12670);
and U13359 (N_13359,N_12755,N_12700);
and U13360 (N_13360,N_12829,N_12692);
or U13361 (N_13361,N_12649,N_12566);
nor U13362 (N_13362,N_12749,N_12736);
nor U13363 (N_13363,N_12619,N_12528);
and U13364 (N_13364,N_12672,N_12538);
and U13365 (N_13365,N_12542,N_12945);
nand U13366 (N_13366,N_12866,N_12629);
or U13367 (N_13367,N_12761,N_12706);
or U13368 (N_13368,N_12970,N_12823);
nor U13369 (N_13369,N_12723,N_12946);
nor U13370 (N_13370,N_12512,N_12541);
or U13371 (N_13371,N_12663,N_12627);
nand U13372 (N_13372,N_12681,N_12813);
and U13373 (N_13373,N_12837,N_12503);
or U13374 (N_13374,N_12964,N_12649);
nand U13375 (N_13375,N_12504,N_12900);
nor U13376 (N_13376,N_12517,N_12884);
nor U13377 (N_13377,N_12834,N_12601);
and U13378 (N_13378,N_12751,N_12859);
or U13379 (N_13379,N_12966,N_12973);
xor U13380 (N_13380,N_12671,N_12567);
nor U13381 (N_13381,N_12513,N_12686);
or U13382 (N_13382,N_12609,N_12831);
nand U13383 (N_13383,N_12728,N_12977);
or U13384 (N_13384,N_12945,N_12506);
nor U13385 (N_13385,N_12508,N_12901);
and U13386 (N_13386,N_12713,N_12647);
or U13387 (N_13387,N_12785,N_12534);
or U13388 (N_13388,N_12510,N_12942);
or U13389 (N_13389,N_12883,N_12742);
and U13390 (N_13390,N_12822,N_12765);
or U13391 (N_13391,N_12632,N_12969);
nand U13392 (N_13392,N_12745,N_12855);
and U13393 (N_13393,N_12597,N_12819);
and U13394 (N_13394,N_12656,N_12599);
and U13395 (N_13395,N_12639,N_12790);
or U13396 (N_13396,N_12668,N_12701);
or U13397 (N_13397,N_12990,N_12876);
nand U13398 (N_13398,N_12557,N_12720);
nor U13399 (N_13399,N_12577,N_12955);
and U13400 (N_13400,N_12675,N_12998);
or U13401 (N_13401,N_12649,N_12589);
nor U13402 (N_13402,N_12620,N_12972);
nand U13403 (N_13403,N_12958,N_12764);
nand U13404 (N_13404,N_12543,N_12711);
or U13405 (N_13405,N_12719,N_12806);
nand U13406 (N_13406,N_12997,N_12763);
or U13407 (N_13407,N_12546,N_12649);
nand U13408 (N_13408,N_12927,N_12816);
nand U13409 (N_13409,N_12914,N_12728);
or U13410 (N_13410,N_12646,N_12523);
and U13411 (N_13411,N_12744,N_12980);
or U13412 (N_13412,N_12949,N_12739);
nand U13413 (N_13413,N_12694,N_12832);
nor U13414 (N_13414,N_12501,N_12839);
or U13415 (N_13415,N_12857,N_12575);
or U13416 (N_13416,N_12717,N_12733);
nand U13417 (N_13417,N_12742,N_12816);
and U13418 (N_13418,N_12753,N_12674);
nor U13419 (N_13419,N_12524,N_12854);
or U13420 (N_13420,N_12880,N_12790);
and U13421 (N_13421,N_12945,N_12922);
and U13422 (N_13422,N_12979,N_12549);
nand U13423 (N_13423,N_12900,N_12864);
nand U13424 (N_13424,N_12802,N_12523);
xnor U13425 (N_13425,N_12892,N_12574);
and U13426 (N_13426,N_12720,N_12843);
and U13427 (N_13427,N_12890,N_12921);
nand U13428 (N_13428,N_12631,N_12513);
or U13429 (N_13429,N_12857,N_12939);
nor U13430 (N_13430,N_12644,N_12508);
and U13431 (N_13431,N_12694,N_12993);
nor U13432 (N_13432,N_12601,N_12630);
nor U13433 (N_13433,N_12916,N_12612);
nor U13434 (N_13434,N_12653,N_12582);
nor U13435 (N_13435,N_12792,N_12720);
or U13436 (N_13436,N_12864,N_12941);
and U13437 (N_13437,N_12620,N_12569);
or U13438 (N_13438,N_12790,N_12811);
or U13439 (N_13439,N_12565,N_12948);
and U13440 (N_13440,N_12937,N_12540);
and U13441 (N_13441,N_12948,N_12961);
nor U13442 (N_13442,N_12827,N_12976);
nor U13443 (N_13443,N_12889,N_12566);
or U13444 (N_13444,N_12848,N_12869);
or U13445 (N_13445,N_12981,N_12968);
and U13446 (N_13446,N_12647,N_12681);
and U13447 (N_13447,N_12839,N_12983);
nor U13448 (N_13448,N_12720,N_12853);
xor U13449 (N_13449,N_12786,N_12974);
or U13450 (N_13450,N_12526,N_12672);
or U13451 (N_13451,N_12996,N_12886);
and U13452 (N_13452,N_12963,N_12574);
xnor U13453 (N_13453,N_12502,N_12630);
xor U13454 (N_13454,N_12976,N_12782);
nor U13455 (N_13455,N_12741,N_12516);
nor U13456 (N_13456,N_12764,N_12603);
nor U13457 (N_13457,N_12825,N_12775);
nor U13458 (N_13458,N_12617,N_12948);
nand U13459 (N_13459,N_12840,N_12573);
and U13460 (N_13460,N_12581,N_12765);
nor U13461 (N_13461,N_12890,N_12873);
nor U13462 (N_13462,N_12527,N_12774);
nand U13463 (N_13463,N_12749,N_12976);
nand U13464 (N_13464,N_12795,N_12542);
nand U13465 (N_13465,N_12634,N_12729);
and U13466 (N_13466,N_12834,N_12956);
or U13467 (N_13467,N_12544,N_12618);
nor U13468 (N_13468,N_12594,N_12809);
and U13469 (N_13469,N_12805,N_12798);
and U13470 (N_13470,N_12923,N_12646);
or U13471 (N_13471,N_12694,N_12722);
and U13472 (N_13472,N_12515,N_12880);
or U13473 (N_13473,N_12898,N_12874);
nand U13474 (N_13474,N_12627,N_12771);
or U13475 (N_13475,N_12590,N_12893);
or U13476 (N_13476,N_12896,N_12794);
nor U13477 (N_13477,N_12610,N_12661);
and U13478 (N_13478,N_12679,N_12973);
nand U13479 (N_13479,N_12972,N_12527);
nor U13480 (N_13480,N_12981,N_12605);
nor U13481 (N_13481,N_12521,N_12732);
nor U13482 (N_13482,N_12998,N_12852);
nor U13483 (N_13483,N_12784,N_12596);
and U13484 (N_13484,N_12641,N_12946);
or U13485 (N_13485,N_12922,N_12791);
nor U13486 (N_13486,N_12763,N_12646);
and U13487 (N_13487,N_12661,N_12929);
or U13488 (N_13488,N_12635,N_12820);
and U13489 (N_13489,N_12694,N_12876);
and U13490 (N_13490,N_12981,N_12530);
nand U13491 (N_13491,N_12583,N_12569);
nor U13492 (N_13492,N_12942,N_12761);
or U13493 (N_13493,N_12552,N_12546);
or U13494 (N_13494,N_12844,N_12556);
nand U13495 (N_13495,N_12605,N_12970);
nand U13496 (N_13496,N_12963,N_12650);
or U13497 (N_13497,N_12939,N_12711);
nand U13498 (N_13498,N_12912,N_12602);
and U13499 (N_13499,N_12967,N_12610);
nand U13500 (N_13500,N_13039,N_13274);
nor U13501 (N_13501,N_13165,N_13291);
nand U13502 (N_13502,N_13468,N_13390);
nand U13503 (N_13503,N_13445,N_13436);
or U13504 (N_13504,N_13391,N_13011);
nand U13505 (N_13505,N_13371,N_13079);
nor U13506 (N_13506,N_13180,N_13042);
nand U13507 (N_13507,N_13377,N_13097);
or U13508 (N_13508,N_13401,N_13145);
and U13509 (N_13509,N_13238,N_13398);
and U13510 (N_13510,N_13091,N_13077);
and U13511 (N_13511,N_13218,N_13177);
nor U13512 (N_13512,N_13441,N_13214);
and U13513 (N_13513,N_13296,N_13240);
nand U13514 (N_13514,N_13276,N_13063);
or U13515 (N_13515,N_13169,N_13173);
and U13516 (N_13516,N_13175,N_13481);
nand U13517 (N_13517,N_13243,N_13161);
nand U13518 (N_13518,N_13285,N_13379);
xnor U13519 (N_13519,N_13256,N_13029);
and U13520 (N_13520,N_13034,N_13031);
nand U13521 (N_13521,N_13139,N_13208);
nand U13522 (N_13522,N_13216,N_13052);
nor U13523 (N_13523,N_13469,N_13232);
and U13524 (N_13524,N_13115,N_13096);
or U13525 (N_13525,N_13466,N_13373);
nand U13526 (N_13526,N_13267,N_13261);
nor U13527 (N_13527,N_13100,N_13168);
nor U13528 (N_13528,N_13114,N_13176);
or U13529 (N_13529,N_13473,N_13319);
nor U13530 (N_13530,N_13066,N_13086);
and U13531 (N_13531,N_13082,N_13278);
or U13532 (N_13532,N_13056,N_13016);
xnor U13533 (N_13533,N_13032,N_13498);
nor U13534 (N_13534,N_13040,N_13370);
nand U13535 (N_13535,N_13340,N_13084);
nand U13536 (N_13536,N_13041,N_13116);
or U13537 (N_13537,N_13048,N_13435);
and U13538 (N_13538,N_13144,N_13088);
and U13539 (N_13539,N_13230,N_13426);
and U13540 (N_13540,N_13229,N_13123);
nor U13541 (N_13541,N_13212,N_13157);
nor U13542 (N_13542,N_13375,N_13258);
or U13543 (N_13543,N_13292,N_13260);
nand U13544 (N_13544,N_13448,N_13148);
nor U13545 (N_13545,N_13110,N_13252);
and U13546 (N_13546,N_13234,N_13002);
nand U13547 (N_13547,N_13217,N_13492);
and U13548 (N_13548,N_13158,N_13433);
and U13549 (N_13549,N_13223,N_13211);
or U13550 (N_13550,N_13081,N_13221);
nand U13551 (N_13551,N_13428,N_13247);
or U13552 (N_13552,N_13359,N_13366);
or U13553 (N_13553,N_13486,N_13017);
and U13554 (N_13554,N_13010,N_13156);
or U13555 (N_13555,N_13182,N_13287);
or U13556 (N_13556,N_13461,N_13255);
or U13557 (N_13557,N_13494,N_13027);
or U13558 (N_13558,N_13421,N_13194);
nor U13559 (N_13559,N_13417,N_13474);
nor U13560 (N_13560,N_13045,N_13286);
xor U13561 (N_13561,N_13279,N_13204);
or U13562 (N_13562,N_13118,N_13069);
nand U13563 (N_13563,N_13351,N_13430);
or U13564 (N_13564,N_13272,N_13119);
and U13565 (N_13565,N_13389,N_13477);
xnor U13566 (N_13566,N_13480,N_13416);
or U13567 (N_13567,N_13344,N_13135);
nand U13568 (N_13568,N_13320,N_13423);
and U13569 (N_13569,N_13155,N_13478);
or U13570 (N_13570,N_13326,N_13284);
or U13571 (N_13571,N_13363,N_13248);
or U13572 (N_13572,N_13227,N_13308);
and U13573 (N_13573,N_13266,N_13269);
nor U13574 (N_13574,N_13209,N_13452);
and U13575 (N_13575,N_13089,N_13178);
nand U13576 (N_13576,N_13313,N_13304);
nor U13577 (N_13577,N_13275,N_13489);
nor U13578 (N_13578,N_13050,N_13338);
and U13579 (N_13579,N_13087,N_13303);
or U13580 (N_13580,N_13244,N_13397);
or U13581 (N_13581,N_13254,N_13321);
and U13582 (N_13582,N_13044,N_13183);
and U13583 (N_13583,N_13455,N_13404);
and U13584 (N_13584,N_13021,N_13413);
or U13585 (N_13585,N_13402,N_13093);
or U13586 (N_13586,N_13141,N_13008);
nand U13587 (N_13587,N_13309,N_13047);
nand U13588 (N_13588,N_13219,N_13072);
nor U13589 (N_13589,N_13190,N_13378);
or U13590 (N_13590,N_13293,N_13064);
nand U13591 (N_13591,N_13387,N_13405);
nor U13592 (N_13592,N_13264,N_13277);
nand U13593 (N_13593,N_13488,N_13393);
and U13594 (N_13594,N_13015,N_13483);
and U13595 (N_13595,N_13409,N_13419);
nand U13596 (N_13596,N_13470,N_13280);
nor U13597 (N_13597,N_13347,N_13497);
or U13598 (N_13598,N_13224,N_13271);
nand U13599 (N_13599,N_13418,N_13174);
or U13600 (N_13600,N_13225,N_13111);
or U13601 (N_13601,N_13080,N_13289);
or U13602 (N_13602,N_13228,N_13226);
nand U13603 (N_13603,N_13410,N_13236);
and U13604 (N_13604,N_13137,N_13130);
nand U13605 (N_13605,N_13472,N_13235);
or U13606 (N_13606,N_13198,N_13439);
nand U13607 (N_13607,N_13490,N_13432);
nand U13608 (N_13608,N_13476,N_13457);
or U13609 (N_13609,N_13000,N_13411);
nor U13610 (N_13610,N_13210,N_13049);
and U13611 (N_13611,N_13188,N_13202);
nand U13612 (N_13612,N_13171,N_13364);
nand U13613 (N_13613,N_13456,N_13342);
nand U13614 (N_13614,N_13310,N_13067);
nand U13615 (N_13615,N_13388,N_13153);
nand U13616 (N_13616,N_13160,N_13143);
nand U13617 (N_13617,N_13462,N_13443);
nand U13618 (N_13618,N_13330,N_13458);
and U13619 (N_13619,N_13181,N_13055);
or U13620 (N_13620,N_13120,N_13147);
nand U13621 (N_13621,N_13140,N_13288);
nand U13622 (N_13622,N_13249,N_13193);
xor U13623 (N_13623,N_13323,N_13295);
and U13624 (N_13624,N_13487,N_13365);
nor U13625 (N_13625,N_13463,N_13427);
nand U13626 (N_13626,N_13242,N_13400);
and U13627 (N_13627,N_13440,N_13369);
nand U13628 (N_13628,N_13422,N_13028);
or U13629 (N_13629,N_13268,N_13142);
nor U13630 (N_13630,N_13170,N_13335);
nor U13631 (N_13631,N_13134,N_13282);
nor U13632 (N_13632,N_13043,N_13349);
nand U13633 (N_13633,N_13128,N_13030);
nor U13634 (N_13634,N_13071,N_13172);
nand U13635 (N_13635,N_13009,N_13166);
or U13636 (N_13636,N_13192,N_13438);
nor U13637 (N_13637,N_13262,N_13058);
nand U13638 (N_13638,N_13345,N_13380);
nand U13639 (N_13639,N_13053,N_13263);
nand U13640 (N_13640,N_13425,N_13197);
nor U13641 (N_13641,N_13451,N_13003);
xor U13642 (N_13642,N_13203,N_13300);
nor U13643 (N_13643,N_13311,N_13103);
nor U13644 (N_13644,N_13434,N_13241);
nor U13645 (N_13645,N_13367,N_13499);
nor U13646 (N_13646,N_13297,N_13206);
or U13647 (N_13647,N_13414,N_13429);
or U13648 (N_13648,N_13121,N_13394);
nor U13649 (N_13649,N_13151,N_13060);
and U13650 (N_13650,N_13459,N_13339);
nor U13651 (N_13651,N_13374,N_13454);
or U13652 (N_13652,N_13117,N_13083);
or U13653 (N_13653,N_13301,N_13307);
and U13654 (N_13654,N_13471,N_13383);
or U13655 (N_13655,N_13122,N_13104);
or U13656 (N_13656,N_13290,N_13162);
nand U13657 (N_13657,N_13036,N_13105);
nand U13658 (N_13658,N_13037,N_13065);
nand U13659 (N_13659,N_13001,N_13150);
and U13660 (N_13660,N_13315,N_13098);
nor U13661 (N_13661,N_13403,N_13154);
or U13662 (N_13662,N_13057,N_13446);
and U13663 (N_13663,N_13251,N_13493);
nand U13664 (N_13664,N_13306,N_13314);
or U13665 (N_13665,N_13442,N_13195);
or U13666 (N_13666,N_13350,N_13189);
or U13667 (N_13667,N_13132,N_13012);
nand U13668 (N_13668,N_13025,N_13412);
nor U13669 (N_13669,N_13113,N_13129);
nand U13670 (N_13670,N_13179,N_13450);
nand U13671 (N_13671,N_13281,N_13099);
nand U13672 (N_13672,N_13059,N_13343);
or U13673 (N_13673,N_13386,N_13207);
nor U13674 (N_13674,N_13465,N_13112);
and U13675 (N_13675,N_13026,N_13213);
or U13676 (N_13676,N_13259,N_13149);
nand U13677 (N_13677,N_13333,N_13233);
nor U13678 (N_13678,N_13362,N_13231);
nor U13679 (N_13679,N_13075,N_13331);
nor U13680 (N_13680,N_13341,N_13384);
nand U13681 (N_13681,N_13250,N_13201);
and U13682 (N_13682,N_13205,N_13020);
nor U13683 (N_13683,N_13068,N_13396);
nor U13684 (N_13684,N_13273,N_13222);
and U13685 (N_13685,N_13361,N_13395);
or U13686 (N_13686,N_13239,N_13152);
or U13687 (N_13687,N_13453,N_13392);
nor U13688 (N_13688,N_13354,N_13073);
or U13689 (N_13689,N_13246,N_13299);
and U13690 (N_13690,N_13046,N_13336);
nor U13691 (N_13691,N_13054,N_13424);
nor U13692 (N_13692,N_13187,N_13191);
nand U13693 (N_13693,N_13467,N_13167);
nor U13694 (N_13694,N_13186,N_13159);
nand U13695 (N_13695,N_13479,N_13327);
nor U13696 (N_13696,N_13334,N_13108);
or U13697 (N_13697,N_13399,N_13022);
nand U13698 (N_13698,N_13092,N_13136);
nor U13699 (N_13699,N_13051,N_13265);
nand U13700 (N_13700,N_13196,N_13024);
or U13701 (N_13701,N_13127,N_13408);
nor U13702 (N_13702,N_13245,N_13184);
nand U13703 (N_13703,N_13076,N_13106);
nor U13704 (N_13704,N_13382,N_13360);
nor U13705 (N_13705,N_13305,N_13270);
nor U13706 (N_13706,N_13346,N_13163);
nand U13707 (N_13707,N_13356,N_13355);
xnor U13708 (N_13708,N_13283,N_13131);
and U13709 (N_13709,N_13294,N_13023);
and U13710 (N_13710,N_13407,N_13447);
nor U13711 (N_13711,N_13325,N_13038);
or U13712 (N_13712,N_13164,N_13107);
or U13713 (N_13713,N_13101,N_13317);
xor U13714 (N_13714,N_13484,N_13199);
nand U13715 (N_13715,N_13406,N_13316);
nand U13716 (N_13716,N_13094,N_13328);
nor U13717 (N_13717,N_13125,N_13352);
nand U13718 (N_13718,N_13337,N_13482);
xnor U13719 (N_13719,N_13253,N_13298);
or U13720 (N_13720,N_13376,N_13491);
nand U13721 (N_13721,N_13070,N_13085);
and U13722 (N_13722,N_13485,N_13431);
nor U13723 (N_13723,N_13074,N_13014);
nor U13724 (N_13724,N_13449,N_13138);
or U13725 (N_13725,N_13348,N_13257);
or U13726 (N_13726,N_13133,N_13220);
and U13727 (N_13727,N_13035,N_13078);
or U13728 (N_13728,N_13124,N_13126);
nand U13729 (N_13729,N_13007,N_13332);
nor U13730 (N_13730,N_13353,N_13358);
nand U13731 (N_13731,N_13005,N_13215);
xor U13732 (N_13732,N_13109,N_13496);
and U13733 (N_13733,N_13004,N_13420);
and U13734 (N_13734,N_13324,N_13302);
or U13735 (N_13735,N_13475,N_13013);
or U13736 (N_13736,N_13357,N_13033);
nor U13737 (N_13737,N_13464,N_13095);
and U13738 (N_13738,N_13460,N_13061);
nor U13739 (N_13739,N_13368,N_13006);
and U13740 (N_13740,N_13381,N_13237);
and U13741 (N_13741,N_13415,N_13090);
or U13742 (N_13742,N_13018,N_13385);
or U13743 (N_13743,N_13318,N_13312);
nand U13744 (N_13744,N_13329,N_13200);
and U13745 (N_13745,N_13495,N_13062);
xnor U13746 (N_13746,N_13185,N_13102);
xnor U13747 (N_13747,N_13146,N_13019);
nor U13748 (N_13748,N_13372,N_13444);
nor U13749 (N_13749,N_13322,N_13437);
nand U13750 (N_13750,N_13225,N_13093);
or U13751 (N_13751,N_13409,N_13405);
or U13752 (N_13752,N_13466,N_13204);
nand U13753 (N_13753,N_13250,N_13433);
or U13754 (N_13754,N_13295,N_13189);
or U13755 (N_13755,N_13075,N_13189);
nand U13756 (N_13756,N_13126,N_13142);
nor U13757 (N_13757,N_13416,N_13007);
or U13758 (N_13758,N_13310,N_13468);
or U13759 (N_13759,N_13419,N_13009);
nor U13760 (N_13760,N_13135,N_13384);
nor U13761 (N_13761,N_13190,N_13329);
nand U13762 (N_13762,N_13346,N_13360);
or U13763 (N_13763,N_13263,N_13018);
or U13764 (N_13764,N_13070,N_13020);
or U13765 (N_13765,N_13421,N_13252);
or U13766 (N_13766,N_13126,N_13132);
nor U13767 (N_13767,N_13453,N_13376);
or U13768 (N_13768,N_13302,N_13279);
nor U13769 (N_13769,N_13314,N_13464);
nor U13770 (N_13770,N_13495,N_13094);
nand U13771 (N_13771,N_13170,N_13478);
or U13772 (N_13772,N_13317,N_13319);
nand U13773 (N_13773,N_13448,N_13399);
nand U13774 (N_13774,N_13488,N_13037);
and U13775 (N_13775,N_13356,N_13440);
nand U13776 (N_13776,N_13087,N_13324);
and U13777 (N_13777,N_13275,N_13007);
or U13778 (N_13778,N_13492,N_13430);
or U13779 (N_13779,N_13230,N_13317);
or U13780 (N_13780,N_13294,N_13420);
nand U13781 (N_13781,N_13062,N_13233);
nand U13782 (N_13782,N_13428,N_13457);
nand U13783 (N_13783,N_13466,N_13407);
nor U13784 (N_13784,N_13406,N_13263);
and U13785 (N_13785,N_13042,N_13299);
nand U13786 (N_13786,N_13374,N_13183);
or U13787 (N_13787,N_13179,N_13181);
nand U13788 (N_13788,N_13112,N_13446);
nand U13789 (N_13789,N_13454,N_13266);
nor U13790 (N_13790,N_13070,N_13182);
or U13791 (N_13791,N_13210,N_13165);
and U13792 (N_13792,N_13380,N_13189);
or U13793 (N_13793,N_13147,N_13409);
nor U13794 (N_13794,N_13267,N_13037);
or U13795 (N_13795,N_13132,N_13266);
or U13796 (N_13796,N_13309,N_13446);
or U13797 (N_13797,N_13136,N_13239);
nor U13798 (N_13798,N_13318,N_13028);
nand U13799 (N_13799,N_13455,N_13008);
nand U13800 (N_13800,N_13032,N_13003);
and U13801 (N_13801,N_13142,N_13197);
nand U13802 (N_13802,N_13139,N_13317);
nand U13803 (N_13803,N_13017,N_13244);
nor U13804 (N_13804,N_13459,N_13069);
xor U13805 (N_13805,N_13287,N_13323);
or U13806 (N_13806,N_13448,N_13300);
nand U13807 (N_13807,N_13263,N_13181);
and U13808 (N_13808,N_13455,N_13106);
nor U13809 (N_13809,N_13319,N_13040);
nor U13810 (N_13810,N_13026,N_13467);
nor U13811 (N_13811,N_13034,N_13055);
nand U13812 (N_13812,N_13491,N_13240);
and U13813 (N_13813,N_13108,N_13093);
and U13814 (N_13814,N_13273,N_13029);
or U13815 (N_13815,N_13232,N_13399);
and U13816 (N_13816,N_13448,N_13262);
or U13817 (N_13817,N_13141,N_13137);
nand U13818 (N_13818,N_13318,N_13426);
and U13819 (N_13819,N_13355,N_13077);
or U13820 (N_13820,N_13319,N_13182);
nor U13821 (N_13821,N_13077,N_13460);
nor U13822 (N_13822,N_13064,N_13253);
nand U13823 (N_13823,N_13039,N_13028);
or U13824 (N_13824,N_13451,N_13149);
or U13825 (N_13825,N_13360,N_13259);
nor U13826 (N_13826,N_13323,N_13145);
or U13827 (N_13827,N_13251,N_13331);
nand U13828 (N_13828,N_13437,N_13321);
nand U13829 (N_13829,N_13195,N_13130);
xnor U13830 (N_13830,N_13138,N_13071);
or U13831 (N_13831,N_13313,N_13192);
nand U13832 (N_13832,N_13214,N_13225);
nor U13833 (N_13833,N_13161,N_13039);
xnor U13834 (N_13834,N_13351,N_13012);
and U13835 (N_13835,N_13064,N_13214);
nand U13836 (N_13836,N_13165,N_13243);
nand U13837 (N_13837,N_13465,N_13227);
nor U13838 (N_13838,N_13488,N_13198);
and U13839 (N_13839,N_13003,N_13184);
or U13840 (N_13840,N_13396,N_13370);
and U13841 (N_13841,N_13023,N_13354);
nor U13842 (N_13842,N_13362,N_13021);
nand U13843 (N_13843,N_13026,N_13121);
or U13844 (N_13844,N_13389,N_13181);
nand U13845 (N_13845,N_13168,N_13390);
or U13846 (N_13846,N_13197,N_13252);
or U13847 (N_13847,N_13463,N_13093);
and U13848 (N_13848,N_13192,N_13207);
nand U13849 (N_13849,N_13259,N_13222);
nor U13850 (N_13850,N_13287,N_13172);
or U13851 (N_13851,N_13002,N_13249);
or U13852 (N_13852,N_13088,N_13196);
nor U13853 (N_13853,N_13243,N_13306);
and U13854 (N_13854,N_13090,N_13014);
and U13855 (N_13855,N_13406,N_13285);
nor U13856 (N_13856,N_13225,N_13205);
nor U13857 (N_13857,N_13495,N_13306);
and U13858 (N_13858,N_13232,N_13390);
nor U13859 (N_13859,N_13470,N_13434);
or U13860 (N_13860,N_13170,N_13047);
nand U13861 (N_13861,N_13392,N_13248);
or U13862 (N_13862,N_13023,N_13429);
nand U13863 (N_13863,N_13323,N_13380);
nor U13864 (N_13864,N_13311,N_13160);
and U13865 (N_13865,N_13064,N_13195);
nand U13866 (N_13866,N_13477,N_13451);
xnor U13867 (N_13867,N_13143,N_13264);
or U13868 (N_13868,N_13328,N_13382);
nor U13869 (N_13869,N_13377,N_13236);
nand U13870 (N_13870,N_13457,N_13219);
nor U13871 (N_13871,N_13213,N_13051);
or U13872 (N_13872,N_13292,N_13250);
or U13873 (N_13873,N_13370,N_13312);
and U13874 (N_13874,N_13162,N_13248);
nor U13875 (N_13875,N_13123,N_13279);
or U13876 (N_13876,N_13095,N_13347);
and U13877 (N_13877,N_13193,N_13323);
or U13878 (N_13878,N_13225,N_13154);
and U13879 (N_13879,N_13095,N_13297);
nand U13880 (N_13880,N_13111,N_13362);
nand U13881 (N_13881,N_13241,N_13169);
nor U13882 (N_13882,N_13496,N_13363);
nor U13883 (N_13883,N_13377,N_13062);
and U13884 (N_13884,N_13381,N_13418);
or U13885 (N_13885,N_13198,N_13209);
xor U13886 (N_13886,N_13201,N_13424);
nor U13887 (N_13887,N_13341,N_13170);
nand U13888 (N_13888,N_13455,N_13213);
or U13889 (N_13889,N_13380,N_13235);
nor U13890 (N_13890,N_13027,N_13401);
nor U13891 (N_13891,N_13182,N_13461);
or U13892 (N_13892,N_13262,N_13426);
nor U13893 (N_13893,N_13249,N_13359);
nor U13894 (N_13894,N_13360,N_13121);
or U13895 (N_13895,N_13228,N_13141);
nor U13896 (N_13896,N_13299,N_13372);
nor U13897 (N_13897,N_13268,N_13308);
nor U13898 (N_13898,N_13470,N_13131);
nor U13899 (N_13899,N_13390,N_13304);
nand U13900 (N_13900,N_13289,N_13024);
or U13901 (N_13901,N_13093,N_13456);
and U13902 (N_13902,N_13466,N_13450);
or U13903 (N_13903,N_13151,N_13197);
nand U13904 (N_13904,N_13356,N_13371);
or U13905 (N_13905,N_13312,N_13199);
or U13906 (N_13906,N_13158,N_13027);
nor U13907 (N_13907,N_13436,N_13272);
nand U13908 (N_13908,N_13054,N_13210);
nand U13909 (N_13909,N_13322,N_13398);
nand U13910 (N_13910,N_13185,N_13444);
nor U13911 (N_13911,N_13447,N_13459);
nor U13912 (N_13912,N_13363,N_13119);
and U13913 (N_13913,N_13249,N_13340);
or U13914 (N_13914,N_13174,N_13244);
nor U13915 (N_13915,N_13362,N_13492);
nor U13916 (N_13916,N_13306,N_13198);
nand U13917 (N_13917,N_13403,N_13453);
nor U13918 (N_13918,N_13114,N_13448);
nor U13919 (N_13919,N_13380,N_13283);
or U13920 (N_13920,N_13284,N_13224);
and U13921 (N_13921,N_13465,N_13392);
nand U13922 (N_13922,N_13345,N_13174);
and U13923 (N_13923,N_13043,N_13325);
nand U13924 (N_13924,N_13166,N_13178);
nor U13925 (N_13925,N_13075,N_13027);
or U13926 (N_13926,N_13473,N_13002);
nand U13927 (N_13927,N_13436,N_13361);
or U13928 (N_13928,N_13467,N_13366);
and U13929 (N_13929,N_13317,N_13487);
nor U13930 (N_13930,N_13415,N_13186);
and U13931 (N_13931,N_13248,N_13146);
and U13932 (N_13932,N_13469,N_13435);
and U13933 (N_13933,N_13134,N_13104);
or U13934 (N_13934,N_13473,N_13008);
and U13935 (N_13935,N_13019,N_13172);
and U13936 (N_13936,N_13148,N_13190);
and U13937 (N_13937,N_13030,N_13127);
nor U13938 (N_13938,N_13431,N_13296);
or U13939 (N_13939,N_13298,N_13471);
and U13940 (N_13940,N_13127,N_13063);
and U13941 (N_13941,N_13217,N_13124);
and U13942 (N_13942,N_13059,N_13095);
and U13943 (N_13943,N_13206,N_13107);
nor U13944 (N_13944,N_13422,N_13024);
or U13945 (N_13945,N_13128,N_13056);
or U13946 (N_13946,N_13105,N_13426);
and U13947 (N_13947,N_13061,N_13040);
and U13948 (N_13948,N_13226,N_13244);
nor U13949 (N_13949,N_13129,N_13346);
and U13950 (N_13950,N_13128,N_13298);
and U13951 (N_13951,N_13311,N_13484);
or U13952 (N_13952,N_13243,N_13436);
and U13953 (N_13953,N_13294,N_13476);
or U13954 (N_13954,N_13289,N_13127);
xnor U13955 (N_13955,N_13021,N_13080);
nor U13956 (N_13956,N_13404,N_13474);
nand U13957 (N_13957,N_13398,N_13455);
or U13958 (N_13958,N_13473,N_13028);
and U13959 (N_13959,N_13144,N_13022);
nand U13960 (N_13960,N_13457,N_13243);
nor U13961 (N_13961,N_13429,N_13025);
nor U13962 (N_13962,N_13156,N_13147);
nor U13963 (N_13963,N_13155,N_13204);
and U13964 (N_13964,N_13141,N_13334);
or U13965 (N_13965,N_13189,N_13117);
or U13966 (N_13966,N_13172,N_13312);
nor U13967 (N_13967,N_13071,N_13233);
nand U13968 (N_13968,N_13121,N_13372);
or U13969 (N_13969,N_13081,N_13027);
xnor U13970 (N_13970,N_13049,N_13420);
or U13971 (N_13971,N_13279,N_13353);
and U13972 (N_13972,N_13366,N_13336);
nand U13973 (N_13973,N_13264,N_13262);
nand U13974 (N_13974,N_13212,N_13007);
nand U13975 (N_13975,N_13429,N_13440);
or U13976 (N_13976,N_13087,N_13420);
nor U13977 (N_13977,N_13054,N_13121);
nand U13978 (N_13978,N_13453,N_13274);
nand U13979 (N_13979,N_13151,N_13329);
nand U13980 (N_13980,N_13236,N_13114);
nand U13981 (N_13981,N_13217,N_13062);
xnor U13982 (N_13982,N_13375,N_13363);
and U13983 (N_13983,N_13133,N_13192);
nor U13984 (N_13984,N_13489,N_13465);
nor U13985 (N_13985,N_13043,N_13495);
nor U13986 (N_13986,N_13265,N_13498);
nor U13987 (N_13987,N_13473,N_13426);
nand U13988 (N_13988,N_13310,N_13222);
nand U13989 (N_13989,N_13291,N_13220);
nor U13990 (N_13990,N_13059,N_13215);
nand U13991 (N_13991,N_13383,N_13120);
nand U13992 (N_13992,N_13344,N_13425);
nor U13993 (N_13993,N_13023,N_13447);
nand U13994 (N_13994,N_13295,N_13047);
nor U13995 (N_13995,N_13421,N_13275);
and U13996 (N_13996,N_13109,N_13165);
or U13997 (N_13997,N_13190,N_13452);
and U13998 (N_13998,N_13419,N_13159);
or U13999 (N_13999,N_13361,N_13421);
and U14000 (N_14000,N_13877,N_13510);
nor U14001 (N_14001,N_13947,N_13934);
nand U14002 (N_14002,N_13693,N_13633);
nand U14003 (N_14003,N_13787,N_13678);
nor U14004 (N_14004,N_13970,N_13672);
nor U14005 (N_14005,N_13817,N_13533);
and U14006 (N_14006,N_13881,N_13614);
nand U14007 (N_14007,N_13968,N_13680);
or U14008 (N_14008,N_13631,N_13894);
and U14009 (N_14009,N_13760,N_13880);
nor U14010 (N_14010,N_13807,N_13886);
or U14011 (N_14011,N_13524,N_13851);
nor U14012 (N_14012,N_13517,N_13897);
nor U14013 (N_14013,N_13858,N_13771);
and U14014 (N_14014,N_13662,N_13889);
and U14015 (N_14015,N_13827,N_13818);
nand U14016 (N_14016,N_13679,N_13879);
or U14017 (N_14017,N_13557,N_13520);
and U14018 (N_14018,N_13608,N_13863);
and U14019 (N_14019,N_13625,N_13561);
and U14020 (N_14020,N_13584,N_13830);
nand U14021 (N_14021,N_13790,N_13500);
and U14022 (N_14022,N_13930,N_13700);
and U14023 (N_14023,N_13865,N_13891);
nand U14024 (N_14024,N_13786,N_13748);
or U14025 (N_14025,N_13546,N_13715);
and U14026 (N_14026,N_13536,N_13742);
nor U14027 (N_14027,N_13929,N_13802);
nor U14028 (N_14028,N_13980,N_13683);
nor U14029 (N_14029,N_13942,N_13728);
or U14030 (N_14030,N_13972,N_13888);
nor U14031 (N_14031,N_13567,N_13819);
or U14032 (N_14032,N_13768,N_13842);
nor U14033 (N_14033,N_13637,N_13754);
nor U14034 (N_14034,N_13724,N_13843);
nand U14035 (N_14035,N_13767,N_13931);
and U14036 (N_14036,N_13593,N_13822);
or U14037 (N_14037,N_13563,N_13624);
nand U14038 (N_14038,N_13738,N_13961);
nand U14039 (N_14039,N_13752,N_13749);
or U14040 (N_14040,N_13706,N_13909);
nand U14041 (N_14041,N_13795,N_13993);
or U14042 (N_14042,N_13745,N_13639);
nand U14043 (N_14043,N_13620,N_13750);
or U14044 (N_14044,N_13873,N_13659);
nor U14045 (N_14045,N_13606,N_13723);
or U14046 (N_14046,N_13591,N_13765);
nor U14047 (N_14047,N_13984,N_13804);
and U14048 (N_14048,N_13833,N_13844);
nor U14049 (N_14049,N_13840,N_13987);
xnor U14050 (N_14050,N_13784,N_13834);
nor U14051 (N_14051,N_13585,N_13655);
and U14052 (N_14052,N_13609,N_13741);
nor U14053 (N_14053,N_13660,N_13986);
nor U14054 (N_14054,N_13799,N_13674);
nor U14055 (N_14055,N_13564,N_13667);
nand U14056 (N_14056,N_13649,N_13726);
or U14057 (N_14057,N_13725,N_13869);
and U14058 (N_14058,N_13922,N_13789);
and U14059 (N_14059,N_13868,N_13645);
nand U14060 (N_14060,N_13872,N_13664);
or U14061 (N_14061,N_13601,N_13617);
nand U14062 (N_14062,N_13534,N_13730);
or U14063 (N_14063,N_13974,N_13707);
or U14064 (N_14064,N_13963,N_13918);
or U14065 (N_14065,N_13945,N_13692);
or U14066 (N_14066,N_13914,N_13526);
nand U14067 (N_14067,N_13924,N_13927);
nand U14068 (N_14068,N_13530,N_13831);
nand U14069 (N_14069,N_13857,N_13686);
or U14070 (N_14070,N_13782,N_13702);
nor U14071 (N_14071,N_13973,N_13568);
nand U14072 (N_14072,N_13991,N_13944);
nand U14073 (N_14073,N_13850,N_13965);
nand U14074 (N_14074,N_13501,N_13525);
nor U14075 (N_14075,N_13673,N_13710);
or U14076 (N_14076,N_13531,N_13855);
or U14077 (N_14077,N_13920,N_13569);
nor U14078 (N_14078,N_13856,N_13607);
nor U14079 (N_14079,N_13718,N_13956);
or U14080 (N_14080,N_13537,N_13647);
nor U14081 (N_14081,N_13504,N_13737);
nor U14082 (N_14082,N_13511,N_13936);
nand U14083 (N_14083,N_13657,N_13992);
nand U14084 (N_14084,N_13803,N_13717);
and U14085 (N_14085,N_13740,N_13713);
or U14086 (N_14086,N_13592,N_13556);
and U14087 (N_14087,N_13836,N_13732);
nand U14088 (N_14088,N_13554,N_13602);
and U14089 (N_14089,N_13763,N_13957);
nor U14090 (N_14090,N_13917,N_13506);
nor U14091 (N_14091,N_13755,N_13597);
and U14092 (N_14092,N_13849,N_13788);
nand U14093 (N_14093,N_13845,N_13578);
and U14094 (N_14094,N_13923,N_13698);
and U14095 (N_14095,N_13908,N_13959);
nand U14096 (N_14096,N_13995,N_13998);
and U14097 (N_14097,N_13539,N_13703);
and U14098 (N_14098,N_13780,N_13636);
or U14099 (N_14099,N_13684,N_13596);
nor U14100 (N_14100,N_13976,N_13581);
nor U14101 (N_14101,N_13800,N_13926);
and U14102 (N_14102,N_13635,N_13600);
or U14103 (N_14103,N_13604,N_13971);
nor U14104 (N_14104,N_13716,N_13935);
nor U14105 (N_14105,N_13816,N_13798);
or U14106 (N_14106,N_13874,N_13793);
or U14107 (N_14107,N_13846,N_13773);
and U14108 (N_14108,N_13670,N_13669);
xnor U14109 (N_14109,N_13646,N_13764);
and U14110 (N_14110,N_13985,N_13518);
and U14111 (N_14111,N_13582,N_13859);
nand U14112 (N_14112,N_13954,N_13919);
nand U14113 (N_14113,N_13792,N_13777);
nand U14114 (N_14114,N_13829,N_13630);
nand U14115 (N_14115,N_13576,N_13502);
nor U14116 (N_14116,N_13676,N_13528);
or U14117 (N_14117,N_13515,N_13523);
nand U14118 (N_14118,N_13785,N_13878);
nor U14119 (N_14119,N_13967,N_13911);
or U14120 (N_14120,N_13529,N_13562);
nand U14121 (N_14121,N_13677,N_13907);
nor U14122 (N_14122,N_13598,N_13571);
nand U14123 (N_14123,N_13644,N_13915);
nand U14124 (N_14124,N_13729,N_13847);
and U14125 (N_14125,N_13699,N_13514);
or U14126 (N_14126,N_13812,N_13590);
nor U14127 (N_14127,N_13952,N_13721);
nand U14128 (N_14128,N_13558,N_13746);
nand U14129 (N_14129,N_13550,N_13542);
or U14130 (N_14130,N_13675,N_13762);
or U14131 (N_14131,N_13666,N_13513);
nand U14132 (N_14132,N_13797,N_13938);
and U14133 (N_14133,N_13811,N_13714);
nand U14134 (N_14134,N_13808,N_13825);
and U14135 (N_14135,N_13731,N_13876);
nand U14136 (N_14136,N_13652,N_13977);
or U14137 (N_14137,N_13940,N_13629);
xor U14138 (N_14138,N_13982,N_13941);
and U14139 (N_14139,N_13555,N_13621);
nand U14140 (N_14140,N_13925,N_13663);
nand U14141 (N_14141,N_13573,N_13580);
or U14142 (N_14142,N_13769,N_13766);
or U14143 (N_14143,N_13705,N_13966);
and U14144 (N_14144,N_13905,N_13559);
and U14145 (N_14145,N_13835,N_13711);
xor U14146 (N_14146,N_13892,N_13516);
nand U14147 (N_14147,N_13508,N_13574);
nor U14148 (N_14148,N_13871,N_13906);
nand U14149 (N_14149,N_13653,N_13512);
and U14150 (N_14150,N_13722,N_13588);
or U14151 (N_14151,N_13988,N_13572);
and U14152 (N_14152,N_13913,N_13866);
or U14153 (N_14153,N_13996,N_13902);
or U14154 (N_14154,N_13575,N_13778);
nor U14155 (N_14155,N_13734,N_13813);
nand U14156 (N_14156,N_13781,N_13656);
and U14157 (N_14157,N_13688,N_13904);
and U14158 (N_14158,N_13743,N_13538);
nand U14159 (N_14159,N_13616,N_13640);
and U14160 (N_14160,N_13566,N_13634);
or U14161 (N_14161,N_13951,N_13937);
or U14162 (N_14162,N_13695,N_13544);
or U14163 (N_14163,N_13898,N_13691);
nand U14164 (N_14164,N_13791,N_13503);
or U14165 (N_14165,N_13747,N_13687);
nor U14166 (N_14166,N_13757,N_13739);
or U14167 (N_14167,N_13964,N_13583);
or U14168 (N_14168,N_13779,N_13933);
nor U14169 (N_14169,N_13658,N_13643);
nor U14170 (N_14170,N_13541,N_13838);
nor U14171 (N_14171,N_13610,N_13650);
nor U14172 (N_14172,N_13823,N_13595);
and U14173 (N_14173,N_13638,N_13751);
and U14174 (N_14174,N_13783,N_13577);
or U14175 (N_14175,N_13837,N_13668);
nand U14176 (N_14176,N_13651,N_13547);
nor U14177 (N_14177,N_13758,N_13854);
and U14178 (N_14178,N_13615,N_13841);
nor U14179 (N_14179,N_13611,N_13776);
nand U14180 (N_14180,N_13978,N_13552);
nand U14181 (N_14181,N_13532,N_13627);
nor U14182 (N_14182,N_13989,N_13540);
nand U14183 (N_14183,N_13895,N_13862);
or U14184 (N_14184,N_13543,N_13619);
and U14185 (N_14185,N_13912,N_13623);
nand U14186 (N_14186,N_13682,N_13551);
or U14187 (N_14187,N_13744,N_13613);
nor U14188 (N_14188,N_13587,N_13654);
nor U14189 (N_14189,N_13548,N_13860);
nor U14190 (N_14190,N_13887,N_13948);
and U14191 (N_14191,N_13916,N_13527);
or U14192 (N_14192,N_13522,N_13709);
nand U14193 (N_14193,N_13960,N_13852);
or U14194 (N_14194,N_13910,N_13735);
nor U14195 (N_14195,N_13832,N_13736);
and U14196 (N_14196,N_13507,N_13999);
nor U14197 (N_14197,N_13618,N_13893);
nand U14198 (N_14198,N_13505,N_13853);
nor U14199 (N_14199,N_13928,N_13545);
xor U14200 (N_14200,N_13824,N_13809);
or U14201 (N_14201,N_13519,N_13805);
nand U14202 (N_14202,N_13774,N_13896);
and U14203 (N_14203,N_13796,N_13826);
nand U14204 (N_14204,N_13884,N_13815);
and U14205 (N_14205,N_13570,N_13761);
nor U14206 (N_14206,N_13794,N_13969);
or U14207 (N_14207,N_13821,N_13612);
nor U14208 (N_14208,N_13870,N_13733);
nor U14209 (N_14209,N_13939,N_13641);
or U14210 (N_14210,N_13983,N_13839);
nand U14211 (N_14211,N_13950,N_13990);
nor U14212 (N_14212,N_13861,N_13708);
and U14213 (N_14213,N_13599,N_13770);
nand U14214 (N_14214,N_13586,N_13622);
or U14215 (N_14215,N_13594,N_13632);
nand U14216 (N_14216,N_13720,N_13560);
and U14217 (N_14217,N_13697,N_13810);
or U14218 (N_14218,N_13828,N_13981);
and U14219 (N_14219,N_13565,N_13704);
and U14220 (N_14220,N_13900,N_13867);
or U14221 (N_14221,N_13901,N_13759);
and U14222 (N_14222,N_13642,N_13753);
nand U14223 (N_14223,N_13975,N_13890);
nand U14224 (N_14224,N_13775,N_13535);
or U14225 (N_14225,N_13921,N_13814);
nand U14226 (N_14226,N_13932,N_13997);
or U14227 (N_14227,N_13943,N_13756);
or U14228 (N_14228,N_13953,N_13605);
or U14229 (N_14229,N_13628,N_13521);
or U14230 (N_14230,N_13661,N_13696);
or U14231 (N_14231,N_13962,N_13712);
or U14232 (N_14232,N_13579,N_13694);
or U14233 (N_14233,N_13958,N_13820);
or U14234 (N_14234,N_13883,N_13885);
or U14235 (N_14235,N_13685,N_13681);
and U14236 (N_14236,N_13553,N_13648);
nor U14237 (N_14237,N_13701,N_13549);
nand U14238 (N_14238,N_13903,N_13875);
or U14239 (N_14239,N_13882,N_13949);
nor U14240 (N_14240,N_13626,N_13946);
xor U14241 (N_14241,N_13689,N_13665);
and U14242 (N_14242,N_13690,N_13772);
nand U14243 (N_14243,N_13603,N_13589);
nor U14244 (N_14244,N_13994,N_13979);
nand U14245 (N_14245,N_13509,N_13727);
nor U14246 (N_14246,N_13671,N_13719);
nor U14247 (N_14247,N_13801,N_13955);
or U14248 (N_14248,N_13806,N_13899);
or U14249 (N_14249,N_13864,N_13848);
nor U14250 (N_14250,N_13829,N_13736);
nand U14251 (N_14251,N_13669,N_13924);
or U14252 (N_14252,N_13518,N_13897);
nor U14253 (N_14253,N_13796,N_13932);
or U14254 (N_14254,N_13847,N_13782);
nor U14255 (N_14255,N_13853,N_13681);
nand U14256 (N_14256,N_13956,N_13996);
or U14257 (N_14257,N_13643,N_13672);
and U14258 (N_14258,N_13985,N_13622);
and U14259 (N_14259,N_13828,N_13705);
and U14260 (N_14260,N_13563,N_13663);
or U14261 (N_14261,N_13944,N_13705);
nand U14262 (N_14262,N_13862,N_13651);
and U14263 (N_14263,N_13800,N_13706);
and U14264 (N_14264,N_13545,N_13874);
and U14265 (N_14265,N_13565,N_13652);
nor U14266 (N_14266,N_13596,N_13638);
or U14267 (N_14267,N_13689,N_13787);
and U14268 (N_14268,N_13658,N_13551);
nand U14269 (N_14269,N_13777,N_13737);
and U14270 (N_14270,N_13992,N_13619);
nor U14271 (N_14271,N_13813,N_13552);
nor U14272 (N_14272,N_13967,N_13955);
and U14273 (N_14273,N_13672,N_13772);
or U14274 (N_14274,N_13825,N_13740);
or U14275 (N_14275,N_13704,N_13860);
nand U14276 (N_14276,N_13623,N_13748);
nor U14277 (N_14277,N_13779,N_13761);
and U14278 (N_14278,N_13888,N_13590);
nand U14279 (N_14279,N_13651,N_13921);
nor U14280 (N_14280,N_13678,N_13709);
nor U14281 (N_14281,N_13852,N_13706);
or U14282 (N_14282,N_13893,N_13816);
or U14283 (N_14283,N_13822,N_13746);
and U14284 (N_14284,N_13857,N_13773);
and U14285 (N_14285,N_13949,N_13507);
nand U14286 (N_14286,N_13737,N_13810);
or U14287 (N_14287,N_13907,N_13604);
nand U14288 (N_14288,N_13838,N_13564);
nand U14289 (N_14289,N_13801,N_13796);
nor U14290 (N_14290,N_13593,N_13576);
nand U14291 (N_14291,N_13914,N_13767);
nor U14292 (N_14292,N_13813,N_13692);
nor U14293 (N_14293,N_13763,N_13587);
or U14294 (N_14294,N_13829,N_13957);
and U14295 (N_14295,N_13927,N_13562);
nand U14296 (N_14296,N_13990,N_13789);
or U14297 (N_14297,N_13982,N_13551);
or U14298 (N_14298,N_13942,N_13794);
nand U14299 (N_14299,N_13684,N_13725);
nand U14300 (N_14300,N_13807,N_13908);
and U14301 (N_14301,N_13934,N_13952);
nand U14302 (N_14302,N_13911,N_13585);
nand U14303 (N_14303,N_13684,N_13911);
and U14304 (N_14304,N_13739,N_13509);
or U14305 (N_14305,N_13571,N_13781);
and U14306 (N_14306,N_13751,N_13857);
nand U14307 (N_14307,N_13952,N_13760);
xnor U14308 (N_14308,N_13746,N_13565);
or U14309 (N_14309,N_13549,N_13903);
nor U14310 (N_14310,N_13666,N_13627);
or U14311 (N_14311,N_13623,N_13509);
nand U14312 (N_14312,N_13826,N_13617);
nor U14313 (N_14313,N_13783,N_13687);
or U14314 (N_14314,N_13548,N_13951);
nor U14315 (N_14315,N_13939,N_13871);
or U14316 (N_14316,N_13686,N_13783);
and U14317 (N_14317,N_13936,N_13920);
nand U14318 (N_14318,N_13855,N_13791);
and U14319 (N_14319,N_13585,N_13692);
and U14320 (N_14320,N_13741,N_13729);
nor U14321 (N_14321,N_13592,N_13924);
nand U14322 (N_14322,N_13838,N_13917);
and U14323 (N_14323,N_13852,N_13771);
or U14324 (N_14324,N_13887,N_13627);
and U14325 (N_14325,N_13836,N_13821);
or U14326 (N_14326,N_13588,N_13814);
nor U14327 (N_14327,N_13544,N_13982);
nor U14328 (N_14328,N_13693,N_13615);
xor U14329 (N_14329,N_13737,N_13664);
and U14330 (N_14330,N_13987,N_13744);
or U14331 (N_14331,N_13542,N_13961);
nand U14332 (N_14332,N_13692,N_13631);
nor U14333 (N_14333,N_13803,N_13727);
nor U14334 (N_14334,N_13745,N_13584);
and U14335 (N_14335,N_13535,N_13640);
or U14336 (N_14336,N_13644,N_13547);
and U14337 (N_14337,N_13992,N_13788);
nor U14338 (N_14338,N_13816,N_13900);
and U14339 (N_14339,N_13779,N_13643);
nand U14340 (N_14340,N_13716,N_13799);
xor U14341 (N_14341,N_13537,N_13791);
or U14342 (N_14342,N_13534,N_13672);
or U14343 (N_14343,N_13606,N_13578);
nor U14344 (N_14344,N_13504,N_13884);
nand U14345 (N_14345,N_13775,N_13826);
nand U14346 (N_14346,N_13977,N_13547);
and U14347 (N_14347,N_13512,N_13978);
nand U14348 (N_14348,N_13700,N_13969);
and U14349 (N_14349,N_13697,N_13552);
or U14350 (N_14350,N_13589,N_13733);
and U14351 (N_14351,N_13568,N_13986);
and U14352 (N_14352,N_13580,N_13752);
nand U14353 (N_14353,N_13949,N_13965);
and U14354 (N_14354,N_13526,N_13880);
or U14355 (N_14355,N_13717,N_13828);
and U14356 (N_14356,N_13714,N_13843);
nor U14357 (N_14357,N_13708,N_13777);
nand U14358 (N_14358,N_13714,N_13886);
nor U14359 (N_14359,N_13830,N_13711);
nand U14360 (N_14360,N_13624,N_13534);
or U14361 (N_14361,N_13674,N_13723);
and U14362 (N_14362,N_13750,N_13635);
nand U14363 (N_14363,N_13752,N_13744);
or U14364 (N_14364,N_13559,N_13976);
nor U14365 (N_14365,N_13682,N_13712);
nor U14366 (N_14366,N_13958,N_13892);
nand U14367 (N_14367,N_13572,N_13925);
nand U14368 (N_14368,N_13577,N_13653);
nor U14369 (N_14369,N_13612,N_13615);
and U14370 (N_14370,N_13759,N_13953);
nor U14371 (N_14371,N_13753,N_13736);
and U14372 (N_14372,N_13647,N_13633);
xnor U14373 (N_14373,N_13549,N_13745);
and U14374 (N_14374,N_13632,N_13976);
xnor U14375 (N_14375,N_13920,N_13956);
and U14376 (N_14376,N_13735,N_13540);
nor U14377 (N_14377,N_13961,N_13577);
or U14378 (N_14378,N_13710,N_13814);
nor U14379 (N_14379,N_13970,N_13977);
nand U14380 (N_14380,N_13559,N_13653);
nor U14381 (N_14381,N_13961,N_13971);
and U14382 (N_14382,N_13844,N_13984);
nor U14383 (N_14383,N_13813,N_13926);
or U14384 (N_14384,N_13642,N_13617);
xor U14385 (N_14385,N_13570,N_13532);
and U14386 (N_14386,N_13638,N_13637);
nor U14387 (N_14387,N_13551,N_13790);
nor U14388 (N_14388,N_13562,N_13864);
or U14389 (N_14389,N_13786,N_13507);
nor U14390 (N_14390,N_13950,N_13628);
nand U14391 (N_14391,N_13703,N_13994);
nand U14392 (N_14392,N_13762,N_13971);
or U14393 (N_14393,N_13522,N_13668);
nand U14394 (N_14394,N_13861,N_13828);
nand U14395 (N_14395,N_13559,N_13931);
nor U14396 (N_14396,N_13759,N_13853);
and U14397 (N_14397,N_13890,N_13779);
nor U14398 (N_14398,N_13894,N_13735);
and U14399 (N_14399,N_13671,N_13539);
or U14400 (N_14400,N_13519,N_13602);
or U14401 (N_14401,N_13874,N_13843);
nor U14402 (N_14402,N_13743,N_13824);
nand U14403 (N_14403,N_13544,N_13592);
nand U14404 (N_14404,N_13877,N_13502);
or U14405 (N_14405,N_13699,N_13678);
nor U14406 (N_14406,N_13868,N_13574);
nor U14407 (N_14407,N_13739,N_13791);
and U14408 (N_14408,N_13895,N_13758);
and U14409 (N_14409,N_13532,N_13752);
nand U14410 (N_14410,N_13525,N_13915);
nor U14411 (N_14411,N_13691,N_13611);
nand U14412 (N_14412,N_13908,N_13697);
nand U14413 (N_14413,N_13574,N_13840);
nand U14414 (N_14414,N_13833,N_13859);
and U14415 (N_14415,N_13792,N_13534);
and U14416 (N_14416,N_13874,N_13753);
nor U14417 (N_14417,N_13772,N_13968);
and U14418 (N_14418,N_13895,N_13680);
nor U14419 (N_14419,N_13923,N_13936);
nand U14420 (N_14420,N_13584,N_13848);
and U14421 (N_14421,N_13648,N_13804);
or U14422 (N_14422,N_13776,N_13507);
nand U14423 (N_14423,N_13732,N_13709);
or U14424 (N_14424,N_13511,N_13748);
nand U14425 (N_14425,N_13510,N_13544);
and U14426 (N_14426,N_13961,N_13635);
nor U14427 (N_14427,N_13832,N_13667);
or U14428 (N_14428,N_13718,N_13886);
or U14429 (N_14429,N_13501,N_13565);
or U14430 (N_14430,N_13557,N_13769);
and U14431 (N_14431,N_13928,N_13883);
or U14432 (N_14432,N_13626,N_13771);
nor U14433 (N_14433,N_13581,N_13944);
and U14434 (N_14434,N_13612,N_13730);
nand U14435 (N_14435,N_13898,N_13501);
nor U14436 (N_14436,N_13905,N_13539);
nand U14437 (N_14437,N_13770,N_13805);
and U14438 (N_14438,N_13658,N_13566);
nand U14439 (N_14439,N_13708,N_13732);
or U14440 (N_14440,N_13916,N_13728);
or U14441 (N_14441,N_13923,N_13696);
nand U14442 (N_14442,N_13530,N_13644);
nor U14443 (N_14443,N_13692,N_13954);
nor U14444 (N_14444,N_13746,N_13982);
xnor U14445 (N_14445,N_13867,N_13538);
nor U14446 (N_14446,N_13975,N_13502);
nor U14447 (N_14447,N_13666,N_13977);
or U14448 (N_14448,N_13677,N_13933);
and U14449 (N_14449,N_13842,N_13559);
and U14450 (N_14450,N_13908,N_13979);
nand U14451 (N_14451,N_13808,N_13736);
or U14452 (N_14452,N_13959,N_13890);
and U14453 (N_14453,N_13979,N_13530);
and U14454 (N_14454,N_13601,N_13828);
nor U14455 (N_14455,N_13709,N_13578);
nor U14456 (N_14456,N_13888,N_13547);
nor U14457 (N_14457,N_13914,N_13850);
nand U14458 (N_14458,N_13655,N_13590);
nand U14459 (N_14459,N_13771,N_13836);
or U14460 (N_14460,N_13535,N_13835);
nand U14461 (N_14461,N_13543,N_13871);
nor U14462 (N_14462,N_13930,N_13829);
or U14463 (N_14463,N_13730,N_13874);
or U14464 (N_14464,N_13874,N_13933);
nor U14465 (N_14465,N_13782,N_13765);
nand U14466 (N_14466,N_13920,N_13768);
and U14467 (N_14467,N_13544,N_13772);
nand U14468 (N_14468,N_13750,N_13621);
nor U14469 (N_14469,N_13747,N_13753);
or U14470 (N_14470,N_13871,N_13789);
nor U14471 (N_14471,N_13524,N_13518);
nor U14472 (N_14472,N_13587,N_13724);
or U14473 (N_14473,N_13833,N_13847);
or U14474 (N_14474,N_13833,N_13650);
or U14475 (N_14475,N_13912,N_13542);
nor U14476 (N_14476,N_13752,N_13993);
and U14477 (N_14477,N_13974,N_13701);
nand U14478 (N_14478,N_13761,N_13641);
nor U14479 (N_14479,N_13648,N_13667);
nor U14480 (N_14480,N_13550,N_13507);
and U14481 (N_14481,N_13547,N_13735);
nor U14482 (N_14482,N_13572,N_13866);
and U14483 (N_14483,N_13674,N_13973);
and U14484 (N_14484,N_13625,N_13976);
or U14485 (N_14485,N_13771,N_13955);
nand U14486 (N_14486,N_13916,N_13560);
and U14487 (N_14487,N_13928,N_13777);
and U14488 (N_14488,N_13712,N_13831);
nor U14489 (N_14489,N_13675,N_13535);
and U14490 (N_14490,N_13852,N_13988);
nor U14491 (N_14491,N_13862,N_13943);
and U14492 (N_14492,N_13655,N_13739);
nor U14493 (N_14493,N_13646,N_13750);
nand U14494 (N_14494,N_13828,N_13984);
nor U14495 (N_14495,N_13773,N_13651);
or U14496 (N_14496,N_13712,N_13716);
nand U14497 (N_14497,N_13986,N_13844);
nor U14498 (N_14498,N_13639,N_13550);
nand U14499 (N_14499,N_13887,N_13579);
and U14500 (N_14500,N_14069,N_14473);
nor U14501 (N_14501,N_14470,N_14268);
or U14502 (N_14502,N_14189,N_14456);
or U14503 (N_14503,N_14402,N_14392);
nor U14504 (N_14504,N_14321,N_14007);
nand U14505 (N_14505,N_14166,N_14480);
nor U14506 (N_14506,N_14050,N_14218);
and U14507 (N_14507,N_14284,N_14110);
nand U14508 (N_14508,N_14361,N_14495);
nand U14509 (N_14509,N_14187,N_14451);
and U14510 (N_14510,N_14333,N_14012);
nand U14511 (N_14511,N_14244,N_14198);
or U14512 (N_14512,N_14000,N_14222);
nor U14513 (N_14513,N_14227,N_14107);
and U14514 (N_14514,N_14475,N_14086);
and U14515 (N_14515,N_14250,N_14108);
nand U14516 (N_14516,N_14140,N_14448);
nand U14517 (N_14517,N_14347,N_14421);
xnor U14518 (N_14518,N_14300,N_14292);
nor U14519 (N_14519,N_14038,N_14494);
and U14520 (N_14520,N_14242,N_14306);
or U14521 (N_14521,N_14183,N_14433);
nor U14522 (N_14522,N_14450,N_14149);
nand U14523 (N_14523,N_14194,N_14207);
or U14524 (N_14524,N_14482,N_14235);
nor U14525 (N_14525,N_14053,N_14279);
and U14526 (N_14526,N_14133,N_14178);
nor U14527 (N_14527,N_14098,N_14365);
and U14528 (N_14528,N_14464,N_14371);
xnor U14529 (N_14529,N_14021,N_14415);
and U14530 (N_14530,N_14144,N_14177);
or U14531 (N_14531,N_14376,N_14136);
nand U14532 (N_14532,N_14124,N_14233);
or U14533 (N_14533,N_14134,N_14182);
nor U14534 (N_14534,N_14083,N_14370);
or U14535 (N_14535,N_14161,N_14383);
or U14536 (N_14536,N_14385,N_14212);
nand U14537 (N_14537,N_14153,N_14315);
and U14538 (N_14538,N_14018,N_14199);
and U14539 (N_14539,N_14301,N_14229);
nor U14540 (N_14540,N_14224,N_14163);
nand U14541 (N_14541,N_14232,N_14428);
or U14542 (N_14542,N_14310,N_14299);
or U14543 (N_14543,N_14334,N_14303);
and U14544 (N_14544,N_14266,N_14155);
nand U14545 (N_14545,N_14010,N_14308);
nand U14546 (N_14546,N_14080,N_14011);
or U14547 (N_14547,N_14491,N_14109);
or U14548 (N_14548,N_14208,N_14346);
or U14549 (N_14549,N_14390,N_14372);
or U14550 (N_14550,N_14019,N_14492);
nand U14551 (N_14551,N_14202,N_14430);
nand U14552 (N_14552,N_14079,N_14230);
nor U14553 (N_14553,N_14049,N_14287);
nand U14554 (N_14554,N_14269,N_14078);
and U14555 (N_14555,N_14017,N_14096);
xnor U14556 (N_14556,N_14200,N_14245);
nand U14557 (N_14557,N_14400,N_14264);
nor U14558 (N_14558,N_14132,N_14258);
and U14559 (N_14559,N_14173,N_14403);
or U14560 (N_14560,N_14138,N_14351);
or U14561 (N_14561,N_14337,N_14023);
nor U14562 (N_14562,N_14131,N_14204);
or U14563 (N_14563,N_14190,N_14197);
nor U14564 (N_14564,N_14239,N_14338);
or U14565 (N_14565,N_14317,N_14395);
nor U14566 (N_14566,N_14236,N_14089);
nor U14567 (N_14567,N_14348,N_14209);
and U14568 (N_14568,N_14324,N_14476);
and U14569 (N_14569,N_14001,N_14498);
and U14570 (N_14570,N_14458,N_14090);
nand U14571 (N_14571,N_14062,N_14459);
and U14572 (N_14572,N_14063,N_14359);
and U14573 (N_14573,N_14322,N_14085);
nand U14574 (N_14574,N_14093,N_14024);
nand U14575 (N_14575,N_14467,N_14151);
nand U14576 (N_14576,N_14247,N_14101);
xnor U14577 (N_14577,N_14339,N_14353);
and U14578 (N_14578,N_14367,N_14422);
or U14579 (N_14579,N_14123,N_14099);
and U14580 (N_14580,N_14489,N_14465);
nand U14581 (N_14581,N_14249,N_14168);
and U14582 (N_14582,N_14267,N_14397);
and U14583 (N_14583,N_14041,N_14461);
nor U14584 (N_14584,N_14102,N_14288);
or U14585 (N_14585,N_14468,N_14210);
or U14586 (N_14586,N_14398,N_14343);
nor U14587 (N_14587,N_14323,N_14426);
nand U14588 (N_14588,N_14309,N_14354);
nand U14589 (N_14589,N_14329,N_14429);
and U14590 (N_14590,N_14399,N_14028);
nand U14591 (N_14591,N_14439,N_14216);
nand U14592 (N_14592,N_14130,N_14052);
or U14593 (N_14593,N_14157,N_14274);
or U14594 (N_14594,N_14142,N_14170);
and U14595 (N_14595,N_14100,N_14191);
nor U14596 (N_14596,N_14418,N_14466);
nand U14597 (N_14597,N_14427,N_14095);
nand U14598 (N_14598,N_14034,N_14016);
and U14599 (N_14599,N_14253,N_14304);
or U14600 (N_14600,N_14278,N_14262);
and U14601 (N_14601,N_14005,N_14006);
or U14602 (N_14602,N_14043,N_14077);
nand U14603 (N_14603,N_14330,N_14174);
and U14604 (N_14604,N_14217,N_14206);
nand U14605 (N_14605,N_14445,N_14496);
or U14606 (N_14606,N_14412,N_14203);
nor U14607 (N_14607,N_14328,N_14270);
or U14608 (N_14608,N_14298,N_14103);
nor U14609 (N_14609,N_14160,N_14004);
and U14610 (N_14610,N_14296,N_14366);
nor U14611 (N_14611,N_14081,N_14350);
nand U14612 (N_14612,N_14039,N_14345);
nand U14613 (N_14613,N_14251,N_14405);
nand U14614 (N_14614,N_14460,N_14030);
and U14615 (N_14615,N_14380,N_14457);
or U14616 (N_14616,N_14419,N_14072);
and U14617 (N_14617,N_14478,N_14033);
nor U14618 (N_14618,N_14368,N_14228);
and U14619 (N_14619,N_14434,N_14356);
nor U14620 (N_14620,N_14145,N_14424);
or U14621 (N_14621,N_14313,N_14293);
nand U14622 (N_14622,N_14221,N_14488);
and U14623 (N_14623,N_14186,N_14487);
and U14624 (N_14624,N_14407,N_14349);
or U14625 (N_14625,N_14425,N_14499);
nor U14626 (N_14626,N_14435,N_14291);
nor U14627 (N_14627,N_14286,N_14116);
and U14628 (N_14628,N_14256,N_14382);
nand U14629 (N_14629,N_14087,N_14469);
nand U14630 (N_14630,N_14243,N_14146);
nor U14631 (N_14631,N_14234,N_14048);
or U14632 (N_14632,N_14335,N_14357);
and U14633 (N_14633,N_14074,N_14226);
xnor U14634 (N_14634,N_14181,N_14088);
nor U14635 (N_14635,N_14137,N_14396);
nand U14636 (N_14636,N_14193,N_14128);
or U14637 (N_14637,N_14027,N_14238);
and U14638 (N_14638,N_14112,N_14290);
nor U14639 (N_14639,N_14248,N_14097);
and U14640 (N_14640,N_14342,N_14332);
and U14641 (N_14641,N_14477,N_14119);
xor U14642 (N_14642,N_14073,N_14076);
or U14643 (N_14643,N_14273,N_14046);
and U14644 (N_14644,N_14281,N_14386);
nand U14645 (N_14645,N_14423,N_14289);
nand U14646 (N_14646,N_14294,N_14272);
or U14647 (N_14647,N_14118,N_14020);
nor U14648 (N_14648,N_14352,N_14295);
and U14649 (N_14649,N_14064,N_14070);
xnor U14650 (N_14650,N_14241,N_14486);
or U14651 (N_14651,N_14051,N_14462);
nor U14652 (N_14652,N_14285,N_14413);
or U14653 (N_14653,N_14472,N_14331);
nand U14654 (N_14654,N_14388,N_14220);
or U14655 (N_14655,N_14065,N_14214);
or U14656 (N_14656,N_14355,N_14364);
nand U14657 (N_14657,N_14044,N_14246);
nor U14658 (N_14658,N_14122,N_14393);
and U14659 (N_14659,N_14493,N_14008);
nor U14660 (N_14660,N_14114,N_14252);
nand U14661 (N_14661,N_14179,N_14431);
xor U14662 (N_14662,N_14381,N_14307);
nor U14663 (N_14663,N_14254,N_14165);
and U14664 (N_14664,N_14143,N_14061);
or U14665 (N_14665,N_14404,N_14029);
nor U14666 (N_14666,N_14319,N_14013);
or U14667 (N_14667,N_14259,N_14416);
xor U14668 (N_14668,N_14326,N_14261);
or U14669 (N_14669,N_14032,N_14058);
nand U14670 (N_14670,N_14444,N_14271);
nand U14671 (N_14671,N_14180,N_14205);
or U14672 (N_14672,N_14164,N_14237);
nand U14673 (N_14673,N_14188,N_14113);
nor U14674 (N_14674,N_14022,N_14373);
nor U14675 (N_14675,N_14378,N_14040);
nand U14676 (N_14676,N_14185,N_14409);
or U14677 (N_14677,N_14071,N_14255);
or U14678 (N_14678,N_14379,N_14126);
nand U14679 (N_14679,N_14172,N_14117);
nand U14680 (N_14680,N_14213,N_14129);
nand U14681 (N_14681,N_14169,N_14369);
nor U14682 (N_14682,N_14340,N_14260);
or U14683 (N_14683,N_14374,N_14384);
nor U14684 (N_14684,N_14389,N_14201);
nor U14685 (N_14685,N_14042,N_14497);
xor U14686 (N_14686,N_14105,N_14455);
and U14687 (N_14687,N_14036,N_14184);
or U14688 (N_14688,N_14115,N_14167);
and U14689 (N_14689,N_14490,N_14148);
nand U14690 (N_14690,N_14219,N_14015);
nor U14691 (N_14691,N_14263,N_14192);
nor U14692 (N_14692,N_14320,N_14441);
xor U14693 (N_14693,N_14363,N_14452);
nand U14694 (N_14694,N_14014,N_14362);
or U14695 (N_14695,N_14454,N_14276);
and U14696 (N_14696,N_14327,N_14120);
and U14697 (N_14697,N_14394,N_14067);
or U14698 (N_14698,N_14196,N_14104);
and U14699 (N_14699,N_14387,N_14377);
nor U14700 (N_14700,N_14302,N_14344);
or U14701 (N_14701,N_14055,N_14410);
or U14702 (N_14702,N_14047,N_14231);
nand U14703 (N_14703,N_14297,N_14432);
and U14704 (N_14704,N_14280,N_14316);
nor U14705 (N_14705,N_14336,N_14474);
nand U14706 (N_14706,N_14318,N_14401);
nor U14707 (N_14707,N_14141,N_14275);
and U14708 (N_14708,N_14438,N_14240);
or U14709 (N_14709,N_14125,N_14442);
and U14710 (N_14710,N_14437,N_14066);
or U14711 (N_14711,N_14084,N_14175);
xor U14712 (N_14712,N_14481,N_14360);
and U14713 (N_14713,N_14025,N_14283);
or U14714 (N_14714,N_14154,N_14106);
nand U14715 (N_14715,N_14002,N_14037);
nor U14716 (N_14716,N_14406,N_14056);
or U14717 (N_14717,N_14211,N_14453);
and U14718 (N_14718,N_14225,N_14341);
nand U14719 (N_14719,N_14265,N_14162);
or U14720 (N_14720,N_14003,N_14026);
nand U14721 (N_14721,N_14358,N_14150);
xor U14722 (N_14722,N_14156,N_14436);
nand U14723 (N_14723,N_14139,N_14127);
and U14724 (N_14724,N_14059,N_14111);
xor U14725 (N_14725,N_14159,N_14479);
and U14726 (N_14726,N_14215,N_14282);
nor U14727 (N_14727,N_14060,N_14440);
and U14728 (N_14728,N_14054,N_14057);
nor U14729 (N_14729,N_14305,N_14075);
or U14730 (N_14730,N_14420,N_14414);
nor U14731 (N_14731,N_14408,N_14082);
nor U14732 (N_14732,N_14158,N_14068);
nor U14733 (N_14733,N_14031,N_14091);
or U14734 (N_14734,N_14171,N_14484);
or U14735 (N_14735,N_14312,N_14121);
nand U14736 (N_14736,N_14411,N_14443);
or U14737 (N_14737,N_14257,N_14009);
or U14738 (N_14738,N_14176,N_14277);
or U14739 (N_14739,N_14483,N_14314);
and U14740 (N_14740,N_14147,N_14447);
or U14741 (N_14741,N_14375,N_14195);
and U14742 (N_14742,N_14045,N_14446);
or U14743 (N_14743,N_14092,N_14311);
or U14744 (N_14744,N_14223,N_14391);
nor U14745 (N_14745,N_14485,N_14417);
nand U14746 (N_14746,N_14449,N_14325);
nand U14747 (N_14747,N_14471,N_14094);
nand U14748 (N_14748,N_14463,N_14135);
nor U14749 (N_14749,N_14152,N_14035);
or U14750 (N_14750,N_14389,N_14379);
or U14751 (N_14751,N_14039,N_14232);
nand U14752 (N_14752,N_14469,N_14399);
xor U14753 (N_14753,N_14369,N_14229);
nor U14754 (N_14754,N_14315,N_14122);
or U14755 (N_14755,N_14444,N_14397);
and U14756 (N_14756,N_14077,N_14111);
nand U14757 (N_14757,N_14103,N_14260);
or U14758 (N_14758,N_14420,N_14280);
or U14759 (N_14759,N_14274,N_14192);
or U14760 (N_14760,N_14258,N_14334);
nand U14761 (N_14761,N_14125,N_14204);
nor U14762 (N_14762,N_14293,N_14083);
nor U14763 (N_14763,N_14280,N_14063);
nand U14764 (N_14764,N_14402,N_14285);
nand U14765 (N_14765,N_14063,N_14095);
nand U14766 (N_14766,N_14470,N_14261);
or U14767 (N_14767,N_14226,N_14297);
or U14768 (N_14768,N_14178,N_14081);
nor U14769 (N_14769,N_14117,N_14310);
nor U14770 (N_14770,N_14336,N_14353);
nand U14771 (N_14771,N_14166,N_14110);
or U14772 (N_14772,N_14419,N_14324);
or U14773 (N_14773,N_14475,N_14497);
or U14774 (N_14774,N_14103,N_14402);
and U14775 (N_14775,N_14293,N_14155);
or U14776 (N_14776,N_14479,N_14413);
nor U14777 (N_14777,N_14149,N_14288);
or U14778 (N_14778,N_14213,N_14251);
or U14779 (N_14779,N_14278,N_14041);
and U14780 (N_14780,N_14221,N_14312);
nor U14781 (N_14781,N_14437,N_14463);
nand U14782 (N_14782,N_14216,N_14382);
or U14783 (N_14783,N_14041,N_14098);
nand U14784 (N_14784,N_14152,N_14470);
and U14785 (N_14785,N_14020,N_14416);
nor U14786 (N_14786,N_14290,N_14159);
and U14787 (N_14787,N_14245,N_14144);
and U14788 (N_14788,N_14186,N_14429);
nor U14789 (N_14789,N_14105,N_14475);
nand U14790 (N_14790,N_14289,N_14153);
and U14791 (N_14791,N_14363,N_14035);
and U14792 (N_14792,N_14374,N_14057);
nor U14793 (N_14793,N_14335,N_14435);
or U14794 (N_14794,N_14384,N_14198);
and U14795 (N_14795,N_14388,N_14268);
nor U14796 (N_14796,N_14222,N_14011);
nor U14797 (N_14797,N_14329,N_14213);
nand U14798 (N_14798,N_14405,N_14079);
and U14799 (N_14799,N_14074,N_14259);
xnor U14800 (N_14800,N_14263,N_14291);
nor U14801 (N_14801,N_14329,N_14060);
nor U14802 (N_14802,N_14463,N_14462);
nor U14803 (N_14803,N_14495,N_14039);
nand U14804 (N_14804,N_14212,N_14057);
and U14805 (N_14805,N_14301,N_14360);
nand U14806 (N_14806,N_14450,N_14133);
nand U14807 (N_14807,N_14023,N_14340);
nand U14808 (N_14808,N_14483,N_14311);
nor U14809 (N_14809,N_14174,N_14254);
nand U14810 (N_14810,N_14404,N_14060);
and U14811 (N_14811,N_14353,N_14405);
or U14812 (N_14812,N_14271,N_14331);
nand U14813 (N_14813,N_14310,N_14102);
and U14814 (N_14814,N_14028,N_14383);
and U14815 (N_14815,N_14182,N_14258);
nor U14816 (N_14816,N_14077,N_14037);
or U14817 (N_14817,N_14174,N_14473);
nand U14818 (N_14818,N_14070,N_14472);
and U14819 (N_14819,N_14217,N_14031);
nor U14820 (N_14820,N_14336,N_14035);
nor U14821 (N_14821,N_14262,N_14031);
and U14822 (N_14822,N_14451,N_14496);
nand U14823 (N_14823,N_14129,N_14262);
and U14824 (N_14824,N_14289,N_14287);
and U14825 (N_14825,N_14418,N_14382);
nand U14826 (N_14826,N_14267,N_14224);
or U14827 (N_14827,N_14193,N_14484);
nor U14828 (N_14828,N_14022,N_14279);
nand U14829 (N_14829,N_14311,N_14495);
or U14830 (N_14830,N_14401,N_14281);
or U14831 (N_14831,N_14450,N_14356);
or U14832 (N_14832,N_14230,N_14294);
nor U14833 (N_14833,N_14279,N_14125);
or U14834 (N_14834,N_14278,N_14005);
or U14835 (N_14835,N_14051,N_14295);
nand U14836 (N_14836,N_14213,N_14202);
or U14837 (N_14837,N_14075,N_14269);
or U14838 (N_14838,N_14457,N_14123);
nor U14839 (N_14839,N_14413,N_14308);
or U14840 (N_14840,N_14194,N_14017);
nand U14841 (N_14841,N_14282,N_14491);
nand U14842 (N_14842,N_14486,N_14168);
nor U14843 (N_14843,N_14025,N_14169);
nor U14844 (N_14844,N_14169,N_14364);
nor U14845 (N_14845,N_14121,N_14265);
or U14846 (N_14846,N_14178,N_14372);
or U14847 (N_14847,N_14138,N_14435);
and U14848 (N_14848,N_14266,N_14096);
or U14849 (N_14849,N_14139,N_14074);
or U14850 (N_14850,N_14449,N_14435);
and U14851 (N_14851,N_14234,N_14188);
nand U14852 (N_14852,N_14097,N_14133);
nor U14853 (N_14853,N_14338,N_14059);
or U14854 (N_14854,N_14366,N_14205);
nor U14855 (N_14855,N_14110,N_14382);
xor U14856 (N_14856,N_14023,N_14127);
and U14857 (N_14857,N_14403,N_14428);
or U14858 (N_14858,N_14330,N_14483);
and U14859 (N_14859,N_14324,N_14298);
or U14860 (N_14860,N_14175,N_14437);
and U14861 (N_14861,N_14310,N_14003);
nand U14862 (N_14862,N_14205,N_14378);
nand U14863 (N_14863,N_14464,N_14153);
nor U14864 (N_14864,N_14182,N_14059);
and U14865 (N_14865,N_14205,N_14240);
nor U14866 (N_14866,N_14324,N_14491);
and U14867 (N_14867,N_14497,N_14150);
nand U14868 (N_14868,N_14247,N_14316);
and U14869 (N_14869,N_14090,N_14443);
nand U14870 (N_14870,N_14214,N_14033);
or U14871 (N_14871,N_14394,N_14119);
or U14872 (N_14872,N_14117,N_14321);
nor U14873 (N_14873,N_14168,N_14145);
nor U14874 (N_14874,N_14176,N_14383);
nor U14875 (N_14875,N_14371,N_14236);
and U14876 (N_14876,N_14337,N_14169);
or U14877 (N_14877,N_14046,N_14009);
or U14878 (N_14878,N_14285,N_14469);
and U14879 (N_14879,N_14253,N_14001);
xnor U14880 (N_14880,N_14199,N_14126);
nor U14881 (N_14881,N_14267,N_14177);
nor U14882 (N_14882,N_14249,N_14195);
nor U14883 (N_14883,N_14132,N_14144);
nor U14884 (N_14884,N_14080,N_14169);
or U14885 (N_14885,N_14166,N_14010);
and U14886 (N_14886,N_14481,N_14149);
or U14887 (N_14887,N_14141,N_14285);
nand U14888 (N_14888,N_14422,N_14440);
and U14889 (N_14889,N_14328,N_14097);
nand U14890 (N_14890,N_14332,N_14167);
nand U14891 (N_14891,N_14002,N_14359);
and U14892 (N_14892,N_14425,N_14344);
nand U14893 (N_14893,N_14234,N_14462);
and U14894 (N_14894,N_14411,N_14473);
and U14895 (N_14895,N_14236,N_14434);
nand U14896 (N_14896,N_14231,N_14428);
xor U14897 (N_14897,N_14289,N_14319);
nor U14898 (N_14898,N_14292,N_14184);
or U14899 (N_14899,N_14190,N_14369);
xor U14900 (N_14900,N_14034,N_14452);
or U14901 (N_14901,N_14420,N_14386);
and U14902 (N_14902,N_14310,N_14435);
or U14903 (N_14903,N_14098,N_14219);
nor U14904 (N_14904,N_14157,N_14145);
and U14905 (N_14905,N_14274,N_14465);
nor U14906 (N_14906,N_14119,N_14227);
nor U14907 (N_14907,N_14388,N_14469);
nand U14908 (N_14908,N_14328,N_14026);
nand U14909 (N_14909,N_14171,N_14440);
or U14910 (N_14910,N_14420,N_14203);
and U14911 (N_14911,N_14404,N_14163);
and U14912 (N_14912,N_14069,N_14238);
or U14913 (N_14913,N_14270,N_14001);
nand U14914 (N_14914,N_14420,N_14325);
or U14915 (N_14915,N_14217,N_14332);
nor U14916 (N_14916,N_14420,N_14432);
nor U14917 (N_14917,N_14355,N_14379);
nand U14918 (N_14918,N_14214,N_14284);
and U14919 (N_14919,N_14329,N_14001);
nand U14920 (N_14920,N_14297,N_14470);
nand U14921 (N_14921,N_14129,N_14190);
nand U14922 (N_14922,N_14267,N_14076);
nand U14923 (N_14923,N_14014,N_14443);
xor U14924 (N_14924,N_14207,N_14467);
and U14925 (N_14925,N_14121,N_14098);
and U14926 (N_14926,N_14083,N_14230);
nor U14927 (N_14927,N_14229,N_14044);
and U14928 (N_14928,N_14012,N_14042);
and U14929 (N_14929,N_14253,N_14259);
nand U14930 (N_14930,N_14402,N_14101);
nand U14931 (N_14931,N_14399,N_14337);
nand U14932 (N_14932,N_14087,N_14069);
or U14933 (N_14933,N_14263,N_14389);
and U14934 (N_14934,N_14456,N_14454);
nor U14935 (N_14935,N_14197,N_14173);
and U14936 (N_14936,N_14379,N_14277);
nor U14937 (N_14937,N_14303,N_14473);
nor U14938 (N_14938,N_14071,N_14246);
nand U14939 (N_14939,N_14227,N_14322);
nor U14940 (N_14940,N_14248,N_14130);
and U14941 (N_14941,N_14114,N_14140);
and U14942 (N_14942,N_14371,N_14419);
or U14943 (N_14943,N_14004,N_14103);
and U14944 (N_14944,N_14411,N_14165);
or U14945 (N_14945,N_14240,N_14057);
and U14946 (N_14946,N_14059,N_14212);
nand U14947 (N_14947,N_14176,N_14152);
or U14948 (N_14948,N_14465,N_14172);
nand U14949 (N_14949,N_14489,N_14256);
or U14950 (N_14950,N_14137,N_14009);
and U14951 (N_14951,N_14134,N_14391);
or U14952 (N_14952,N_14435,N_14141);
or U14953 (N_14953,N_14146,N_14390);
nand U14954 (N_14954,N_14450,N_14065);
nor U14955 (N_14955,N_14432,N_14144);
or U14956 (N_14956,N_14226,N_14461);
nor U14957 (N_14957,N_14138,N_14306);
nand U14958 (N_14958,N_14467,N_14342);
and U14959 (N_14959,N_14120,N_14248);
nand U14960 (N_14960,N_14003,N_14246);
nand U14961 (N_14961,N_14414,N_14158);
and U14962 (N_14962,N_14346,N_14141);
nand U14963 (N_14963,N_14445,N_14368);
nand U14964 (N_14964,N_14438,N_14157);
or U14965 (N_14965,N_14214,N_14377);
nor U14966 (N_14966,N_14254,N_14424);
or U14967 (N_14967,N_14049,N_14251);
and U14968 (N_14968,N_14204,N_14460);
or U14969 (N_14969,N_14446,N_14405);
and U14970 (N_14970,N_14196,N_14404);
and U14971 (N_14971,N_14146,N_14038);
nand U14972 (N_14972,N_14259,N_14087);
and U14973 (N_14973,N_14043,N_14384);
xnor U14974 (N_14974,N_14214,N_14274);
and U14975 (N_14975,N_14405,N_14167);
nor U14976 (N_14976,N_14009,N_14152);
and U14977 (N_14977,N_14188,N_14282);
and U14978 (N_14978,N_14307,N_14339);
or U14979 (N_14979,N_14374,N_14016);
nand U14980 (N_14980,N_14472,N_14306);
and U14981 (N_14981,N_14200,N_14473);
and U14982 (N_14982,N_14136,N_14366);
or U14983 (N_14983,N_14198,N_14308);
or U14984 (N_14984,N_14012,N_14159);
or U14985 (N_14985,N_14404,N_14479);
or U14986 (N_14986,N_14206,N_14198);
xor U14987 (N_14987,N_14073,N_14062);
and U14988 (N_14988,N_14374,N_14178);
and U14989 (N_14989,N_14426,N_14335);
and U14990 (N_14990,N_14247,N_14136);
nor U14991 (N_14991,N_14004,N_14152);
nand U14992 (N_14992,N_14348,N_14044);
nor U14993 (N_14993,N_14194,N_14334);
nand U14994 (N_14994,N_14355,N_14229);
and U14995 (N_14995,N_14424,N_14130);
nor U14996 (N_14996,N_14085,N_14364);
nand U14997 (N_14997,N_14491,N_14439);
or U14998 (N_14998,N_14210,N_14331);
nand U14999 (N_14999,N_14276,N_14156);
xor U15000 (N_15000,N_14950,N_14984);
nand U15001 (N_15001,N_14542,N_14605);
nand U15002 (N_15002,N_14664,N_14949);
or U15003 (N_15003,N_14595,N_14970);
or U15004 (N_15004,N_14942,N_14543);
and U15005 (N_15005,N_14990,N_14904);
or U15006 (N_15006,N_14886,N_14860);
nor U15007 (N_15007,N_14686,N_14819);
nand U15008 (N_15008,N_14853,N_14678);
nand U15009 (N_15009,N_14934,N_14926);
nor U15010 (N_15010,N_14539,N_14932);
and U15011 (N_15011,N_14612,N_14710);
nor U15012 (N_15012,N_14703,N_14712);
nor U15013 (N_15013,N_14848,N_14788);
nor U15014 (N_15014,N_14776,N_14622);
and U15015 (N_15015,N_14696,N_14509);
or U15016 (N_15016,N_14545,N_14842);
or U15017 (N_15017,N_14979,N_14514);
or U15018 (N_15018,N_14974,N_14516);
nand U15019 (N_15019,N_14709,N_14851);
nor U15020 (N_15020,N_14689,N_14895);
or U15021 (N_15021,N_14897,N_14981);
and U15022 (N_15022,N_14881,N_14646);
and U15023 (N_15023,N_14922,N_14898);
and U15024 (N_15024,N_14796,N_14896);
and U15025 (N_15025,N_14517,N_14994);
and U15026 (N_15026,N_14617,N_14915);
nand U15027 (N_15027,N_14794,N_14580);
nand U15028 (N_15028,N_14911,N_14756);
or U15029 (N_15029,N_14618,N_14875);
xnor U15030 (N_15030,N_14912,N_14791);
and U15031 (N_15031,N_14939,N_14888);
or U15032 (N_15032,N_14845,N_14682);
nand U15033 (N_15033,N_14836,N_14634);
and U15034 (N_15034,N_14874,N_14597);
or U15035 (N_15035,N_14620,N_14591);
nand U15036 (N_15036,N_14892,N_14577);
and U15037 (N_15037,N_14565,N_14831);
or U15038 (N_15038,N_14906,N_14744);
or U15039 (N_15039,N_14515,N_14790);
nand U15040 (N_15040,N_14699,N_14698);
nand U15041 (N_15041,N_14977,N_14708);
xor U15042 (N_15042,N_14769,N_14735);
or U15043 (N_15043,N_14601,N_14960);
nand U15044 (N_15044,N_14623,N_14676);
nand U15045 (N_15045,N_14792,N_14723);
nand U15046 (N_15046,N_14571,N_14876);
nor U15047 (N_15047,N_14726,N_14508);
or U15048 (N_15048,N_14971,N_14887);
or U15049 (N_15049,N_14656,N_14611);
and U15050 (N_15050,N_14606,N_14745);
and U15051 (N_15051,N_14841,N_14732);
nand U15052 (N_15052,N_14569,N_14899);
and U15053 (N_15053,N_14529,N_14551);
nand U15054 (N_15054,N_14574,N_14501);
or U15055 (N_15055,N_14777,N_14650);
or U15056 (N_15056,N_14525,N_14833);
and U15057 (N_15057,N_14568,N_14614);
or U15058 (N_15058,N_14955,N_14958);
nor U15059 (N_15059,N_14628,N_14588);
or U15060 (N_15060,N_14714,N_14763);
and U15061 (N_15061,N_14590,N_14579);
and U15062 (N_15062,N_14780,N_14827);
and U15063 (N_15063,N_14558,N_14526);
or U15064 (N_15064,N_14805,N_14843);
xnor U15065 (N_15065,N_14826,N_14690);
or U15066 (N_15066,N_14559,N_14787);
or U15067 (N_15067,N_14861,N_14866);
nand U15068 (N_15068,N_14627,N_14941);
or U15069 (N_15069,N_14644,N_14933);
or U15070 (N_15070,N_14505,N_14662);
and U15071 (N_15071,N_14832,N_14547);
or U15072 (N_15072,N_14901,N_14661);
or U15073 (N_15073,N_14809,N_14964);
nor U15074 (N_15074,N_14625,N_14671);
or U15075 (N_15075,N_14862,N_14931);
and U15076 (N_15076,N_14695,N_14564);
and U15077 (N_15077,N_14867,N_14968);
and U15078 (N_15078,N_14540,N_14534);
and U15079 (N_15079,N_14997,N_14582);
and U15080 (N_15080,N_14637,N_14679);
nand U15081 (N_15081,N_14996,N_14834);
or U15082 (N_15082,N_14655,N_14600);
and U15083 (N_15083,N_14716,N_14761);
xnor U15084 (N_15084,N_14885,N_14718);
nand U15085 (N_15085,N_14585,N_14755);
or U15086 (N_15086,N_14506,N_14803);
nor U15087 (N_15087,N_14513,N_14518);
nor U15088 (N_15088,N_14621,N_14511);
nand U15089 (N_15089,N_14793,N_14795);
nand U15090 (N_15090,N_14757,N_14880);
nor U15091 (N_15091,N_14555,N_14884);
or U15092 (N_15092,N_14654,N_14573);
and U15093 (N_15093,N_14663,N_14594);
nand U15094 (N_15094,N_14976,N_14812);
and U15095 (N_15095,N_14639,N_14632);
or U15096 (N_15096,N_14658,N_14677);
and U15097 (N_15097,N_14570,N_14972);
or U15098 (N_15098,N_14849,N_14672);
or U15099 (N_15099,N_14648,N_14584);
and U15100 (N_15100,N_14856,N_14747);
nand U15101 (N_15101,N_14989,N_14925);
nand U15102 (N_15102,N_14711,N_14552);
and U15103 (N_15103,N_14838,N_14967);
or U15104 (N_15104,N_14855,N_14905);
and U15105 (N_15105,N_14903,N_14801);
or U15106 (N_15106,N_14765,N_14828);
and U15107 (N_15107,N_14993,N_14754);
and U15108 (N_15108,N_14742,N_14953);
nor U15109 (N_15109,N_14798,N_14642);
nand U15110 (N_15110,N_14500,N_14963);
nor U15111 (N_15111,N_14909,N_14956);
and U15112 (N_15112,N_14604,N_14613);
and U15113 (N_15113,N_14669,N_14523);
nor U15114 (N_15114,N_14507,N_14969);
and U15115 (N_15115,N_14846,N_14715);
and U15116 (N_15116,N_14923,N_14945);
and U15117 (N_15117,N_14973,N_14952);
and U15118 (N_15118,N_14921,N_14748);
xnor U15119 (N_15119,N_14725,N_14512);
nor U15120 (N_15120,N_14734,N_14636);
or U15121 (N_15121,N_14946,N_14847);
nor U15122 (N_15122,N_14766,N_14645);
or U15123 (N_15123,N_14857,N_14771);
xnor U15124 (N_15124,N_14630,N_14889);
nand U15125 (N_15125,N_14821,N_14865);
nand U15126 (N_15126,N_14774,N_14680);
nor U15127 (N_15127,N_14802,N_14635);
or U15128 (N_15128,N_14685,N_14626);
and U15129 (N_15129,N_14729,N_14930);
and U15130 (N_15130,N_14998,N_14666);
nor U15131 (N_15131,N_14687,N_14739);
nor U15132 (N_15132,N_14631,N_14829);
or U15133 (N_15133,N_14649,N_14693);
and U15134 (N_15134,N_14948,N_14770);
or U15135 (N_15135,N_14657,N_14550);
nand U15136 (N_15136,N_14879,N_14728);
nand U15137 (N_15137,N_14562,N_14781);
nand U15138 (N_15138,N_14837,N_14786);
nor U15139 (N_15139,N_14814,N_14920);
nor U15140 (N_15140,N_14951,N_14528);
nand U15141 (N_15141,N_14872,N_14720);
nand U15142 (N_15142,N_14741,N_14882);
or U15143 (N_15143,N_14944,N_14587);
or U15144 (N_15144,N_14520,N_14918);
nor U15145 (N_15145,N_14576,N_14760);
nor U15146 (N_15146,N_14916,N_14927);
nand U15147 (N_15147,N_14667,N_14533);
or U15148 (N_15148,N_14894,N_14554);
or U15149 (N_15149,N_14980,N_14844);
nand U15150 (N_15150,N_14924,N_14936);
or U15151 (N_15151,N_14722,N_14929);
or U15152 (N_15152,N_14633,N_14919);
nor U15153 (N_15153,N_14531,N_14959);
or U15154 (N_15154,N_14753,N_14768);
nand U15155 (N_15155,N_14987,N_14638);
nand U15156 (N_15156,N_14779,N_14991);
or U15157 (N_15157,N_14675,N_14799);
or U15158 (N_15158,N_14624,N_14824);
xor U15159 (N_15159,N_14684,N_14615);
or U15160 (N_15160,N_14940,N_14581);
nor U15161 (N_15161,N_14785,N_14806);
or U15162 (N_15162,N_14810,N_14691);
or U15163 (N_15163,N_14752,N_14983);
nor U15164 (N_15164,N_14784,N_14530);
nor U15165 (N_15165,N_14891,N_14608);
and U15166 (N_15166,N_14640,N_14907);
or U15167 (N_15167,N_14999,N_14789);
nand U15168 (N_15168,N_14557,N_14721);
or U15169 (N_15169,N_14902,N_14823);
or U15170 (N_15170,N_14840,N_14816);
or U15171 (N_15171,N_14578,N_14572);
and U15172 (N_15172,N_14536,N_14750);
nor U15173 (N_15173,N_14730,N_14727);
nand U15174 (N_15174,N_14521,N_14811);
and U15175 (N_15175,N_14982,N_14873);
or U15176 (N_15176,N_14758,N_14546);
and U15177 (N_15177,N_14705,N_14743);
nand U15178 (N_15178,N_14825,N_14870);
nor U15179 (N_15179,N_14878,N_14702);
or U15180 (N_15180,N_14704,N_14673);
nor U15181 (N_15181,N_14804,N_14719);
and U15182 (N_15182,N_14852,N_14775);
nand U15183 (N_15183,N_14822,N_14913);
and U15184 (N_15184,N_14544,N_14817);
and U15185 (N_15185,N_14589,N_14619);
and U15186 (N_15186,N_14566,N_14778);
nand U15187 (N_15187,N_14858,N_14800);
nor U15188 (N_15188,N_14808,N_14773);
nand U15189 (N_15189,N_14724,N_14935);
nand U15190 (N_15190,N_14556,N_14736);
nor U15191 (N_15191,N_14890,N_14504);
or U15192 (N_15192,N_14864,N_14740);
or U15193 (N_15193,N_14586,N_14641);
xnor U15194 (N_15194,N_14561,N_14647);
and U15195 (N_15195,N_14681,N_14807);
nor U15196 (N_15196,N_14535,N_14797);
nand U15197 (N_15197,N_14522,N_14975);
and U15198 (N_15198,N_14563,N_14575);
and U15199 (N_15199,N_14524,N_14961);
nor U15200 (N_15200,N_14995,N_14532);
and U15201 (N_15201,N_14707,N_14553);
nand U15202 (N_15202,N_14937,N_14697);
or U15203 (N_15203,N_14603,N_14610);
or U15204 (N_15204,N_14717,N_14954);
or U15205 (N_15205,N_14738,N_14830);
xor U15206 (N_15206,N_14985,N_14914);
or U15207 (N_15207,N_14660,N_14527);
and U15208 (N_15208,N_14883,N_14674);
or U15209 (N_15209,N_14598,N_14772);
or U15210 (N_15210,N_14746,N_14868);
nand U15211 (N_15211,N_14762,N_14957);
nor U15212 (N_15212,N_14652,N_14908);
nand U15213 (N_15213,N_14694,N_14668);
nor U15214 (N_15214,N_14541,N_14502);
and U15215 (N_15215,N_14503,N_14871);
nor U15216 (N_15216,N_14938,N_14859);
nor U15217 (N_15217,N_14629,N_14992);
nor U15218 (N_15218,N_14737,N_14583);
or U15219 (N_15219,N_14820,N_14659);
nor U15220 (N_15220,N_14607,N_14602);
nor U15221 (N_15221,N_14665,N_14733);
nand U15222 (N_15222,N_14700,N_14813);
nand U15223 (N_15223,N_14643,N_14850);
nand U15224 (N_15224,N_14962,N_14567);
nand U15225 (N_15225,N_14548,N_14749);
nor U15226 (N_15226,N_14943,N_14653);
nor U15227 (N_15227,N_14713,N_14988);
nor U15228 (N_15228,N_14818,N_14701);
and U15229 (N_15229,N_14549,N_14978);
nand U15230 (N_15230,N_14835,N_14965);
and U15231 (N_15231,N_14609,N_14966);
and U15232 (N_15232,N_14616,N_14782);
and U15233 (N_15233,N_14537,N_14519);
or U15234 (N_15234,N_14731,N_14910);
nor U15235 (N_15235,N_14764,N_14706);
or U15236 (N_15236,N_14869,N_14593);
xor U15237 (N_15237,N_14596,N_14683);
xor U15238 (N_15238,N_14592,N_14751);
nand U15239 (N_15239,N_14560,N_14893);
and U15240 (N_15240,N_14815,N_14767);
nor U15241 (N_15241,N_14759,N_14877);
nand U15242 (N_15242,N_14986,N_14510);
nand U15243 (N_15243,N_14538,N_14900);
nand U15244 (N_15244,N_14670,N_14688);
and U15245 (N_15245,N_14928,N_14947);
and U15246 (N_15246,N_14783,N_14917);
nor U15247 (N_15247,N_14692,N_14854);
nand U15248 (N_15248,N_14839,N_14599);
or U15249 (N_15249,N_14863,N_14651);
or U15250 (N_15250,N_14657,N_14710);
nor U15251 (N_15251,N_14539,N_14695);
nor U15252 (N_15252,N_14884,N_14784);
nor U15253 (N_15253,N_14984,N_14591);
nor U15254 (N_15254,N_14937,N_14851);
or U15255 (N_15255,N_14687,N_14851);
or U15256 (N_15256,N_14605,N_14798);
nor U15257 (N_15257,N_14821,N_14603);
nand U15258 (N_15258,N_14771,N_14740);
nor U15259 (N_15259,N_14759,N_14826);
and U15260 (N_15260,N_14510,N_14719);
nor U15261 (N_15261,N_14878,N_14916);
or U15262 (N_15262,N_14675,N_14673);
and U15263 (N_15263,N_14910,N_14933);
and U15264 (N_15264,N_14783,N_14644);
or U15265 (N_15265,N_14665,N_14512);
nand U15266 (N_15266,N_14549,N_14765);
nand U15267 (N_15267,N_14895,N_14825);
nor U15268 (N_15268,N_14503,N_14598);
nand U15269 (N_15269,N_14799,N_14601);
and U15270 (N_15270,N_14516,N_14795);
or U15271 (N_15271,N_14729,N_14909);
nand U15272 (N_15272,N_14580,N_14840);
nor U15273 (N_15273,N_14607,N_14950);
or U15274 (N_15274,N_14518,N_14963);
or U15275 (N_15275,N_14669,N_14788);
or U15276 (N_15276,N_14501,N_14978);
and U15277 (N_15277,N_14573,N_14568);
and U15278 (N_15278,N_14756,N_14945);
or U15279 (N_15279,N_14742,N_14611);
or U15280 (N_15280,N_14681,N_14512);
nand U15281 (N_15281,N_14630,N_14633);
xor U15282 (N_15282,N_14793,N_14699);
and U15283 (N_15283,N_14536,N_14955);
nand U15284 (N_15284,N_14841,N_14810);
nand U15285 (N_15285,N_14503,N_14767);
and U15286 (N_15286,N_14511,N_14709);
xor U15287 (N_15287,N_14849,N_14628);
nor U15288 (N_15288,N_14645,N_14661);
nand U15289 (N_15289,N_14603,N_14754);
or U15290 (N_15290,N_14984,N_14602);
and U15291 (N_15291,N_14947,N_14783);
and U15292 (N_15292,N_14639,N_14726);
or U15293 (N_15293,N_14697,N_14705);
and U15294 (N_15294,N_14689,N_14760);
or U15295 (N_15295,N_14747,N_14799);
or U15296 (N_15296,N_14609,N_14686);
nand U15297 (N_15297,N_14705,N_14511);
nor U15298 (N_15298,N_14849,N_14949);
and U15299 (N_15299,N_14585,N_14797);
or U15300 (N_15300,N_14599,N_14979);
and U15301 (N_15301,N_14546,N_14542);
nand U15302 (N_15302,N_14697,N_14534);
nand U15303 (N_15303,N_14971,N_14661);
and U15304 (N_15304,N_14639,N_14513);
nand U15305 (N_15305,N_14679,N_14815);
nand U15306 (N_15306,N_14652,N_14968);
xnor U15307 (N_15307,N_14569,N_14993);
nand U15308 (N_15308,N_14504,N_14775);
nand U15309 (N_15309,N_14924,N_14897);
or U15310 (N_15310,N_14835,N_14522);
nor U15311 (N_15311,N_14589,N_14889);
or U15312 (N_15312,N_14750,N_14634);
and U15313 (N_15313,N_14949,N_14926);
or U15314 (N_15314,N_14870,N_14761);
or U15315 (N_15315,N_14701,N_14794);
nor U15316 (N_15316,N_14637,N_14962);
and U15317 (N_15317,N_14631,N_14731);
or U15318 (N_15318,N_14899,N_14881);
nand U15319 (N_15319,N_14844,N_14946);
or U15320 (N_15320,N_14603,N_14852);
nor U15321 (N_15321,N_14626,N_14977);
nor U15322 (N_15322,N_14599,N_14687);
and U15323 (N_15323,N_14918,N_14504);
nand U15324 (N_15324,N_14606,N_14954);
and U15325 (N_15325,N_14994,N_14513);
nor U15326 (N_15326,N_14515,N_14963);
nand U15327 (N_15327,N_14589,N_14793);
nand U15328 (N_15328,N_14589,N_14626);
nand U15329 (N_15329,N_14819,N_14853);
and U15330 (N_15330,N_14889,N_14569);
or U15331 (N_15331,N_14797,N_14736);
or U15332 (N_15332,N_14663,N_14509);
xor U15333 (N_15333,N_14709,N_14540);
or U15334 (N_15334,N_14712,N_14523);
or U15335 (N_15335,N_14623,N_14831);
and U15336 (N_15336,N_14844,N_14957);
or U15337 (N_15337,N_14569,N_14872);
and U15338 (N_15338,N_14934,N_14553);
and U15339 (N_15339,N_14613,N_14829);
and U15340 (N_15340,N_14750,N_14779);
or U15341 (N_15341,N_14780,N_14679);
or U15342 (N_15342,N_14792,N_14746);
and U15343 (N_15343,N_14547,N_14613);
nand U15344 (N_15344,N_14740,N_14943);
and U15345 (N_15345,N_14778,N_14759);
nand U15346 (N_15346,N_14828,N_14838);
nand U15347 (N_15347,N_14972,N_14860);
and U15348 (N_15348,N_14635,N_14964);
or U15349 (N_15349,N_14784,N_14819);
or U15350 (N_15350,N_14504,N_14980);
or U15351 (N_15351,N_14810,N_14898);
nand U15352 (N_15352,N_14782,N_14603);
nand U15353 (N_15353,N_14546,N_14912);
nor U15354 (N_15354,N_14615,N_14680);
nor U15355 (N_15355,N_14967,N_14855);
nor U15356 (N_15356,N_14963,N_14638);
nand U15357 (N_15357,N_14909,N_14742);
or U15358 (N_15358,N_14591,N_14906);
xnor U15359 (N_15359,N_14704,N_14964);
and U15360 (N_15360,N_14575,N_14826);
and U15361 (N_15361,N_14933,N_14745);
nor U15362 (N_15362,N_14922,N_14579);
and U15363 (N_15363,N_14542,N_14524);
nand U15364 (N_15364,N_14598,N_14727);
or U15365 (N_15365,N_14789,N_14588);
nand U15366 (N_15366,N_14681,N_14827);
and U15367 (N_15367,N_14648,N_14775);
nor U15368 (N_15368,N_14509,N_14659);
and U15369 (N_15369,N_14681,N_14771);
nor U15370 (N_15370,N_14646,N_14551);
and U15371 (N_15371,N_14508,N_14586);
nand U15372 (N_15372,N_14657,N_14908);
and U15373 (N_15373,N_14715,N_14568);
or U15374 (N_15374,N_14594,N_14646);
and U15375 (N_15375,N_14765,N_14699);
or U15376 (N_15376,N_14713,N_14686);
and U15377 (N_15377,N_14507,N_14977);
nand U15378 (N_15378,N_14989,N_14505);
and U15379 (N_15379,N_14686,N_14975);
nor U15380 (N_15380,N_14860,N_14642);
nand U15381 (N_15381,N_14570,N_14617);
and U15382 (N_15382,N_14956,N_14830);
or U15383 (N_15383,N_14693,N_14520);
nor U15384 (N_15384,N_14813,N_14921);
nor U15385 (N_15385,N_14682,N_14589);
and U15386 (N_15386,N_14738,N_14979);
nor U15387 (N_15387,N_14762,N_14909);
and U15388 (N_15388,N_14547,N_14918);
nand U15389 (N_15389,N_14914,N_14818);
and U15390 (N_15390,N_14633,N_14522);
and U15391 (N_15391,N_14958,N_14828);
nor U15392 (N_15392,N_14611,N_14567);
or U15393 (N_15393,N_14872,N_14788);
or U15394 (N_15394,N_14888,N_14982);
nand U15395 (N_15395,N_14549,N_14685);
nor U15396 (N_15396,N_14759,N_14912);
nand U15397 (N_15397,N_14957,N_14772);
nor U15398 (N_15398,N_14816,N_14649);
and U15399 (N_15399,N_14706,N_14827);
nand U15400 (N_15400,N_14885,N_14872);
nand U15401 (N_15401,N_14639,N_14906);
and U15402 (N_15402,N_14737,N_14764);
or U15403 (N_15403,N_14844,N_14620);
or U15404 (N_15404,N_14907,N_14762);
nand U15405 (N_15405,N_14693,N_14656);
nand U15406 (N_15406,N_14837,N_14934);
nor U15407 (N_15407,N_14873,N_14608);
nor U15408 (N_15408,N_14569,N_14589);
or U15409 (N_15409,N_14567,N_14759);
nor U15410 (N_15410,N_14870,N_14886);
nor U15411 (N_15411,N_14537,N_14562);
or U15412 (N_15412,N_14773,N_14811);
nor U15413 (N_15413,N_14813,N_14997);
or U15414 (N_15414,N_14657,N_14585);
and U15415 (N_15415,N_14553,N_14866);
and U15416 (N_15416,N_14929,N_14992);
nand U15417 (N_15417,N_14531,N_14854);
nand U15418 (N_15418,N_14926,N_14854);
nor U15419 (N_15419,N_14758,N_14507);
or U15420 (N_15420,N_14834,N_14646);
and U15421 (N_15421,N_14790,N_14740);
or U15422 (N_15422,N_14989,N_14911);
or U15423 (N_15423,N_14530,N_14611);
nand U15424 (N_15424,N_14650,N_14665);
or U15425 (N_15425,N_14854,N_14979);
nand U15426 (N_15426,N_14991,N_14656);
nor U15427 (N_15427,N_14775,N_14510);
nor U15428 (N_15428,N_14994,N_14614);
nand U15429 (N_15429,N_14953,N_14847);
nand U15430 (N_15430,N_14779,N_14928);
or U15431 (N_15431,N_14597,N_14540);
or U15432 (N_15432,N_14761,N_14885);
nor U15433 (N_15433,N_14687,N_14538);
or U15434 (N_15434,N_14982,N_14771);
nand U15435 (N_15435,N_14531,N_14947);
nand U15436 (N_15436,N_14649,N_14793);
or U15437 (N_15437,N_14989,N_14763);
nand U15438 (N_15438,N_14870,N_14996);
and U15439 (N_15439,N_14932,N_14976);
nand U15440 (N_15440,N_14562,N_14518);
nor U15441 (N_15441,N_14763,N_14675);
nor U15442 (N_15442,N_14580,N_14662);
nor U15443 (N_15443,N_14659,N_14651);
or U15444 (N_15444,N_14882,N_14937);
nand U15445 (N_15445,N_14800,N_14566);
nor U15446 (N_15446,N_14771,N_14832);
nand U15447 (N_15447,N_14981,N_14854);
and U15448 (N_15448,N_14801,N_14713);
nand U15449 (N_15449,N_14533,N_14625);
and U15450 (N_15450,N_14896,N_14694);
and U15451 (N_15451,N_14822,N_14619);
nand U15452 (N_15452,N_14825,N_14703);
nand U15453 (N_15453,N_14898,N_14572);
or U15454 (N_15454,N_14516,N_14701);
nor U15455 (N_15455,N_14872,N_14849);
or U15456 (N_15456,N_14735,N_14603);
and U15457 (N_15457,N_14944,N_14824);
nand U15458 (N_15458,N_14928,N_14870);
nor U15459 (N_15459,N_14998,N_14895);
and U15460 (N_15460,N_14987,N_14632);
nor U15461 (N_15461,N_14667,N_14883);
nor U15462 (N_15462,N_14661,N_14948);
and U15463 (N_15463,N_14820,N_14689);
nor U15464 (N_15464,N_14928,N_14804);
and U15465 (N_15465,N_14503,N_14679);
nand U15466 (N_15466,N_14661,N_14805);
or U15467 (N_15467,N_14544,N_14970);
nor U15468 (N_15468,N_14919,N_14531);
and U15469 (N_15469,N_14995,N_14592);
nor U15470 (N_15470,N_14990,N_14841);
and U15471 (N_15471,N_14685,N_14773);
nor U15472 (N_15472,N_14730,N_14801);
and U15473 (N_15473,N_14912,N_14992);
and U15474 (N_15474,N_14846,N_14594);
nand U15475 (N_15475,N_14708,N_14958);
and U15476 (N_15476,N_14895,N_14623);
nand U15477 (N_15477,N_14592,N_14700);
nand U15478 (N_15478,N_14707,N_14617);
nand U15479 (N_15479,N_14901,N_14586);
xor U15480 (N_15480,N_14656,N_14856);
nand U15481 (N_15481,N_14590,N_14955);
or U15482 (N_15482,N_14917,N_14647);
and U15483 (N_15483,N_14600,N_14512);
or U15484 (N_15484,N_14548,N_14508);
nand U15485 (N_15485,N_14737,N_14778);
nand U15486 (N_15486,N_14628,N_14805);
nand U15487 (N_15487,N_14646,N_14696);
xor U15488 (N_15488,N_14773,N_14551);
nor U15489 (N_15489,N_14766,N_14799);
nand U15490 (N_15490,N_14652,N_14826);
and U15491 (N_15491,N_14831,N_14971);
nand U15492 (N_15492,N_14836,N_14713);
or U15493 (N_15493,N_14594,N_14620);
nand U15494 (N_15494,N_14590,N_14880);
and U15495 (N_15495,N_14662,N_14802);
nor U15496 (N_15496,N_14612,N_14598);
nand U15497 (N_15497,N_14736,N_14514);
or U15498 (N_15498,N_14685,N_14571);
nor U15499 (N_15499,N_14507,N_14940);
or U15500 (N_15500,N_15325,N_15196);
nand U15501 (N_15501,N_15225,N_15040);
or U15502 (N_15502,N_15224,N_15339);
and U15503 (N_15503,N_15303,N_15242);
nor U15504 (N_15504,N_15289,N_15266);
nor U15505 (N_15505,N_15489,N_15376);
nor U15506 (N_15506,N_15055,N_15485);
and U15507 (N_15507,N_15497,N_15286);
nor U15508 (N_15508,N_15424,N_15195);
nand U15509 (N_15509,N_15361,N_15282);
nand U15510 (N_15510,N_15301,N_15235);
nor U15511 (N_15511,N_15134,N_15052);
or U15512 (N_15512,N_15063,N_15096);
nor U15513 (N_15513,N_15486,N_15093);
and U15514 (N_15514,N_15437,N_15365);
or U15515 (N_15515,N_15280,N_15244);
and U15516 (N_15516,N_15024,N_15336);
nand U15517 (N_15517,N_15122,N_15086);
nor U15518 (N_15518,N_15165,N_15205);
or U15519 (N_15519,N_15124,N_15239);
xnor U15520 (N_15520,N_15105,N_15413);
and U15521 (N_15521,N_15221,N_15284);
nor U15522 (N_15522,N_15396,N_15227);
nand U15523 (N_15523,N_15322,N_15341);
or U15524 (N_15524,N_15395,N_15329);
nand U15525 (N_15525,N_15050,N_15032);
and U15526 (N_15526,N_15245,N_15030);
or U15527 (N_15527,N_15130,N_15180);
xor U15528 (N_15528,N_15384,N_15042);
xor U15529 (N_15529,N_15360,N_15057);
or U15530 (N_15530,N_15209,N_15213);
nand U15531 (N_15531,N_15185,N_15025);
and U15532 (N_15532,N_15228,N_15248);
or U15533 (N_15533,N_15255,N_15297);
or U15534 (N_15534,N_15327,N_15385);
nand U15535 (N_15535,N_15357,N_15406);
nor U15536 (N_15536,N_15456,N_15265);
or U15537 (N_15537,N_15471,N_15309);
nand U15538 (N_15538,N_15495,N_15436);
nand U15539 (N_15539,N_15342,N_15249);
or U15540 (N_15540,N_15064,N_15117);
or U15541 (N_15541,N_15007,N_15299);
nand U15542 (N_15542,N_15252,N_15317);
or U15543 (N_15543,N_15141,N_15380);
and U15544 (N_15544,N_15474,N_15375);
or U15545 (N_15545,N_15462,N_15412);
nand U15546 (N_15546,N_15171,N_15021);
xnor U15547 (N_15547,N_15022,N_15150);
nand U15548 (N_15548,N_15074,N_15060);
or U15549 (N_15549,N_15381,N_15210);
nor U15550 (N_15550,N_15427,N_15388);
or U15551 (N_15551,N_15447,N_15005);
nand U15552 (N_15552,N_15354,N_15182);
or U15553 (N_15553,N_15291,N_15222);
nor U15554 (N_15554,N_15496,N_15145);
and U15555 (N_15555,N_15401,N_15493);
and U15556 (N_15556,N_15374,N_15149);
or U15557 (N_15557,N_15008,N_15218);
nor U15558 (N_15558,N_15020,N_15109);
and U15559 (N_15559,N_15431,N_15494);
or U15560 (N_15560,N_15318,N_15203);
and U15561 (N_15561,N_15461,N_15107);
nor U15562 (N_15562,N_15217,N_15369);
or U15563 (N_15563,N_15448,N_15283);
and U15564 (N_15564,N_15389,N_15438);
or U15565 (N_15565,N_15464,N_15029);
nor U15566 (N_15566,N_15099,N_15332);
nand U15567 (N_15567,N_15321,N_15194);
nor U15568 (N_15568,N_15451,N_15056);
nor U15569 (N_15569,N_15428,N_15162);
nand U15570 (N_15570,N_15095,N_15103);
nand U15571 (N_15571,N_15405,N_15215);
and U15572 (N_15572,N_15144,N_15373);
nor U15573 (N_15573,N_15425,N_15310);
or U15574 (N_15574,N_15426,N_15142);
and U15575 (N_15575,N_15068,N_15308);
and U15576 (N_15576,N_15295,N_15220);
and U15577 (N_15577,N_15006,N_15268);
and U15578 (N_15578,N_15331,N_15250);
and U15579 (N_15579,N_15017,N_15113);
nor U15580 (N_15580,N_15367,N_15372);
nand U15581 (N_15581,N_15458,N_15212);
nor U15582 (N_15582,N_15070,N_15368);
and U15583 (N_15583,N_15479,N_15123);
or U15584 (N_15584,N_15200,N_15163);
nor U15585 (N_15585,N_15168,N_15264);
or U15586 (N_15586,N_15112,N_15137);
nand U15587 (N_15587,N_15466,N_15053);
and U15588 (N_15588,N_15079,N_15257);
and U15589 (N_15589,N_15358,N_15313);
nor U15590 (N_15590,N_15167,N_15118);
nand U15591 (N_15591,N_15154,N_15298);
nand U15592 (N_15592,N_15128,N_15039);
and U15593 (N_15593,N_15108,N_15326);
or U15594 (N_15594,N_15492,N_15034);
nand U15595 (N_15595,N_15433,N_15261);
nand U15596 (N_15596,N_15197,N_15409);
nand U15597 (N_15597,N_15482,N_15316);
and U15598 (N_15598,N_15363,N_15411);
and U15599 (N_15599,N_15186,N_15347);
nand U15600 (N_15600,N_15232,N_15088);
xor U15601 (N_15601,N_15353,N_15345);
and U15602 (N_15602,N_15417,N_15275);
and U15603 (N_15603,N_15161,N_15340);
xor U15604 (N_15604,N_15419,N_15273);
nor U15605 (N_15605,N_15164,N_15491);
nor U15606 (N_15606,N_15391,N_15083);
or U15607 (N_15607,N_15234,N_15080);
or U15608 (N_15608,N_15430,N_15281);
and U15609 (N_15609,N_15382,N_15364);
or U15610 (N_15610,N_15013,N_15027);
or U15611 (N_15611,N_15238,N_15192);
nand U15612 (N_15612,N_15000,N_15176);
nor U15613 (N_15613,N_15293,N_15175);
nor U15614 (N_15614,N_15460,N_15440);
nor U15615 (N_15615,N_15211,N_15014);
or U15616 (N_15616,N_15119,N_15153);
nand U15617 (N_15617,N_15432,N_15028);
nand U15618 (N_15618,N_15467,N_15259);
nor U15619 (N_15619,N_15151,N_15287);
nor U15620 (N_15620,N_15352,N_15087);
and U15621 (N_15621,N_15454,N_15469);
and U15622 (N_15622,N_15279,N_15306);
and U15623 (N_15623,N_15045,N_15499);
or U15624 (N_15624,N_15035,N_15267);
xor U15625 (N_15625,N_15251,N_15094);
and U15626 (N_15626,N_15136,N_15077);
xor U15627 (N_15627,N_15468,N_15319);
nor U15628 (N_15628,N_15156,N_15429);
or U15629 (N_15629,N_15140,N_15247);
or U15630 (N_15630,N_15243,N_15481);
or U15631 (N_15631,N_15059,N_15246);
or U15632 (N_15632,N_15002,N_15237);
xnor U15633 (N_15633,N_15009,N_15061);
and U15634 (N_15634,N_15018,N_15044);
or U15635 (N_15635,N_15393,N_15110);
nor U15636 (N_15636,N_15387,N_15449);
nand U15637 (N_15637,N_15157,N_15229);
nor U15638 (N_15638,N_15477,N_15473);
or U15639 (N_15639,N_15386,N_15048);
or U15640 (N_15640,N_15072,N_15148);
or U15641 (N_15641,N_15160,N_15120);
and U15642 (N_15642,N_15410,N_15392);
or U15643 (N_15643,N_15397,N_15138);
nand U15644 (N_15644,N_15398,N_15423);
nor U15645 (N_15645,N_15478,N_15133);
and U15646 (N_15646,N_15135,N_15075);
nor U15647 (N_15647,N_15260,N_15101);
nand U15648 (N_15648,N_15498,N_15198);
or U15649 (N_15649,N_15344,N_15125);
nor U15650 (N_15650,N_15285,N_15253);
nor U15651 (N_15651,N_15177,N_15004);
nand U15652 (N_15652,N_15178,N_15484);
nand U15653 (N_15653,N_15199,N_15115);
nor U15654 (N_15654,N_15324,N_15179);
nor U15655 (N_15655,N_15434,N_15031);
xor U15656 (N_15656,N_15294,N_15051);
nand U15657 (N_15657,N_15403,N_15445);
nand U15658 (N_15658,N_15288,N_15443);
nand U15659 (N_15659,N_15292,N_15277);
or U15660 (N_15660,N_15183,N_15240);
and U15661 (N_15661,N_15335,N_15082);
or U15662 (N_15662,N_15187,N_15166);
nand U15663 (N_15663,N_15349,N_15241);
and U15664 (N_15664,N_15129,N_15037);
or U15665 (N_15665,N_15330,N_15097);
or U15666 (N_15666,N_15450,N_15256);
nand U15667 (N_15667,N_15001,N_15269);
or U15668 (N_15668,N_15089,N_15254);
and U15669 (N_15669,N_15147,N_15204);
and U15670 (N_15670,N_15311,N_15091);
nand U15671 (N_15671,N_15062,N_15312);
or U15672 (N_15672,N_15219,N_15366);
and U15673 (N_15673,N_15362,N_15226);
or U15674 (N_15674,N_15414,N_15402);
or U15675 (N_15675,N_15290,N_15069);
and U15676 (N_15676,N_15333,N_15016);
and U15677 (N_15677,N_15370,N_15067);
and U15678 (N_15678,N_15158,N_15026);
and U15679 (N_15679,N_15262,N_15202);
or U15680 (N_15680,N_15003,N_15476);
nand U15681 (N_15681,N_15407,N_15463);
nand U15682 (N_15682,N_15404,N_15033);
nor U15683 (N_15683,N_15049,N_15258);
nand U15684 (N_15684,N_15173,N_15400);
nand U15685 (N_15685,N_15098,N_15296);
or U15686 (N_15686,N_15155,N_15421);
or U15687 (N_15687,N_15488,N_15416);
or U15688 (N_15688,N_15399,N_15208);
and U15689 (N_15689,N_15439,N_15092);
or U15690 (N_15690,N_15216,N_15371);
nor U15691 (N_15691,N_15278,N_15076);
xnor U15692 (N_15692,N_15106,N_15274);
or U15693 (N_15693,N_15146,N_15015);
nor U15694 (N_15694,N_15348,N_15159);
xnor U15695 (N_15695,N_15054,N_15104);
and U15696 (N_15696,N_15090,N_15441);
and U15697 (N_15697,N_15172,N_15444);
nand U15698 (N_15698,N_15011,N_15422);
nand U15699 (N_15699,N_15420,N_15415);
and U15700 (N_15700,N_15487,N_15207);
and U15701 (N_15701,N_15206,N_15270);
or U15702 (N_15702,N_15356,N_15383);
nor U15703 (N_15703,N_15276,N_15272);
or U15704 (N_15704,N_15408,N_15066);
nor U15705 (N_15705,N_15390,N_15453);
and U15706 (N_15706,N_15346,N_15189);
nor U15707 (N_15707,N_15169,N_15305);
nor U15708 (N_15708,N_15435,N_15233);
nand U15709 (N_15709,N_15377,N_15036);
nand U15710 (N_15710,N_15043,N_15442);
or U15711 (N_15711,N_15012,N_15271);
xor U15712 (N_15712,N_15126,N_15320);
nand U15713 (N_15713,N_15046,N_15190);
and U15714 (N_15714,N_15201,N_15010);
and U15715 (N_15715,N_15121,N_15193);
or U15716 (N_15716,N_15457,N_15188);
nand U15717 (N_15717,N_15334,N_15465);
and U15718 (N_15718,N_15302,N_15470);
nand U15719 (N_15719,N_15214,N_15181);
and U15720 (N_15720,N_15023,N_15139);
nor U15721 (N_15721,N_15170,N_15078);
and U15722 (N_15722,N_15081,N_15314);
nor U15723 (N_15723,N_15174,N_15459);
and U15724 (N_15724,N_15058,N_15114);
nand U15725 (N_15725,N_15111,N_15452);
and U15726 (N_15726,N_15315,N_15131);
nor U15727 (N_15727,N_15337,N_15084);
nand U15728 (N_15728,N_15355,N_15127);
nor U15729 (N_15729,N_15071,N_15446);
nor U15730 (N_15730,N_15338,N_15116);
nand U15731 (N_15731,N_15073,N_15231);
or U15732 (N_15732,N_15191,N_15047);
nor U15733 (N_15733,N_15230,N_15307);
xnor U15734 (N_15734,N_15304,N_15455);
nand U15735 (N_15735,N_15378,N_15019);
and U15736 (N_15736,N_15472,N_15418);
nand U15737 (N_15737,N_15263,N_15490);
or U15738 (N_15738,N_15343,N_15132);
or U15739 (N_15739,N_15184,N_15323);
nor U15740 (N_15740,N_15475,N_15100);
nor U15741 (N_15741,N_15480,N_15394);
nor U15742 (N_15742,N_15041,N_15065);
or U15743 (N_15743,N_15379,N_15038);
and U15744 (N_15744,N_15102,N_15236);
nor U15745 (N_15745,N_15350,N_15085);
nand U15746 (N_15746,N_15351,N_15143);
xnor U15747 (N_15747,N_15328,N_15359);
nor U15748 (N_15748,N_15483,N_15152);
xor U15749 (N_15749,N_15223,N_15300);
or U15750 (N_15750,N_15443,N_15477);
nor U15751 (N_15751,N_15099,N_15188);
or U15752 (N_15752,N_15055,N_15157);
or U15753 (N_15753,N_15488,N_15119);
or U15754 (N_15754,N_15038,N_15039);
nand U15755 (N_15755,N_15102,N_15390);
nand U15756 (N_15756,N_15034,N_15380);
nand U15757 (N_15757,N_15416,N_15295);
or U15758 (N_15758,N_15104,N_15488);
nor U15759 (N_15759,N_15008,N_15176);
xor U15760 (N_15760,N_15392,N_15137);
nor U15761 (N_15761,N_15489,N_15488);
nor U15762 (N_15762,N_15356,N_15438);
and U15763 (N_15763,N_15482,N_15069);
xor U15764 (N_15764,N_15268,N_15284);
nor U15765 (N_15765,N_15390,N_15281);
and U15766 (N_15766,N_15480,N_15272);
or U15767 (N_15767,N_15138,N_15336);
or U15768 (N_15768,N_15057,N_15285);
nor U15769 (N_15769,N_15251,N_15246);
nor U15770 (N_15770,N_15302,N_15277);
or U15771 (N_15771,N_15221,N_15176);
nor U15772 (N_15772,N_15122,N_15001);
or U15773 (N_15773,N_15475,N_15354);
nor U15774 (N_15774,N_15224,N_15422);
or U15775 (N_15775,N_15138,N_15202);
nor U15776 (N_15776,N_15255,N_15386);
and U15777 (N_15777,N_15041,N_15333);
nand U15778 (N_15778,N_15248,N_15201);
nor U15779 (N_15779,N_15287,N_15199);
or U15780 (N_15780,N_15379,N_15363);
or U15781 (N_15781,N_15026,N_15001);
nand U15782 (N_15782,N_15360,N_15277);
nor U15783 (N_15783,N_15406,N_15011);
or U15784 (N_15784,N_15085,N_15329);
nand U15785 (N_15785,N_15093,N_15277);
and U15786 (N_15786,N_15201,N_15273);
nor U15787 (N_15787,N_15081,N_15260);
nor U15788 (N_15788,N_15488,N_15040);
or U15789 (N_15789,N_15272,N_15381);
nand U15790 (N_15790,N_15066,N_15290);
nand U15791 (N_15791,N_15007,N_15098);
nand U15792 (N_15792,N_15036,N_15068);
or U15793 (N_15793,N_15483,N_15059);
or U15794 (N_15794,N_15308,N_15217);
nor U15795 (N_15795,N_15250,N_15267);
nor U15796 (N_15796,N_15495,N_15155);
or U15797 (N_15797,N_15429,N_15043);
and U15798 (N_15798,N_15160,N_15155);
nand U15799 (N_15799,N_15177,N_15140);
nand U15800 (N_15800,N_15437,N_15089);
nand U15801 (N_15801,N_15287,N_15031);
or U15802 (N_15802,N_15197,N_15335);
nand U15803 (N_15803,N_15471,N_15406);
or U15804 (N_15804,N_15247,N_15237);
nand U15805 (N_15805,N_15348,N_15397);
nor U15806 (N_15806,N_15096,N_15029);
or U15807 (N_15807,N_15007,N_15442);
or U15808 (N_15808,N_15218,N_15328);
nor U15809 (N_15809,N_15325,N_15482);
nand U15810 (N_15810,N_15073,N_15483);
and U15811 (N_15811,N_15133,N_15119);
nor U15812 (N_15812,N_15279,N_15195);
nor U15813 (N_15813,N_15388,N_15291);
nand U15814 (N_15814,N_15293,N_15259);
nand U15815 (N_15815,N_15254,N_15385);
xnor U15816 (N_15816,N_15461,N_15142);
and U15817 (N_15817,N_15192,N_15106);
nor U15818 (N_15818,N_15263,N_15194);
or U15819 (N_15819,N_15315,N_15312);
nor U15820 (N_15820,N_15034,N_15260);
nor U15821 (N_15821,N_15075,N_15109);
or U15822 (N_15822,N_15209,N_15486);
xor U15823 (N_15823,N_15127,N_15017);
xor U15824 (N_15824,N_15279,N_15331);
and U15825 (N_15825,N_15424,N_15024);
nor U15826 (N_15826,N_15354,N_15323);
or U15827 (N_15827,N_15402,N_15200);
and U15828 (N_15828,N_15279,N_15176);
nand U15829 (N_15829,N_15205,N_15128);
nor U15830 (N_15830,N_15454,N_15239);
nor U15831 (N_15831,N_15463,N_15342);
nand U15832 (N_15832,N_15373,N_15338);
and U15833 (N_15833,N_15171,N_15486);
and U15834 (N_15834,N_15135,N_15129);
nand U15835 (N_15835,N_15058,N_15230);
or U15836 (N_15836,N_15272,N_15043);
or U15837 (N_15837,N_15244,N_15083);
or U15838 (N_15838,N_15328,N_15035);
or U15839 (N_15839,N_15024,N_15052);
and U15840 (N_15840,N_15048,N_15389);
nor U15841 (N_15841,N_15267,N_15060);
and U15842 (N_15842,N_15164,N_15349);
and U15843 (N_15843,N_15092,N_15207);
and U15844 (N_15844,N_15138,N_15038);
or U15845 (N_15845,N_15362,N_15493);
nand U15846 (N_15846,N_15405,N_15446);
nand U15847 (N_15847,N_15409,N_15269);
nor U15848 (N_15848,N_15100,N_15104);
nand U15849 (N_15849,N_15060,N_15070);
nand U15850 (N_15850,N_15221,N_15428);
and U15851 (N_15851,N_15192,N_15182);
and U15852 (N_15852,N_15269,N_15153);
or U15853 (N_15853,N_15309,N_15079);
nand U15854 (N_15854,N_15083,N_15315);
and U15855 (N_15855,N_15040,N_15364);
nand U15856 (N_15856,N_15411,N_15446);
nand U15857 (N_15857,N_15469,N_15257);
nor U15858 (N_15858,N_15254,N_15391);
nor U15859 (N_15859,N_15408,N_15445);
and U15860 (N_15860,N_15219,N_15163);
nor U15861 (N_15861,N_15074,N_15379);
or U15862 (N_15862,N_15388,N_15042);
nand U15863 (N_15863,N_15382,N_15271);
nor U15864 (N_15864,N_15338,N_15265);
or U15865 (N_15865,N_15138,N_15434);
or U15866 (N_15866,N_15107,N_15021);
and U15867 (N_15867,N_15324,N_15418);
or U15868 (N_15868,N_15476,N_15442);
or U15869 (N_15869,N_15315,N_15467);
and U15870 (N_15870,N_15110,N_15247);
or U15871 (N_15871,N_15354,N_15472);
nand U15872 (N_15872,N_15233,N_15134);
nor U15873 (N_15873,N_15294,N_15310);
nor U15874 (N_15874,N_15088,N_15460);
or U15875 (N_15875,N_15003,N_15075);
nor U15876 (N_15876,N_15098,N_15235);
nor U15877 (N_15877,N_15287,N_15392);
or U15878 (N_15878,N_15280,N_15277);
nor U15879 (N_15879,N_15344,N_15161);
nor U15880 (N_15880,N_15438,N_15314);
nor U15881 (N_15881,N_15140,N_15135);
nor U15882 (N_15882,N_15189,N_15104);
and U15883 (N_15883,N_15068,N_15254);
or U15884 (N_15884,N_15206,N_15392);
nand U15885 (N_15885,N_15447,N_15146);
nand U15886 (N_15886,N_15108,N_15194);
or U15887 (N_15887,N_15341,N_15489);
nand U15888 (N_15888,N_15164,N_15051);
and U15889 (N_15889,N_15482,N_15121);
or U15890 (N_15890,N_15350,N_15436);
and U15891 (N_15891,N_15227,N_15306);
xor U15892 (N_15892,N_15185,N_15067);
nand U15893 (N_15893,N_15179,N_15468);
and U15894 (N_15894,N_15016,N_15435);
or U15895 (N_15895,N_15067,N_15218);
or U15896 (N_15896,N_15410,N_15295);
nand U15897 (N_15897,N_15142,N_15045);
nor U15898 (N_15898,N_15355,N_15143);
nand U15899 (N_15899,N_15267,N_15279);
and U15900 (N_15900,N_15392,N_15473);
and U15901 (N_15901,N_15019,N_15039);
and U15902 (N_15902,N_15278,N_15450);
nor U15903 (N_15903,N_15463,N_15162);
nor U15904 (N_15904,N_15188,N_15032);
or U15905 (N_15905,N_15315,N_15225);
nor U15906 (N_15906,N_15140,N_15497);
nor U15907 (N_15907,N_15258,N_15461);
nand U15908 (N_15908,N_15031,N_15243);
and U15909 (N_15909,N_15343,N_15390);
and U15910 (N_15910,N_15445,N_15273);
nor U15911 (N_15911,N_15431,N_15069);
nor U15912 (N_15912,N_15484,N_15226);
nand U15913 (N_15913,N_15378,N_15138);
and U15914 (N_15914,N_15144,N_15278);
xnor U15915 (N_15915,N_15190,N_15007);
or U15916 (N_15916,N_15011,N_15298);
nor U15917 (N_15917,N_15114,N_15226);
nor U15918 (N_15918,N_15396,N_15050);
nor U15919 (N_15919,N_15282,N_15045);
and U15920 (N_15920,N_15151,N_15235);
or U15921 (N_15921,N_15070,N_15133);
nand U15922 (N_15922,N_15285,N_15052);
nor U15923 (N_15923,N_15303,N_15189);
or U15924 (N_15924,N_15093,N_15367);
xnor U15925 (N_15925,N_15230,N_15397);
or U15926 (N_15926,N_15314,N_15006);
or U15927 (N_15927,N_15273,N_15172);
nor U15928 (N_15928,N_15256,N_15027);
nor U15929 (N_15929,N_15265,N_15249);
and U15930 (N_15930,N_15212,N_15174);
nand U15931 (N_15931,N_15151,N_15001);
and U15932 (N_15932,N_15038,N_15287);
nand U15933 (N_15933,N_15047,N_15005);
nand U15934 (N_15934,N_15027,N_15065);
and U15935 (N_15935,N_15179,N_15413);
nand U15936 (N_15936,N_15026,N_15329);
and U15937 (N_15937,N_15170,N_15466);
or U15938 (N_15938,N_15243,N_15156);
or U15939 (N_15939,N_15111,N_15356);
and U15940 (N_15940,N_15492,N_15160);
and U15941 (N_15941,N_15410,N_15441);
and U15942 (N_15942,N_15185,N_15150);
and U15943 (N_15943,N_15006,N_15443);
or U15944 (N_15944,N_15462,N_15349);
nor U15945 (N_15945,N_15189,N_15047);
and U15946 (N_15946,N_15379,N_15419);
or U15947 (N_15947,N_15380,N_15453);
nand U15948 (N_15948,N_15103,N_15029);
nor U15949 (N_15949,N_15101,N_15195);
nor U15950 (N_15950,N_15262,N_15494);
nand U15951 (N_15951,N_15439,N_15367);
nor U15952 (N_15952,N_15447,N_15370);
and U15953 (N_15953,N_15262,N_15191);
nand U15954 (N_15954,N_15406,N_15161);
or U15955 (N_15955,N_15119,N_15408);
nor U15956 (N_15956,N_15207,N_15056);
xor U15957 (N_15957,N_15147,N_15282);
nand U15958 (N_15958,N_15152,N_15352);
or U15959 (N_15959,N_15282,N_15378);
or U15960 (N_15960,N_15360,N_15073);
and U15961 (N_15961,N_15184,N_15472);
or U15962 (N_15962,N_15124,N_15182);
nand U15963 (N_15963,N_15294,N_15129);
nor U15964 (N_15964,N_15179,N_15325);
or U15965 (N_15965,N_15363,N_15184);
and U15966 (N_15966,N_15154,N_15146);
nand U15967 (N_15967,N_15153,N_15046);
nor U15968 (N_15968,N_15236,N_15169);
nor U15969 (N_15969,N_15066,N_15412);
and U15970 (N_15970,N_15053,N_15094);
and U15971 (N_15971,N_15112,N_15432);
or U15972 (N_15972,N_15436,N_15287);
xnor U15973 (N_15973,N_15180,N_15079);
or U15974 (N_15974,N_15004,N_15262);
or U15975 (N_15975,N_15251,N_15041);
xnor U15976 (N_15976,N_15135,N_15195);
xnor U15977 (N_15977,N_15051,N_15486);
or U15978 (N_15978,N_15283,N_15241);
xnor U15979 (N_15979,N_15293,N_15273);
nor U15980 (N_15980,N_15067,N_15271);
or U15981 (N_15981,N_15095,N_15255);
and U15982 (N_15982,N_15135,N_15413);
nor U15983 (N_15983,N_15254,N_15173);
and U15984 (N_15984,N_15010,N_15405);
nor U15985 (N_15985,N_15130,N_15404);
nor U15986 (N_15986,N_15063,N_15159);
nor U15987 (N_15987,N_15477,N_15368);
and U15988 (N_15988,N_15095,N_15000);
and U15989 (N_15989,N_15448,N_15161);
nor U15990 (N_15990,N_15328,N_15471);
nand U15991 (N_15991,N_15186,N_15497);
nor U15992 (N_15992,N_15126,N_15325);
nor U15993 (N_15993,N_15335,N_15443);
or U15994 (N_15994,N_15104,N_15252);
nor U15995 (N_15995,N_15112,N_15239);
or U15996 (N_15996,N_15160,N_15178);
nand U15997 (N_15997,N_15398,N_15408);
or U15998 (N_15998,N_15087,N_15467);
nor U15999 (N_15999,N_15151,N_15297);
and U16000 (N_16000,N_15629,N_15958);
nand U16001 (N_16001,N_15835,N_15661);
and U16002 (N_16002,N_15969,N_15543);
nor U16003 (N_16003,N_15867,N_15587);
or U16004 (N_16004,N_15895,N_15648);
or U16005 (N_16005,N_15740,N_15711);
and U16006 (N_16006,N_15727,N_15715);
and U16007 (N_16007,N_15870,N_15521);
nand U16008 (N_16008,N_15858,N_15618);
or U16009 (N_16009,N_15600,N_15731);
or U16010 (N_16010,N_15941,N_15555);
nand U16011 (N_16011,N_15844,N_15642);
or U16012 (N_16012,N_15755,N_15896);
or U16013 (N_16013,N_15964,N_15585);
nand U16014 (N_16014,N_15726,N_15691);
nand U16015 (N_16015,N_15548,N_15967);
nand U16016 (N_16016,N_15553,N_15977);
nor U16017 (N_16017,N_15512,N_15809);
nor U16018 (N_16018,N_15817,N_15529);
and U16019 (N_16019,N_15938,N_15743);
nand U16020 (N_16020,N_15811,N_15614);
nor U16021 (N_16021,N_15792,N_15537);
or U16022 (N_16022,N_15762,N_15576);
or U16023 (N_16023,N_15959,N_15586);
nor U16024 (N_16024,N_15992,N_15852);
nand U16025 (N_16025,N_15664,N_15903);
and U16026 (N_16026,N_15683,N_15594);
and U16027 (N_16027,N_15693,N_15517);
nor U16028 (N_16028,N_15504,N_15502);
and U16029 (N_16029,N_15939,N_15577);
and U16030 (N_16030,N_15682,N_15772);
nand U16031 (N_16031,N_15847,N_15957);
nand U16032 (N_16032,N_15805,N_15886);
nor U16033 (N_16033,N_15595,N_15632);
or U16034 (N_16034,N_15652,N_15936);
nand U16035 (N_16035,N_15606,N_15803);
and U16036 (N_16036,N_15589,N_15701);
or U16037 (N_16037,N_15604,N_15819);
nor U16038 (N_16038,N_15651,N_15611);
nor U16039 (N_16039,N_15593,N_15556);
and U16040 (N_16040,N_15946,N_15793);
nand U16041 (N_16041,N_15873,N_15884);
and U16042 (N_16042,N_15729,N_15524);
nor U16043 (N_16043,N_15826,N_15754);
or U16044 (N_16044,N_15963,N_15893);
and U16045 (N_16045,N_15944,N_15808);
or U16046 (N_16046,N_15782,N_15891);
nand U16047 (N_16047,N_15931,N_15721);
and U16048 (N_16048,N_15995,N_15676);
nand U16049 (N_16049,N_15568,N_15528);
nor U16050 (N_16050,N_15500,N_15771);
and U16051 (N_16051,N_15636,N_15850);
or U16052 (N_16052,N_15766,N_15872);
and U16053 (N_16053,N_15597,N_15518);
nor U16054 (N_16054,N_15877,N_15552);
nor U16055 (N_16055,N_15843,N_15745);
or U16056 (N_16056,N_15566,N_15523);
nand U16057 (N_16057,N_15695,N_15789);
and U16058 (N_16058,N_15708,N_15562);
nor U16059 (N_16059,N_15821,N_15666);
and U16060 (N_16060,N_15706,N_15685);
or U16061 (N_16061,N_15741,N_15725);
or U16062 (N_16062,N_15712,N_15719);
nand U16063 (N_16063,N_15993,N_15833);
and U16064 (N_16064,N_15732,N_15972);
or U16065 (N_16065,N_15783,N_15971);
nand U16066 (N_16066,N_15637,N_15979);
nor U16067 (N_16067,N_15617,N_15526);
xor U16068 (N_16068,N_15961,N_15910);
nor U16069 (N_16069,N_15840,N_15862);
nor U16070 (N_16070,N_15716,N_15613);
nor U16071 (N_16071,N_15780,N_15897);
or U16072 (N_16072,N_15538,N_15807);
nor U16073 (N_16073,N_15994,N_15530);
nor U16074 (N_16074,N_15759,N_15610);
nor U16075 (N_16075,N_15943,N_15573);
nand U16076 (N_16076,N_15883,N_15677);
or U16077 (N_16077,N_15687,N_15778);
and U16078 (N_16078,N_15767,N_15527);
and U16079 (N_16079,N_15810,N_15746);
or U16080 (N_16080,N_15544,N_15848);
and U16081 (N_16081,N_15916,N_15922);
nand U16082 (N_16082,N_15774,N_15569);
nand U16083 (N_16083,N_15752,N_15668);
and U16084 (N_16084,N_15698,N_15907);
and U16085 (N_16085,N_15813,N_15531);
nand U16086 (N_16086,N_15503,N_15737);
nand U16087 (N_16087,N_15832,N_15854);
nor U16088 (N_16088,N_15855,N_15702);
and U16089 (N_16089,N_15650,N_15738);
and U16090 (N_16090,N_15918,N_15709);
or U16091 (N_16091,N_15519,N_15894);
nand U16092 (N_16092,N_15620,N_15881);
nand U16093 (N_16093,N_15559,N_15564);
nor U16094 (N_16094,N_15744,N_15608);
nor U16095 (N_16095,N_15710,N_15558);
and U16096 (N_16096,N_15796,N_15928);
nand U16097 (N_16097,N_15799,N_15734);
nor U16098 (N_16098,N_15624,N_15934);
nor U16099 (N_16099,N_15542,N_15549);
or U16100 (N_16100,N_15889,N_15692);
nor U16101 (N_16101,N_15615,N_15787);
and U16102 (N_16102,N_15601,N_15700);
nand U16103 (N_16103,N_15545,N_15742);
or U16104 (N_16104,N_15863,N_15827);
and U16105 (N_16105,N_15968,N_15839);
or U16106 (N_16106,N_15937,N_15776);
nor U16107 (N_16107,N_15975,N_15717);
or U16108 (N_16108,N_15550,N_15980);
nor U16109 (N_16109,N_15565,N_15983);
and U16110 (N_16110,N_15921,N_15535);
and U16111 (N_16111,N_15663,N_15658);
nor U16112 (N_16112,N_15665,N_15997);
and U16113 (N_16113,N_15641,N_15800);
or U16114 (N_16114,N_15536,N_15984);
nand U16115 (N_16115,N_15869,N_15806);
or U16116 (N_16116,N_15962,N_15768);
or U16117 (N_16117,N_15675,N_15546);
and U16118 (N_16118,N_15859,N_15728);
nor U16119 (N_16119,N_15525,N_15798);
nand U16120 (N_16120,N_15976,N_15582);
or U16121 (N_16121,N_15824,N_15973);
nand U16122 (N_16122,N_15563,N_15747);
and U16123 (N_16123,N_15511,N_15765);
nor U16124 (N_16124,N_15953,N_15689);
nand U16125 (N_16125,N_15670,N_15705);
or U16126 (N_16126,N_15667,N_15534);
nand U16127 (N_16127,N_15707,N_15876);
and U16128 (N_16128,N_15913,N_15630);
or U16129 (N_16129,N_15690,N_15764);
and U16130 (N_16130,N_15951,N_15812);
nor U16131 (N_16131,N_15818,N_15911);
nor U16132 (N_16132,N_15671,N_15802);
or U16133 (N_16133,N_15501,N_15533);
or U16134 (N_16134,N_15507,N_15539);
and U16135 (N_16135,N_15591,N_15924);
and U16136 (N_16136,N_15834,N_15860);
nor U16137 (N_16137,N_15914,N_15655);
nor U16138 (N_16138,N_15887,N_15786);
nor U16139 (N_16139,N_15837,N_15758);
nor U16140 (N_16140,N_15982,N_15804);
and U16141 (N_16141,N_15784,N_15570);
or U16142 (N_16142,N_15761,N_15952);
nand U16143 (N_16143,N_15919,N_15628);
and U16144 (N_16144,N_15956,N_15763);
and U16145 (N_16145,N_15830,N_15880);
or U16146 (N_16146,N_15927,N_15541);
nand U16147 (N_16147,N_15888,N_15815);
nand U16148 (N_16148,N_15505,N_15781);
or U16149 (N_16149,N_15684,N_15627);
or U16150 (N_16150,N_15584,N_15688);
nor U16151 (N_16151,N_15836,N_15633);
nor U16152 (N_16152,N_15875,N_15602);
nor U16153 (N_16153,N_15510,N_15756);
nand U16154 (N_16154,N_15753,N_15902);
or U16155 (N_16155,N_15865,N_15704);
or U16156 (N_16156,N_15609,N_15596);
or U16157 (N_16157,N_15659,N_15920);
xnor U16158 (N_16158,N_15828,N_15788);
xor U16159 (N_16159,N_15857,N_15933);
nor U16160 (N_16160,N_15795,N_15669);
nor U16161 (N_16161,N_15878,N_15578);
or U16162 (N_16162,N_15508,N_15657);
and U16163 (N_16163,N_15739,N_15987);
nand U16164 (N_16164,N_15966,N_15592);
or U16165 (N_16165,N_15736,N_15714);
nor U16166 (N_16166,N_15686,N_15643);
nand U16167 (N_16167,N_15634,N_15890);
nand U16168 (N_16168,N_15965,N_15769);
nor U16169 (N_16169,N_15681,N_15791);
and U16170 (N_16170,N_15703,N_15879);
and U16171 (N_16171,N_15723,N_15645);
and U16172 (N_16172,N_15574,N_15926);
nor U16173 (N_16173,N_15599,N_15978);
nor U16174 (N_16174,N_15674,N_15751);
nor U16175 (N_16175,N_15750,N_15583);
nor U16176 (N_16176,N_15845,N_15989);
and U16177 (N_16177,N_15955,N_15842);
or U16178 (N_16178,N_15654,N_15849);
or U16179 (N_16179,N_15861,N_15697);
nor U16180 (N_16180,N_15724,N_15930);
and U16181 (N_16181,N_15998,N_15942);
or U16182 (N_16182,N_15797,N_15540);
nor U16183 (N_16183,N_15901,N_15825);
or U16184 (N_16184,N_15612,N_15838);
or U16185 (N_16185,N_15514,N_15988);
nor U16186 (N_16186,N_15581,N_15794);
or U16187 (N_16187,N_15874,N_15991);
nand U16188 (N_16188,N_15892,N_15621);
nand U16189 (N_16189,N_15622,N_15678);
or U16190 (N_16190,N_15770,N_15831);
xor U16191 (N_16191,N_15954,N_15713);
nand U16192 (N_16192,N_15720,N_15516);
xor U16193 (N_16193,N_15580,N_15760);
and U16194 (N_16194,N_15900,N_15853);
or U16195 (N_16195,N_15801,N_15699);
or U16196 (N_16196,N_15572,N_15730);
nor U16197 (N_16197,N_15898,N_15579);
nor U16198 (N_16198,N_15822,N_15912);
nand U16199 (N_16199,N_15814,N_15626);
and U16200 (N_16200,N_15649,N_15945);
nand U16201 (N_16201,N_15588,N_15868);
and U16202 (N_16202,N_15974,N_15619);
and U16203 (N_16203,N_15935,N_15950);
nor U16204 (N_16204,N_15616,N_15605);
and U16205 (N_16205,N_15785,N_15673);
or U16206 (N_16206,N_15639,N_15749);
nor U16207 (N_16207,N_15718,N_15680);
or U16208 (N_16208,N_15773,N_15899);
and U16209 (N_16209,N_15990,N_15885);
and U16210 (N_16210,N_15679,N_15777);
and U16211 (N_16211,N_15672,N_15635);
and U16212 (N_16212,N_15513,N_15623);
and U16213 (N_16213,N_15647,N_15947);
nor U16214 (N_16214,N_15551,N_15905);
nor U16215 (N_16215,N_15925,N_15640);
nor U16216 (N_16216,N_15557,N_15607);
nor U16217 (N_16217,N_15561,N_15917);
and U16218 (N_16218,N_15970,N_15923);
nor U16219 (N_16219,N_15638,N_15625);
nand U16220 (N_16220,N_15735,N_15871);
or U16221 (N_16221,N_15757,N_15866);
or U16222 (N_16222,N_15948,N_15554);
xor U16223 (N_16223,N_15915,N_15520);
and U16224 (N_16224,N_15999,N_15851);
nand U16225 (N_16225,N_15694,N_15509);
nand U16226 (N_16226,N_15940,N_15748);
nand U16227 (N_16227,N_15909,N_15660);
nor U16228 (N_16228,N_15571,N_15653);
and U16229 (N_16229,N_15908,N_15515);
nor U16230 (N_16230,N_15906,N_15986);
and U16231 (N_16231,N_15996,N_15864);
or U16232 (N_16232,N_15775,N_15506);
and U16233 (N_16233,N_15547,N_15696);
or U16234 (N_16234,N_15904,N_15662);
nor U16235 (N_16235,N_15598,N_15816);
and U16236 (N_16236,N_15656,N_15646);
or U16237 (N_16237,N_15929,N_15829);
nand U16238 (N_16238,N_15981,N_15560);
nor U16239 (N_16239,N_15841,N_15603);
or U16240 (N_16240,N_15823,N_15856);
nor U16241 (N_16241,N_15722,N_15779);
nand U16242 (N_16242,N_15846,N_15631);
nand U16243 (N_16243,N_15733,N_15949);
nand U16244 (N_16244,N_15882,N_15567);
or U16245 (N_16245,N_15575,N_15932);
or U16246 (N_16246,N_15590,N_15790);
nor U16247 (N_16247,N_15644,N_15522);
or U16248 (N_16248,N_15532,N_15820);
and U16249 (N_16249,N_15960,N_15985);
nand U16250 (N_16250,N_15812,N_15613);
and U16251 (N_16251,N_15794,N_15924);
nand U16252 (N_16252,N_15694,N_15608);
nand U16253 (N_16253,N_15832,N_15684);
or U16254 (N_16254,N_15725,N_15686);
nand U16255 (N_16255,N_15790,N_15523);
nand U16256 (N_16256,N_15983,N_15558);
and U16257 (N_16257,N_15826,N_15856);
nand U16258 (N_16258,N_15756,N_15571);
nand U16259 (N_16259,N_15614,N_15793);
nand U16260 (N_16260,N_15508,N_15975);
or U16261 (N_16261,N_15754,N_15555);
and U16262 (N_16262,N_15633,N_15881);
or U16263 (N_16263,N_15810,N_15745);
nand U16264 (N_16264,N_15958,N_15650);
and U16265 (N_16265,N_15600,N_15872);
nand U16266 (N_16266,N_15815,N_15639);
and U16267 (N_16267,N_15707,N_15700);
and U16268 (N_16268,N_15885,N_15868);
and U16269 (N_16269,N_15580,N_15866);
and U16270 (N_16270,N_15541,N_15956);
nor U16271 (N_16271,N_15514,N_15607);
and U16272 (N_16272,N_15720,N_15716);
and U16273 (N_16273,N_15857,N_15998);
nor U16274 (N_16274,N_15674,N_15627);
nor U16275 (N_16275,N_15513,N_15822);
nand U16276 (N_16276,N_15943,N_15909);
nand U16277 (N_16277,N_15624,N_15659);
and U16278 (N_16278,N_15822,N_15764);
and U16279 (N_16279,N_15745,N_15708);
nand U16280 (N_16280,N_15866,N_15958);
nor U16281 (N_16281,N_15618,N_15513);
and U16282 (N_16282,N_15549,N_15512);
or U16283 (N_16283,N_15719,N_15961);
and U16284 (N_16284,N_15644,N_15637);
nor U16285 (N_16285,N_15820,N_15535);
nand U16286 (N_16286,N_15664,N_15531);
and U16287 (N_16287,N_15866,N_15761);
nand U16288 (N_16288,N_15806,N_15858);
nand U16289 (N_16289,N_15916,N_15529);
or U16290 (N_16290,N_15514,N_15587);
and U16291 (N_16291,N_15878,N_15931);
nand U16292 (N_16292,N_15551,N_15903);
and U16293 (N_16293,N_15650,N_15821);
and U16294 (N_16294,N_15535,N_15828);
and U16295 (N_16295,N_15574,N_15807);
nand U16296 (N_16296,N_15818,N_15976);
nand U16297 (N_16297,N_15938,N_15608);
nand U16298 (N_16298,N_15740,N_15934);
and U16299 (N_16299,N_15525,N_15758);
nor U16300 (N_16300,N_15907,N_15943);
or U16301 (N_16301,N_15960,N_15949);
nand U16302 (N_16302,N_15918,N_15533);
nand U16303 (N_16303,N_15793,N_15780);
and U16304 (N_16304,N_15839,N_15501);
nor U16305 (N_16305,N_15541,N_15513);
nor U16306 (N_16306,N_15926,N_15786);
nor U16307 (N_16307,N_15514,N_15538);
nor U16308 (N_16308,N_15675,N_15572);
nand U16309 (N_16309,N_15550,N_15973);
nor U16310 (N_16310,N_15962,N_15594);
nor U16311 (N_16311,N_15707,N_15621);
or U16312 (N_16312,N_15834,N_15952);
nor U16313 (N_16313,N_15769,N_15887);
nor U16314 (N_16314,N_15659,N_15906);
or U16315 (N_16315,N_15664,N_15919);
nand U16316 (N_16316,N_15786,N_15844);
nor U16317 (N_16317,N_15992,N_15563);
nor U16318 (N_16318,N_15918,N_15954);
nor U16319 (N_16319,N_15577,N_15740);
nor U16320 (N_16320,N_15617,N_15597);
and U16321 (N_16321,N_15670,N_15678);
nand U16322 (N_16322,N_15688,N_15966);
or U16323 (N_16323,N_15614,N_15516);
nor U16324 (N_16324,N_15736,N_15552);
nor U16325 (N_16325,N_15883,N_15957);
nand U16326 (N_16326,N_15632,N_15515);
nand U16327 (N_16327,N_15688,N_15589);
nor U16328 (N_16328,N_15601,N_15785);
nand U16329 (N_16329,N_15953,N_15945);
xnor U16330 (N_16330,N_15600,N_15578);
or U16331 (N_16331,N_15945,N_15760);
nand U16332 (N_16332,N_15653,N_15600);
nand U16333 (N_16333,N_15806,N_15542);
nand U16334 (N_16334,N_15586,N_15871);
nand U16335 (N_16335,N_15963,N_15800);
or U16336 (N_16336,N_15934,N_15568);
nand U16337 (N_16337,N_15866,N_15649);
nand U16338 (N_16338,N_15913,N_15785);
nor U16339 (N_16339,N_15793,N_15887);
nand U16340 (N_16340,N_15981,N_15948);
nand U16341 (N_16341,N_15818,N_15752);
nand U16342 (N_16342,N_15917,N_15914);
nand U16343 (N_16343,N_15707,N_15906);
nor U16344 (N_16344,N_15767,N_15966);
or U16345 (N_16345,N_15761,N_15907);
and U16346 (N_16346,N_15638,N_15788);
and U16347 (N_16347,N_15685,N_15862);
nor U16348 (N_16348,N_15554,N_15785);
xnor U16349 (N_16349,N_15763,N_15645);
nor U16350 (N_16350,N_15547,N_15652);
and U16351 (N_16351,N_15710,N_15577);
and U16352 (N_16352,N_15750,N_15792);
or U16353 (N_16353,N_15546,N_15505);
or U16354 (N_16354,N_15715,N_15585);
nor U16355 (N_16355,N_15698,N_15533);
and U16356 (N_16356,N_15563,N_15554);
nand U16357 (N_16357,N_15530,N_15815);
nor U16358 (N_16358,N_15922,N_15584);
and U16359 (N_16359,N_15602,N_15616);
nand U16360 (N_16360,N_15903,N_15510);
or U16361 (N_16361,N_15753,N_15707);
and U16362 (N_16362,N_15565,N_15523);
and U16363 (N_16363,N_15853,N_15885);
or U16364 (N_16364,N_15576,N_15892);
nand U16365 (N_16365,N_15926,N_15869);
or U16366 (N_16366,N_15579,N_15619);
or U16367 (N_16367,N_15742,N_15526);
nor U16368 (N_16368,N_15800,N_15732);
nor U16369 (N_16369,N_15669,N_15733);
nor U16370 (N_16370,N_15861,N_15827);
nand U16371 (N_16371,N_15512,N_15831);
or U16372 (N_16372,N_15722,N_15861);
nand U16373 (N_16373,N_15744,N_15569);
nand U16374 (N_16374,N_15615,N_15541);
nand U16375 (N_16375,N_15791,N_15637);
nand U16376 (N_16376,N_15730,N_15964);
and U16377 (N_16377,N_15532,N_15841);
or U16378 (N_16378,N_15706,N_15979);
nor U16379 (N_16379,N_15565,N_15622);
or U16380 (N_16380,N_15807,N_15520);
nand U16381 (N_16381,N_15701,N_15544);
nor U16382 (N_16382,N_15614,N_15692);
nor U16383 (N_16383,N_15791,N_15707);
nor U16384 (N_16384,N_15956,N_15979);
or U16385 (N_16385,N_15963,N_15563);
nand U16386 (N_16386,N_15743,N_15526);
or U16387 (N_16387,N_15848,N_15665);
and U16388 (N_16388,N_15672,N_15666);
nor U16389 (N_16389,N_15700,N_15631);
nand U16390 (N_16390,N_15771,N_15887);
or U16391 (N_16391,N_15665,N_15516);
nor U16392 (N_16392,N_15616,N_15927);
and U16393 (N_16393,N_15565,N_15925);
nand U16394 (N_16394,N_15567,N_15607);
nor U16395 (N_16395,N_15526,N_15875);
nand U16396 (N_16396,N_15620,N_15637);
and U16397 (N_16397,N_15991,N_15508);
and U16398 (N_16398,N_15812,N_15528);
nand U16399 (N_16399,N_15865,N_15929);
nand U16400 (N_16400,N_15852,N_15778);
or U16401 (N_16401,N_15765,N_15615);
nor U16402 (N_16402,N_15502,N_15514);
and U16403 (N_16403,N_15781,N_15885);
nand U16404 (N_16404,N_15676,N_15674);
nand U16405 (N_16405,N_15766,N_15811);
nand U16406 (N_16406,N_15583,N_15735);
nor U16407 (N_16407,N_15942,N_15784);
nor U16408 (N_16408,N_15543,N_15836);
or U16409 (N_16409,N_15939,N_15616);
nor U16410 (N_16410,N_15818,N_15567);
or U16411 (N_16411,N_15550,N_15533);
nand U16412 (N_16412,N_15615,N_15888);
nand U16413 (N_16413,N_15657,N_15517);
nand U16414 (N_16414,N_15527,N_15609);
and U16415 (N_16415,N_15855,N_15691);
nor U16416 (N_16416,N_15756,N_15549);
nor U16417 (N_16417,N_15867,N_15756);
nand U16418 (N_16418,N_15976,N_15864);
or U16419 (N_16419,N_15845,N_15549);
and U16420 (N_16420,N_15520,N_15677);
nand U16421 (N_16421,N_15805,N_15766);
nand U16422 (N_16422,N_15536,N_15771);
nor U16423 (N_16423,N_15727,N_15757);
xor U16424 (N_16424,N_15632,N_15743);
or U16425 (N_16425,N_15847,N_15587);
nand U16426 (N_16426,N_15680,N_15782);
nor U16427 (N_16427,N_15838,N_15901);
and U16428 (N_16428,N_15684,N_15797);
and U16429 (N_16429,N_15784,N_15768);
nand U16430 (N_16430,N_15890,N_15757);
or U16431 (N_16431,N_15591,N_15792);
and U16432 (N_16432,N_15642,N_15684);
nand U16433 (N_16433,N_15711,N_15863);
nor U16434 (N_16434,N_15850,N_15852);
or U16435 (N_16435,N_15808,N_15855);
or U16436 (N_16436,N_15947,N_15769);
and U16437 (N_16437,N_15588,N_15698);
or U16438 (N_16438,N_15748,N_15513);
nor U16439 (N_16439,N_15922,N_15585);
nor U16440 (N_16440,N_15857,N_15656);
and U16441 (N_16441,N_15797,N_15822);
and U16442 (N_16442,N_15727,N_15558);
nor U16443 (N_16443,N_15663,N_15776);
nor U16444 (N_16444,N_15532,N_15770);
nor U16445 (N_16445,N_15676,N_15619);
nand U16446 (N_16446,N_15599,N_15554);
and U16447 (N_16447,N_15587,N_15575);
or U16448 (N_16448,N_15890,N_15970);
and U16449 (N_16449,N_15696,N_15701);
or U16450 (N_16450,N_15748,N_15936);
and U16451 (N_16451,N_15562,N_15710);
nor U16452 (N_16452,N_15631,N_15841);
xnor U16453 (N_16453,N_15874,N_15832);
or U16454 (N_16454,N_15759,N_15828);
and U16455 (N_16455,N_15690,N_15594);
nor U16456 (N_16456,N_15717,N_15779);
or U16457 (N_16457,N_15623,N_15823);
nor U16458 (N_16458,N_15907,N_15855);
nor U16459 (N_16459,N_15911,N_15532);
nor U16460 (N_16460,N_15827,N_15705);
or U16461 (N_16461,N_15778,N_15653);
and U16462 (N_16462,N_15869,N_15726);
nor U16463 (N_16463,N_15899,N_15942);
nor U16464 (N_16464,N_15921,N_15566);
nand U16465 (N_16465,N_15674,N_15930);
nand U16466 (N_16466,N_15571,N_15910);
and U16467 (N_16467,N_15583,N_15559);
nand U16468 (N_16468,N_15720,N_15732);
and U16469 (N_16469,N_15865,N_15967);
or U16470 (N_16470,N_15663,N_15906);
nor U16471 (N_16471,N_15814,N_15831);
or U16472 (N_16472,N_15930,N_15699);
nor U16473 (N_16473,N_15760,N_15713);
nand U16474 (N_16474,N_15883,N_15635);
nand U16475 (N_16475,N_15814,N_15832);
nor U16476 (N_16476,N_15854,N_15694);
nor U16477 (N_16477,N_15628,N_15897);
nand U16478 (N_16478,N_15888,N_15851);
and U16479 (N_16479,N_15668,N_15674);
and U16480 (N_16480,N_15693,N_15766);
or U16481 (N_16481,N_15714,N_15971);
and U16482 (N_16482,N_15974,N_15631);
nor U16483 (N_16483,N_15913,N_15654);
or U16484 (N_16484,N_15978,N_15982);
or U16485 (N_16485,N_15813,N_15503);
or U16486 (N_16486,N_15519,N_15577);
nand U16487 (N_16487,N_15980,N_15545);
and U16488 (N_16488,N_15630,N_15869);
and U16489 (N_16489,N_15863,N_15550);
nor U16490 (N_16490,N_15713,N_15651);
nor U16491 (N_16491,N_15582,N_15978);
nand U16492 (N_16492,N_15705,N_15871);
and U16493 (N_16493,N_15513,N_15954);
xor U16494 (N_16494,N_15687,N_15732);
and U16495 (N_16495,N_15968,N_15866);
xor U16496 (N_16496,N_15798,N_15687);
nor U16497 (N_16497,N_15803,N_15906);
or U16498 (N_16498,N_15585,N_15541);
nand U16499 (N_16499,N_15917,N_15544);
nor U16500 (N_16500,N_16428,N_16383);
and U16501 (N_16501,N_16238,N_16433);
and U16502 (N_16502,N_16464,N_16386);
or U16503 (N_16503,N_16171,N_16218);
nor U16504 (N_16504,N_16212,N_16313);
or U16505 (N_16505,N_16442,N_16052);
nor U16506 (N_16506,N_16271,N_16364);
nand U16507 (N_16507,N_16497,N_16480);
nor U16508 (N_16508,N_16165,N_16429);
nand U16509 (N_16509,N_16077,N_16153);
nor U16510 (N_16510,N_16270,N_16340);
nor U16511 (N_16511,N_16359,N_16177);
nor U16512 (N_16512,N_16179,N_16185);
or U16513 (N_16513,N_16457,N_16363);
nor U16514 (N_16514,N_16229,N_16056);
nand U16515 (N_16515,N_16059,N_16007);
and U16516 (N_16516,N_16256,N_16242);
nand U16517 (N_16517,N_16411,N_16085);
nand U16518 (N_16518,N_16342,N_16083);
and U16519 (N_16519,N_16087,N_16304);
nand U16520 (N_16520,N_16322,N_16157);
nor U16521 (N_16521,N_16160,N_16444);
and U16522 (N_16522,N_16125,N_16152);
nand U16523 (N_16523,N_16408,N_16425);
and U16524 (N_16524,N_16244,N_16335);
nand U16525 (N_16525,N_16134,N_16004);
nand U16526 (N_16526,N_16044,N_16172);
or U16527 (N_16527,N_16217,N_16448);
nand U16528 (N_16528,N_16431,N_16490);
nand U16529 (N_16529,N_16100,N_16112);
and U16530 (N_16530,N_16113,N_16397);
xnor U16531 (N_16531,N_16226,N_16272);
and U16532 (N_16532,N_16065,N_16277);
or U16533 (N_16533,N_16137,N_16224);
and U16534 (N_16534,N_16144,N_16042);
and U16535 (N_16535,N_16417,N_16024);
xnor U16536 (N_16536,N_16390,N_16158);
nand U16537 (N_16537,N_16231,N_16063);
nand U16538 (N_16538,N_16170,N_16365);
nand U16539 (N_16539,N_16298,N_16026);
and U16540 (N_16540,N_16126,N_16110);
and U16541 (N_16541,N_16409,N_16093);
and U16542 (N_16542,N_16205,N_16067);
and U16543 (N_16543,N_16117,N_16379);
or U16544 (N_16544,N_16141,N_16202);
and U16545 (N_16545,N_16459,N_16263);
or U16546 (N_16546,N_16209,N_16441);
or U16547 (N_16547,N_16233,N_16176);
nor U16548 (N_16548,N_16255,N_16316);
or U16549 (N_16549,N_16039,N_16465);
and U16550 (N_16550,N_16296,N_16210);
nand U16551 (N_16551,N_16345,N_16275);
nand U16552 (N_16552,N_16415,N_16033);
and U16553 (N_16553,N_16062,N_16373);
and U16554 (N_16554,N_16037,N_16199);
nand U16555 (N_16555,N_16147,N_16114);
or U16556 (N_16556,N_16047,N_16173);
nand U16557 (N_16557,N_16181,N_16162);
and U16558 (N_16558,N_16201,N_16483);
or U16559 (N_16559,N_16090,N_16370);
nor U16560 (N_16560,N_16399,N_16168);
or U16561 (N_16561,N_16161,N_16167);
and U16562 (N_16562,N_16462,N_16387);
and U16563 (N_16563,N_16422,N_16427);
nor U16564 (N_16564,N_16315,N_16355);
nor U16565 (N_16565,N_16143,N_16198);
nor U16566 (N_16566,N_16469,N_16104);
and U16567 (N_16567,N_16394,N_16048);
and U16568 (N_16568,N_16347,N_16252);
and U16569 (N_16569,N_16010,N_16333);
and U16570 (N_16570,N_16352,N_16071);
or U16571 (N_16571,N_16265,N_16262);
nand U16572 (N_16572,N_16487,N_16456);
nor U16573 (N_16573,N_16301,N_16377);
xnor U16574 (N_16574,N_16380,N_16159);
or U16575 (N_16575,N_16107,N_16474);
nand U16576 (N_16576,N_16261,N_16232);
or U16577 (N_16577,N_16346,N_16412);
nand U16578 (N_16578,N_16268,N_16097);
or U16579 (N_16579,N_16020,N_16248);
and U16580 (N_16580,N_16368,N_16068);
nand U16581 (N_16581,N_16495,N_16401);
nand U16582 (N_16582,N_16361,N_16180);
nand U16583 (N_16583,N_16016,N_16019);
nor U16584 (N_16584,N_16021,N_16192);
nor U16585 (N_16585,N_16310,N_16151);
nor U16586 (N_16586,N_16269,N_16317);
nor U16587 (N_16587,N_16496,N_16050);
and U16588 (N_16588,N_16372,N_16384);
nand U16589 (N_16589,N_16430,N_16498);
nor U16590 (N_16590,N_16030,N_16109);
nand U16591 (N_16591,N_16282,N_16400);
nor U16592 (N_16592,N_16145,N_16150);
and U16593 (N_16593,N_16253,N_16435);
nand U16594 (N_16594,N_16403,N_16139);
and U16595 (N_16595,N_16002,N_16289);
nor U16596 (N_16596,N_16036,N_16075);
nand U16597 (N_16597,N_16041,N_16453);
nor U16598 (N_16598,N_16178,N_16029);
nor U16599 (N_16599,N_16091,N_16321);
nand U16600 (N_16600,N_16341,N_16294);
and U16601 (N_16601,N_16481,N_16475);
nand U16602 (N_16602,N_16102,N_16095);
and U16603 (N_16603,N_16455,N_16472);
or U16604 (N_16604,N_16008,N_16283);
nand U16605 (N_16605,N_16308,N_16274);
nor U16606 (N_16606,N_16076,N_16385);
nor U16607 (N_16607,N_16482,N_16392);
and U16608 (N_16608,N_16299,N_16461);
nor U16609 (N_16609,N_16329,N_16437);
nand U16610 (N_16610,N_16418,N_16108);
nor U16611 (N_16611,N_16343,N_16471);
nand U16612 (N_16612,N_16225,N_16051);
and U16613 (N_16613,N_16318,N_16058);
xor U16614 (N_16614,N_16351,N_16327);
nor U16615 (N_16615,N_16066,N_16358);
or U16616 (N_16616,N_16494,N_16436);
or U16617 (N_16617,N_16410,N_16486);
and U16618 (N_16618,N_16404,N_16079);
and U16619 (N_16619,N_16196,N_16072);
and U16620 (N_16620,N_16460,N_16458);
or U16621 (N_16621,N_16046,N_16200);
nor U16622 (N_16622,N_16064,N_16362);
nor U16623 (N_16623,N_16367,N_16115);
nand U16624 (N_16624,N_16419,N_16499);
nor U16625 (N_16625,N_16396,N_16307);
and U16626 (N_16626,N_16366,N_16260);
or U16627 (N_16627,N_16088,N_16006);
or U16628 (N_16628,N_16291,N_16309);
or U16629 (N_16629,N_16395,N_16003);
and U16630 (N_16630,N_16440,N_16191);
and U16631 (N_16631,N_16290,N_16023);
and U16632 (N_16632,N_16257,N_16353);
and U16633 (N_16633,N_16193,N_16204);
and U16634 (N_16634,N_16339,N_16197);
nor U16635 (N_16635,N_16479,N_16045);
or U16636 (N_16636,N_16325,N_16406);
or U16637 (N_16637,N_16413,N_16454);
xnor U16638 (N_16638,N_16426,N_16297);
nand U16639 (N_16639,N_16300,N_16214);
nand U16640 (N_16640,N_16203,N_16451);
and U16641 (N_16641,N_16124,N_16184);
xor U16642 (N_16642,N_16398,N_16287);
and U16643 (N_16643,N_16120,N_16069);
nor U16644 (N_16644,N_16240,N_16488);
nor U16645 (N_16645,N_16211,N_16468);
or U16646 (N_16646,N_16149,N_16049);
nor U16647 (N_16647,N_16086,N_16070);
and U16648 (N_16648,N_16215,N_16247);
nand U16649 (N_16649,N_16190,N_16078);
nand U16650 (N_16650,N_16273,N_16133);
nand U16651 (N_16651,N_16101,N_16138);
nand U16652 (N_16652,N_16103,N_16323);
or U16653 (N_16653,N_16130,N_16374);
nand U16654 (N_16654,N_16350,N_16434);
nor U16655 (N_16655,N_16131,N_16241);
and U16656 (N_16656,N_16280,N_16420);
nand U16657 (N_16657,N_16140,N_16493);
nor U16658 (N_16658,N_16094,N_16227);
nor U16659 (N_16659,N_16080,N_16009);
nand U16660 (N_16660,N_16013,N_16014);
nor U16661 (N_16661,N_16354,N_16450);
or U16662 (N_16662,N_16254,N_16337);
and U16663 (N_16663,N_16182,N_16393);
nand U16664 (N_16664,N_16098,N_16338);
and U16665 (N_16665,N_16073,N_16348);
and U16666 (N_16666,N_16040,N_16278);
nor U16667 (N_16667,N_16228,N_16328);
nand U16668 (N_16668,N_16326,N_16319);
nand U16669 (N_16669,N_16470,N_16446);
and U16670 (N_16670,N_16332,N_16135);
and U16671 (N_16671,N_16034,N_16236);
nand U16672 (N_16672,N_16074,N_16312);
or U16673 (N_16673,N_16320,N_16249);
nor U16674 (N_16674,N_16473,N_16416);
nor U16675 (N_16675,N_16424,N_16443);
and U16676 (N_16676,N_16142,N_16027);
and U16677 (N_16677,N_16447,N_16292);
nand U16678 (N_16678,N_16356,N_16127);
nor U16679 (N_16679,N_16038,N_16402);
and U16680 (N_16680,N_16357,N_16295);
nand U16681 (N_16681,N_16285,N_16466);
or U16682 (N_16682,N_16432,N_16264);
or U16683 (N_16683,N_16061,N_16208);
or U16684 (N_16684,N_16251,N_16467);
or U16685 (N_16685,N_16035,N_16188);
nand U16686 (N_16686,N_16005,N_16258);
and U16687 (N_16687,N_16243,N_16237);
and U16688 (N_16688,N_16279,N_16166);
and U16689 (N_16689,N_16018,N_16000);
or U16690 (N_16690,N_16476,N_16206);
or U16691 (N_16691,N_16491,N_16223);
or U16692 (N_16692,N_16175,N_16389);
and U16693 (N_16693,N_16414,N_16477);
nor U16694 (N_16694,N_16331,N_16055);
nand U16695 (N_16695,N_16119,N_16043);
nand U16696 (N_16696,N_16025,N_16311);
or U16697 (N_16697,N_16452,N_16111);
nand U16698 (N_16698,N_16266,N_16154);
and U16699 (N_16699,N_16187,N_16084);
nand U16700 (N_16700,N_16017,N_16489);
xor U16701 (N_16701,N_16445,N_16303);
and U16702 (N_16702,N_16123,N_16246);
or U16703 (N_16703,N_16221,N_16360);
or U16704 (N_16704,N_16118,N_16250);
and U16705 (N_16705,N_16314,N_16028);
nand U16706 (N_16706,N_16219,N_16156);
or U16707 (N_16707,N_16281,N_16492);
nand U16708 (N_16708,N_16106,N_16189);
and U16709 (N_16709,N_16349,N_16092);
nand U16710 (N_16710,N_16267,N_16132);
or U16711 (N_16711,N_16060,N_16245);
or U16712 (N_16712,N_16146,N_16421);
and U16713 (N_16713,N_16239,N_16082);
xnor U16714 (N_16714,N_16423,N_16382);
nand U16715 (N_16715,N_16405,N_16121);
or U16716 (N_16716,N_16183,N_16449);
nand U16717 (N_16717,N_16302,N_16288);
or U16718 (N_16718,N_16089,N_16334);
nand U16719 (N_16719,N_16293,N_16330);
nor U16720 (N_16720,N_16286,N_16324);
nand U16721 (N_16721,N_16012,N_16439);
nand U16722 (N_16722,N_16381,N_16186);
or U16723 (N_16723,N_16031,N_16478);
nand U16724 (N_16724,N_16195,N_16015);
nor U16725 (N_16725,N_16463,N_16163);
or U16726 (N_16726,N_16378,N_16053);
and U16727 (N_16727,N_16081,N_16011);
or U16728 (N_16728,N_16174,N_16485);
nor U16729 (N_16729,N_16222,N_16054);
and U16730 (N_16730,N_16369,N_16438);
nand U16731 (N_16731,N_16207,N_16344);
nor U16732 (N_16732,N_16336,N_16057);
or U16733 (N_16733,N_16306,N_16001);
or U16734 (N_16734,N_16128,N_16213);
or U16735 (N_16735,N_16032,N_16375);
or U16736 (N_16736,N_16259,N_16230);
nor U16737 (N_16737,N_16099,N_16096);
and U16738 (N_16738,N_16194,N_16371);
and U16739 (N_16739,N_16105,N_16305);
nor U16740 (N_16740,N_16136,N_16235);
and U16741 (N_16741,N_16234,N_16388);
and U16742 (N_16742,N_16407,N_16116);
nand U16743 (N_16743,N_16164,N_16376);
and U16744 (N_16744,N_16148,N_16216);
and U16745 (N_16745,N_16122,N_16276);
nor U16746 (N_16746,N_16022,N_16220);
nor U16747 (N_16747,N_16155,N_16391);
and U16748 (N_16748,N_16169,N_16484);
nand U16749 (N_16749,N_16284,N_16129);
xor U16750 (N_16750,N_16160,N_16074);
or U16751 (N_16751,N_16407,N_16217);
nand U16752 (N_16752,N_16102,N_16182);
and U16753 (N_16753,N_16131,N_16310);
or U16754 (N_16754,N_16354,N_16223);
nor U16755 (N_16755,N_16367,N_16423);
or U16756 (N_16756,N_16325,N_16293);
nor U16757 (N_16757,N_16300,N_16437);
nand U16758 (N_16758,N_16260,N_16484);
nor U16759 (N_16759,N_16351,N_16365);
or U16760 (N_16760,N_16401,N_16226);
nor U16761 (N_16761,N_16416,N_16162);
nor U16762 (N_16762,N_16026,N_16248);
nand U16763 (N_16763,N_16275,N_16460);
nor U16764 (N_16764,N_16107,N_16359);
or U16765 (N_16765,N_16271,N_16165);
or U16766 (N_16766,N_16239,N_16306);
or U16767 (N_16767,N_16427,N_16047);
nand U16768 (N_16768,N_16474,N_16179);
xor U16769 (N_16769,N_16280,N_16403);
and U16770 (N_16770,N_16169,N_16029);
nand U16771 (N_16771,N_16082,N_16148);
nor U16772 (N_16772,N_16041,N_16378);
and U16773 (N_16773,N_16244,N_16121);
nand U16774 (N_16774,N_16096,N_16404);
xnor U16775 (N_16775,N_16475,N_16347);
or U16776 (N_16776,N_16392,N_16165);
nor U16777 (N_16777,N_16073,N_16448);
and U16778 (N_16778,N_16472,N_16080);
nand U16779 (N_16779,N_16058,N_16314);
and U16780 (N_16780,N_16485,N_16115);
nor U16781 (N_16781,N_16468,N_16396);
or U16782 (N_16782,N_16401,N_16203);
or U16783 (N_16783,N_16215,N_16043);
or U16784 (N_16784,N_16041,N_16165);
nor U16785 (N_16785,N_16055,N_16110);
and U16786 (N_16786,N_16016,N_16407);
or U16787 (N_16787,N_16181,N_16189);
or U16788 (N_16788,N_16085,N_16313);
nor U16789 (N_16789,N_16117,N_16041);
nor U16790 (N_16790,N_16193,N_16404);
nand U16791 (N_16791,N_16453,N_16405);
or U16792 (N_16792,N_16423,N_16343);
or U16793 (N_16793,N_16268,N_16055);
nand U16794 (N_16794,N_16310,N_16279);
nand U16795 (N_16795,N_16146,N_16121);
nor U16796 (N_16796,N_16073,N_16039);
or U16797 (N_16797,N_16312,N_16112);
or U16798 (N_16798,N_16360,N_16170);
nand U16799 (N_16799,N_16468,N_16155);
nand U16800 (N_16800,N_16261,N_16350);
nand U16801 (N_16801,N_16189,N_16316);
nand U16802 (N_16802,N_16045,N_16299);
or U16803 (N_16803,N_16202,N_16443);
nand U16804 (N_16804,N_16314,N_16202);
or U16805 (N_16805,N_16311,N_16493);
nand U16806 (N_16806,N_16214,N_16430);
nand U16807 (N_16807,N_16306,N_16363);
nor U16808 (N_16808,N_16287,N_16233);
or U16809 (N_16809,N_16276,N_16395);
nand U16810 (N_16810,N_16399,N_16277);
nor U16811 (N_16811,N_16118,N_16002);
nor U16812 (N_16812,N_16372,N_16217);
nor U16813 (N_16813,N_16336,N_16022);
and U16814 (N_16814,N_16167,N_16124);
or U16815 (N_16815,N_16149,N_16182);
and U16816 (N_16816,N_16222,N_16462);
nand U16817 (N_16817,N_16483,N_16495);
nor U16818 (N_16818,N_16458,N_16102);
nand U16819 (N_16819,N_16147,N_16143);
and U16820 (N_16820,N_16324,N_16362);
or U16821 (N_16821,N_16164,N_16324);
and U16822 (N_16822,N_16266,N_16228);
nor U16823 (N_16823,N_16018,N_16423);
nand U16824 (N_16824,N_16189,N_16312);
and U16825 (N_16825,N_16388,N_16264);
or U16826 (N_16826,N_16197,N_16160);
and U16827 (N_16827,N_16217,N_16378);
nor U16828 (N_16828,N_16199,N_16473);
or U16829 (N_16829,N_16041,N_16020);
and U16830 (N_16830,N_16253,N_16295);
or U16831 (N_16831,N_16274,N_16014);
and U16832 (N_16832,N_16146,N_16083);
or U16833 (N_16833,N_16389,N_16440);
and U16834 (N_16834,N_16340,N_16199);
nand U16835 (N_16835,N_16270,N_16110);
and U16836 (N_16836,N_16197,N_16403);
or U16837 (N_16837,N_16183,N_16324);
and U16838 (N_16838,N_16153,N_16256);
nand U16839 (N_16839,N_16186,N_16125);
and U16840 (N_16840,N_16363,N_16100);
nand U16841 (N_16841,N_16278,N_16334);
nand U16842 (N_16842,N_16269,N_16081);
nand U16843 (N_16843,N_16434,N_16157);
nand U16844 (N_16844,N_16087,N_16013);
nand U16845 (N_16845,N_16116,N_16107);
xnor U16846 (N_16846,N_16408,N_16294);
or U16847 (N_16847,N_16043,N_16442);
nor U16848 (N_16848,N_16148,N_16429);
nand U16849 (N_16849,N_16194,N_16440);
and U16850 (N_16850,N_16423,N_16069);
or U16851 (N_16851,N_16396,N_16215);
nand U16852 (N_16852,N_16495,N_16327);
nand U16853 (N_16853,N_16355,N_16479);
nor U16854 (N_16854,N_16298,N_16140);
and U16855 (N_16855,N_16099,N_16216);
or U16856 (N_16856,N_16362,N_16204);
nand U16857 (N_16857,N_16410,N_16258);
and U16858 (N_16858,N_16368,N_16456);
and U16859 (N_16859,N_16472,N_16106);
and U16860 (N_16860,N_16437,N_16473);
nand U16861 (N_16861,N_16309,N_16474);
nor U16862 (N_16862,N_16219,N_16083);
and U16863 (N_16863,N_16403,N_16010);
and U16864 (N_16864,N_16108,N_16220);
nand U16865 (N_16865,N_16341,N_16003);
or U16866 (N_16866,N_16478,N_16392);
nand U16867 (N_16867,N_16273,N_16428);
nand U16868 (N_16868,N_16126,N_16021);
or U16869 (N_16869,N_16478,N_16363);
or U16870 (N_16870,N_16361,N_16415);
or U16871 (N_16871,N_16016,N_16493);
nor U16872 (N_16872,N_16414,N_16021);
nor U16873 (N_16873,N_16493,N_16300);
xnor U16874 (N_16874,N_16494,N_16143);
or U16875 (N_16875,N_16073,N_16205);
nand U16876 (N_16876,N_16387,N_16452);
nand U16877 (N_16877,N_16327,N_16461);
and U16878 (N_16878,N_16158,N_16485);
nor U16879 (N_16879,N_16420,N_16232);
nor U16880 (N_16880,N_16316,N_16387);
or U16881 (N_16881,N_16327,N_16396);
nor U16882 (N_16882,N_16177,N_16017);
nor U16883 (N_16883,N_16190,N_16090);
nor U16884 (N_16884,N_16111,N_16481);
nand U16885 (N_16885,N_16188,N_16016);
nor U16886 (N_16886,N_16292,N_16031);
or U16887 (N_16887,N_16420,N_16245);
nand U16888 (N_16888,N_16432,N_16426);
or U16889 (N_16889,N_16150,N_16037);
or U16890 (N_16890,N_16420,N_16175);
and U16891 (N_16891,N_16344,N_16238);
nor U16892 (N_16892,N_16123,N_16185);
or U16893 (N_16893,N_16420,N_16192);
or U16894 (N_16894,N_16140,N_16134);
and U16895 (N_16895,N_16221,N_16442);
or U16896 (N_16896,N_16228,N_16390);
nand U16897 (N_16897,N_16379,N_16255);
or U16898 (N_16898,N_16379,N_16429);
nand U16899 (N_16899,N_16166,N_16136);
nor U16900 (N_16900,N_16485,N_16082);
or U16901 (N_16901,N_16483,N_16278);
and U16902 (N_16902,N_16076,N_16133);
nor U16903 (N_16903,N_16092,N_16305);
or U16904 (N_16904,N_16277,N_16468);
and U16905 (N_16905,N_16353,N_16252);
and U16906 (N_16906,N_16292,N_16430);
or U16907 (N_16907,N_16186,N_16493);
nand U16908 (N_16908,N_16349,N_16176);
and U16909 (N_16909,N_16306,N_16110);
or U16910 (N_16910,N_16299,N_16078);
nand U16911 (N_16911,N_16486,N_16237);
nand U16912 (N_16912,N_16014,N_16404);
and U16913 (N_16913,N_16234,N_16087);
or U16914 (N_16914,N_16412,N_16098);
and U16915 (N_16915,N_16359,N_16439);
nor U16916 (N_16916,N_16462,N_16316);
or U16917 (N_16917,N_16413,N_16335);
and U16918 (N_16918,N_16098,N_16129);
and U16919 (N_16919,N_16002,N_16364);
and U16920 (N_16920,N_16113,N_16420);
and U16921 (N_16921,N_16381,N_16382);
nor U16922 (N_16922,N_16459,N_16420);
or U16923 (N_16923,N_16084,N_16296);
nand U16924 (N_16924,N_16412,N_16393);
nand U16925 (N_16925,N_16195,N_16310);
or U16926 (N_16926,N_16207,N_16131);
or U16927 (N_16927,N_16283,N_16298);
and U16928 (N_16928,N_16368,N_16411);
nand U16929 (N_16929,N_16111,N_16377);
nor U16930 (N_16930,N_16172,N_16336);
nor U16931 (N_16931,N_16161,N_16226);
and U16932 (N_16932,N_16138,N_16477);
nand U16933 (N_16933,N_16355,N_16175);
or U16934 (N_16934,N_16123,N_16091);
nand U16935 (N_16935,N_16333,N_16006);
nand U16936 (N_16936,N_16295,N_16131);
nor U16937 (N_16937,N_16360,N_16050);
nand U16938 (N_16938,N_16227,N_16487);
nor U16939 (N_16939,N_16072,N_16404);
nor U16940 (N_16940,N_16178,N_16309);
and U16941 (N_16941,N_16096,N_16087);
xnor U16942 (N_16942,N_16429,N_16413);
nand U16943 (N_16943,N_16063,N_16290);
and U16944 (N_16944,N_16198,N_16462);
and U16945 (N_16945,N_16440,N_16189);
nor U16946 (N_16946,N_16463,N_16272);
nor U16947 (N_16947,N_16235,N_16317);
or U16948 (N_16948,N_16173,N_16096);
or U16949 (N_16949,N_16069,N_16412);
nand U16950 (N_16950,N_16473,N_16305);
or U16951 (N_16951,N_16474,N_16259);
nand U16952 (N_16952,N_16298,N_16153);
nand U16953 (N_16953,N_16475,N_16484);
nor U16954 (N_16954,N_16459,N_16247);
nand U16955 (N_16955,N_16470,N_16396);
and U16956 (N_16956,N_16465,N_16414);
nor U16957 (N_16957,N_16011,N_16149);
or U16958 (N_16958,N_16268,N_16499);
and U16959 (N_16959,N_16299,N_16032);
and U16960 (N_16960,N_16410,N_16042);
nor U16961 (N_16961,N_16062,N_16405);
nand U16962 (N_16962,N_16010,N_16377);
or U16963 (N_16963,N_16033,N_16304);
nor U16964 (N_16964,N_16245,N_16039);
nand U16965 (N_16965,N_16372,N_16274);
nand U16966 (N_16966,N_16147,N_16044);
and U16967 (N_16967,N_16058,N_16131);
or U16968 (N_16968,N_16421,N_16003);
nor U16969 (N_16969,N_16421,N_16445);
nand U16970 (N_16970,N_16336,N_16391);
or U16971 (N_16971,N_16485,N_16305);
or U16972 (N_16972,N_16195,N_16436);
or U16973 (N_16973,N_16295,N_16182);
nor U16974 (N_16974,N_16204,N_16427);
or U16975 (N_16975,N_16242,N_16275);
and U16976 (N_16976,N_16328,N_16378);
and U16977 (N_16977,N_16480,N_16362);
nor U16978 (N_16978,N_16122,N_16314);
or U16979 (N_16979,N_16308,N_16303);
nand U16980 (N_16980,N_16239,N_16414);
nor U16981 (N_16981,N_16417,N_16498);
nand U16982 (N_16982,N_16386,N_16161);
or U16983 (N_16983,N_16262,N_16141);
or U16984 (N_16984,N_16295,N_16390);
and U16985 (N_16985,N_16276,N_16499);
or U16986 (N_16986,N_16061,N_16143);
nand U16987 (N_16987,N_16306,N_16170);
xor U16988 (N_16988,N_16108,N_16409);
nor U16989 (N_16989,N_16130,N_16430);
and U16990 (N_16990,N_16049,N_16227);
and U16991 (N_16991,N_16296,N_16101);
nor U16992 (N_16992,N_16154,N_16225);
or U16993 (N_16993,N_16095,N_16126);
and U16994 (N_16994,N_16096,N_16462);
xor U16995 (N_16995,N_16178,N_16315);
nand U16996 (N_16996,N_16304,N_16009);
and U16997 (N_16997,N_16411,N_16286);
or U16998 (N_16998,N_16417,N_16349);
xnor U16999 (N_16999,N_16275,N_16086);
nor U17000 (N_17000,N_16880,N_16557);
nand U17001 (N_17001,N_16886,N_16785);
and U17002 (N_17002,N_16995,N_16946);
nand U17003 (N_17003,N_16893,N_16959);
and U17004 (N_17004,N_16826,N_16737);
and U17005 (N_17005,N_16521,N_16824);
or U17006 (N_17006,N_16853,N_16718);
nand U17007 (N_17007,N_16874,N_16822);
and U17008 (N_17008,N_16912,N_16601);
and U17009 (N_17009,N_16520,N_16794);
nand U17010 (N_17010,N_16745,N_16799);
and U17011 (N_17011,N_16855,N_16990);
or U17012 (N_17012,N_16631,N_16622);
nor U17013 (N_17013,N_16905,N_16936);
nand U17014 (N_17014,N_16660,N_16613);
or U17015 (N_17015,N_16689,N_16892);
nor U17016 (N_17016,N_16906,N_16781);
or U17017 (N_17017,N_16612,N_16553);
and U17018 (N_17018,N_16791,N_16569);
nor U17019 (N_17019,N_16506,N_16789);
nand U17020 (N_17020,N_16820,N_16604);
nand U17021 (N_17021,N_16808,N_16558);
and U17022 (N_17022,N_16917,N_16694);
or U17023 (N_17023,N_16716,N_16502);
nor U17024 (N_17024,N_16866,N_16840);
nand U17025 (N_17025,N_16541,N_16652);
or U17026 (N_17026,N_16849,N_16878);
and U17027 (N_17027,N_16938,N_16534);
nand U17028 (N_17028,N_16698,N_16910);
or U17029 (N_17029,N_16589,N_16619);
or U17030 (N_17030,N_16548,N_16725);
or U17031 (N_17031,N_16816,N_16516);
and U17032 (N_17032,N_16638,N_16828);
or U17033 (N_17033,N_16634,N_16764);
or U17034 (N_17034,N_16955,N_16721);
nor U17035 (N_17035,N_16903,N_16830);
and U17036 (N_17036,N_16802,N_16796);
and U17037 (N_17037,N_16658,N_16738);
and U17038 (N_17038,N_16611,N_16811);
or U17039 (N_17039,N_16549,N_16571);
and U17040 (N_17040,N_16605,N_16897);
nand U17041 (N_17041,N_16735,N_16944);
or U17042 (N_17042,N_16544,N_16530);
nor U17043 (N_17043,N_16931,N_16713);
nand U17044 (N_17044,N_16957,N_16760);
and U17045 (N_17045,N_16927,N_16607);
or U17046 (N_17046,N_16679,N_16630);
and U17047 (N_17047,N_16835,N_16812);
nor U17048 (N_17048,N_16527,N_16709);
and U17049 (N_17049,N_16674,N_16772);
or U17050 (N_17050,N_16987,N_16720);
or U17051 (N_17051,N_16695,N_16861);
nor U17052 (N_17052,N_16623,N_16814);
nor U17053 (N_17053,N_16675,N_16645);
nand U17054 (N_17054,N_16700,N_16710);
nor U17055 (N_17055,N_16852,N_16921);
or U17056 (N_17056,N_16865,N_16692);
nand U17057 (N_17057,N_16625,N_16975);
nor U17058 (N_17058,N_16673,N_16860);
and U17059 (N_17059,N_16948,N_16896);
nor U17060 (N_17060,N_16732,N_16503);
nand U17061 (N_17061,N_16726,N_16514);
nand U17062 (N_17062,N_16668,N_16884);
nand U17063 (N_17063,N_16617,N_16641);
xnor U17064 (N_17064,N_16554,N_16647);
nor U17065 (N_17065,N_16699,N_16600);
nor U17066 (N_17066,N_16810,N_16629);
and U17067 (N_17067,N_16743,N_16986);
or U17068 (N_17068,N_16951,N_16817);
nor U17069 (N_17069,N_16838,N_16529);
nand U17070 (N_17070,N_16627,N_16654);
and U17071 (N_17071,N_16572,N_16934);
or U17072 (N_17072,N_16671,N_16872);
nand U17073 (N_17073,N_16770,N_16940);
nor U17074 (N_17074,N_16680,N_16644);
nor U17075 (N_17075,N_16528,N_16784);
or U17076 (N_17076,N_16797,N_16815);
or U17077 (N_17077,N_16924,N_16588);
or U17078 (N_17078,N_16985,N_16915);
nor U17079 (N_17079,N_16819,N_16564);
and U17080 (N_17080,N_16597,N_16561);
or U17081 (N_17081,N_16596,N_16531);
and U17082 (N_17082,N_16967,N_16583);
nand U17083 (N_17083,N_16578,N_16804);
nand U17084 (N_17084,N_16515,N_16888);
or U17085 (N_17085,N_16657,N_16992);
or U17086 (N_17086,N_16672,N_16926);
xnor U17087 (N_17087,N_16902,N_16733);
and U17088 (N_17088,N_16937,N_16842);
and U17089 (N_17089,N_16535,N_16839);
and U17090 (N_17090,N_16923,N_16730);
xnor U17091 (N_17091,N_16945,N_16859);
xnor U17092 (N_17092,N_16963,N_16961);
and U17093 (N_17093,N_16688,N_16524);
nand U17094 (N_17094,N_16523,N_16996);
nand U17095 (N_17095,N_16882,N_16773);
nand U17096 (N_17096,N_16669,N_16591);
nand U17097 (N_17097,N_16640,N_16593);
nand U17098 (N_17098,N_16509,N_16580);
or U17099 (N_17099,N_16685,N_16599);
nand U17100 (N_17100,N_16821,N_16505);
or U17101 (N_17101,N_16598,N_16576);
and U17102 (N_17102,N_16895,N_16960);
or U17103 (N_17103,N_16707,N_16546);
nand U17104 (N_17104,N_16939,N_16847);
or U17105 (N_17105,N_16751,N_16532);
or U17106 (N_17106,N_16898,N_16649);
and U17107 (N_17107,N_16703,N_16574);
nand U17108 (N_17108,N_16543,N_16740);
nor U17109 (N_17109,N_16628,N_16925);
or U17110 (N_17110,N_16786,N_16891);
nor U17111 (N_17111,N_16782,N_16662);
nand U17112 (N_17112,N_16517,N_16508);
or U17113 (N_17113,N_16650,N_16941);
or U17114 (N_17114,N_16550,N_16954);
or U17115 (N_17115,N_16979,N_16877);
nand U17116 (N_17116,N_16510,N_16603);
nor U17117 (N_17117,N_16953,N_16994);
nor U17118 (N_17118,N_16736,N_16862);
nand U17119 (N_17119,N_16587,N_16901);
nand U17120 (N_17120,N_16846,N_16581);
or U17121 (N_17121,N_16854,N_16761);
nand U17122 (N_17122,N_16916,N_16648);
nor U17123 (N_17123,N_16519,N_16755);
or U17124 (N_17124,N_16827,N_16632);
or U17125 (N_17125,N_16837,N_16970);
and U17126 (N_17126,N_16507,N_16551);
nand U17127 (N_17127,N_16690,N_16741);
and U17128 (N_17128,N_16633,N_16920);
and U17129 (N_17129,N_16869,N_16907);
or U17130 (N_17130,N_16973,N_16919);
or U17131 (N_17131,N_16614,N_16766);
and U17132 (N_17132,N_16731,N_16972);
or U17133 (N_17133,N_16542,N_16806);
or U17134 (N_17134,N_16590,N_16818);
nand U17135 (N_17135,N_16900,N_16547);
or U17136 (N_17136,N_16845,N_16559);
and U17137 (N_17137,N_16798,N_16608);
nand U17138 (N_17138,N_16678,N_16964);
nor U17139 (N_17139,N_16594,N_16702);
nor U17140 (N_17140,N_16778,N_16930);
nor U17141 (N_17141,N_16722,N_16929);
nor U17142 (N_17142,N_16800,N_16750);
nor U17143 (N_17143,N_16579,N_16780);
or U17144 (N_17144,N_16592,N_16705);
nor U17145 (N_17145,N_16833,N_16881);
and U17146 (N_17146,N_16844,N_16663);
and U17147 (N_17147,N_16670,N_16932);
nor U17148 (N_17148,N_16762,N_16701);
nor U17149 (N_17149,N_16918,N_16928);
nor U17150 (N_17150,N_16803,N_16585);
and U17151 (N_17151,N_16795,N_16834);
and U17152 (N_17152,N_16697,N_16825);
and U17153 (N_17153,N_16914,N_16533);
nand U17154 (N_17154,N_16727,N_16922);
and U17155 (N_17155,N_16942,N_16746);
or U17156 (N_17156,N_16752,N_16949);
nand U17157 (N_17157,N_16651,N_16643);
xor U17158 (N_17158,N_16609,N_16909);
and U17159 (N_17159,N_16693,N_16704);
nand U17160 (N_17160,N_16586,N_16974);
nor U17161 (N_17161,N_16763,N_16950);
nand U17162 (N_17162,N_16618,N_16624);
nand U17163 (N_17163,N_16687,N_16536);
or U17164 (N_17164,N_16655,N_16863);
nand U17165 (N_17165,N_16904,N_16653);
nor U17166 (N_17166,N_16984,N_16570);
or U17167 (N_17167,N_16988,N_16767);
or U17168 (N_17168,N_16696,N_16841);
nand U17169 (N_17169,N_16753,N_16538);
or U17170 (N_17170,N_16676,N_16894);
nand U17171 (N_17171,N_16962,N_16666);
nor U17172 (N_17172,N_16754,N_16620);
nor U17173 (N_17173,N_16978,N_16562);
nand U17174 (N_17174,N_16991,N_16626);
nor U17175 (N_17175,N_16980,N_16723);
or U17176 (N_17176,N_16525,N_16777);
or U17177 (N_17177,N_16768,N_16686);
or U17178 (N_17178,N_16565,N_16998);
xor U17179 (N_17179,N_16993,N_16749);
nand U17180 (N_17180,N_16708,N_16775);
nand U17181 (N_17181,N_16968,N_16969);
or U17182 (N_17182,N_16684,N_16511);
or U17183 (N_17183,N_16813,N_16756);
and U17184 (N_17184,N_16563,N_16876);
and U17185 (N_17185,N_16691,N_16513);
or U17186 (N_17186,N_16717,N_16560);
nand U17187 (N_17187,N_16602,N_16724);
nor U17188 (N_17188,N_16729,N_16831);
nand U17189 (N_17189,N_16913,N_16765);
or U17190 (N_17190,N_16889,N_16883);
and U17191 (N_17191,N_16646,N_16879);
or U17192 (N_17192,N_16575,N_16997);
or U17193 (N_17193,N_16867,N_16779);
and U17194 (N_17194,N_16537,N_16555);
nor U17195 (N_17195,N_16790,N_16665);
or U17196 (N_17196,N_16769,N_16595);
nand U17197 (N_17197,N_16843,N_16656);
or U17198 (N_17198,N_16864,N_16805);
or U17199 (N_17199,N_16667,N_16989);
nand U17200 (N_17200,N_16848,N_16832);
and U17201 (N_17201,N_16636,N_16540);
nor U17202 (N_17202,N_16965,N_16635);
and U17203 (N_17203,N_16911,N_16734);
and U17204 (N_17204,N_16664,N_16661);
nand U17205 (N_17205,N_16606,N_16783);
nand U17206 (N_17206,N_16711,N_16801);
nand U17207 (N_17207,N_16871,N_16759);
and U17208 (N_17208,N_16744,N_16850);
and U17209 (N_17209,N_16642,N_16823);
and U17210 (N_17210,N_16504,N_16512);
or U17211 (N_17211,N_16577,N_16682);
nor U17212 (N_17212,N_16719,N_16947);
nor U17213 (N_17213,N_16573,N_16681);
and U17214 (N_17214,N_16639,N_16857);
or U17215 (N_17215,N_16539,N_16836);
nand U17216 (N_17216,N_16758,N_16966);
nand U17217 (N_17217,N_16899,N_16933);
nor U17218 (N_17218,N_16976,N_16977);
and U17219 (N_17219,N_16518,N_16757);
and U17220 (N_17220,N_16582,N_16868);
or U17221 (N_17221,N_16856,N_16637);
or U17222 (N_17222,N_16875,N_16567);
and U17223 (N_17223,N_16870,N_16771);
and U17224 (N_17224,N_16776,N_16873);
or U17225 (N_17225,N_16792,N_16935);
nor U17226 (N_17226,N_16952,N_16615);
or U17227 (N_17227,N_16793,N_16728);
or U17228 (N_17228,N_16712,N_16500);
nor U17229 (N_17229,N_16621,N_16677);
and U17230 (N_17230,N_16568,N_16742);
nor U17231 (N_17231,N_16748,N_16706);
nor U17232 (N_17232,N_16982,N_16616);
or U17233 (N_17233,N_16526,N_16683);
and U17234 (N_17234,N_16858,N_16552);
nand U17235 (N_17235,N_16545,N_16659);
or U17236 (N_17236,N_16943,N_16774);
or U17237 (N_17237,N_16983,N_16809);
nand U17238 (N_17238,N_16887,N_16788);
or U17239 (N_17239,N_16584,N_16885);
and U17240 (N_17240,N_16890,N_16908);
nand U17241 (N_17241,N_16566,N_16971);
nor U17242 (N_17242,N_16747,N_16851);
and U17243 (N_17243,N_16739,N_16956);
nor U17244 (N_17244,N_16958,N_16714);
nand U17245 (N_17245,N_16556,N_16501);
and U17246 (N_17246,N_16981,N_16715);
and U17247 (N_17247,N_16610,N_16787);
nor U17248 (N_17248,N_16807,N_16999);
and U17249 (N_17249,N_16522,N_16829);
or U17250 (N_17250,N_16835,N_16907);
and U17251 (N_17251,N_16862,N_16976);
nand U17252 (N_17252,N_16934,N_16948);
nand U17253 (N_17253,N_16513,N_16731);
nand U17254 (N_17254,N_16713,N_16781);
or U17255 (N_17255,N_16883,N_16723);
or U17256 (N_17256,N_16670,N_16856);
xor U17257 (N_17257,N_16665,N_16514);
nor U17258 (N_17258,N_16919,N_16834);
nor U17259 (N_17259,N_16715,N_16716);
and U17260 (N_17260,N_16572,N_16662);
and U17261 (N_17261,N_16873,N_16828);
nand U17262 (N_17262,N_16886,N_16863);
xnor U17263 (N_17263,N_16608,N_16923);
or U17264 (N_17264,N_16735,N_16911);
nand U17265 (N_17265,N_16920,N_16688);
and U17266 (N_17266,N_16838,N_16612);
nand U17267 (N_17267,N_16818,N_16889);
and U17268 (N_17268,N_16528,N_16854);
or U17269 (N_17269,N_16864,N_16856);
or U17270 (N_17270,N_16713,N_16569);
or U17271 (N_17271,N_16525,N_16663);
or U17272 (N_17272,N_16961,N_16541);
or U17273 (N_17273,N_16599,N_16870);
or U17274 (N_17274,N_16966,N_16915);
nand U17275 (N_17275,N_16890,N_16601);
and U17276 (N_17276,N_16732,N_16743);
nand U17277 (N_17277,N_16893,N_16617);
nand U17278 (N_17278,N_16705,N_16601);
nand U17279 (N_17279,N_16582,N_16724);
nor U17280 (N_17280,N_16745,N_16919);
nor U17281 (N_17281,N_16711,N_16531);
nand U17282 (N_17282,N_16590,N_16797);
or U17283 (N_17283,N_16610,N_16995);
nor U17284 (N_17284,N_16988,N_16647);
or U17285 (N_17285,N_16548,N_16882);
nand U17286 (N_17286,N_16528,N_16998);
and U17287 (N_17287,N_16800,N_16629);
nand U17288 (N_17288,N_16766,N_16891);
or U17289 (N_17289,N_16918,N_16547);
and U17290 (N_17290,N_16810,N_16991);
and U17291 (N_17291,N_16772,N_16987);
nand U17292 (N_17292,N_16843,N_16546);
or U17293 (N_17293,N_16811,N_16606);
and U17294 (N_17294,N_16852,N_16540);
nor U17295 (N_17295,N_16531,N_16557);
or U17296 (N_17296,N_16706,N_16820);
nand U17297 (N_17297,N_16745,N_16623);
and U17298 (N_17298,N_16835,N_16776);
nand U17299 (N_17299,N_16601,N_16832);
or U17300 (N_17300,N_16539,N_16549);
and U17301 (N_17301,N_16775,N_16809);
or U17302 (N_17302,N_16637,N_16645);
nand U17303 (N_17303,N_16951,N_16733);
and U17304 (N_17304,N_16801,N_16929);
nor U17305 (N_17305,N_16903,N_16865);
and U17306 (N_17306,N_16650,N_16767);
nor U17307 (N_17307,N_16540,N_16585);
nor U17308 (N_17308,N_16687,N_16659);
nor U17309 (N_17309,N_16636,N_16846);
or U17310 (N_17310,N_16531,N_16972);
or U17311 (N_17311,N_16707,N_16581);
and U17312 (N_17312,N_16583,N_16778);
nand U17313 (N_17313,N_16666,N_16716);
and U17314 (N_17314,N_16587,N_16637);
or U17315 (N_17315,N_16864,N_16784);
or U17316 (N_17316,N_16979,N_16686);
nor U17317 (N_17317,N_16528,N_16992);
nor U17318 (N_17318,N_16961,N_16955);
nor U17319 (N_17319,N_16613,N_16576);
and U17320 (N_17320,N_16932,N_16974);
and U17321 (N_17321,N_16538,N_16915);
or U17322 (N_17322,N_16603,N_16515);
nand U17323 (N_17323,N_16948,N_16749);
and U17324 (N_17324,N_16901,N_16575);
or U17325 (N_17325,N_16508,N_16779);
nor U17326 (N_17326,N_16575,N_16958);
or U17327 (N_17327,N_16551,N_16982);
nor U17328 (N_17328,N_16789,N_16911);
and U17329 (N_17329,N_16577,N_16857);
nand U17330 (N_17330,N_16645,N_16671);
nand U17331 (N_17331,N_16565,N_16540);
nand U17332 (N_17332,N_16569,N_16520);
or U17333 (N_17333,N_16568,N_16804);
nand U17334 (N_17334,N_16910,N_16849);
nor U17335 (N_17335,N_16986,N_16849);
nand U17336 (N_17336,N_16613,N_16524);
nand U17337 (N_17337,N_16713,N_16907);
nand U17338 (N_17338,N_16602,N_16950);
or U17339 (N_17339,N_16659,N_16718);
nand U17340 (N_17340,N_16572,N_16836);
or U17341 (N_17341,N_16751,N_16776);
nor U17342 (N_17342,N_16718,N_16621);
and U17343 (N_17343,N_16548,N_16582);
and U17344 (N_17344,N_16976,N_16896);
nand U17345 (N_17345,N_16617,N_16583);
and U17346 (N_17346,N_16619,N_16552);
or U17347 (N_17347,N_16992,N_16845);
and U17348 (N_17348,N_16515,N_16880);
nor U17349 (N_17349,N_16505,N_16876);
and U17350 (N_17350,N_16636,N_16677);
nand U17351 (N_17351,N_16810,N_16586);
or U17352 (N_17352,N_16798,N_16866);
nor U17353 (N_17353,N_16685,N_16891);
nand U17354 (N_17354,N_16766,N_16895);
nor U17355 (N_17355,N_16985,N_16943);
and U17356 (N_17356,N_16638,N_16855);
nand U17357 (N_17357,N_16561,N_16721);
nor U17358 (N_17358,N_16838,N_16982);
nand U17359 (N_17359,N_16730,N_16617);
or U17360 (N_17360,N_16782,N_16703);
nor U17361 (N_17361,N_16784,N_16688);
nand U17362 (N_17362,N_16571,N_16846);
nor U17363 (N_17363,N_16855,N_16648);
and U17364 (N_17364,N_16990,N_16902);
nor U17365 (N_17365,N_16556,N_16994);
nor U17366 (N_17366,N_16953,N_16726);
and U17367 (N_17367,N_16907,N_16576);
or U17368 (N_17368,N_16842,N_16584);
nor U17369 (N_17369,N_16713,N_16675);
nand U17370 (N_17370,N_16544,N_16578);
nor U17371 (N_17371,N_16899,N_16793);
and U17372 (N_17372,N_16605,N_16744);
nand U17373 (N_17373,N_16904,N_16785);
nor U17374 (N_17374,N_16580,N_16796);
and U17375 (N_17375,N_16538,N_16907);
and U17376 (N_17376,N_16961,N_16747);
and U17377 (N_17377,N_16616,N_16779);
nand U17378 (N_17378,N_16544,N_16942);
nor U17379 (N_17379,N_16609,N_16554);
nor U17380 (N_17380,N_16552,N_16526);
nand U17381 (N_17381,N_16965,N_16542);
or U17382 (N_17382,N_16757,N_16907);
nor U17383 (N_17383,N_16821,N_16598);
and U17384 (N_17384,N_16660,N_16732);
and U17385 (N_17385,N_16761,N_16802);
nor U17386 (N_17386,N_16864,N_16673);
or U17387 (N_17387,N_16525,N_16619);
or U17388 (N_17388,N_16870,N_16516);
or U17389 (N_17389,N_16531,N_16983);
nand U17390 (N_17390,N_16630,N_16702);
xor U17391 (N_17391,N_16981,N_16602);
and U17392 (N_17392,N_16916,N_16966);
nand U17393 (N_17393,N_16891,N_16789);
nand U17394 (N_17394,N_16822,N_16552);
nor U17395 (N_17395,N_16965,N_16575);
or U17396 (N_17396,N_16612,N_16949);
and U17397 (N_17397,N_16927,N_16500);
nor U17398 (N_17398,N_16826,N_16695);
nor U17399 (N_17399,N_16617,N_16992);
nor U17400 (N_17400,N_16708,N_16531);
nand U17401 (N_17401,N_16754,N_16846);
nand U17402 (N_17402,N_16690,N_16961);
or U17403 (N_17403,N_16741,N_16771);
nand U17404 (N_17404,N_16874,N_16800);
nor U17405 (N_17405,N_16572,N_16855);
and U17406 (N_17406,N_16657,N_16748);
nand U17407 (N_17407,N_16799,N_16587);
and U17408 (N_17408,N_16536,N_16723);
and U17409 (N_17409,N_16781,N_16544);
or U17410 (N_17410,N_16984,N_16883);
xnor U17411 (N_17411,N_16662,N_16809);
and U17412 (N_17412,N_16881,N_16616);
or U17413 (N_17413,N_16923,N_16605);
or U17414 (N_17414,N_16794,N_16502);
or U17415 (N_17415,N_16938,N_16526);
nand U17416 (N_17416,N_16894,N_16925);
and U17417 (N_17417,N_16865,N_16895);
nand U17418 (N_17418,N_16760,N_16877);
and U17419 (N_17419,N_16592,N_16513);
nor U17420 (N_17420,N_16807,N_16791);
and U17421 (N_17421,N_16677,N_16680);
and U17422 (N_17422,N_16734,N_16838);
and U17423 (N_17423,N_16684,N_16930);
and U17424 (N_17424,N_16945,N_16796);
nand U17425 (N_17425,N_16755,N_16961);
nor U17426 (N_17426,N_16805,N_16712);
nand U17427 (N_17427,N_16808,N_16583);
nand U17428 (N_17428,N_16696,N_16976);
or U17429 (N_17429,N_16878,N_16823);
nor U17430 (N_17430,N_16721,N_16956);
and U17431 (N_17431,N_16755,N_16511);
or U17432 (N_17432,N_16753,N_16726);
nand U17433 (N_17433,N_16654,N_16691);
or U17434 (N_17434,N_16544,N_16880);
and U17435 (N_17435,N_16885,N_16744);
nor U17436 (N_17436,N_16867,N_16536);
nand U17437 (N_17437,N_16733,N_16823);
nand U17438 (N_17438,N_16807,N_16830);
nand U17439 (N_17439,N_16800,N_16717);
nor U17440 (N_17440,N_16828,N_16917);
and U17441 (N_17441,N_16718,N_16557);
nor U17442 (N_17442,N_16586,N_16752);
nor U17443 (N_17443,N_16970,N_16611);
and U17444 (N_17444,N_16646,N_16704);
or U17445 (N_17445,N_16635,N_16953);
nor U17446 (N_17446,N_16955,N_16964);
nor U17447 (N_17447,N_16542,N_16839);
nand U17448 (N_17448,N_16726,N_16916);
nor U17449 (N_17449,N_16954,N_16841);
nor U17450 (N_17450,N_16809,N_16897);
nor U17451 (N_17451,N_16728,N_16872);
or U17452 (N_17452,N_16893,N_16718);
and U17453 (N_17453,N_16942,N_16540);
and U17454 (N_17454,N_16804,N_16726);
or U17455 (N_17455,N_16606,N_16597);
or U17456 (N_17456,N_16801,N_16808);
or U17457 (N_17457,N_16825,N_16815);
and U17458 (N_17458,N_16621,N_16661);
and U17459 (N_17459,N_16799,N_16594);
and U17460 (N_17460,N_16595,N_16857);
nand U17461 (N_17461,N_16517,N_16868);
or U17462 (N_17462,N_16710,N_16603);
nor U17463 (N_17463,N_16627,N_16901);
nand U17464 (N_17464,N_16622,N_16910);
nor U17465 (N_17465,N_16876,N_16628);
and U17466 (N_17466,N_16607,N_16665);
nand U17467 (N_17467,N_16992,N_16700);
nor U17468 (N_17468,N_16742,N_16695);
nor U17469 (N_17469,N_16517,N_16668);
or U17470 (N_17470,N_16653,N_16903);
and U17471 (N_17471,N_16932,N_16789);
or U17472 (N_17472,N_16892,N_16557);
or U17473 (N_17473,N_16619,N_16721);
or U17474 (N_17474,N_16987,N_16918);
nor U17475 (N_17475,N_16883,N_16771);
and U17476 (N_17476,N_16576,N_16993);
nor U17477 (N_17477,N_16655,N_16536);
or U17478 (N_17478,N_16565,N_16846);
nand U17479 (N_17479,N_16557,N_16757);
nor U17480 (N_17480,N_16820,N_16942);
nand U17481 (N_17481,N_16741,N_16755);
nand U17482 (N_17482,N_16664,N_16964);
nor U17483 (N_17483,N_16588,N_16806);
or U17484 (N_17484,N_16613,N_16898);
nor U17485 (N_17485,N_16872,N_16696);
nand U17486 (N_17486,N_16779,N_16711);
nor U17487 (N_17487,N_16902,N_16808);
nor U17488 (N_17488,N_16507,N_16830);
nor U17489 (N_17489,N_16957,N_16695);
and U17490 (N_17490,N_16699,N_16584);
and U17491 (N_17491,N_16968,N_16508);
or U17492 (N_17492,N_16553,N_16720);
xnor U17493 (N_17493,N_16656,N_16659);
or U17494 (N_17494,N_16896,N_16881);
or U17495 (N_17495,N_16968,N_16535);
nand U17496 (N_17496,N_16956,N_16732);
and U17497 (N_17497,N_16728,N_16932);
and U17498 (N_17498,N_16755,N_16943);
nor U17499 (N_17499,N_16639,N_16908);
nor U17500 (N_17500,N_17181,N_17213);
nor U17501 (N_17501,N_17452,N_17384);
and U17502 (N_17502,N_17416,N_17197);
or U17503 (N_17503,N_17393,N_17426);
nand U17504 (N_17504,N_17327,N_17085);
xor U17505 (N_17505,N_17039,N_17270);
nand U17506 (N_17506,N_17277,N_17128);
and U17507 (N_17507,N_17492,N_17383);
nand U17508 (N_17508,N_17049,N_17402);
or U17509 (N_17509,N_17314,N_17227);
and U17510 (N_17510,N_17468,N_17407);
or U17511 (N_17511,N_17204,N_17088);
nand U17512 (N_17512,N_17359,N_17486);
and U17513 (N_17513,N_17048,N_17023);
nand U17514 (N_17514,N_17196,N_17487);
nor U17515 (N_17515,N_17377,N_17150);
nor U17516 (N_17516,N_17084,N_17086);
nor U17517 (N_17517,N_17073,N_17001);
and U17518 (N_17518,N_17463,N_17059);
nand U17519 (N_17519,N_17067,N_17311);
nor U17520 (N_17520,N_17089,N_17496);
or U17521 (N_17521,N_17046,N_17449);
or U17522 (N_17522,N_17349,N_17003);
nand U17523 (N_17523,N_17279,N_17470);
nor U17524 (N_17524,N_17348,N_17082);
nor U17525 (N_17525,N_17040,N_17062);
nor U17526 (N_17526,N_17388,N_17098);
and U17527 (N_17527,N_17281,N_17199);
and U17528 (N_17528,N_17378,N_17251);
and U17529 (N_17529,N_17057,N_17207);
or U17530 (N_17530,N_17136,N_17029);
or U17531 (N_17531,N_17410,N_17341);
or U17532 (N_17532,N_17269,N_17072);
xnor U17533 (N_17533,N_17068,N_17322);
nor U17534 (N_17534,N_17376,N_17351);
and U17535 (N_17535,N_17119,N_17493);
nor U17536 (N_17536,N_17484,N_17256);
xnor U17537 (N_17537,N_17032,N_17024);
nor U17538 (N_17538,N_17053,N_17333);
nand U17539 (N_17539,N_17090,N_17236);
nor U17540 (N_17540,N_17448,N_17299);
nor U17541 (N_17541,N_17389,N_17397);
nor U17542 (N_17542,N_17056,N_17058);
nor U17543 (N_17543,N_17478,N_17229);
and U17544 (N_17544,N_17160,N_17362);
and U17545 (N_17545,N_17353,N_17329);
and U17546 (N_17546,N_17273,N_17079);
or U17547 (N_17547,N_17445,N_17016);
or U17548 (N_17548,N_17316,N_17392);
or U17549 (N_17549,N_17069,N_17144);
nor U17550 (N_17550,N_17159,N_17363);
or U17551 (N_17551,N_17497,N_17409);
nand U17552 (N_17552,N_17284,N_17011);
nor U17553 (N_17553,N_17276,N_17442);
nor U17554 (N_17554,N_17390,N_17203);
xor U17555 (N_17555,N_17296,N_17044);
or U17556 (N_17556,N_17163,N_17356);
nor U17557 (N_17557,N_17161,N_17176);
xor U17558 (N_17558,N_17135,N_17050);
and U17559 (N_17559,N_17274,N_17483);
nor U17560 (N_17560,N_17330,N_17495);
and U17561 (N_17561,N_17433,N_17107);
or U17562 (N_17562,N_17000,N_17194);
and U17563 (N_17563,N_17450,N_17177);
nor U17564 (N_17564,N_17360,N_17352);
or U17565 (N_17565,N_17216,N_17428);
or U17566 (N_17566,N_17110,N_17182);
and U17567 (N_17567,N_17052,N_17342);
and U17568 (N_17568,N_17337,N_17071);
nand U17569 (N_17569,N_17063,N_17117);
nor U17570 (N_17570,N_17241,N_17343);
or U17571 (N_17571,N_17244,N_17443);
and U17572 (N_17572,N_17317,N_17162);
nor U17573 (N_17573,N_17247,N_17315);
and U17574 (N_17574,N_17122,N_17007);
or U17575 (N_17575,N_17141,N_17218);
or U17576 (N_17576,N_17025,N_17231);
nor U17577 (N_17577,N_17020,N_17455);
or U17578 (N_17578,N_17149,N_17419);
nor U17579 (N_17579,N_17192,N_17103);
nand U17580 (N_17580,N_17260,N_17168);
or U17581 (N_17581,N_17254,N_17152);
or U17582 (N_17582,N_17457,N_17259);
nand U17583 (N_17583,N_17258,N_17075);
nor U17584 (N_17584,N_17013,N_17239);
or U17585 (N_17585,N_17386,N_17193);
nor U17586 (N_17586,N_17081,N_17187);
nand U17587 (N_17587,N_17441,N_17275);
or U17588 (N_17588,N_17369,N_17232);
nor U17589 (N_17589,N_17083,N_17022);
nand U17590 (N_17590,N_17105,N_17051);
xnor U17591 (N_17591,N_17476,N_17195);
nand U17592 (N_17592,N_17403,N_17070);
nor U17593 (N_17593,N_17220,N_17094);
nand U17594 (N_17594,N_17246,N_17235);
nor U17595 (N_17595,N_17158,N_17268);
or U17596 (N_17596,N_17139,N_17435);
nor U17597 (N_17597,N_17242,N_17401);
nor U17598 (N_17598,N_17221,N_17190);
nand U17599 (N_17599,N_17233,N_17146);
nor U17600 (N_17600,N_17200,N_17347);
nor U17601 (N_17601,N_17436,N_17173);
xor U17602 (N_17602,N_17300,N_17164);
and U17603 (N_17603,N_17208,N_17026);
and U17604 (N_17604,N_17382,N_17148);
nand U17605 (N_17605,N_17261,N_17250);
or U17606 (N_17606,N_17368,N_17267);
or U17607 (N_17607,N_17425,N_17042);
nand U17608 (N_17608,N_17485,N_17114);
nand U17609 (N_17609,N_17255,N_17466);
xnor U17610 (N_17610,N_17321,N_17350);
or U17611 (N_17611,N_17074,N_17406);
nand U17612 (N_17612,N_17033,N_17440);
and U17613 (N_17613,N_17120,N_17278);
nand U17614 (N_17614,N_17472,N_17249);
and U17615 (N_17615,N_17238,N_17215);
nand U17616 (N_17616,N_17184,N_17320);
or U17617 (N_17617,N_17453,N_17087);
or U17618 (N_17618,N_17325,N_17400);
and U17619 (N_17619,N_17387,N_17465);
and U17620 (N_17620,N_17475,N_17118);
or U17621 (N_17621,N_17340,N_17174);
and U17622 (N_17622,N_17143,N_17209);
or U17623 (N_17623,N_17396,N_17112);
or U17624 (N_17624,N_17202,N_17418);
and U17625 (N_17625,N_17447,N_17096);
and U17626 (N_17626,N_17093,N_17432);
or U17627 (N_17627,N_17293,N_17129);
nor U17628 (N_17628,N_17041,N_17291);
nor U17629 (N_17629,N_17272,N_17477);
or U17630 (N_17630,N_17106,N_17155);
and U17631 (N_17631,N_17345,N_17423);
nand U17632 (N_17632,N_17456,N_17123);
nand U17633 (N_17633,N_17370,N_17469);
nand U17634 (N_17634,N_17212,N_17334);
and U17635 (N_17635,N_17134,N_17482);
nand U17636 (N_17636,N_17346,N_17055);
and U17637 (N_17637,N_17228,N_17338);
or U17638 (N_17638,N_17132,N_17313);
nor U17639 (N_17639,N_17367,N_17344);
and U17640 (N_17640,N_17121,N_17294);
or U17641 (N_17641,N_17131,N_17262);
nor U17642 (N_17642,N_17210,N_17153);
and U17643 (N_17643,N_17065,N_17439);
nand U17644 (N_17644,N_17361,N_17167);
nand U17645 (N_17645,N_17318,N_17461);
nand U17646 (N_17646,N_17230,N_17223);
nand U17647 (N_17647,N_17156,N_17133);
or U17648 (N_17648,N_17422,N_17140);
or U17649 (N_17649,N_17336,N_17028);
nor U17650 (N_17650,N_17429,N_17288);
and U17651 (N_17651,N_17111,N_17489);
nor U17652 (N_17652,N_17004,N_17287);
and U17653 (N_17653,N_17467,N_17171);
and U17654 (N_17654,N_17038,N_17339);
and U17655 (N_17655,N_17286,N_17295);
or U17656 (N_17656,N_17289,N_17283);
nand U17657 (N_17657,N_17309,N_17408);
nand U17658 (N_17658,N_17101,N_17175);
nor U17659 (N_17659,N_17104,N_17198);
or U17660 (N_17660,N_17054,N_17014);
and U17661 (N_17661,N_17091,N_17394);
or U17662 (N_17662,N_17460,N_17189);
nor U17663 (N_17663,N_17464,N_17126);
or U17664 (N_17664,N_17109,N_17335);
or U17665 (N_17665,N_17015,N_17061);
or U17666 (N_17666,N_17324,N_17328);
and U17667 (N_17667,N_17302,N_17290);
nand U17668 (N_17668,N_17264,N_17405);
or U17669 (N_17669,N_17364,N_17166);
nor U17670 (N_17670,N_17234,N_17301);
nor U17671 (N_17671,N_17430,N_17374);
nor U17672 (N_17672,N_17180,N_17080);
nand U17673 (N_17673,N_17248,N_17027);
or U17674 (N_17674,N_17375,N_17115);
nor U17675 (N_17675,N_17017,N_17127);
and U17676 (N_17676,N_17271,N_17308);
and U17677 (N_17677,N_17357,N_17266);
nor U17678 (N_17678,N_17043,N_17037);
xnor U17679 (N_17679,N_17446,N_17404);
or U17680 (N_17680,N_17380,N_17355);
or U17681 (N_17681,N_17481,N_17245);
nor U17682 (N_17682,N_17124,N_17462);
and U17683 (N_17683,N_17205,N_17490);
nor U17684 (N_17684,N_17045,N_17391);
nand U17685 (N_17685,N_17398,N_17219);
nor U17686 (N_17686,N_17385,N_17169);
or U17687 (N_17687,N_17373,N_17165);
xor U17688 (N_17688,N_17005,N_17417);
and U17689 (N_17689,N_17036,N_17185);
and U17690 (N_17690,N_17395,N_17225);
nand U17691 (N_17691,N_17444,N_17310);
and U17692 (N_17692,N_17331,N_17116);
nand U17693 (N_17693,N_17030,N_17459);
nand U17694 (N_17694,N_17170,N_17280);
or U17695 (N_17695,N_17031,N_17018);
nor U17696 (N_17696,N_17237,N_17008);
nor U17697 (N_17697,N_17130,N_17222);
nand U17698 (N_17698,N_17421,N_17147);
nand U17699 (N_17699,N_17240,N_17113);
and U17700 (N_17700,N_17186,N_17191);
nor U17701 (N_17701,N_17066,N_17097);
and U17702 (N_17702,N_17172,N_17019);
or U17703 (N_17703,N_17252,N_17076);
or U17704 (N_17704,N_17413,N_17437);
nand U17705 (N_17705,N_17379,N_17060);
nor U17706 (N_17706,N_17479,N_17499);
nor U17707 (N_17707,N_17206,N_17035);
nand U17708 (N_17708,N_17471,N_17095);
or U17709 (N_17709,N_17157,N_17078);
and U17710 (N_17710,N_17145,N_17306);
or U17711 (N_17711,N_17491,N_17381);
and U17712 (N_17712,N_17188,N_17179);
and U17713 (N_17713,N_17354,N_17473);
or U17714 (N_17714,N_17323,N_17285);
or U17715 (N_17715,N_17399,N_17319);
nand U17716 (N_17716,N_17420,N_17297);
and U17717 (N_17717,N_17138,N_17125);
and U17718 (N_17718,N_17458,N_17292);
or U17719 (N_17719,N_17102,N_17411);
or U17720 (N_17720,N_17108,N_17312);
nor U17721 (N_17721,N_17332,N_17498);
nor U17722 (N_17722,N_17434,N_17431);
or U17723 (N_17723,N_17021,N_17365);
and U17724 (N_17724,N_17183,N_17454);
and U17725 (N_17725,N_17488,N_17034);
or U17726 (N_17726,N_17414,N_17253);
or U17727 (N_17727,N_17142,N_17263);
nand U17728 (N_17728,N_17077,N_17047);
nor U17729 (N_17729,N_17154,N_17372);
and U17730 (N_17730,N_17178,N_17438);
and U17731 (N_17731,N_17282,N_17427);
nor U17732 (N_17732,N_17100,N_17366);
or U17733 (N_17733,N_17064,N_17243);
nor U17734 (N_17734,N_17305,N_17415);
and U17735 (N_17735,N_17257,N_17137);
or U17736 (N_17736,N_17010,N_17211);
nand U17737 (N_17737,N_17412,N_17009);
and U17738 (N_17738,N_17358,N_17298);
nand U17739 (N_17739,N_17151,N_17265);
or U17740 (N_17740,N_17012,N_17099);
and U17741 (N_17741,N_17304,N_17480);
nand U17742 (N_17742,N_17226,N_17303);
and U17743 (N_17743,N_17002,N_17326);
or U17744 (N_17744,N_17217,N_17307);
and U17745 (N_17745,N_17224,N_17371);
or U17746 (N_17746,N_17092,N_17474);
nor U17747 (N_17747,N_17494,N_17451);
nor U17748 (N_17748,N_17424,N_17201);
or U17749 (N_17749,N_17006,N_17214);
or U17750 (N_17750,N_17398,N_17061);
and U17751 (N_17751,N_17390,N_17010);
nand U17752 (N_17752,N_17161,N_17135);
nor U17753 (N_17753,N_17130,N_17389);
nand U17754 (N_17754,N_17365,N_17008);
nor U17755 (N_17755,N_17328,N_17472);
xnor U17756 (N_17756,N_17324,N_17353);
nor U17757 (N_17757,N_17309,N_17220);
nand U17758 (N_17758,N_17348,N_17476);
and U17759 (N_17759,N_17355,N_17426);
nand U17760 (N_17760,N_17296,N_17325);
nand U17761 (N_17761,N_17405,N_17360);
or U17762 (N_17762,N_17208,N_17055);
or U17763 (N_17763,N_17257,N_17031);
nand U17764 (N_17764,N_17393,N_17029);
or U17765 (N_17765,N_17293,N_17212);
nor U17766 (N_17766,N_17012,N_17111);
nor U17767 (N_17767,N_17090,N_17115);
nor U17768 (N_17768,N_17021,N_17371);
or U17769 (N_17769,N_17313,N_17424);
or U17770 (N_17770,N_17365,N_17292);
and U17771 (N_17771,N_17317,N_17226);
nand U17772 (N_17772,N_17006,N_17216);
nand U17773 (N_17773,N_17458,N_17417);
and U17774 (N_17774,N_17418,N_17218);
nand U17775 (N_17775,N_17366,N_17189);
or U17776 (N_17776,N_17063,N_17382);
nand U17777 (N_17777,N_17205,N_17090);
and U17778 (N_17778,N_17091,N_17492);
and U17779 (N_17779,N_17019,N_17259);
and U17780 (N_17780,N_17244,N_17223);
or U17781 (N_17781,N_17466,N_17097);
nand U17782 (N_17782,N_17158,N_17035);
and U17783 (N_17783,N_17327,N_17136);
nor U17784 (N_17784,N_17231,N_17391);
and U17785 (N_17785,N_17255,N_17246);
and U17786 (N_17786,N_17262,N_17409);
nor U17787 (N_17787,N_17044,N_17479);
and U17788 (N_17788,N_17158,N_17063);
nand U17789 (N_17789,N_17307,N_17197);
nand U17790 (N_17790,N_17349,N_17207);
or U17791 (N_17791,N_17063,N_17099);
or U17792 (N_17792,N_17297,N_17216);
and U17793 (N_17793,N_17165,N_17112);
xor U17794 (N_17794,N_17057,N_17164);
and U17795 (N_17795,N_17472,N_17149);
and U17796 (N_17796,N_17140,N_17448);
or U17797 (N_17797,N_17053,N_17447);
and U17798 (N_17798,N_17478,N_17158);
or U17799 (N_17799,N_17490,N_17053);
nor U17800 (N_17800,N_17363,N_17271);
and U17801 (N_17801,N_17399,N_17422);
or U17802 (N_17802,N_17285,N_17282);
or U17803 (N_17803,N_17298,N_17302);
xor U17804 (N_17804,N_17133,N_17285);
and U17805 (N_17805,N_17327,N_17288);
nor U17806 (N_17806,N_17426,N_17219);
nand U17807 (N_17807,N_17032,N_17442);
nor U17808 (N_17808,N_17397,N_17328);
and U17809 (N_17809,N_17164,N_17000);
or U17810 (N_17810,N_17118,N_17200);
nand U17811 (N_17811,N_17035,N_17237);
or U17812 (N_17812,N_17324,N_17498);
nor U17813 (N_17813,N_17248,N_17315);
nand U17814 (N_17814,N_17190,N_17231);
and U17815 (N_17815,N_17200,N_17262);
nand U17816 (N_17816,N_17200,N_17150);
or U17817 (N_17817,N_17210,N_17020);
nand U17818 (N_17818,N_17237,N_17081);
or U17819 (N_17819,N_17345,N_17104);
and U17820 (N_17820,N_17192,N_17077);
nand U17821 (N_17821,N_17076,N_17355);
nor U17822 (N_17822,N_17305,N_17241);
xor U17823 (N_17823,N_17435,N_17073);
nor U17824 (N_17824,N_17450,N_17271);
nor U17825 (N_17825,N_17185,N_17306);
xnor U17826 (N_17826,N_17143,N_17190);
or U17827 (N_17827,N_17472,N_17343);
nor U17828 (N_17828,N_17086,N_17369);
nand U17829 (N_17829,N_17019,N_17189);
nand U17830 (N_17830,N_17126,N_17023);
or U17831 (N_17831,N_17196,N_17178);
and U17832 (N_17832,N_17042,N_17432);
or U17833 (N_17833,N_17244,N_17156);
nor U17834 (N_17834,N_17386,N_17269);
nand U17835 (N_17835,N_17137,N_17151);
and U17836 (N_17836,N_17258,N_17291);
nor U17837 (N_17837,N_17410,N_17372);
and U17838 (N_17838,N_17208,N_17172);
nor U17839 (N_17839,N_17090,N_17050);
nand U17840 (N_17840,N_17014,N_17021);
nand U17841 (N_17841,N_17111,N_17251);
nand U17842 (N_17842,N_17095,N_17110);
and U17843 (N_17843,N_17457,N_17347);
nor U17844 (N_17844,N_17487,N_17331);
nor U17845 (N_17845,N_17240,N_17122);
nand U17846 (N_17846,N_17232,N_17471);
nand U17847 (N_17847,N_17134,N_17281);
nor U17848 (N_17848,N_17401,N_17239);
nand U17849 (N_17849,N_17271,N_17068);
nand U17850 (N_17850,N_17042,N_17256);
nand U17851 (N_17851,N_17117,N_17287);
or U17852 (N_17852,N_17455,N_17115);
and U17853 (N_17853,N_17353,N_17330);
nand U17854 (N_17854,N_17125,N_17041);
nor U17855 (N_17855,N_17169,N_17139);
nor U17856 (N_17856,N_17299,N_17088);
or U17857 (N_17857,N_17149,N_17026);
nand U17858 (N_17858,N_17416,N_17015);
or U17859 (N_17859,N_17178,N_17398);
xnor U17860 (N_17860,N_17112,N_17419);
nand U17861 (N_17861,N_17077,N_17418);
nand U17862 (N_17862,N_17414,N_17176);
nand U17863 (N_17863,N_17123,N_17264);
nor U17864 (N_17864,N_17188,N_17041);
and U17865 (N_17865,N_17077,N_17031);
nand U17866 (N_17866,N_17333,N_17216);
nand U17867 (N_17867,N_17411,N_17038);
nor U17868 (N_17868,N_17434,N_17406);
nand U17869 (N_17869,N_17320,N_17366);
nand U17870 (N_17870,N_17171,N_17141);
nand U17871 (N_17871,N_17273,N_17059);
xnor U17872 (N_17872,N_17438,N_17150);
or U17873 (N_17873,N_17499,N_17412);
or U17874 (N_17874,N_17227,N_17201);
nand U17875 (N_17875,N_17447,N_17173);
nand U17876 (N_17876,N_17169,N_17221);
nor U17877 (N_17877,N_17081,N_17363);
and U17878 (N_17878,N_17471,N_17248);
and U17879 (N_17879,N_17361,N_17457);
nand U17880 (N_17880,N_17199,N_17381);
nor U17881 (N_17881,N_17362,N_17374);
nor U17882 (N_17882,N_17085,N_17400);
and U17883 (N_17883,N_17101,N_17489);
or U17884 (N_17884,N_17400,N_17225);
or U17885 (N_17885,N_17248,N_17271);
and U17886 (N_17886,N_17452,N_17146);
and U17887 (N_17887,N_17211,N_17153);
or U17888 (N_17888,N_17326,N_17186);
or U17889 (N_17889,N_17372,N_17490);
and U17890 (N_17890,N_17249,N_17284);
nand U17891 (N_17891,N_17213,N_17227);
nor U17892 (N_17892,N_17176,N_17035);
nor U17893 (N_17893,N_17403,N_17301);
or U17894 (N_17894,N_17052,N_17123);
nand U17895 (N_17895,N_17082,N_17332);
nor U17896 (N_17896,N_17106,N_17243);
nand U17897 (N_17897,N_17409,N_17088);
nor U17898 (N_17898,N_17404,N_17464);
nand U17899 (N_17899,N_17005,N_17485);
nand U17900 (N_17900,N_17045,N_17348);
or U17901 (N_17901,N_17357,N_17442);
nor U17902 (N_17902,N_17043,N_17357);
nor U17903 (N_17903,N_17252,N_17077);
nor U17904 (N_17904,N_17312,N_17362);
and U17905 (N_17905,N_17289,N_17290);
or U17906 (N_17906,N_17479,N_17282);
and U17907 (N_17907,N_17466,N_17452);
and U17908 (N_17908,N_17110,N_17070);
nand U17909 (N_17909,N_17080,N_17435);
and U17910 (N_17910,N_17348,N_17321);
and U17911 (N_17911,N_17296,N_17197);
or U17912 (N_17912,N_17329,N_17073);
nand U17913 (N_17913,N_17000,N_17392);
nor U17914 (N_17914,N_17156,N_17059);
or U17915 (N_17915,N_17035,N_17342);
xor U17916 (N_17916,N_17159,N_17224);
nor U17917 (N_17917,N_17046,N_17175);
or U17918 (N_17918,N_17193,N_17230);
nand U17919 (N_17919,N_17395,N_17423);
nand U17920 (N_17920,N_17472,N_17032);
nand U17921 (N_17921,N_17125,N_17235);
nand U17922 (N_17922,N_17488,N_17072);
nor U17923 (N_17923,N_17031,N_17459);
xnor U17924 (N_17924,N_17489,N_17091);
nand U17925 (N_17925,N_17336,N_17153);
nor U17926 (N_17926,N_17268,N_17151);
nand U17927 (N_17927,N_17200,N_17082);
nand U17928 (N_17928,N_17351,N_17479);
or U17929 (N_17929,N_17047,N_17229);
nand U17930 (N_17930,N_17051,N_17156);
nor U17931 (N_17931,N_17210,N_17187);
nor U17932 (N_17932,N_17085,N_17032);
or U17933 (N_17933,N_17197,N_17023);
nor U17934 (N_17934,N_17324,N_17006);
and U17935 (N_17935,N_17147,N_17410);
or U17936 (N_17936,N_17103,N_17024);
or U17937 (N_17937,N_17228,N_17083);
and U17938 (N_17938,N_17376,N_17112);
or U17939 (N_17939,N_17399,N_17050);
and U17940 (N_17940,N_17405,N_17173);
or U17941 (N_17941,N_17042,N_17096);
nand U17942 (N_17942,N_17024,N_17283);
and U17943 (N_17943,N_17424,N_17274);
and U17944 (N_17944,N_17436,N_17046);
nor U17945 (N_17945,N_17196,N_17198);
and U17946 (N_17946,N_17424,N_17418);
nor U17947 (N_17947,N_17309,N_17136);
nor U17948 (N_17948,N_17498,N_17263);
and U17949 (N_17949,N_17434,N_17250);
nand U17950 (N_17950,N_17211,N_17041);
nand U17951 (N_17951,N_17492,N_17486);
and U17952 (N_17952,N_17114,N_17041);
or U17953 (N_17953,N_17002,N_17197);
and U17954 (N_17954,N_17437,N_17108);
and U17955 (N_17955,N_17205,N_17437);
nand U17956 (N_17956,N_17304,N_17106);
nand U17957 (N_17957,N_17019,N_17303);
nand U17958 (N_17958,N_17374,N_17161);
xnor U17959 (N_17959,N_17158,N_17329);
nand U17960 (N_17960,N_17414,N_17357);
nor U17961 (N_17961,N_17066,N_17078);
nor U17962 (N_17962,N_17431,N_17476);
or U17963 (N_17963,N_17019,N_17087);
or U17964 (N_17964,N_17224,N_17412);
xnor U17965 (N_17965,N_17410,N_17111);
and U17966 (N_17966,N_17417,N_17474);
nand U17967 (N_17967,N_17440,N_17086);
nand U17968 (N_17968,N_17330,N_17115);
or U17969 (N_17969,N_17037,N_17253);
nand U17970 (N_17970,N_17033,N_17159);
and U17971 (N_17971,N_17444,N_17486);
or U17972 (N_17972,N_17452,N_17030);
nor U17973 (N_17973,N_17253,N_17492);
or U17974 (N_17974,N_17442,N_17110);
nor U17975 (N_17975,N_17247,N_17312);
nand U17976 (N_17976,N_17368,N_17301);
nor U17977 (N_17977,N_17409,N_17456);
or U17978 (N_17978,N_17061,N_17402);
or U17979 (N_17979,N_17188,N_17121);
or U17980 (N_17980,N_17449,N_17467);
nand U17981 (N_17981,N_17458,N_17067);
nand U17982 (N_17982,N_17215,N_17320);
and U17983 (N_17983,N_17099,N_17289);
nor U17984 (N_17984,N_17237,N_17142);
or U17985 (N_17985,N_17024,N_17034);
nor U17986 (N_17986,N_17484,N_17226);
nor U17987 (N_17987,N_17169,N_17238);
nor U17988 (N_17988,N_17086,N_17407);
and U17989 (N_17989,N_17380,N_17351);
or U17990 (N_17990,N_17285,N_17239);
and U17991 (N_17991,N_17024,N_17118);
and U17992 (N_17992,N_17321,N_17248);
nor U17993 (N_17993,N_17047,N_17382);
and U17994 (N_17994,N_17447,N_17305);
nor U17995 (N_17995,N_17341,N_17355);
or U17996 (N_17996,N_17218,N_17039);
nand U17997 (N_17997,N_17490,N_17200);
nand U17998 (N_17998,N_17444,N_17496);
nand U17999 (N_17999,N_17041,N_17055);
or U18000 (N_18000,N_17979,N_17647);
nor U18001 (N_18001,N_17856,N_17952);
and U18002 (N_18002,N_17871,N_17673);
or U18003 (N_18003,N_17506,N_17783);
and U18004 (N_18004,N_17615,N_17646);
or U18005 (N_18005,N_17635,N_17714);
nor U18006 (N_18006,N_17942,N_17622);
and U18007 (N_18007,N_17529,N_17521);
nor U18008 (N_18008,N_17539,N_17924);
nand U18009 (N_18009,N_17965,N_17758);
and U18010 (N_18010,N_17860,N_17730);
xnor U18011 (N_18011,N_17610,N_17722);
nand U18012 (N_18012,N_17763,N_17697);
nand U18013 (N_18013,N_17626,N_17684);
or U18014 (N_18014,N_17654,N_17584);
nand U18015 (N_18015,N_17900,N_17962);
nand U18016 (N_18016,N_17837,N_17875);
or U18017 (N_18017,N_17554,N_17855);
and U18018 (N_18018,N_17543,N_17891);
and U18019 (N_18019,N_17825,N_17806);
nand U18020 (N_18020,N_17883,N_17970);
xor U18021 (N_18021,N_17811,N_17940);
or U18022 (N_18022,N_17538,N_17822);
or U18023 (N_18023,N_17953,N_17872);
nor U18024 (N_18024,N_17606,N_17939);
xnor U18025 (N_18025,N_17810,N_17551);
and U18026 (N_18026,N_17963,N_17674);
nand U18027 (N_18027,N_17641,N_17898);
nand U18028 (N_18028,N_17914,N_17896);
or U18029 (N_18029,N_17852,N_17735);
nand U18030 (N_18030,N_17514,N_17612);
and U18031 (N_18031,N_17808,N_17794);
and U18032 (N_18032,N_17907,N_17677);
or U18033 (N_18033,N_17733,N_17755);
nor U18034 (N_18034,N_17642,N_17704);
and U18035 (N_18035,N_17645,N_17519);
or U18036 (N_18036,N_17936,N_17785);
nor U18037 (N_18037,N_17887,N_17574);
or U18038 (N_18038,N_17540,N_17873);
or U18039 (N_18039,N_17548,N_17536);
and U18040 (N_18040,N_17602,N_17816);
and U18041 (N_18041,N_17868,N_17839);
and U18042 (N_18042,N_17870,N_17959);
nor U18043 (N_18043,N_17503,N_17636);
or U18044 (N_18044,N_17997,N_17788);
and U18045 (N_18045,N_17618,N_17964);
nor U18046 (N_18046,N_17706,N_17643);
and U18047 (N_18047,N_17966,N_17848);
nor U18048 (N_18048,N_17805,N_17798);
nand U18049 (N_18049,N_17754,N_17687);
or U18050 (N_18050,N_17931,N_17784);
nor U18051 (N_18051,N_17520,N_17975);
nor U18052 (N_18052,N_17571,N_17524);
and U18053 (N_18053,N_17680,N_17599);
or U18054 (N_18054,N_17669,N_17851);
nor U18055 (N_18055,N_17671,N_17594);
nor U18056 (N_18056,N_17889,N_17841);
or U18057 (N_18057,N_17617,N_17682);
or U18058 (N_18058,N_17561,N_17728);
or U18059 (N_18059,N_17661,N_17732);
and U18060 (N_18060,N_17766,N_17570);
xor U18061 (N_18061,N_17830,N_17588);
nand U18062 (N_18062,N_17779,N_17933);
and U18063 (N_18063,N_17879,N_17869);
and U18064 (N_18064,N_17718,N_17526);
or U18065 (N_18065,N_17619,N_17532);
and U18066 (N_18066,N_17700,N_17566);
and U18067 (N_18067,N_17917,N_17653);
nor U18068 (N_18068,N_17972,N_17648);
nor U18069 (N_18069,N_17938,N_17991);
nor U18070 (N_18070,N_17818,N_17545);
nand U18071 (N_18071,N_17862,N_17590);
and U18072 (N_18072,N_17791,N_17683);
and U18073 (N_18073,N_17707,N_17668);
nor U18074 (N_18074,N_17659,N_17639);
nand U18075 (N_18075,N_17880,N_17552);
nor U18076 (N_18076,N_17899,N_17723);
and U18077 (N_18077,N_17840,N_17712);
xnor U18078 (N_18078,N_17751,N_17738);
nand U18079 (N_18079,N_17729,N_17650);
and U18080 (N_18080,N_17500,N_17627);
or U18081 (N_18081,N_17861,N_17748);
or U18082 (N_18082,N_17736,N_17695);
nand U18083 (N_18083,N_17821,N_17507);
and U18084 (N_18084,N_17854,N_17947);
or U18085 (N_18085,N_17663,N_17672);
and U18086 (N_18086,N_17592,N_17937);
nand U18087 (N_18087,N_17874,N_17813);
nand U18088 (N_18088,N_17760,N_17960);
nor U18089 (N_18089,N_17859,N_17579);
or U18090 (N_18090,N_17774,N_17757);
or U18091 (N_18091,N_17787,N_17903);
nand U18092 (N_18092,N_17789,N_17587);
or U18093 (N_18093,N_17812,N_17844);
nand U18094 (N_18094,N_17709,N_17591);
and U18095 (N_18095,N_17995,N_17958);
nand U18096 (N_18096,N_17752,N_17842);
and U18097 (N_18097,N_17781,N_17901);
or U18098 (N_18098,N_17716,N_17982);
and U18099 (N_18099,N_17885,N_17795);
nor U18100 (N_18100,N_17525,N_17527);
and U18101 (N_18101,N_17858,N_17780);
nor U18102 (N_18102,N_17616,N_17656);
or U18103 (N_18103,N_17511,N_17932);
nor U18104 (N_18104,N_17604,N_17989);
nand U18105 (N_18105,N_17853,N_17913);
and U18106 (N_18106,N_17831,N_17739);
nand U18107 (N_18107,N_17568,N_17589);
or U18108 (N_18108,N_17586,N_17513);
and U18109 (N_18109,N_17578,N_17686);
nor U18110 (N_18110,N_17928,N_17814);
and U18111 (N_18111,N_17908,N_17544);
nand U18112 (N_18112,N_17768,N_17703);
nand U18113 (N_18113,N_17542,N_17534);
nand U18114 (N_18114,N_17771,N_17973);
nor U18115 (N_18115,N_17775,N_17782);
nor U18116 (N_18116,N_17807,N_17644);
and U18117 (N_18117,N_17943,N_17691);
nand U18118 (N_18118,N_17727,N_17895);
nor U18119 (N_18119,N_17762,N_17922);
nand U18120 (N_18120,N_17847,N_17567);
or U18121 (N_18121,N_17793,N_17881);
nand U18122 (N_18122,N_17750,N_17621);
nor U18123 (N_18123,N_17944,N_17863);
and U18124 (N_18124,N_17918,N_17849);
and U18125 (N_18125,N_17976,N_17925);
nor U18126 (N_18126,N_17530,N_17804);
and U18127 (N_18127,N_17611,N_17633);
and U18128 (N_18128,N_17778,N_17977);
or U18129 (N_18129,N_17670,N_17609);
or U18130 (N_18130,N_17662,N_17523);
nor U18131 (N_18131,N_17572,N_17710);
and U18132 (N_18132,N_17508,N_17776);
and U18133 (N_18133,N_17559,N_17877);
and U18134 (N_18134,N_17585,N_17876);
nand U18135 (N_18135,N_17528,N_17535);
nand U18136 (N_18136,N_17846,N_17580);
or U18137 (N_18137,N_17769,N_17819);
nor U18138 (N_18138,N_17773,N_17603);
and U18139 (N_18139,N_17509,N_17660);
or U18140 (N_18140,N_17665,N_17721);
and U18141 (N_18141,N_17927,N_17745);
and U18142 (N_18142,N_17517,N_17607);
or U18143 (N_18143,N_17613,N_17546);
and U18144 (N_18144,N_17838,N_17878);
nand U18145 (N_18145,N_17749,N_17950);
and U18146 (N_18146,N_17817,N_17630);
nand U18147 (N_18147,N_17921,N_17558);
or U18148 (N_18148,N_17857,N_17713);
nor U18149 (N_18149,N_17676,N_17725);
nand U18150 (N_18150,N_17951,N_17505);
or U18151 (N_18151,N_17930,N_17957);
or U18152 (N_18152,N_17985,N_17850);
nand U18153 (N_18153,N_17595,N_17608);
or U18154 (N_18154,N_17549,N_17833);
or U18155 (N_18155,N_17990,N_17614);
nand U18156 (N_18156,N_17689,N_17967);
or U18157 (N_18157,N_17888,N_17598);
nand U18158 (N_18158,N_17702,N_17563);
and U18159 (N_18159,N_17890,N_17577);
nor U18160 (N_18160,N_17770,N_17583);
nor U18161 (N_18161,N_17634,N_17971);
nand U18162 (N_18162,N_17945,N_17553);
and U18163 (N_18163,N_17845,N_17946);
nand U18164 (N_18164,N_17919,N_17912);
or U18165 (N_18165,N_17726,N_17777);
or U18166 (N_18166,N_17765,N_17988);
nand U18167 (N_18167,N_17601,N_17693);
nor U18168 (N_18168,N_17620,N_17655);
and U18169 (N_18169,N_17911,N_17694);
or U18170 (N_18170,N_17832,N_17843);
or U18171 (N_18171,N_17623,N_17799);
nor U18172 (N_18172,N_17910,N_17664);
and U18173 (N_18173,N_17756,N_17564);
and U18174 (N_18174,N_17993,N_17600);
or U18175 (N_18175,N_17699,N_17666);
or U18176 (N_18176,N_17741,N_17685);
and U18177 (N_18177,N_17904,N_17893);
or U18178 (N_18178,N_17605,N_17892);
nor U18179 (N_18179,N_17698,N_17987);
and U18180 (N_18180,N_17941,N_17929);
or U18181 (N_18181,N_17675,N_17550);
or U18182 (N_18182,N_17955,N_17565);
nor U18183 (N_18183,N_17984,N_17961);
nor U18184 (N_18184,N_17701,N_17581);
and U18185 (N_18185,N_17688,N_17518);
or U18186 (N_18186,N_17696,N_17681);
and U18187 (N_18187,N_17596,N_17974);
and U18188 (N_18188,N_17835,N_17935);
nor U18189 (N_18189,N_17746,N_17510);
or U18190 (N_18190,N_17954,N_17555);
nand U18191 (N_18191,N_17826,N_17516);
nor U18192 (N_18192,N_17593,N_17753);
nand U18193 (N_18193,N_17690,N_17720);
xnor U18194 (N_18194,N_17836,N_17560);
nor U18195 (N_18195,N_17999,N_17562);
or U18196 (N_18196,N_17575,N_17502);
nor U18197 (N_18197,N_17827,N_17864);
and U18198 (N_18198,N_17692,N_17740);
and U18199 (N_18199,N_17969,N_17926);
xor U18200 (N_18200,N_17992,N_17824);
and U18201 (N_18201,N_17978,N_17533);
and U18202 (N_18202,N_17537,N_17800);
or U18203 (N_18203,N_17717,N_17708);
nand U18204 (N_18204,N_17867,N_17923);
nand U18205 (N_18205,N_17796,N_17998);
or U18206 (N_18206,N_17980,N_17920);
nand U18207 (N_18207,N_17801,N_17994);
nor U18208 (N_18208,N_17886,N_17547);
or U18209 (N_18209,N_17815,N_17678);
nand U18210 (N_18210,N_17759,N_17576);
nand U18211 (N_18211,N_17638,N_17522);
and U18212 (N_18212,N_17996,N_17790);
nand U18213 (N_18213,N_17557,N_17981);
and U18214 (N_18214,N_17829,N_17724);
nor U18215 (N_18215,N_17802,N_17823);
xor U18216 (N_18216,N_17747,N_17632);
nand U18217 (N_18217,N_17744,N_17764);
or U18218 (N_18218,N_17651,N_17905);
nand U18219 (N_18219,N_17531,N_17742);
nor U18220 (N_18220,N_17631,N_17916);
or U18221 (N_18221,N_17652,N_17948);
nand U18222 (N_18222,N_17786,N_17640);
nand U18223 (N_18223,N_17956,N_17865);
nand U18224 (N_18224,N_17515,N_17711);
or U18225 (N_18225,N_17731,N_17934);
nor U18226 (N_18226,N_17820,N_17983);
nor U18227 (N_18227,N_17986,N_17637);
nor U18228 (N_18228,N_17556,N_17897);
and U18229 (N_18229,N_17828,N_17582);
or U18230 (N_18230,N_17809,N_17569);
or U18231 (N_18231,N_17882,N_17909);
nor U18232 (N_18232,N_17541,N_17649);
and U18233 (N_18233,N_17792,N_17657);
and U18234 (N_18234,N_17625,N_17772);
or U18235 (N_18235,N_17501,N_17884);
nand U18236 (N_18236,N_17968,N_17658);
or U18237 (N_18237,N_17597,N_17628);
or U18238 (N_18238,N_17715,N_17902);
nand U18239 (N_18239,N_17512,N_17906);
xor U18240 (N_18240,N_17624,N_17803);
nand U18241 (N_18241,N_17949,N_17737);
and U18242 (N_18242,N_17767,N_17797);
and U18243 (N_18243,N_17629,N_17667);
nor U18244 (N_18244,N_17504,N_17894);
and U18245 (N_18245,N_17719,N_17866);
nand U18246 (N_18246,N_17679,N_17834);
and U18247 (N_18247,N_17705,N_17915);
nand U18248 (N_18248,N_17743,N_17573);
xnor U18249 (N_18249,N_17734,N_17761);
and U18250 (N_18250,N_17865,N_17694);
and U18251 (N_18251,N_17591,N_17726);
and U18252 (N_18252,N_17949,N_17819);
or U18253 (N_18253,N_17601,N_17604);
and U18254 (N_18254,N_17563,N_17673);
or U18255 (N_18255,N_17540,N_17557);
nor U18256 (N_18256,N_17811,N_17886);
nor U18257 (N_18257,N_17868,N_17942);
nor U18258 (N_18258,N_17600,N_17512);
or U18259 (N_18259,N_17800,N_17613);
nand U18260 (N_18260,N_17582,N_17818);
and U18261 (N_18261,N_17829,N_17590);
or U18262 (N_18262,N_17853,N_17530);
and U18263 (N_18263,N_17723,N_17678);
nand U18264 (N_18264,N_17706,N_17740);
and U18265 (N_18265,N_17506,N_17924);
nand U18266 (N_18266,N_17881,N_17544);
or U18267 (N_18267,N_17561,N_17888);
xnor U18268 (N_18268,N_17709,N_17527);
nand U18269 (N_18269,N_17996,N_17757);
nor U18270 (N_18270,N_17722,N_17810);
or U18271 (N_18271,N_17915,N_17653);
nand U18272 (N_18272,N_17976,N_17922);
nand U18273 (N_18273,N_17693,N_17985);
or U18274 (N_18274,N_17741,N_17682);
nor U18275 (N_18275,N_17555,N_17972);
nor U18276 (N_18276,N_17924,N_17699);
nand U18277 (N_18277,N_17608,N_17562);
and U18278 (N_18278,N_17842,N_17899);
xnor U18279 (N_18279,N_17512,N_17752);
nand U18280 (N_18280,N_17977,N_17667);
nor U18281 (N_18281,N_17508,N_17920);
or U18282 (N_18282,N_17598,N_17536);
nand U18283 (N_18283,N_17627,N_17932);
or U18284 (N_18284,N_17959,N_17614);
or U18285 (N_18285,N_17935,N_17797);
nor U18286 (N_18286,N_17831,N_17755);
or U18287 (N_18287,N_17609,N_17595);
nand U18288 (N_18288,N_17888,N_17630);
nor U18289 (N_18289,N_17625,N_17909);
or U18290 (N_18290,N_17812,N_17673);
nand U18291 (N_18291,N_17678,N_17840);
and U18292 (N_18292,N_17658,N_17678);
and U18293 (N_18293,N_17847,N_17621);
or U18294 (N_18294,N_17968,N_17595);
and U18295 (N_18295,N_17503,N_17612);
xnor U18296 (N_18296,N_17854,N_17531);
and U18297 (N_18297,N_17760,N_17502);
nor U18298 (N_18298,N_17736,N_17613);
or U18299 (N_18299,N_17504,N_17960);
nor U18300 (N_18300,N_17807,N_17716);
or U18301 (N_18301,N_17581,N_17845);
nor U18302 (N_18302,N_17628,N_17519);
nand U18303 (N_18303,N_17969,N_17837);
or U18304 (N_18304,N_17569,N_17852);
or U18305 (N_18305,N_17543,N_17673);
nand U18306 (N_18306,N_17937,N_17916);
or U18307 (N_18307,N_17645,N_17832);
nand U18308 (N_18308,N_17618,N_17707);
nor U18309 (N_18309,N_17832,N_17745);
or U18310 (N_18310,N_17707,N_17660);
nand U18311 (N_18311,N_17932,N_17531);
or U18312 (N_18312,N_17965,N_17941);
or U18313 (N_18313,N_17740,N_17863);
nand U18314 (N_18314,N_17877,N_17911);
nor U18315 (N_18315,N_17706,N_17789);
or U18316 (N_18316,N_17915,N_17767);
or U18317 (N_18317,N_17899,N_17705);
nand U18318 (N_18318,N_17940,N_17531);
nor U18319 (N_18319,N_17582,N_17957);
or U18320 (N_18320,N_17997,N_17922);
and U18321 (N_18321,N_17807,N_17704);
and U18322 (N_18322,N_17501,N_17823);
nor U18323 (N_18323,N_17806,N_17997);
or U18324 (N_18324,N_17613,N_17607);
and U18325 (N_18325,N_17578,N_17667);
nor U18326 (N_18326,N_17580,N_17548);
nand U18327 (N_18327,N_17744,N_17545);
and U18328 (N_18328,N_17583,N_17799);
or U18329 (N_18329,N_17884,N_17563);
and U18330 (N_18330,N_17563,N_17959);
or U18331 (N_18331,N_17528,N_17975);
and U18332 (N_18332,N_17535,N_17917);
nor U18333 (N_18333,N_17933,N_17620);
nand U18334 (N_18334,N_17692,N_17661);
and U18335 (N_18335,N_17935,N_17890);
nand U18336 (N_18336,N_17676,N_17986);
nor U18337 (N_18337,N_17602,N_17954);
nor U18338 (N_18338,N_17766,N_17921);
nand U18339 (N_18339,N_17555,N_17615);
or U18340 (N_18340,N_17910,N_17788);
xor U18341 (N_18341,N_17803,N_17656);
nand U18342 (N_18342,N_17979,N_17554);
nand U18343 (N_18343,N_17579,N_17640);
or U18344 (N_18344,N_17604,N_17577);
nand U18345 (N_18345,N_17776,N_17553);
nor U18346 (N_18346,N_17601,N_17598);
nand U18347 (N_18347,N_17923,N_17763);
nor U18348 (N_18348,N_17736,N_17842);
or U18349 (N_18349,N_17865,N_17671);
or U18350 (N_18350,N_17800,N_17502);
nand U18351 (N_18351,N_17987,N_17695);
nor U18352 (N_18352,N_17948,N_17620);
nand U18353 (N_18353,N_17809,N_17851);
or U18354 (N_18354,N_17740,N_17624);
or U18355 (N_18355,N_17811,N_17561);
or U18356 (N_18356,N_17917,N_17512);
and U18357 (N_18357,N_17656,N_17669);
or U18358 (N_18358,N_17680,N_17792);
or U18359 (N_18359,N_17821,N_17765);
and U18360 (N_18360,N_17845,N_17851);
or U18361 (N_18361,N_17841,N_17871);
and U18362 (N_18362,N_17872,N_17977);
and U18363 (N_18363,N_17934,N_17581);
nor U18364 (N_18364,N_17788,N_17730);
nand U18365 (N_18365,N_17821,N_17651);
nor U18366 (N_18366,N_17523,N_17982);
nor U18367 (N_18367,N_17875,N_17996);
and U18368 (N_18368,N_17870,N_17869);
or U18369 (N_18369,N_17902,N_17913);
nand U18370 (N_18370,N_17722,N_17863);
nand U18371 (N_18371,N_17701,N_17578);
nor U18372 (N_18372,N_17851,N_17711);
and U18373 (N_18373,N_17766,N_17572);
nor U18374 (N_18374,N_17817,N_17852);
and U18375 (N_18375,N_17841,N_17610);
nor U18376 (N_18376,N_17646,N_17845);
and U18377 (N_18377,N_17506,N_17888);
or U18378 (N_18378,N_17680,N_17566);
or U18379 (N_18379,N_17901,N_17515);
and U18380 (N_18380,N_17644,N_17811);
or U18381 (N_18381,N_17726,N_17886);
or U18382 (N_18382,N_17715,N_17916);
nor U18383 (N_18383,N_17790,N_17574);
or U18384 (N_18384,N_17579,N_17869);
nand U18385 (N_18385,N_17970,N_17943);
nand U18386 (N_18386,N_17784,N_17792);
nand U18387 (N_18387,N_17870,N_17700);
or U18388 (N_18388,N_17866,N_17705);
nand U18389 (N_18389,N_17749,N_17916);
nand U18390 (N_18390,N_17699,N_17909);
nor U18391 (N_18391,N_17624,N_17688);
nor U18392 (N_18392,N_17567,N_17884);
or U18393 (N_18393,N_17974,N_17542);
and U18394 (N_18394,N_17867,N_17684);
and U18395 (N_18395,N_17547,N_17695);
nor U18396 (N_18396,N_17601,N_17611);
and U18397 (N_18397,N_17889,N_17661);
or U18398 (N_18398,N_17759,N_17832);
or U18399 (N_18399,N_17779,N_17822);
nand U18400 (N_18400,N_17826,N_17525);
nor U18401 (N_18401,N_17957,N_17768);
nor U18402 (N_18402,N_17827,N_17998);
nor U18403 (N_18403,N_17636,N_17765);
nor U18404 (N_18404,N_17665,N_17511);
and U18405 (N_18405,N_17617,N_17797);
nor U18406 (N_18406,N_17733,N_17585);
nor U18407 (N_18407,N_17857,N_17994);
or U18408 (N_18408,N_17783,N_17684);
or U18409 (N_18409,N_17702,N_17788);
or U18410 (N_18410,N_17930,N_17810);
and U18411 (N_18411,N_17898,N_17796);
or U18412 (N_18412,N_17510,N_17625);
nor U18413 (N_18413,N_17819,N_17501);
and U18414 (N_18414,N_17743,N_17547);
or U18415 (N_18415,N_17629,N_17943);
nor U18416 (N_18416,N_17542,N_17729);
or U18417 (N_18417,N_17876,N_17598);
or U18418 (N_18418,N_17831,N_17933);
nor U18419 (N_18419,N_17737,N_17873);
or U18420 (N_18420,N_17859,N_17668);
nand U18421 (N_18421,N_17948,N_17964);
and U18422 (N_18422,N_17530,N_17857);
nor U18423 (N_18423,N_17708,N_17880);
nor U18424 (N_18424,N_17543,N_17634);
nor U18425 (N_18425,N_17902,N_17806);
or U18426 (N_18426,N_17710,N_17638);
or U18427 (N_18427,N_17984,N_17752);
or U18428 (N_18428,N_17948,N_17722);
nand U18429 (N_18429,N_17796,N_17517);
nand U18430 (N_18430,N_17898,N_17786);
nand U18431 (N_18431,N_17860,N_17631);
nor U18432 (N_18432,N_17651,N_17817);
nand U18433 (N_18433,N_17528,N_17611);
and U18434 (N_18434,N_17888,N_17986);
nor U18435 (N_18435,N_17930,N_17615);
nor U18436 (N_18436,N_17879,N_17589);
or U18437 (N_18437,N_17505,N_17548);
or U18438 (N_18438,N_17779,N_17550);
nor U18439 (N_18439,N_17831,N_17662);
or U18440 (N_18440,N_17839,N_17580);
and U18441 (N_18441,N_17608,N_17812);
nor U18442 (N_18442,N_17736,N_17679);
nor U18443 (N_18443,N_17589,N_17751);
nor U18444 (N_18444,N_17806,N_17941);
and U18445 (N_18445,N_17837,N_17710);
nor U18446 (N_18446,N_17731,N_17680);
or U18447 (N_18447,N_17720,N_17643);
and U18448 (N_18448,N_17886,N_17737);
and U18449 (N_18449,N_17816,N_17856);
and U18450 (N_18450,N_17991,N_17687);
nor U18451 (N_18451,N_17552,N_17820);
nor U18452 (N_18452,N_17871,N_17522);
or U18453 (N_18453,N_17964,N_17665);
xnor U18454 (N_18454,N_17824,N_17619);
nand U18455 (N_18455,N_17710,N_17897);
nand U18456 (N_18456,N_17910,N_17613);
nor U18457 (N_18457,N_17673,N_17500);
nor U18458 (N_18458,N_17666,N_17776);
and U18459 (N_18459,N_17598,N_17725);
nand U18460 (N_18460,N_17754,N_17677);
or U18461 (N_18461,N_17705,N_17968);
or U18462 (N_18462,N_17583,N_17800);
nand U18463 (N_18463,N_17931,N_17513);
or U18464 (N_18464,N_17530,N_17861);
nand U18465 (N_18465,N_17650,N_17891);
and U18466 (N_18466,N_17797,N_17782);
and U18467 (N_18467,N_17583,N_17632);
nand U18468 (N_18468,N_17569,N_17667);
nand U18469 (N_18469,N_17884,N_17801);
or U18470 (N_18470,N_17564,N_17969);
or U18471 (N_18471,N_17683,N_17634);
nand U18472 (N_18472,N_17617,N_17536);
and U18473 (N_18473,N_17866,N_17758);
nand U18474 (N_18474,N_17790,N_17837);
nand U18475 (N_18475,N_17793,N_17707);
or U18476 (N_18476,N_17894,N_17557);
nor U18477 (N_18477,N_17720,N_17896);
and U18478 (N_18478,N_17813,N_17508);
nand U18479 (N_18479,N_17738,N_17861);
nor U18480 (N_18480,N_17977,N_17583);
xor U18481 (N_18481,N_17783,N_17582);
and U18482 (N_18482,N_17542,N_17838);
nor U18483 (N_18483,N_17731,N_17864);
or U18484 (N_18484,N_17596,N_17793);
and U18485 (N_18485,N_17950,N_17719);
and U18486 (N_18486,N_17720,N_17911);
nor U18487 (N_18487,N_17509,N_17770);
nor U18488 (N_18488,N_17607,N_17822);
nand U18489 (N_18489,N_17506,N_17711);
or U18490 (N_18490,N_17974,N_17614);
nand U18491 (N_18491,N_17635,N_17846);
and U18492 (N_18492,N_17917,N_17962);
and U18493 (N_18493,N_17525,N_17896);
and U18494 (N_18494,N_17737,N_17938);
or U18495 (N_18495,N_17655,N_17887);
and U18496 (N_18496,N_17678,N_17637);
nand U18497 (N_18497,N_17809,N_17807);
nor U18498 (N_18498,N_17699,N_17713);
and U18499 (N_18499,N_17925,N_17790);
or U18500 (N_18500,N_18138,N_18338);
or U18501 (N_18501,N_18284,N_18375);
or U18502 (N_18502,N_18341,N_18012);
nand U18503 (N_18503,N_18156,N_18494);
and U18504 (N_18504,N_18498,N_18277);
nor U18505 (N_18505,N_18109,N_18293);
or U18506 (N_18506,N_18459,N_18419);
nor U18507 (N_18507,N_18401,N_18060);
nor U18508 (N_18508,N_18052,N_18224);
nand U18509 (N_18509,N_18182,N_18235);
or U18510 (N_18510,N_18145,N_18026);
or U18511 (N_18511,N_18171,N_18003);
and U18512 (N_18512,N_18472,N_18349);
and U18513 (N_18513,N_18080,N_18385);
or U18514 (N_18514,N_18257,N_18131);
nor U18515 (N_18515,N_18312,N_18367);
and U18516 (N_18516,N_18247,N_18076);
and U18517 (N_18517,N_18212,N_18017);
nand U18518 (N_18518,N_18057,N_18326);
or U18519 (N_18519,N_18451,N_18369);
nand U18520 (N_18520,N_18380,N_18322);
or U18521 (N_18521,N_18496,N_18086);
nor U18522 (N_18522,N_18254,N_18155);
or U18523 (N_18523,N_18475,N_18409);
and U18524 (N_18524,N_18105,N_18097);
nand U18525 (N_18525,N_18303,N_18337);
xor U18526 (N_18526,N_18191,N_18243);
and U18527 (N_18527,N_18092,N_18177);
or U18528 (N_18528,N_18455,N_18088);
nor U18529 (N_18529,N_18020,N_18393);
xor U18530 (N_18530,N_18067,N_18485);
or U18531 (N_18531,N_18445,N_18468);
nand U18532 (N_18532,N_18222,N_18002);
xnor U18533 (N_18533,N_18272,N_18311);
or U18534 (N_18534,N_18252,N_18169);
and U18535 (N_18535,N_18175,N_18047);
and U18536 (N_18536,N_18343,N_18208);
nand U18537 (N_18537,N_18362,N_18134);
or U18538 (N_18538,N_18411,N_18195);
and U18539 (N_18539,N_18050,N_18116);
nor U18540 (N_18540,N_18123,N_18150);
or U18541 (N_18541,N_18427,N_18416);
nand U18542 (N_18542,N_18495,N_18351);
nand U18543 (N_18543,N_18245,N_18077);
nand U18544 (N_18544,N_18137,N_18009);
and U18545 (N_18545,N_18096,N_18314);
and U18546 (N_18546,N_18049,N_18454);
nor U18547 (N_18547,N_18068,N_18471);
or U18548 (N_18548,N_18377,N_18296);
or U18549 (N_18549,N_18480,N_18347);
xor U18550 (N_18550,N_18093,N_18011);
or U18551 (N_18551,N_18373,N_18233);
nand U18552 (N_18552,N_18364,N_18108);
and U18553 (N_18553,N_18430,N_18408);
nor U18554 (N_18554,N_18227,N_18414);
or U18555 (N_18555,N_18170,N_18216);
nor U18556 (N_18556,N_18280,N_18446);
or U18557 (N_18557,N_18354,N_18128);
nor U18558 (N_18558,N_18213,N_18388);
nor U18559 (N_18559,N_18164,N_18141);
or U18560 (N_18560,N_18042,N_18033);
or U18561 (N_18561,N_18100,N_18319);
or U18562 (N_18562,N_18074,N_18342);
nor U18563 (N_18563,N_18111,N_18196);
nand U18564 (N_18564,N_18114,N_18434);
nor U18565 (N_18565,N_18163,N_18010);
or U18566 (N_18566,N_18199,N_18263);
and U18567 (N_18567,N_18302,N_18365);
nor U18568 (N_18568,N_18313,N_18479);
nand U18569 (N_18569,N_18300,N_18045);
and U18570 (N_18570,N_18439,N_18465);
nor U18571 (N_18571,N_18307,N_18085);
and U18572 (N_18572,N_18028,N_18335);
nand U18573 (N_18573,N_18087,N_18320);
and U18574 (N_18574,N_18442,N_18053);
or U18575 (N_18575,N_18112,N_18464);
nor U18576 (N_18576,N_18133,N_18197);
nand U18577 (N_18577,N_18019,N_18031);
nor U18578 (N_18578,N_18330,N_18237);
nor U18579 (N_18579,N_18417,N_18265);
nor U18580 (N_18580,N_18168,N_18415);
or U18581 (N_18581,N_18201,N_18161);
and U18582 (N_18582,N_18249,N_18378);
nor U18583 (N_18583,N_18066,N_18036);
xnor U18584 (N_18584,N_18463,N_18406);
nand U18585 (N_18585,N_18046,N_18497);
xor U18586 (N_18586,N_18193,N_18298);
nand U18587 (N_18587,N_18228,N_18038);
nor U18588 (N_18588,N_18054,N_18185);
nor U18589 (N_18589,N_18437,N_18321);
or U18590 (N_18590,N_18309,N_18223);
nand U18591 (N_18591,N_18005,N_18402);
nor U18592 (N_18592,N_18207,N_18062);
nor U18593 (N_18593,N_18259,N_18018);
nor U18594 (N_18594,N_18355,N_18352);
nor U18595 (N_18595,N_18460,N_18368);
nand U18596 (N_18596,N_18014,N_18157);
xor U18597 (N_18597,N_18139,N_18147);
nand U18598 (N_18598,N_18172,N_18332);
or U18599 (N_18599,N_18246,N_18395);
or U18600 (N_18600,N_18240,N_18482);
or U18601 (N_18601,N_18366,N_18048);
or U18602 (N_18602,N_18275,N_18144);
and U18603 (N_18603,N_18236,N_18413);
or U18604 (N_18604,N_18301,N_18381);
xnor U18605 (N_18605,N_18359,N_18435);
or U18606 (N_18606,N_18032,N_18113);
and U18607 (N_18607,N_18219,N_18286);
nand U18608 (N_18608,N_18059,N_18187);
nand U18609 (N_18609,N_18452,N_18090);
and U18610 (N_18610,N_18082,N_18271);
nand U18611 (N_18611,N_18394,N_18044);
nor U18612 (N_18612,N_18262,N_18340);
nor U18613 (N_18613,N_18421,N_18440);
nand U18614 (N_18614,N_18357,N_18239);
nor U18615 (N_18615,N_18418,N_18013);
or U18616 (N_18616,N_18238,N_18397);
nor U18617 (N_18617,N_18021,N_18390);
nor U18618 (N_18618,N_18255,N_18391);
nor U18619 (N_18619,N_18318,N_18361);
and U18620 (N_18620,N_18091,N_18499);
nand U18621 (N_18621,N_18190,N_18306);
and U18622 (N_18622,N_18467,N_18292);
and U18623 (N_18623,N_18165,N_18051);
nor U18624 (N_18624,N_18407,N_18488);
or U18625 (N_18625,N_18225,N_18140);
nor U18626 (N_18626,N_18184,N_18457);
and U18627 (N_18627,N_18215,N_18094);
nor U18628 (N_18628,N_18030,N_18299);
nand U18629 (N_18629,N_18015,N_18022);
and U18630 (N_18630,N_18428,N_18220);
nand U18631 (N_18631,N_18403,N_18120);
and U18632 (N_18632,N_18056,N_18205);
nor U18633 (N_18633,N_18198,N_18078);
or U18634 (N_18634,N_18115,N_18104);
or U18635 (N_18635,N_18221,N_18143);
nand U18636 (N_18636,N_18248,N_18095);
nand U18637 (N_18637,N_18055,N_18040);
and U18638 (N_18638,N_18209,N_18192);
nor U18639 (N_18639,N_18029,N_18304);
or U18640 (N_18640,N_18079,N_18106);
and U18641 (N_18641,N_18382,N_18126);
and U18642 (N_18642,N_18350,N_18334);
xor U18643 (N_18643,N_18136,N_18173);
or U18644 (N_18644,N_18167,N_18160);
or U18645 (N_18645,N_18384,N_18204);
nand U18646 (N_18646,N_18426,N_18436);
or U18647 (N_18647,N_18148,N_18324);
nand U18648 (N_18648,N_18258,N_18176);
nor U18649 (N_18649,N_18308,N_18400);
nand U18650 (N_18650,N_18289,N_18478);
nand U18651 (N_18651,N_18069,N_18461);
or U18652 (N_18652,N_18230,N_18449);
or U18653 (N_18653,N_18273,N_18119);
nor U18654 (N_18654,N_18244,N_18423);
nand U18655 (N_18655,N_18462,N_18283);
or U18656 (N_18656,N_18486,N_18410);
or U18657 (N_18657,N_18389,N_18231);
nor U18658 (N_18658,N_18226,N_18004);
nor U18659 (N_18659,N_18285,N_18278);
nor U18660 (N_18660,N_18125,N_18360);
or U18661 (N_18661,N_18305,N_18450);
nor U18662 (N_18662,N_18064,N_18178);
and U18663 (N_18663,N_18251,N_18256);
or U18664 (N_18664,N_18466,N_18132);
and U18665 (N_18665,N_18039,N_18279);
nor U18666 (N_18666,N_18179,N_18072);
or U18667 (N_18667,N_18099,N_18058);
nand U18668 (N_18668,N_18084,N_18290);
and U18669 (N_18669,N_18061,N_18353);
nor U18670 (N_18670,N_18037,N_18102);
or U18671 (N_18671,N_18339,N_18081);
and U18672 (N_18672,N_18491,N_18431);
or U18673 (N_18673,N_18127,N_18316);
nor U18674 (N_18674,N_18276,N_18448);
or U18675 (N_18675,N_18383,N_18492);
and U18676 (N_18676,N_18281,N_18315);
and U18677 (N_18677,N_18270,N_18387);
and U18678 (N_18678,N_18124,N_18433);
nor U18679 (N_18679,N_18474,N_18098);
or U18680 (N_18680,N_18470,N_18035);
or U18681 (N_18681,N_18121,N_18000);
and U18682 (N_18682,N_18405,N_18432);
nor U18683 (N_18683,N_18396,N_18268);
nand U18684 (N_18684,N_18203,N_18158);
nor U18685 (N_18685,N_18107,N_18146);
or U18686 (N_18686,N_18376,N_18206);
and U18687 (N_18687,N_18260,N_18101);
nand U18688 (N_18688,N_18398,N_18386);
and U18689 (N_18689,N_18297,N_18487);
nand U18690 (N_18690,N_18149,N_18473);
and U18691 (N_18691,N_18476,N_18073);
and U18692 (N_18692,N_18372,N_18229);
nor U18693 (N_18693,N_18345,N_18489);
or U18694 (N_18694,N_18183,N_18288);
nor U18695 (N_18695,N_18186,N_18024);
nor U18696 (N_18696,N_18370,N_18008);
or U18697 (N_18697,N_18180,N_18135);
nor U18698 (N_18698,N_18202,N_18110);
nand U18699 (N_18699,N_18117,N_18174);
or U18700 (N_18700,N_18344,N_18034);
and U18701 (N_18701,N_18214,N_18118);
nor U18702 (N_18702,N_18453,N_18331);
and U18703 (N_18703,N_18328,N_18234);
or U18704 (N_18704,N_18065,N_18329);
or U18705 (N_18705,N_18481,N_18083);
nand U18706 (N_18706,N_18269,N_18159);
and U18707 (N_18707,N_18162,N_18379);
nand U18708 (N_18708,N_18122,N_18490);
nand U18709 (N_18709,N_18291,N_18264);
and U18710 (N_18710,N_18493,N_18404);
nand U18711 (N_18711,N_18189,N_18211);
nor U18712 (N_18712,N_18154,N_18142);
nand U18713 (N_18713,N_18089,N_18075);
or U18714 (N_18714,N_18358,N_18266);
nand U18715 (N_18715,N_18399,N_18210);
nor U18716 (N_18716,N_18027,N_18250);
or U18717 (N_18717,N_18438,N_18153);
nand U18718 (N_18718,N_18267,N_18310);
or U18719 (N_18719,N_18130,N_18441);
and U18720 (N_18720,N_18043,N_18295);
xor U18721 (N_18721,N_18484,N_18241);
or U18722 (N_18722,N_18242,N_18023);
nor U18723 (N_18723,N_18483,N_18103);
and U18724 (N_18724,N_18363,N_18333);
xor U18725 (N_18725,N_18007,N_18166);
nand U18726 (N_18726,N_18458,N_18129);
and U18727 (N_18727,N_18188,N_18477);
nand U18728 (N_18728,N_18261,N_18317);
and U18729 (N_18729,N_18336,N_18181);
and U18730 (N_18730,N_18217,N_18274);
nor U18731 (N_18731,N_18253,N_18447);
nand U18732 (N_18732,N_18282,N_18456);
nand U18733 (N_18733,N_18348,N_18041);
nor U18734 (N_18734,N_18194,N_18412);
nand U18735 (N_18735,N_18325,N_18327);
or U18736 (N_18736,N_18151,N_18232);
nor U18737 (N_18737,N_18016,N_18006);
nand U18738 (N_18738,N_18443,N_18200);
nor U18739 (N_18739,N_18323,N_18001);
and U18740 (N_18740,N_18420,N_18444);
and U18741 (N_18741,N_18218,N_18424);
and U18742 (N_18742,N_18025,N_18422);
or U18743 (N_18743,N_18063,N_18287);
nand U18744 (N_18744,N_18152,N_18429);
nor U18745 (N_18745,N_18294,N_18469);
nand U18746 (N_18746,N_18425,N_18356);
and U18747 (N_18747,N_18346,N_18392);
or U18748 (N_18748,N_18070,N_18374);
and U18749 (N_18749,N_18071,N_18371);
nand U18750 (N_18750,N_18143,N_18405);
and U18751 (N_18751,N_18135,N_18370);
or U18752 (N_18752,N_18315,N_18421);
and U18753 (N_18753,N_18393,N_18423);
nor U18754 (N_18754,N_18039,N_18004);
or U18755 (N_18755,N_18281,N_18010);
or U18756 (N_18756,N_18115,N_18455);
nor U18757 (N_18757,N_18138,N_18457);
or U18758 (N_18758,N_18175,N_18395);
and U18759 (N_18759,N_18044,N_18049);
nand U18760 (N_18760,N_18071,N_18268);
nor U18761 (N_18761,N_18164,N_18258);
or U18762 (N_18762,N_18473,N_18330);
nand U18763 (N_18763,N_18009,N_18437);
and U18764 (N_18764,N_18305,N_18358);
nor U18765 (N_18765,N_18431,N_18304);
nand U18766 (N_18766,N_18266,N_18110);
nand U18767 (N_18767,N_18358,N_18203);
nand U18768 (N_18768,N_18319,N_18259);
or U18769 (N_18769,N_18103,N_18325);
and U18770 (N_18770,N_18257,N_18223);
or U18771 (N_18771,N_18026,N_18250);
nand U18772 (N_18772,N_18234,N_18316);
and U18773 (N_18773,N_18443,N_18015);
or U18774 (N_18774,N_18295,N_18209);
and U18775 (N_18775,N_18360,N_18122);
and U18776 (N_18776,N_18150,N_18324);
nor U18777 (N_18777,N_18159,N_18158);
nand U18778 (N_18778,N_18141,N_18012);
or U18779 (N_18779,N_18051,N_18094);
or U18780 (N_18780,N_18205,N_18252);
nand U18781 (N_18781,N_18447,N_18042);
or U18782 (N_18782,N_18228,N_18245);
and U18783 (N_18783,N_18052,N_18223);
xor U18784 (N_18784,N_18488,N_18183);
nand U18785 (N_18785,N_18120,N_18337);
nor U18786 (N_18786,N_18494,N_18364);
and U18787 (N_18787,N_18322,N_18115);
nor U18788 (N_18788,N_18081,N_18131);
nand U18789 (N_18789,N_18393,N_18030);
and U18790 (N_18790,N_18257,N_18444);
nor U18791 (N_18791,N_18155,N_18382);
nor U18792 (N_18792,N_18352,N_18094);
nand U18793 (N_18793,N_18182,N_18422);
xor U18794 (N_18794,N_18403,N_18436);
and U18795 (N_18795,N_18226,N_18489);
or U18796 (N_18796,N_18020,N_18487);
and U18797 (N_18797,N_18478,N_18476);
xnor U18798 (N_18798,N_18377,N_18018);
or U18799 (N_18799,N_18366,N_18237);
nor U18800 (N_18800,N_18137,N_18235);
nand U18801 (N_18801,N_18233,N_18075);
and U18802 (N_18802,N_18169,N_18120);
nand U18803 (N_18803,N_18349,N_18015);
or U18804 (N_18804,N_18084,N_18294);
nor U18805 (N_18805,N_18292,N_18102);
and U18806 (N_18806,N_18202,N_18121);
or U18807 (N_18807,N_18406,N_18190);
and U18808 (N_18808,N_18239,N_18303);
nand U18809 (N_18809,N_18426,N_18296);
and U18810 (N_18810,N_18052,N_18255);
or U18811 (N_18811,N_18282,N_18412);
nand U18812 (N_18812,N_18147,N_18203);
or U18813 (N_18813,N_18291,N_18345);
nor U18814 (N_18814,N_18060,N_18416);
nand U18815 (N_18815,N_18156,N_18111);
and U18816 (N_18816,N_18045,N_18355);
or U18817 (N_18817,N_18296,N_18086);
or U18818 (N_18818,N_18496,N_18303);
and U18819 (N_18819,N_18190,N_18362);
nand U18820 (N_18820,N_18002,N_18188);
and U18821 (N_18821,N_18124,N_18409);
nor U18822 (N_18822,N_18097,N_18068);
nand U18823 (N_18823,N_18045,N_18396);
nor U18824 (N_18824,N_18228,N_18030);
nor U18825 (N_18825,N_18178,N_18024);
nor U18826 (N_18826,N_18006,N_18391);
or U18827 (N_18827,N_18292,N_18150);
nor U18828 (N_18828,N_18193,N_18350);
nor U18829 (N_18829,N_18251,N_18116);
xor U18830 (N_18830,N_18453,N_18477);
and U18831 (N_18831,N_18067,N_18192);
or U18832 (N_18832,N_18006,N_18440);
and U18833 (N_18833,N_18058,N_18476);
and U18834 (N_18834,N_18425,N_18290);
and U18835 (N_18835,N_18215,N_18052);
nor U18836 (N_18836,N_18284,N_18416);
and U18837 (N_18837,N_18264,N_18089);
and U18838 (N_18838,N_18080,N_18204);
and U18839 (N_18839,N_18441,N_18477);
or U18840 (N_18840,N_18178,N_18377);
or U18841 (N_18841,N_18295,N_18429);
nand U18842 (N_18842,N_18317,N_18311);
nand U18843 (N_18843,N_18307,N_18146);
or U18844 (N_18844,N_18022,N_18316);
and U18845 (N_18845,N_18099,N_18484);
and U18846 (N_18846,N_18105,N_18111);
or U18847 (N_18847,N_18419,N_18329);
xor U18848 (N_18848,N_18279,N_18455);
and U18849 (N_18849,N_18423,N_18198);
and U18850 (N_18850,N_18302,N_18374);
nand U18851 (N_18851,N_18460,N_18260);
nor U18852 (N_18852,N_18277,N_18428);
or U18853 (N_18853,N_18458,N_18372);
nand U18854 (N_18854,N_18464,N_18423);
nor U18855 (N_18855,N_18425,N_18379);
nand U18856 (N_18856,N_18052,N_18402);
and U18857 (N_18857,N_18234,N_18237);
or U18858 (N_18858,N_18468,N_18096);
or U18859 (N_18859,N_18015,N_18114);
or U18860 (N_18860,N_18119,N_18437);
or U18861 (N_18861,N_18314,N_18335);
nor U18862 (N_18862,N_18499,N_18362);
and U18863 (N_18863,N_18401,N_18081);
and U18864 (N_18864,N_18134,N_18233);
or U18865 (N_18865,N_18018,N_18318);
xor U18866 (N_18866,N_18465,N_18306);
nand U18867 (N_18867,N_18315,N_18055);
nor U18868 (N_18868,N_18367,N_18073);
nor U18869 (N_18869,N_18447,N_18474);
or U18870 (N_18870,N_18439,N_18331);
nor U18871 (N_18871,N_18420,N_18217);
nor U18872 (N_18872,N_18016,N_18075);
or U18873 (N_18873,N_18027,N_18425);
and U18874 (N_18874,N_18490,N_18103);
nor U18875 (N_18875,N_18155,N_18314);
and U18876 (N_18876,N_18101,N_18217);
or U18877 (N_18877,N_18373,N_18145);
and U18878 (N_18878,N_18436,N_18213);
and U18879 (N_18879,N_18182,N_18035);
or U18880 (N_18880,N_18320,N_18299);
nor U18881 (N_18881,N_18074,N_18338);
or U18882 (N_18882,N_18137,N_18350);
or U18883 (N_18883,N_18471,N_18444);
nand U18884 (N_18884,N_18439,N_18015);
nor U18885 (N_18885,N_18089,N_18160);
nand U18886 (N_18886,N_18485,N_18183);
and U18887 (N_18887,N_18240,N_18049);
nand U18888 (N_18888,N_18129,N_18210);
nor U18889 (N_18889,N_18396,N_18254);
nand U18890 (N_18890,N_18155,N_18128);
nor U18891 (N_18891,N_18489,N_18103);
and U18892 (N_18892,N_18440,N_18166);
nor U18893 (N_18893,N_18286,N_18178);
nor U18894 (N_18894,N_18471,N_18214);
nor U18895 (N_18895,N_18000,N_18082);
or U18896 (N_18896,N_18125,N_18458);
nor U18897 (N_18897,N_18235,N_18012);
or U18898 (N_18898,N_18032,N_18316);
or U18899 (N_18899,N_18106,N_18096);
and U18900 (N_18900,N_18281,N_18070);
or U18901 (N_18901,N_18142,N_18342);
and U18902 (N_18902,N_18398,N_18203);
and U18903 (N_18903,N_18415,N_18030);
nand U18904 (N_18904,N_18380,N_18143);
nor U18905 (N_18905,N_18115,N_18190);
nand U18906 (N_18906,N_18424,N_18422);
or U18907 (N_18907,N_18003,N_18433);
nor U18908 (N_18908,N_18071,N_18056);
nand U18909 (N_18909,N_18142,N_18049);
nor U18910 (N_18910,N_18165,N_18399);
or U18911 (N_18911,N_18076,N_18363);
nand U18912 (N_18912,N_18169,N_18314);
nor U18913 (N_18913,N_18316,N_18321);
or U18914 (N_18914,N_18147,N_18457);
nand U18915 (N_18915,N_18269,N_18151);
and U18916 (N_18916,N_18194,N_18012);
and U18917 (N_18917,N_18286,N_18461);
and U18918 (N_18918,N_18297,N_18187);
or U18919 (N_18919,N_18268,N_18370);
and U18920 (N_18920,N_18259,N_18403);
nand U18921 (N_18921,N_18151,N_18316);
nand U18922 (N_18922,N_18149,N_18073);
and U18923 (N_18923,N_18281,N_18191);
or U18924 (N_18924,N_18244,N_18087);
nand U18925 (N_18925,N_18198,N_18328);
nor U18926 (N_18926,N_18409,N_18444);
xor U18927 (N_18927,N_18149,N_18084);
or U18928 (N_18928,N_18367,N_18291);
or U18929 (N_18929,N_18115,N_18139);
and U18930 (N_18930,N_18339,N_18044);
and U18931 (N_18931,N_18224,N_18079);
nor U18932 (N_18932,N_18145,N_18462);
and U18933 (N_18933,N_18013,N_18358);
and U18934 (N_18934,N_18217,N_18374);
and U18935 (N_18935,N_18008,N_18321);
nor U18936 (N_18936,N_18187,N_18080);
nand U18937 (N_18937,N_18440,N_18376);
and U18938 (N_18938,N_18021,N_18057);
nor U18939 (N_18939,N_18108,N_18434);
nor U18940 (N_18940,N_18337,N_18172);
and U18941 (N_18941,N_18288,N_18261);
nor U18942 (N_18942,N_18370,N_18152);
nor U18943 (N_18943,N_18355,N_18382);
nor U18944 (N_18944,N_18422,N_18320);
nor U18945 (N_18945,N_18078,N_18437);
xor U18946 (N_18946,N_18143,N_18268);
nand U18947 (N_18947,N_18072,N_18357);
and U18948 (N_18948,N_18254,N_18382);
nand U18949 (N_18949,N_18109,N_18309);
nor U18950 (N_18950,N_18268,N_18044);
nand U18951 (N_18951,N_18085,N_18156);
or U18952 (N_18952,N_18098,N_18475);
nor U18953 (N_18953,N_18410,N_18203);
and U18954 (N_18954,N_18462,N_18230);
nor U18955 (N_18955,N_18420,N_18421);
nand U18956 (N_18956,N_18139,N_18404);
and U18957 (N_18957,N_18101,N_18171);
nor U18958 (N_18958,N_18405,N_18406);
and U18959 (N_18959,N_18486,N_18286);
nor U18960 (N_18960,N_18048,N_18020);
nand U18961 (N_18961,N_18024,N_18268);
and U18962 (N_18962,N_18326,N_18291);
nor U18963 (N_18963,N_18151,N_18184);
or U18964 (N_18964,N_18185,N_18058);
or U18965 (N_18965,N_18016,N_18278);
or U18966 (N_18966,N_18125,N_18023);
or U18967 (N_18967,N_18077,N_18112);
nand U18968 (N_18968,N_18461,N_18314);
and U18969 (N_18969,N_18141,N_18132);
xnor U18970 (N_18970,N_18357,N_18020);
nor U18971 (N_18971,N_18029,N_18084);
or U18972 (N_18972,N_18289,N_18204);
and U18973 (N_18973,N_18291,N_18125);
or U18974 (N_18974,N_18029,N_18432);
and U18975 (N_18975,N_18328,N_18386);
nand U18976 (N_18976,N_18086,N_18282);
nand U18977 (N_18977,N_18483,N_18456);
and U18978 (N_18978,N_18324,N_18395);
and U18979 (N_18979,N_18358,N_18240);
nor U18980 (N_18980,N_18168,N_18419);
nand U18981 (N_18981,N_18022,N_18196);
and U18982 (N_18982,N_18176,N_18424);
or U18983 (N_18983,N_18263,N_18110);
or U18984 (N_18984,N_18396,N_18264);
or U18985 (N_18985,N_18372,N_18194);
or U18986 (N_18986,N_18193,N_18284);
nor U18987 (N_18987,N_18031,N_18329);
and U18988 (N_18988,N_18476,N_18398);
or U18989 (N_18989,N_18217,N_18130);
nand U18990 (N_18990,N_18298,N_18389);
or U18991 (N_18991,N_18270,N_18304);
and U18992 (N_18992,N_18331,N_18212);
and U18993 (N_18993,N_18499,N_18100);
nor U18994 (N_18994,N_18420,N_18395);
nor U18995 (N_18995,N_18222,N_18029);
nor U18996 (N_18996,N_18389,N_18106);
or U18997 (N_18997,N_18427,N_18348);
or U18998 (N_18998,N_18135,N_18185);
or U18999 (N_18999,N_18334,N_18494);
or U19000 (N_19000,N_18683,N_18693);
and U19001 (N_19001,N_18781,N_18816);
nand U19002 (N_19002,N_18702,N_18673);
or U19003 (N_19003,N_18715,N_18775);
and U19004 (N_19004,N_18574,N_18815);
and U19005 (N_19005,N_18818,N_18844);
or U19006 (N_19006,N_18806,N_18835);
nand U19007 (N_19007,N_18593,N_18720);
or U19008 (N_19008,N_18920,N_18779);
nor U19009 (N_19009,N_18944,N_18760);
nor U19010 (N_19010,N_18954,N_18690);
nand U19011 (N_19011,N_18628,N_18773);
or U19012 (N_19012,N_18650,N_18735);
nor U19013 (N_19013,N_18597,N_18562);
nand U19014 (N_19014,N_18919,N_18631);
or U19015 (N_19015,N_18810,N_18968);
nor U19016 (N_19016,N_18997,N_18502);
nand U19017 (N_19017,N_18967,N_18855);
or U19018 (N_19018,N_18868,N_18769);
and U19019 (N_19019,N_18830,N_18639);
or U19020 (N_19020,N_18785,N_18619);
nand U19021 (N_19021,N_18795,N_18667);
xor U19022 (N_19022,N_18821,N_18825);
or U19023 (N_19023,N_18800,N_18978);
and U19024 (N_19024,N_18636,N_18550);
and U19025 (N_19025,N_18762,N_18764);
or U19026 (N_19026,N_18543,N_18851);
and U19027 (N_19027,N_18515,N_18789);
nand U19028 (N_19028,N_18909,N_18588);
nand U19029 (N_19029,N_18642,N_18699);
nand U19030 (N_19030,N_18956,N_18946);
or U19031 (N_19031,N_18974,N_18500);
nor U19032 (N_19032,N_18834,N_18763);
xnor U19033 (N_19033,N_18626,N_18923);
nand U19034 (N_19034,N_18857,N_18756);
and U19035 (N_19035,N_18988,N_18669);
nor U19036 (N_19036,N_18627,N_18655);
and U19037 (N_19037,N_18556,N_18520);
and U19038 (N_19038,N_18982,N_18758);
and U19039 (N_19039,N_18646,N_18659);
and U19040 (N_19040,N_18560,N_18686);
or U19041 (N_19041,N_18587,N_18796);
nor U19042 (N_19042,N_18737,N_18647);
or U19043 (N_19043,N_18506,N_18569);
or U19044 (N_19044,N_18722,N_18525);
nand U19045 (N_19045,N_18869,N_18808);
and U19046 (N_19046,N_18575,N_18805);
or U19047 (N_19047,N_18987,N_18616);
or U19048 (N_19048,N_18952,N_18695);
and U19049 (N_19049,N_18675,N_18989);
nor U19050 (N_19050,N_18605,N_18552);
or U19051 (N_19051,N_18798,N_18558);
nor U19052 (N_19052,N_18547,N_18966);
nor U19053 (N_19053,N_18714,N_18866);
nand U19054 (N_19054,N_18939,N_18738);
and U19055 (N_19055,N_18880,N_18662);
nor U19056 (N_19056,N_18536,N_18514);
nand U19057 (N_19057,N_18841,N_18533);
or U19058 (N_19058,N_18774,N_18538);
and U19059 (N_19059,N_18827,N_18973);
and U19060 (N_19060,N_18895,N_18850);
xnor U19061 (N_19061,N_18567,N_18860);
and U19062 (N_19062,N_18622,N_18656);
nand U19063 (N_19063,N_18826,N_18976);
nor U19064 (N_19064,N_18545,N_18728);
nand U19065 (N_19065,N_18638,N_18910);
or U19066 (N_19066,N_18522,N_18936);
or U19067 (N_19067,N_18518,N_18649);
nor U19068 (N_19068,N_18941,N_18721);
nand U19069 (N_19069,N_18573,N_18685);
nor U19070 (N_19070,N_18768,N_18513);
nand U19071 (N_19071,N_18846,N_18801);
and U19072 (N_19072,N_18599,N_18927);
nand U19073 (N_19073,N_18623,N_18963);
and U19074 (N_19074,N_18965,N_18697);
or U19075 (N_19075,N_18742,N_18791);
nor U19076 (N_19076,N_18561,N_18645);
and U19077 (N_19077,N_18889,N_18688);
nor U19078 (N_19078,N_18904,N_18881);
nor U19079 (N_19079,N_18915,N_18777);
or U19080 (N_19080,N_18677,N_18894);
nand U19081 (N_19081,N_18576,N_18754);
or U19082 (N_19082,N_18906,N_18644);
or U19083 (N_19083,N_18765,N_18739);
nor U19084 (N_19084,N_18814,N_18848);
nand U19085 (N_19085,N_18694,N_18842);
nand U19086 (N_19086,N_18504,N_18600);
and U19087 (N_19087,N_18847,N_18862);
and U19088 (N_19088,N_18517,N_18858);
or U19089 (N_19089,N_18527,N_18565);
nor U19090 (N_19090,N_18918,N_18661);
nor U19091 (N_19091,N_18886,N_18879);
or U19092 (N_19092,N_18679,N_18975);
and U19093 (N_19093,N_18712,N_18937);
and U19094 (N_19094,N_18892,N_18787);
nand U19095 (N_19095,N_18696,N_18829);
and U19096 (N_19096,N_18797,N_18621);
nor U19097 (N_19097,N_18691,N_18951);
and U19098 (N_19098,N_18732,N_18617);
and U19099 (N_19099,N_18511,N_18658);
or U19100 (N_19100,N_18700,N_18955);
nor U19101 (N_19101,N_18865,N_18548);
and U19102 (N_19102,N_18893,N_18709);
or U19103 (N_19103,N_18554,N_18803);
and U19104 (N_19104,N_18563,N_18990);
nor U19105 (N_19105,N_18716,N_18899);
and U19106 (N_19106,N_18993,N_18926);
nand U19107 (N_19107,N_18689,N_18559);
or U19108 (N_19108,N_18674,N_18723);
and U19109 (N_19109,N_18940,N_18744);
nand U19110 (N_19110,N_18969,N_18983);
or U19111 (N_19111,N_18883,N_18708);
nor U19112 (N_19112,N_18749,N_18579);
nor U19113 (N_19113,N_18703,N_18824);
nor U19114 (N_19114,N_18657,N_18970);
nor U19115 (N_19115,N_18555,N_18871);
nor U19116 (N_19116,N_18611,N_18719);
and U19117 (N_19117,N_18986,N_18596);
nor U19118 (N_19118,N_18804,N_18519);
nand U19119 (N_19119,N_18509,N_18510);
or U19120 (N_19120,N_18705,N_18994);
and U19121 (N_19121,N_18828,N_18707);
nand U19122 (N_19122,N_18584,N_18635);
nor U19123 (N_19123,N_18819,N_18831);
and U19124 (N_19124,N_18745,N_18681);
nand U19125 (N_19125,N_18953,N_18640);
or U19126 (N_19126,N_18531,N_18917);
nand U19127 (N_19127,N_18668,N_18692);
nor U19128 (N_19128,N_18783,N_18535);
nor U19129 (N_19129,N_18949,N_18761);
and U19130 (N_19130,N_18529,N_18602);
nand U19131 (N_19131,N_18580,N_18960);
xor U19132 (N_19132,N_18666,N_18985);
nor U19133 (N_19133,N_18660,N_18750);
nor U19134 (N_19134,N_18788,N_18961);
nand U19135 (N_19135,N_18813,N_18925);
nor U19136 (N_19136,N_18741,N_18746);
nor U19137 (N_19137,N_18874,N_18729);
and U19138 (N_19138,N_18943,N_18507);
or U19139 (N_19139,N_18964,N_18641);
nand U19140 (N_19140,N_18603,N_18770);
nand U19141 (N_19141,N_18671,N_18630);
and U19142 (N_19142,N_18875,N_18891);
or U19143 (N_19143,N_18900,N_18701);
nand U19144 (N_19144,N_18604,N_18537);
and U19145 (N_19145,N_18534,N_18687);
nand U19146 (N_19146,N_18678,N_18908);
or U19147 (N_19147,N_18807,N_18592);
nand U19148 (N_19148,N_18888,N_18947);
and U19149 (N_19149,N_18609,N_18608);
or U19150 (N_19150,N_18962,N_18924);
or U19151 (N_19151,N_18822,N_18505);
nand U19152 (N_19152,N_18928,N_18931);
and U19153 (N_19153,N_18902,N_18654);
nor U19154 (N_19154,N_18615,N_18748);
and U19155 (N_19155,N_18809,N_18629);
or U19156 (N_19156,N_18929,N_18887);
nand U19157 (N_19157,N_18792,N_18524);
and U19158 (N_19158,N_18501,N_18595);
nor U19159 (N_19159,N_18778,N_18878);
or U19160 (N_19160,N_18772,N_18632);
nand U19161 (N_19161,N_18736,N_18759);
and U19162 (N_19162,N_18620,N_18546);
or U19163 (N_19163,N_18942,N_18852);
and U19164 (N_19164,N_18718,N_18583);
or U19165 (N_19165,N_18767,N_18832);
or U19166 (N_19166,N_18757,N_18637);
nor U19167 (N_19167,N_18945,N_18704);
and U19168 (N_19168,N_18726,N_18540);
or U19169 (N_19169,N_18933,N_18590);
or U19170 (N_19170,N_18651,N_18734);
or U19171 (N_19171,N_18867,N_18594);
or U19172 (N_19172,N_18624,N_18849);
or U19173 (N_19173,N_18740,N_18753);
or U19174 (N_19174,N_18585,N_18817);
nand U19175 (N_19175,N_18959,N_18725);
or U19176 (N_19176,N_18652,N_18564);
nor U19177 (N_19177,N_18991,N_18812);
nor U19178 (N_19178,N_18676,N_18903);
or U19179 (N_19179,N_18907,N_18771);
nor U19180 (N_19180,N_18843,N_18836);
and U19181 (N_19181,N_18934,N_18672);
or U19182 (N_19182,N_18713,N_18793);
nand U19183 (N_19183,N_18999,N_18950);
nand U19184 (N_19184,N_18872,N_18972);
nor U19185 (N_19185,N_18998,N_18581);
and U19186 (N_19186,N_18633,N_18782);
and U19187 (N_19187,N_18916,N_18684);
and U19188 (N_19188,N_18802,N_18914);
or U19189 (N_19189,N_18508,N_18730);
and U19190 (N_19190,N_18912,N_18711);
nor U19191 (N_19191,N_18523,N_18532);
or U19192 (N_19192,N_18521,N_18980);
or U19193 (N_19193,N_18820,N_18614);
or U19194 (N_19194,N_18551,N_18911);
or U19195 (N_19195,N_18539,N_18863);
or U19196 (N_19196,N_18528,N_18698);
nor U19197 (N_19197,N_18607,N_18755);
xnor U19198 (N_19198,N_18731,N_18577);
and U19199 (N_19199,N_18612,N_18544);
and U19200 (N_19200,N_18526,N_18582);
nand U19201 (N_19201,N_18780,N_18663);
and U19202 (N_19202,N_18799,N_18516);
nand U19203 (N_19203,N_18776,N_18845);
or U19204 (N_19204,N_18625,N_18724);
nand U19205 (N_19205,N_18885,N_18653);
and U19206 (N_19206,N_18549,N_18905);
or U19207 (N_19207,N_18823,N_18727);
xnor U19208 (N_19208,N_18938,N_18864);
and U19209 (N_19209,N_18981,N_18568);
and U19210 (N_19210,N_18837,N_18876);
nor U19211 (N_19211,N_18870,N_18861);
or U19212 (N_19212,N_18897,N_18971);
nor U19213 (N_19213,N_18571,N_18566);
or U19214 (N_19214,N_18706,N_18884);
nor U19215 (N_19215,N_18752,N_18790);
nor U19216 (N_19216,N_18984,N_18578);
or U19217 (N_19217,N_18922,N_18856);
nor U19218 (N_19218,N_18643,N_18751);
or U19219 (N_19219,N_18882,N_18977);
or U19220 (N_19220,N_18935,N_18979);
nand U19221 (N_19221,N_18680,N_18553);
and U19222 (N_19222,N_18591,N_18840);
xnor U19223 (N_19223,N_18747,N_18948);
or U19224 (N_19224,N_18648,N_18877);
nor U19225 (N_19225,N_18992,N_18530);
nor U19226 (N_19226,N_18930,N_18586);
and U19227 (N_19227,N_18601,N_18598);
nand U19228 (N_19228,N_18839,N_18957);
nor U19229 (N_19229,N_18932,N_18854);
and U19230 (N_19230,N_18958,N_18717);
xnor U19231 (N_19231,N_18618,N_18512);
or U19232 (N_19232,N_18613,N_18794);
and U19233 (N_19233,N_18557,N_18570);
and U19234 (N_19234,N_18890,N_18811);
and U19235 (N_19235,N_18606,N_18710);
and U19236 (N_19236,N_18853,N_18541);
or U19237 (N_19237,N_18996,N_18733);
nand U19238 (N_19238,N_18743,N_18589);
or U19239 (N_19239,N_18913,N_18664);
or U19240 (N_19240,N_18572,N_18670);
nor U19241 (N_19241,N_18766,N_18901);
and U19242 (N_19242,N_18833,N_18665);
nand U19243 (N_19243,N_18786,N_18503);
or U19244 (N_19244,N_18898,N_18873);
xnor U19245 (N_19245,N_18634,N_18784);
and U19246 (N_19246,N_18859,N_18921);
and U19247 (N_19247,N_18995,N_18682);
nor U19248 (N_19248,N_18542,N_18838);
and U19249 (N_19249,N_18896,N_18610);
nor U19250 (N_19250,N_18754,N_18871);
or U19251 (N_19251,N_18638,N_18713);
and U19252 (N_19252,N_18749,N_18577);
or U19253 (N_19253,N_18811,N_18527);
and U19254 (N_19254,N_18581,N_18567);
and U19255 (N_19255,N_18674,N_18711);
nor U19256 (N_19256,N_18588,N_18571);
xnor U19257 (N_19257,N_18896,N_18900);
nor U19258 (N_19258,N_18963,N_18912);
nand U19259 (N_19259,N_18766,N_18574);
or U19260 (N_19260,N_18786,N_18935);
nand U19261 (N_19261,N_18796,N_18878);
and U19262 (N_19262,N_18821,N_18564);
nor U19263 (N_19263,N_18546,N_18742);
xnor U19264 (N_19264,N_18553,N_18928);
nand U19265 (N_19265,N_18847,N_18743);
nand U19266 (N_19266,N_18813,N_18761);
nor U19267 (N_19267,N_18840,N_18621);
nor U19268 (N_19268,N_18627,N_18776);
nor U19269 (N_19269,N_18981,N_18910);
nand U19270 (N_19270,N_18870,N_18661);
and U19271 (N_19271,N_18655,N_18915);
nand U19272 (N_19272,N_18758,N_18651);
or U19273 (N_19273,N_18518,N_18642);
nor U19274 (N_19274,N_18767,N_18651);
and U19275 (N_19275,N_18515,N_18796);
nor U19276 (N_19276,N_18999,N_18821);
and U19277 (N_19277,N_18643,N_18911);
or U19278 (N_19278,N_18815,N_18723);
nor U19279 (N_19279,N_18636,N_18705);
nand U19280 (N_19280,N_18933,N_18895);
nand U19281 (N_19281,N_18700,N_18800);
nor U19282 (N_19282,N_18500,N_18770);
nor U19283 (N_19283,N_18556,N_18886);
nor U19284 (N_19284,N_18606,N_18824);
and U19285 (N_19285,N_18835,N_18901);
or U19286 (N_19286,N_18882,N_18958);
or U19287 (N_19287,N_18963,N_18752);
nand U19288 (N_19288,N_18822,N_18602);
nor U19289 (N_19289,N_18769,N_18563);
nor U19290 (N_19290,N_18991,N_18792);
and U19291 (N_19291,N_18894,N_18999);
nor U19292 (N_19292,N_18825,N_18724);
nor U19293 (N_19293,N_18768,N_18570);
and U19294 (N_19294,N_18727,N_18711);
or U19295 (N_19295,N_18858,N_18806);
and U19296 (N_19296,N_18669,N_18964);
nand U19297 (N_19297,N_18916,N_18893);
or U19298 (N_19298,N_18822,N_18880);
nand U19299 (N_19299,N_18743,N_18526);
or U19300 (N_19300,N_18865,N_18677);
and U19301 (N_19301,N_18516,N_18528);
nand U19302 (N_19302,N_18547,N_18516);
and U19303 (N_19303,N_18578,N_18575);
nor U19304 (N_19304,N_18550,N_18989);
or U19305 (N_19305,N_18991,N_18845);
nor U19306 (N_19306,N_18852,N_18517);
or U19307 (N_19307,N_18893,N_18959);
and U19308 (N_19308,N_18861,N_18509);
nor U19309 (N_19309,N_18697,N_18534);
or U19310 (N_19310,N_18715,N_18764);
nor U19311 (N_19311,N_18899,N_18663);
nor U19312 (N_19312,N_18511,N_18761);
xor U19313 (N_19313,N_18693,N_18698);
nand U19314 (N_19314,N_18923,N_18529);
and U19315 (N_19315,N_18619,N_18856);
nand U19316 (N_19316,N_18844,N_18966);
nor U19317 (N_19317,N_18679,N_18934);
and U19318 (N_19318,N_18678,N_18715);
nand U19319 (N_19319,N_18921,N_18539);
or U19320 (N_19320,N_18859,N_18507);
nor U19321 (N_19321,N_18889,N_18598);
and U19322 (N_19322,N_18545,N_18760);
nand U19323 (N_19323,N_18578,N_18655);
xnor U19324 (N_19324,N_18574,N_18573);
nor U19325 (N_19325,N_18605,N_18844);
or U19326 (N_19326,N_18705,N_18999);
and U19327 (N_19327,N_18871,N_18759);
or U19328 (N_19328,N_18777,N_18600);
nand U19329 (N_19329,N_18582,N_18947);
nand U19330 (N_19330,N_18726,N_18942);
nand U19331 (N_19331,N_18781,N_18730);
nor U19332 (N_19332,N_18891,N_18801);
or U19333 (N_19333,N_18504,N_18770);
or U19334 (N_19334,N_18947,N_18611);
nor U19335 (N_19335,N_18737,N_18636);
or U19336 (N_19336,N_18606,N_18652);
xnor U19337 (N_19337,N_18751,N_18788);
nand U19338 (N_19338,N_18682,N_18962);
or U19339 (N_19339,N_18651,N_18778);
nand U19340 (N_19340,N_18773,N_18500);
nor U19341 (N_19341,N_18954,N_18689);
or U19342 (N_19342,N_18528,N_18513);
nor U19343 (N_19343,N_18996,N_18675);
xor U19344 (N_19344,N_18782,N_18950);
nor U19345 (N_19345,N_18941,N_18597);
or U19346 (N_19346,N_18500,N_18895);
nand U19347 (N_19347,N_18788,N_18842);
nor U19348 (N_19348,N_18571,N_18507);
xnor U19349 (N_19349,N_18641,N_18648);
or U19350 (N_19350,N_18569,N_18702);
nand U19351 (N_19351,N_18824,N_18962);
and U19352 (N_19352,N_18659,N_18519);
nor U19353 (N_19353,N_18767,N_18791);
xor U19354 (N_19354,N_18512,N_18948);
nand U19355 (N_19355,N_18593,N_18718);
nand U19356 (N_19356,N_18891,N_18835);
nand U19357 (N_19357,N_18911,N_18674);
xnor U19358 (N_19358,N_18961,N_18949);
nand U19359 (N_19359,N_18968,N_18909);
and U19360 (N_19360,N_18748,N_18533);
and U19361 (N_19361,N_18529,N_18745);
xnor U19362 (N_19362,N_18782,N_18555);
nand U19363 (N_19363,N_18580,N_18632);
or U19364 (N_19364,N_18630,N_18875);
and U19365 (N_19365,N_18781,N_18751);
and U19366 (N_19366,N_18952,N_18872);
nand U19367 (N_19367,N_18544,N_18681);
and U19368 (N_19368,N_18990,N_18516);
or U19369 (N_19369,N_18643,N_18809);
nand U19370 (N_19370,N_18767,N_18793);
or U19371 (N_19371,N_18746,N_18834);
or U19372 (N_19372,N_18606,N_18938);
or U19373 (N_19373,N_18635,N_18742);
or U19374 (N_19374,N_18811,N_18513);
and U19375 (N_19375,N_18599,N_18517);
or U19376 (N_19376,N_18818,N_18693);
nor U19377 (N_19377,N_18765,N_18603);
nor U19378 (N_19378,N_18566,N_18755);
nor U19379 (N_19379,N_18939,N_18746);
or U19380 (N_19380,N_18738,N_18843);
and U19381 (N_19381,N_18982,N_18676);
and U19382 (N_19382,N_18886,N_18768);
nand U19383 (N_19383,N_18826,N_18680);
and U19384 (N_19384,N_18826,N_18690);
nor U19385 (N_19385,N_18732,N_18987);
and U19386 (N_19386,N_18668,N_18689);
and U19387 (N_19387,N_18740,N_18867);
nor U19388 (N_19388,N_18538,N_18768);
nand U19389 (N_19389,N_18821,N_18986);
or U19390 (N_19390,N_18735,N_18753);
and U19391 (N_19391,N_18525,N_18906);
and U19392 (N_19392,N_18747,N_18682);
or U19393 (N_19393,N_18526,N_18522);
nor U19394 (N_19394,N_18641,N_18766);
nand U19395 (N_19395,N_18797,N_18812);
xnor U19396 (N_19396,N_18617,N_18908);
nand U19397 (N_19397,N_18635,N_18732);
and U19398 (N_19398,N_18704,N_18716);
and U19399 (N_19399,N_18847,N_18886);
or U19400 (N_19400,N_18993,N_18535);
nor U19401 (N_19401,N_18575,N_18837);
nand U19402 (N_19402,N_18995,N_18854);
or U19403 (N_19403,N_18980,N_18625);
nor U19404 (N_19404,N_18535,N_18918);
nor U19405 (N_19405,N_18825,N_18845);
nand U19406 (N_19406,N_18992,N_18895);
or U19407 (N_19407,N_18529,N_18805);
nand U19408 (N_19408,N_18843,N_18784);
or U19409 (N_19409,N_18770,N_18739);
nand U19410 (N_19410,N_18960,N_18735);
nor U19411 (N_19411,N_18905,N_18995);
and U19412 (N_19412,N_18915,N_18845);
nand U19413 (N_19413,N_18946,N_18826);
and U19414 (N_19414,N_18996,N_18845);
or U19415 (N_19415,N_18870,N_18514);
and U19416 (N_19416,N_18890,N_18989);
nand U19417 (N_19417,N_18807,N_18800);
and U19418 (N_19418,N_18690,N_18981);
nor U19419 (N_19419,N_18618,N_18910);
nand U19420 (N_19420,N_18589,N_18905);
nor U19421 (N_19421,N_18945,N_18783);
or U19422 (N_19422,N_18873,N_18965);
nor U19423 (N_19423,N_18791,N_18625);
and U19424 (N_19424,N_18642,N_18936);
or U19425 (N_19425,N_18805,N_18789);
nor U19426 (N_19426,N_18673,N_18897);
and U19427 (N_19427,N_18893,N_18622);
and U19428 (N_19428,N_18581,N_18794);
nor U19429 (N_19429,N_18605,N_18658);
nand U19430 (N_19430,N_18813,N_18880);
or U19431 (N_19431,N_18549,N_18673);
or U19432 (N_19432,N_18950,N_18725);
nor U19433 (N_19433,N_18532,N_18915);
xnor U19434 (N_19434,N_18904,N_18626);
and U19435 (N_19435,N_18993,N_18988);
or U19436 (N_19436,N_18820,N_18719);
nor U19437 (N_19437,N_18545,N_18743);
nor U19438 (N_19438,N_18872,N_18626);
nor U19439 (N_19439,N_18765,N_18900);
or U19440 (N_19440,N_18618,N_18587);
or U19441 (N_19441,N_18848,N_18824);
and U19442 (N_19442,N_18927,N_18926);
or U19443 (N_19443,N_18854,N_18568);
and U19444 (N_19444,N_18678,N_18537);
nand U19445 (N_19445,N_18935,N_18730);
and U19446 (N_19446,N_18530,N_18543);
nor U19447 (N_19447,N_18852,N_18636);
xnor U19448 (N_19448,N_18937,N_18654);
nor U19449 (N_19449,N_18559,N_18709);
and U19450 (N_19450,N_18550,N_18619);
or U19451 (N_19451,N_18930,N_18687);
nand U19452 (N_19452,N_18815,N_18589);
or U19453 (N_19453,N_18533,N_18524);
or U19454 (N_19454,N_18877,N_18879);
nand U19455 (N_19455,N_18774,N_18862);
nor U19456 (N_19456,N_18788,N_18618);
and U19457 (N_19457,N_18694,N_18733);
and U19458 (N_19458,N_18661,N_18639);
or U19459 (N_19459,N_18947,N_18741);
nor U19460 (N_19460,N_18885,N_18853);
and U19461 (N_19461,N_18682,N_18589);
or U19462 (N_19462,N_18572,N_18846);
and U19463 (N_19463,N_18733,N_18961);
nand U19464 (N_19464,N_18519,N_18627);
and U19465 (N_19465,N_18692,N_18529);
nand U19466 (N_19466,N_18907,N_18669);
nand U19467 (N_19467,N_18629,N_18570);
and U19468 (N_19468,N_18674,N_18947);
nor U19469 (N_19469,N_18534,N_18897);
or U19470 (N_19470,N_18615,N_18508);
or U19471 (N_19471,N_18892,N_18983);
nor U19472 (N_19472,N_18502,N_18560);
nor U19473 (N_19473,N_18810,N_18714);
and U19474 (N_19474,N_18758,N_18719);
or U19475 (N_19475,N_18647,N_18902);
nor U19476 (N_19476,N_18958,N_18846);
or U19477 (N_19477,N_18945,N_18637);
and U19478 (N_19478,N_18534,N_18901);
nor U19479 (N_19479,N_18549,N_18626);
nor U19480 (N_19480,N_18548,N_18578);
and U19481 (N_19481,N_18987,N_18710);
xor U19482 (N_19482,N_18685,N_18675);
or U19483 (N_19483,N_18546,N_18853);
nand U19484 (N_19484,N_18604,N_18627);
nand U19485 (N_19485,N_18803,N_18696);
and U19486 (N_19486,N_18686,N_18506);
nand U19487 (N_19487,N_18975,N_18632);
nand U19488 (N_19488,N_18708,N_18956);
or U19489 (N_19489,N_18642,N_18973);
nor U19490 (N_19490,N_18783,N_18632);
xor U19491 (N_19491,N_18924,N_18771);
and U19492 (N_19492,N_18725,N_18966);
xnor U19493 (N_19493,N_18639,N_18502);
or U19494 (N_19494,N_18677,N_18723);
or U19495 (N_19495,N_18919,N_18667);
and U19496 (N_19496,N_18763,N_18965);
nand U19497 (N_19497,N_18689,N_18910);
and U19498 (N_19498,N_18808,N_18762);
or U19499 (N_19499,N_18531,N_18977);
nor U19500 (N_19500,N_19353,N_19266);
or U19501 (N_19501,N_19205,N_19332);
nor U19502 (N_19502,N_19317,N_19161);
xor U19503 (N_19503,N_19407,N_19419);
nor U19504 (N_19504,N_19031,N_19399);
nand U19505 (N_19505,N_19046,N_19019);
or U19506 (N_19506,N_19142,N_19440);
nand U19507 (N_19507,N_19413,N_19453);
and U19508 (N_19508,N_19428,N_19193);
and U19509 (N_19509,N_19214,N_19203);
nand U19510 (N_19510,N_19243,N_19000);
nand U19511 (N_19511,N_19138,N_19326);
nor U19512 (N_19512,N_19129,N_19423);
and U19513 (N_19513,N_19213,N_19258);
nand U19514 (N_19514,N_19004,N_19447);
or U19515 (N_19515,N_19387,N_19474);
nand U19516 (N_19516,N_19469,N_19181);
or U19517 (N_19517,N_19371,N_19248);
and U19518 (N_19518,N_19079,N_19246);
nand U19519 (N_19519,N_19064,N_19329);
or U19520 (N_19520,N_19376,N_19273);
and U19521 (N_19521,N_19264,N_19063);
and U19522 (N_19522,N_19035,N_19037);
nor U19523 (N_19523,N_19437,N_19402);
nand U19524 (N_19524,N_19366,N_19251);
or U19525 (N_19525,N_19165,N_19051);
or U19526 (N_19526,N_19049,N_19357);
nand U19527 (N_19527,N_19052,N_19297);
or U19528 (N_19528,N_19128,N_19062);
nand U19529 (N_19529,N_19302,N_19173);
nor U19530 (N_19530,N_19429,N_19348);
or U19531 (N_19531,N_19075,N_19236);
nor U19532 (N_19532,N_19085,N_19185);
and U19533 (N_19533,N_19304,N_19081);
and U19534 (N_19534,N_19150,N_19089);
nor U19535 (N_19535,N_19252,N_19218);
and U19536 (N_19536,N_19333,N_19389);
nand U19537 (N_19537,N_19337,N_19416);
nand U19538 (N_19538,N_19274,N_19253);
and U19539 (N_19539,N_19498,N_19444);
nand U19540 (N_19540,N_19118,N_19272);
or U19541 (N_19541,N_19277,N_19050);
and U19542 (N_19542,N_19146,N_19306);
and U19543 (N_19543,N_19044,N_19137);
nor U19544 (N_19544,N_19270,N_19202);
nor U19545 (N_19545,N_19341,N_19324);
nand U19546 (N_19546,N_19080,N_19382);
nor U19547 (N_19547,N_19462,N_19295);
xnor U19548 (N_19548,N_19372,N_19321);
and U19549 (N_19549,N_19155,N_19268);
nor U19550 (N_19550,N_19254,N_19334);
and U19551 (N_19551,N_19336,N_19397);
or U19552 (N_19552,N_19493,N_19244);
nand U19553 (N_19553,N_19412,N_19293);
or U19554 (N_19554,N_19263,N_19346);
nand U19555 (N_19555,N_19294,N_19014);
nor U19556 (N_19556,N_19340,N_19426);
and U19557 (N_19557,N_19191,N_19163);
nand U19558 (N_19558,N_19471,N_19066);
nor U19559 (N_19559,N_19182,N_19145);
nor U19560 (N_19560,N_19409,N_19406);
nand U19561 (N_19561,N_19093,N_19410);
nor U19562 (N_19562,N_19386,N_19126);
and U19563 (N_19563,N_19188,N_19108);
nand U19564 (N_19564,N_19132,N_19158);
nor U19565 (N_19565,N_19276,N_19076);
nand U19566 (N_19566,N_19058,N_19457);
or U19567 (N_19567,N_19492,N_19026);
or U19568 (N_19568,N_19124,N_19443);
xor U19569 (N_19569,N_19168,N_19384);
and U19570 (N_19570,N_19069,N_19176);
and U19571 (N_19571,N_19458,N_19421);
nand U19572 (N_19572,N_19141,N_19223);
nand U19573 (N_19573,N_19491,N_19178);
nor U19574 (N_19574,N_19180,N_19356);
nand U19575 (N_19575,N_19029,N_19260);
nand U19576 (N_19576,N_19121,N_19083);
and U19577 (N_19577,N_19209,N_19184);
and U19578 (N_19578,N_19327,N_19338);
nand U19579 (N_19579,N_19436,N_19430);
nor U19580 (N_19580,N_19100,N_19149);
nor U19581 (N_19581,N_19082,N_19005);
nand U19582 (N_19582,N_19257,N_19127);
nor U19583 (N_19583,N_19283,N_19284);
nand U19584 (N_19584,N_19060,N_19393);
or U19585 (N_19585,N_19370,N_19422);
and U19586 (N_19586,N_19227,N_19130);
and U19587 (N_19587,N_19009,N_19299);
or U19588 (N_19588,N_19164,N_19090);
nor U19589 (N_19589,N_19278,N_19032);
nand U19590 (N_19590,N_19048,N_19225);
or U19591 (N_19591,N_19388,N_19434);
or U19592 (N_19592,N_19078,N_19136);
nor U19593 (N_19593,N_19194,N_19403);
and U19594 (N_19594,N_19210,N_19343);
nor U19595 (N_19595,N_19224,N_19087);
nand U19596 (N_19596,N_19433,N_19237);
nor U19597 (N_19597,N_19394,N_19255);
and U19598 (N_19598,N_19111,N_19368);
and U19599 (N_19599,N_19139,N_19016);
nand U19600 (N_19600,N_19379,N_19170);
or U19601 (N_19601,N_19449,N_19047);
and U19602 (N_19602,N_19404,N_19098);
or U19603 (N_19603,N_19454,N_19411);
nor U19604 (N_19604,N_19094,N_19424);
and U19605 (N_19605,N_19012,N_19301);
nand U19606 (N_19606,N_19183,N_19310);
and U19607 (N_19607,N_19110,N_19077);
nand U19608 (N_19608,N_19425,N_19204);
and U19609 (N_19609,N_19177,N_19140);
nand U19610 (N_19610,N_19490,N_19119);
nand U19611 (N_19611,N_19380,N_19358);
or U19612 (N_19612,N_19298,N_19355);
nand U19613 (N_19613,N_19347,N_19465);
or U19614 (N_19614,N_19109,N_19486);
nor U19615 (N_19615,N_19296,N_19311);
nand U19616 (N_19616,N_19024,N_19056);
nand U19617 (N_19617,N_19395,N_19431);
nor U19618 (N_19618,N_19418,N_19484);
nor U19619 (N_19619,N_19269,N_19441);
or U19620 (N_19620,N_19286,N_19488);
or U19621 (N_19621,N_19467,N_19420);
and U19622 (N_19622,N_19199,N_19249);
and U19623 (N_19623,N_19006,N_19452);
and U19624 (N_19624,N_19114,N_19192);
nor U19625 (N_19625,N_19360,N_19313);
or U19626 (N_19626,N_19041,N_19095);
nor U19627 (N_19627,N_19435,N_19282);
nand U19628 (N_19628,N_19091,N_19143);
xor U19629 (N_19629,N_19001,N_19461);
and U19630 (N_19630,N_19365,N_19175);
nor U19631 (N_19631,N_19135,N_19215);
nor U19632 (N_19632,N_19456,N_19201);
nor U19633 (N_19633,N_19101,N_19442);
or U19634 (N_19634,N_19445,N_19247);
or U19635 (N_19635,N_19207,N_19065);
and U19636 (N_19636,N_19231,N_19017);
and U19637 (N_19637,N_19305,N_19328);
nor U19638 (N_19638,N_19112,N_19217);
or U19639 (N_19639,N_19446,N_19369);
and U19640 (N_19640,N_19351,N_19289);
nor U19641 (N_19641,N_19314,N_19220);
nand U19642 (N_19642,N_19157,N_19342);
or U19643 (N_19643,N_19238,N_19068);
or U19644 (N_19644,N_19038,N_19007);
or U19645 (N_19645,N_19073,N_19279);
nand U19646 (N_19646,N_19361,N_19107);
nand U19647 (N_19647,N_19468,N_19400);
and U19648 (N_19648,N_19460,N_19401);
nand U19649 (N_19649,N_19497,N_19022);
nor U19650 (N_19650,N_19228,N_19359);
nand U19651 (N_19651,N_19025,N_19042);
nor U19652 (N_19652,N_19450,N_19120);
nand U19653 (N_19653,N_19233,N_19055);
xnor U19654 (N_19654,N_19144,N_19378);
nand U19655 (N_19655,N_19432,N_19349);
and U19656 (N_19656,N_19466,N_19088);
nand U19657 (N_19657,N_19169,N_19148);
nor U19658 (N_19658,N_19216,N_19020);
nor U19659 (N_19659,N_19134,N_19187);
nor U19660 (N_19660,N_19221,N_19325);
nor U19661 (N_19661,N_19285,N_19339);
nor U19662 (N_19662,N_19097,N_19408);
nor U19663 (N_19663,N_19023,N_19463);
nand U19664 (N_19664,N_19195,N_19256);
nand U19665 (N_19665,N_19479,N_19105);
and U19666 (N_19666,N_19487,N_19480);
or U19667 (N_19667,N_19160,N_19464);
or U19668 (N_19668,N_19290,N_19013);
and U19669 (N_19669,N_19417,N_19451);
and U19670 (N_19670,N_19459,N_19222);
and U19671 (N_19671,N_19106,N_19345);
nand U19672 (N_19672,N_19003,N_19167);
and U19673 (N_19673,N_19125,N_19240);
nand U19674 (N_19674,N_19381,N_19316);
or U19675 (N_19675,N_19067,N_19331);
or U19676 (N_19676,N_19239,N_19472);
nand U19677 (N_19677,N_19320,N_19166);
and U19678 (N_19678,N_19259,N_19245);
or U19679 (N_19679,N_19219,N_19485);
or U19680 (N_19680,N_19117,N_19071);
nand U19681 (N_19681,N_19318,N_19212);
nor U19682 (N_19682,N_19092,N_19190);
nor U19683 (N_19683,N_19483,N_19281);
xnor U19684 (N_19684,N_19481,N_19116);
and U19685 (N_19685,N_19053,N_19208);
nor U19686 (N_19686,N_19034,N_19280);
nor U19687 (N_19687,N_19392,N_19131);
and U19688 (N_19688,N_19186,N_19229);
and U19689 (N_19689,N_19102,N_19265);
and U19690 (N_19690,N_19473,N_19174);
and U19691 (N_19691,N_19377,N_19494);
xnor U19692 (N_19692,N_19096,N_19200);
or U19693 (N_19693,N_19405,N_19030);
or U19694 (N_19694,N_19291,N_19061);
or U19695 (N_19695,N_19288,N_19367);
nor U19696 (N_19696,N_19010,N_19335);
nor U19697 (N_19697,N_19039,N_19330);
or U19698 (N_19698,N_19070,N_19439);
nor U19699 (N_19699,N_19002,N_19057);
nand U19700 (N_19700,N_19113,N_19122);
or U19701 (N_19701,N_19364,N_19027);
or U19702 (N_19702,N_19300,N_19262);
and U19703 (N_19703,N_19011,N_19015);
nand U19704 (N_19704,N_19230,N_19028);
and U19705 (N_19705,N_19103,N_19261);
nand U19706 (N_19706,N_19235,N_19390);
or U19707 (N_19707,N_19308,N_19241);
or U19708 (N_19708,N_19344,N_19226);
nor U19709 (N_19709,N_19375,N_19267);
nand U19710 (N_19710,N_19363,N_19396);
nand U19711 (N_19711,N_19043,N_19312);
or U19712 (N_19712,N_19415,N_19499);
nand U19713 (N_19713,N_19072,N_19414);
nand U19714 (N_19714,N_19232,N_19322);
nand U19715 (N_19715,N_19383,N_19319);
and U19716 (N_19716,N_19287,N_19197);
nor U19717 (N_19717,N_19495,N_19156);
nor U19718 (N_19718,N_19292,N_19162);
and U19719 (N_19719,N_19489,N_19309);
or U19720 (N_19720,N_19374,N_19496);
nand U19721 (N_19721,N_19350,N_19352);
and U19722 (N_19722,N_19198,N_19172);
and U19723 (N_19723,N_19159,N_19398);
or U19724 (N_19724,N_19021,N_19234);
nand U19725 (N_19725,N_19086,N_19033);
nand U19726 (N_19726,N_19153,N_19151);
nand U19727 (N_19727,N_19179,N_19385);
or U19728 (N_19728,N_19242,N_19315);
nand U19729 (N_19729,N_19133,N_19478);
and U19730 (N_19730,N_19045,N_19354);
or U19731 (N_19731,N_19373,N_19362);
nor U19732 (N_19732,N_19448,N_19171);
nor U19733 (N_19733,N_19115,N_19206);
and U19734 (N_19734,N_19099,N_19104);
nand U19735 (N_19735,N_19482,N_19196);
or U19736 (N_19736,N_19211,N_19476);
and U19737 (N_19737,N_19455,N_19154);
or U19738 (N_19738,N_19147,N_19018);
nand U19739 (N_19739,N_19427,N_19275);
nor U19740 (N_19740,N_19084,N_19271);
or U19741 (N_19741,N_19074,N_19307);
xor U19742 (N_19742,N_19470,N_19040);
or U19743 (N_19743,N_19250,N_19189);
nand U19744 (N_19744,N_19391,N_19477);
nor U19745 (N_19745,N_19323,N_19303);
or U19746 (N_19746,N_19059,N_19123);
or U19747 (N_19747,N_19036,N_19008);
or U19748 (N_19748,N_19438,N_19054);
nand U19749 (N_19749,N_19475,N_19152);
and U19750 (N_19750,N_19115,N_19242);
nor U19751 (N_19751,N_19120,N_19246);
nand U19752 (N_19752,N_19147,N_19378);
nand U19753 (N_19753,N_19395,N_19204);
nor U19754 (N_19754,N_19469,N_19156);
nand U19755 (N_19755,N_19323,N_19458);
and U19756 (N_19756,N_19068,N_19033);
and U19757 (N_19757,N_19332,N_19210);
and U19758 (N_19758,N_19324,N_19356);
nor U19759 (N_19759,N_19430,N_19045);
nand U19760 (N_19760,N_19180,N_19307);
nor U19761 (N_19761,N_19344,N_19058);
and U19762 (N_19762,N_19354,N_19020);
or U19763 (N_19763,N_19055,N_19353);
or U19764 (N_19764,N_19124,N_19349);
nor U19765 (N_19765,N_19420,N_19181);
or U19766 (N_19766,N_19420,N_19172);
nand U19767 (N_19767,N_19363,N_19122);
or U19768 (N_19768,N_19114,N_19247);
nand U19769 (N_19769,N_19409,N_19217);
and U19770 (N_19770,N_19308,N_19334);
and U19771 (N_19771,N_19059,N_19258);
nand U19772 (N_19772,N_19123,N_19067);
nand U19773 (N_19773,N_19480,N_19069);
nor U19774 (N_19774,N_19201,N_19411);
nand U19775 (N_19775,N_19267,N_19204);
and U19776 (N_19776,N_19312,N_19384);
and U19777 (N_19777,N_19242,N_19368);
or U19778 (N_19778,N_19380,N_19162);
nand U19779 (N_19779,N_19353,N_19157);
and U19780 (N_19780,N_19332,N_19339);
xor U19781 (N_19781,N_19273,N_19000);
nand U19782 (N_19782,N_19129,N_19209);
nand U19783 (N_19783,N_19299,N_19205);
or U19784 (N_19784,N_19166,N_19432);
nand U19785 (N_19785,N_19072,N_19384);
nand U19786 (N_19786,N_19349,N_19412);
nor U19787 (N_19787,N_19200,N_19261);
or U19788 (N_19788,N_19421,N_19180);
or U19789 (N_19789,N_19440,N_19337);
nand U19790 (N_19790,N_19008,N_19497);
xor U19791 (N_19791,N_19124,N_19087);
and U19792 (N_19792,N_19461,N_19239);
or U19793 (N_19793,N_19105,N_19398);
nand U19794 (N_19794,N_19326,N_19479);
or U19795 (N_19795,N_19470,N_19404);
and U19796 (N_19796,N_19394,N_19243);
or U19797 (N_19797,N_19060,N_19343);
or U19798 (N_19798,N_19097,N_19332);
and U19799 (N_19799,N_19340,N_19186);
and U19800 (N_19800,N_19020,N_19369);
nand U19801 (N_19801,N_19471,N_19163);
or U19802 (N_19802,N_19163,N_19118);
and U19803 (N_19803,N_19084,N_19144);
nor U19804 (N_19804,N_19317,N_19461);
xnor U19805 (N_19805,N_19062,N_19168);
and U19806 (N_19806,N_19156,N_19006);
or U19807 (N_19807,N_19031,N_19247);
or U19808 (N_19808,N_19031,N_19441);
nand U19809 (N_19809,N_19119,N_19018);
and U19810 (N_19810,N_19161,N_19302);
and U19811 (N_19811,N_19283,N_19400);
or U19812 (N_19812,N_19089,N_19163);
nor U19813 (N_19813,N_19320,N_19036);
nor U19814 (N_19814,N_19199,N_19128);
nor U19815 (N_19815,N_19248,N_19454);
xor U19816 (N_19816,N_19319,N_19100);
or U19817 (N_19817,N_19226,N_19241);
and U19818 (N_19818,N_19213,N_19265);
or U19819 (N_19819,N_19238,N_19128);
or U19820 (N_19820,N_19426,N_19198);
nor U19821 (N_19821,N_19168,N_19152);
nor U19822 (N_19822,N_19202,N_19214);
and U19823 (N_19823,N_19220,N_19464);
and U19824 (N_19824,N_19289,N_19145);
and U19825 (N_19825,N_19063,N_19042);
and U19826 (N_19826,N_19344,N_19469);
and U19827 (N_19827,N_19333,N_19447);
and U19828 (N_19828,N_19371,N_19285);
or U19829 (N_19829,N_19313,N_19271);
or U19830 (N_19830,N_19259,N_19321);
nor U19831 (N_19831,N_19209,N_19256);
or U19832 (N_19832,N_19396,N_19273);
or U19833 (N_19833,N_19295,N_19050);
and U19834 (N_19834,N_19204,N_19442);
and U19835 (N_19835,N_19196,N_19239);
or U19836 (N_19836,N_19379,N_19112);
and U19837 (N_19837,N_19004,N_19290);
or U19838 (N_19838,N_19305,N_19126);
nor U19839 (N_19839,N_19401,N_19290);
nand U19840 (N_19840,N_19300,N_19437);
or U19841 (N_19841,N_19117,N_19228);
nor U19842 (N_19842,N_19430,N_19427);
nand U19843 (N_19843,N_19203,N_19096);
xor U19844 (N_19844,N_19121,N_19497);
nor U19845 (N_19845,N_19110,N_19341);
or U19846 (N_19846,N_19413,N_19094);
nor U19847 (N_19847,N_19054,N_19424);
nand U19848 (N_19848,N_19317,N_19272);
or U19849 (N_19849,N_19166,N_19005);
and U19850 (N_19850,N_19122,N_19074);
and U19851 (N_19851,N_19437,N_19425);
and U19852 (N_19852,N_19457,N_19137);
or U19853 (N_19853,N_19257,N_19147);
nor U19854 (N_19854,N_19129,N_19096);
nand U19855 (N_19855,N_19175,N_19151);
xnor U19856 (N_19856,N_19421,N_19112);
nor U19857 (N_19857,N_19097,N_19212);
nand U19858 (N_19858,N_19034,N_19444);
and U19859 (N_19859,N_19026,N_19168);
and U19860 (N_19860,N_19457,N_19044);
nor U19861 (N_19861,N_19187,N_19376);
nand U19862 (N_19862,N_19107,N_19019);
and U19863 (N_19863,N_19377,N_19011);
xor U19864 (N_19864,N_19030,N_19100);
and U19865 (N_19865,N_19013,N_19298);
nor U19866 (N_19866,N_19141,N_19037);
or U19867 (N_19867,N_19118,N_19214);
or U19868 (N_19868,N_19106,N_19253);
and U19869 (N_19869,N_19068,N_19128);
and U19870 (N_19870,N_19453,N_19199);
and U19871 (N_19871,N_19074,N_19357);
or U19872 (N_19872,N_19431,N_19284);
or U19873 (N_19873,N_19258,N_19291);
nand U19874 (N_19874,N_19151,N_19286);
or U19875 (N_19875,N_19189,N_19261);
nor U19876 (N_19876,N_19424,N_19097);
nand U19877 (N_19877,N_19127,N_19435);
or U19878 (N_19878,N_19092,N_19056);
and U19879 (N_19879,N_19499,N_19187);
and U19880 (N_19880,N_19052,N_19319);
and U19881 (N_19881,N_19044,N_19475);
nand U19882 (N_19882,N_19253,N_19149);
and U19883 (N_19883,N_19289,N_19361);
or U19884 (N_19884,N_19228,N_19090);
and U19885 (N_19885,N_19028,N_19380);
nand U19886 (N_19886,N_19245,N_19030);
nor U19887 (N_19887,N_19049,N_19439);
or U19888 (N_19888,N_19105,N_19196);
and U19889 (N_19889,N_19106,N_19022);
and U19890 (N_19890,N_19343,N_19102);
nor U19891 (N_19891,N_19340,N_19165);
nor U19892 (N_19892,N_19479,N_19070);
and U19893 (N_19893,N_19256,N_19100);
or U19894 (N_19894,N_19013,N_19190);
nand U19895 (N_19895,N_19296,N_19182);
xor U19896 (N_19896,N_19471,N_19145);
and U19897 (N_19897,N_19185,N_19220);
or U19898 (N_19898,N_19288,N_19253);
or U19899 (N_19899,N_19395,N_19394);
nand U19900 (N_19900,N_19400,N_19366);
nand U19901 (N_19901,N_19488,N_19427);
nor U19902 (N_19902,N_19138,N_19071);
and U19903 (N_19903,N_19388,N_19405);
or U19904 (N_19904,N_19011,N_19170);
nand U19905 (N_19905,N_19072,N_19359);
or U19906 (N_19906,N_19411,N_19394);
nor U19907 (N_19907,N_19098,N_19168);
and U19908 (N_19908,N_19005,N_19258);
or U19909 (N_19909,N_19063,N_19342);
xnor U19910 (N_19910,N_19200,N_19186);
nor U19911 (N_19911,N_19365,N_19094);
and U19912 (N_19912,N_19037,N_19231);
or U19913 (N_19913,N_19400,N_19413);
or U19914 (N_19914,N_19275,N_19459);
nand U19915 (N_19915,N_19219,N_19291);
nand U19916 (N_19916,N_19402,N_19150);
nor U19917 (N_19917,N_19193,N_19025);
xor U19918 (N_19918,N_19425,N_19012);
and U19919 (N_19919,N_19435,N_19378);
and U19920 (N_19920,N_19198,N_19201);
or U19921 (N_19921,N_19257,N_19174);
and U19922 (N_19922,N_19201,N_19169);
and U19923 (N_19923,N_19341,N_19471);
nand U19924 (N_19924,N_19313,N_19201);
and U19925 (N_19925,N_19019,N_19204);
nor U19926 (N_19926,N_19398,N_19409);
xor U19927 (N_19927,N_19376,N_19302);
or U19928 (N_19928,N_19337,N_19212);
nor U19929 (N_19929,N_19052,N_19005);
nor U19930 (N_19930,N_19155,N_19135);
nor U19931 (N_19931,N_19098,N_19159);
nor U19932 (N_19932,N_19470,N_19454);
and U19933 (N_19933,N_19355,N_19269);
nor U19934 (N_19934,N_19030,N_19002);
and U19935 (N_19935,N_19466,N_19290);
xnor U19936 (N_19936,N_19356,N_19215);
nand U19937 (N_19937,N_19118,N_19181);
nor U19938 (N_19938,N_19305,N_19046);
or U19939 (N_19939,N_19167,N_19091);
nand U19940 (N_19940,N_19349,N_19393);
nand U19941 (N_19941,N_19110,N_19204);
nor U19942 (N_19942,N_19352,N_19057);
nand U19943 (N_19943,N_19219,N_19428);
nand U19944 (N_19944,N_19353,N_19403);
and U19945 (N_19945,N_19172,N_19018);
or U19946 (N_19946,N_19354,N_19130);
nor U19947 (N_19947,N_19007,N_19372);
and U19948 (N_19948,N_19287,N_19441);
or U19949 (N_19949,N_19480,N_19374);
or U19950 (N_19950,N_19428,N_19425);
nor U19951 (N_19951,N_19336,N_19213);
or U19952 (N_19952,N_19379,N_19290);
or U19953 (N_19953,N_19059,N_19222);
or U19954 (N_19954,N_19326,N_19258);
nand U19955 (N_19955,N_19300,N_19491);
nor U19956 (N_19956,N_19284,N_19387);
and U19957 (N_19957,N_19070,N_19300);
or U19958 (N_19958,N_19380,N_19389);
nor U19959 (N_19959,N_19304,N_19323);
nor U19960 (N_19960,N_19405,N_19023);
xor U19961 (N_19961,N_19390,N_19110);
nand U19962 (N_19962,N_19451,N_19367);
nor U19963 (N_19963,N_19040,N_19257);
nand U19964 (N_19964,N_19093,N_19012);
or U19965 (N_19965,N_19136,N_19013);
nor U19966 (N_19966,N_19272,N_19491);
nor U19967 (N_19967,N_19466,N_19404);
nor U19968 (N_19968,N_19264,N_19167);
and U19969 (N_19969,N_19239,N_19198);
and U19970 (N_19970,N_19265,N_19456);
and U19971 (N_19971,N_19075,N_19087);
xor U19972 (N_19972,N_19219,N_19377);
nor U19973 (N_19973,N_19122,N_19083);
and U19974 (N_19974,N_19149,N_19398);
and U19975 (N_19975,N_19187,N_19223);
xnor U19976 (N_19976,N_19058,N_19211);
nand U19977 (N_19977,N_19075,N_19235);
and U19978 (N_19978,N_19281,N_19150);
or U19979 (N_19979,N_19038,N_19385);
nor U19980 (N_19980,N_19261,N_19155);
and U19981 (N_19981,N_19123,N_19472);
or U19982 (N_19982,N_19459,N_19001);
and U19983 (N_19983,N_19159,N_19386);
nor U19984 (N_19984,N_19013,N_19361);
or U19985 (N_19985,N_19317,N_19312);
and U19986 (N_19986,N_19231,N_19406);
and U19987 (N_19987,N_19111,N_19390);
nand U19988 (N_19988,N_19004,N_19448);
or U19989 (N_19989,N_19445,N_19398);
or U19990 (N_19990,N_19058,N_19264);
and U19991 (N_19991,N_19407,N_19320);
and U19992 (N_19992,N_19488,N_19463);
nor U19993 (N_19993,N_19142,N_19073);
and U19994 (N_19994,N_19464,N_19324);
and U19995 (N_19995,N_19173,N_19494);
nand U19996 (N_19996,N_19392,N_19385);
nand U19997 (N_19997,N_19194,N_19068);
nor U19998 (N_19998,N_19240,N_19430);
and U19999 (N_19999,N_19074,N_19248);
nand U20000 (N_20000,N_19823,N_19801);
and U20001 (N_20001,N_19615,N_19750);
nor U20002 (N_20002,N_19938,N_19623);
or U20003 (N_20003,N_19928,N_19683);
or U20004 (N_20004,N_19996,N_19632);
or U20005 (N_20005,N_19787,N_19713);
nand U20006 (N_20006,N_19723,N_19877);
nand U20007 (N_20007,N_19789,N_19709);
nor U20008 (N_20008,N_19667,N_19951);
nor U20009 (N_20009,N_19721,N_19532);
nand U20010 (N_20010,N_19715,N_19521);
nand U20011 (N_20011,N_19846,N_19635);
or U20012 (N_20012,N_19813,N_19828);
and U20013 (N_20013,N_19871,N_19754);
nand U20014 (N_20014,N_19971,N_19855);
or U20015 (N_20015,N_19516,N_19980);
nor U20016 (N_20016,N_19740,N_19940);
nor U20017 (N_20017,N_19894,N_19743);
nor U20018 (N_20018,N_19729,N_19926);
nor U20019 (N_20019,N_19874,N_19745);
nor U20020 (N_20020,N_19912,N_19949);
nand U20021 (N_20021,N_19941,N_19773);
nor U20022 (N_20022,N_19512,N_19884);
nand U20023 (N_20023,N_19907,N_19782);
nor U20024 (N_20024,N_19785,N_19654);
nand U20025 (N_20025,N_19503,N_19784);
or U20026 (N_20026,N_19880,N_19794);
or U20027 (N_20027,N_19682,N_19933);
nor U20028 (N_20028,N_19681,N_19541);
nand U20029 (N_20029,N_19526,N_19869);
nand U20030 (N_20030,N_19563,N_19589);
and U20031 (N_20031,N_19583,N_19741);
or U20032 (N_20032,N_19889,N_19560);
nand U20033 (N_20033,N_19790,N_19509);
or U20034 (N_20034,N_19712,N_19694);
nand U20035 (N_20035,N_19927,N_19973);
nand U20036 (N_20036,N_19847,N_19539);
nand U20037 (N_20037,N_19964,N_19867);
or U20038 (N_20038,N_19558,N_19738);
nor U20039 (N_20039,N_19525,N_19859);
nand U20040 (N_20040,N_19991,N_19848);
or U20041 (N_20041,N_19751,N_19752);
and U20042 (N_20042,N_19810,N_19691);
or U20043 (N_20043,N_19827,N_19962);
and U20044 (N_20044,N_19625,N_19722);
nor U20045 (N_20045,N_19984,N_19585);
and U20046 (N_20046,N_19868,N_19590);
nor U20047 (N_20047,N_19711,N_19582);
nand U20048 (N_20048,N_19897,N_19976);
or U20049 (N_20049,N_19915,N_19506);
and U20050 (N_20050,N_19699,N_19760);
nor U20051 (N_20051,N_19830,N_19646);
and U20052 (N_20052,N_19770,N_19698);
and U20053 (N_20053,N_19505,N_19580);
xnor U20054 (N_20054,N_19725,N_19831);
nor U20055 (N_20055,N_19955,N_19781);
or U20056 (N_20056,N_19882,N_19579);
nor U20057 (N_20057,N_19766,N_19645);
or U20058 (N_20058,N_19876,N_19661);
and U20059 (N_20059,N_19960,N_19730);
or U20060 (N_20060,N_19815,N_19961);
nor U20061 (N_20061,N_19858,N_19974);
or U20062 (N_20062,N_19975,N_19598);
or U20063 (N_20063,N_19545,N_19764);
and U20064 (N_20064,N_19936,N_19538);
and U20065 (N_20065,N_19557,N_19651);
and U20066 (N_20066,N_19644,N_19888);
xor U20067 (N_20067,N_19826,N_19788);
nor U20068 (N_20068,N_19909,N_19527);
or U20069 (N_20069,N_19688,N_19524);
or U20070 (N_20070,N_19739,N_19686);
or U20071 (N_20071,N_19865,N_19504);
and U20072 (N_20072,N_19786,N_19501);
nor U20073 (N_20073,N_19531,N_19900);
or U20074 (N_20074,N_19844,N_19954);
or U20075 (N_20075,N_19696,N_19717);
and U20076 (N_20076,N_19779,N_19817);
nor U20077 (N_20077,N_19919,N_19614);
nand U20078 (N_20078,N_19604,N_19736);
or U20079 (N_20079,N_19547,N_19780);
nor U20080 (N_20080,N_19668,N_19576);
nor U20081 (N_20081,N_19612,N_19596);
nand U20082 (N_20082,N_19594,N_19956);
nor U20083 (N_20083,N_19633,N_19553);
nor U20084 (N_20084,N_19600,N_19591);
nand U20085 (N_20085,N_19572,N_19845);
nand U20086 (N_20086,N_19670,N_19957);
or U20087 (N_20087,N_19536,N_19890);
nand U20088 (N_20088,N_19842,N_19966);
nor U20089 (N_20089,N_19514,N_19999);
or U20090 (N_20090,N_19925,N_19673);
nor U20091 (N_20091,N_19837,N_19684);
or U20092 (N_20092,N_19567,N_19692);
nand U20093 (N_20093,N_19613,N_19735);
nor U20094 (N_20094,N_19647,N_19593);
nand U20095 (N_20095,N_19573,N_19737);
or U20096 (N_20096,N_19861,N_19706);
nor U20097 (N_20097,N_19854,N_19948);
and U20098 (N_20098,N_19893,N_19913);
nor U20099 (N_20099,N_19914,N_19978);
nor U20100 (N_20100,N_19908,N_19977);
nand U20101 (N_20101,N_19822,N_19998);
nand U20102 (N_20102,N_19551,N_19638);
nor U20103 (N_20103,N_19758,N_19626);
and U20104 (N_20104,N_19648,N_19838);
and U20105 (N_20105,N_19857,N_19814);
nor U20106 (N_20106,N_19552,N_19548);
nor U20107 (N_20107,N_19641,N_19860);
and U20108 (N_20108,N_19881,N_19771);
or U20109 (N_20109,N_19829,N_19783);
nor U20110 (N_20110,N_19533,N_19762);
nor U20111 (N_20111,N_19719,N_19849);
nand U20112 (N_20112,N_19664,N_19995);
and U20113 (N_20113,N_19796,N_19963);
or U20114 (N_20114,N_19507,N_19929);
and U20115 (N_20115,N_19522,N_19839);
and U20116 (N_20116,N_19776,N_19834);
nor U20117 (N_20117,N_19566,N_19609);
and U20118 (N_20118,N_19875,N_19791);
and U20119 (N_20119,N_19901,N_19989);
nor U20120 (N_20120,N_19918,N_19685);
nand U20121 (N_20121,N_19852,N_19958);
and U20122 (N_20122,N_19990,N_19768);
nor U20123 (N_20123,N_19595,N_19569);
and U20124 (N_20124,N_19879,N_19746);
or U20125 (N_20125,N_19643,N_19680);
and U20126 (N_20126,N_19666,N_19602);
and U20127 (N_20127,N_19800,N_19803);
nor U20128 (N_20128,N_19759,N_19732);
xnor U20129 (N_20129,N_19820,N_19697);
nand U20130 (N_20130,N_19708,N_19693);
nand U20131 (N_20131,N_19904,N_19703);
or U20132 (N_20132,N_19657,N_19825);
xnor U20133 (N_20133,N_19959,N_19924);
or U20134 (N_20134,N_19891,N_19931);
nor U20135 (N_20135,N_19777,N_19588);
nor U20136 (N_20136,N_19578,N_19607);
nor U20137 (N_20137,N_19523,N_19559);
and U20138 (N_20138,N_19610,N_19833);
nand U20139 (N_20139,N_19902,N_19679);
nor U20140 (N_20140,N_19639,N_19898);
nand U20141 (N_20141,N_19674,N_19749);
or U20142 (N_20142,N_19671,N_19608);
or U20143 (N_20143,N_19658,N_19896);
and U20144 (N_20144,N_19716,N_19528);
xnor U20145 (N_20145,N_19795,N_19985);
or U20146 (N_20146,N_19581,N_19793);
and U20147 (N_20147,N_19627,N_19701);
nor U20148 (N_20148,N_19519,N_19618);
and U20149 (N_20149,N_19747,N_19952);
nand U20150 (N_20150,N_19836,N_19887);
or U20151 (N_20151,N_19606,N_19910);
and U20152 (N_20152,N_19630,N_19689);
nor U20153 (N_20153,N_19763,N_19944);
and U20154 (N_20154,N_19702,N_19953);
or U20155 (N_20155,N_19824,N_19932);
or U20156 (N_20156,N_19850,N_19634);
nand U20157 (N_20157,N_19575,N_19744);
nor U20158 (N_20158,N_19895,N_19775);
or U20159 (N_20159,N_19549,N_19637);
or U20160 (N_20160,N_19798,N_19577);
or U20161 (N_20161,N_19508,N_19947);
nand U20162 (N_20162,N_19562,N_19946);
or U20163 (N_20163,N_19676,N_19631);
and U20164 (N_20164,N_19642,N_19731);
and U20165 (N_20165,N_19979,N_19772);
or U20166 (N_20166,N_19917,N_19905);
and U20167 (N_20167,N_19544,N_19565);
nor U20168 (N_20168,N_19540,N_19678);
and U20169 (N_20169,N_19930,N_19943);
nor U20170 (N_20170,N_19568,N_19530);
and U20171 (N_20171,N_19811,N_19864);
xor U20172 (N_20172,N_19601,N_19517);
nand U20173 (N_20173,N_19714,N_19866);
nand U20174 (N_20174,N_19659,N_19767);
or U20175 (N_20175,N_19605,N_19535);
and U20176 (N_20176,N_19804,N_19599);
and U20177 (N_20177,N_19921,N_19862);
or U20178 (N_20178,N_19624,N_19677);
nand U20179 (N_20179,N_19835,N_19856);
or U20180 (N_20180,N_19650,N_19853);
nand U20181 (N_20181,N_19660,N_19537);
nand U20182 (N_20182,N_19863,N_19797);
or U20183 (N_20183,N_19942,N_19570);
nand U20184 (N_20184,N_19808,N_19872);
nor U20185 (N_20185,N_19653,N_19983);
and U20186 (N_20186,N_19704,N_19982);
nand U20187 (N_20187,N_19621,N_19500);
and U20188 (N_20188,N_19748,N_19923);
nor U20189 (N_20189,N_19733,N_19669);
or U20190 (N_20190,N_19756,N_19640);
nor U20191 (N_20191,N_19520,N_19922);
and U20192 (N_20192,N_19807,N_19970);
xor U20193 (N_20193,N_19916,N_19753);
nor U20194 (N_20194,N_19755,N_19769);
xnor U20195 (N_20195,N_19662,N_19886);
or U20196 (N_20196,N_19611,N_19710);
nand U20197 (N_20197,N_19529,N_19665);
nor U20198 (N_20198,N_19988,N_19718);
or U20199 (N_20199,N_19550,N_19802);
nand U20200 (N_20200,N_19792,N_19554);
or U20201 (N_20201,N_19597,N_19812);
or U20202 (N_20202,N_19742,N_19878);
and U20203 (N_20203,N_19841,N_19799);
or U20204 (N_20204,N_19840,N_19816);
and U20205 (N_20205,N_19513,N_19726);
and U20206 (N_20206,N_19720,N_19656);
or U20207 (N_20207,N_19972,N_19851);
and U20208 (N_20208,N_19965,N_19636);
nand U20209 (N_20209,N_19655,N_19761);
nor U20210 (N_20210,N_19906,N_19968);
nand U20211 (N_20211,N_19690,N_19993);
or U20212 (N_20212,N_19546,N_19652);
nand U20213 (N_20213,N_19727,N_19707);
nor U20214 (N_20214,N_19571,N_19700);
or U20215 (N_20215,N_19903,N_19969);
nor U20216 (N_20216,N_19987,N_19832);
nor U20217 (N_20217,N_19778,N_19809);
and U20218 (N_20218,N_19561,N_19883);
or U20219 (N_20219,N_19873,N_19510);
nand U20220 (N_20220,N_19911,N_19518);
and U20221 (N_20221,N_19805,N_19843);
xor U20222 (N_20222,N_19821,N_19728);
nor U20223 (N_20223,N_19672,N_19986);
and U20224 (N_20224,N_19734,N_19534);
nand U20225 (N_20225,N_19620,N_19649);
xor U20226 (N_20226,N_19997,N_19870);
or U20227 (N_20227,N_19586,N_19555);
nor U20228 (N_20228,N_19939,N_19592);
or U20229 (N_20229,N_19935,N_19628);
nand U20230 (N_20230,N_19818,N_19705);
or U20231 (N_20231,N_19967,N_19515);
nor U20232 (N_20232,N_19950,N_19502);
or U20233 (N_20233,N_19695,N_19574);
or U20234 (N_20234,N_19757,N_19603);
and U20235 (N_20235,N_19587,N_19675);
nand U20236 (N_20236,N_19994,N_19806);
and U20237 (N_20237,N_19542,N_19663);
and U20238 (N_20238,N_19937,N_19687);
and U20239 (N_20239,N_19617,N_19934);
xnor U20240 (N_20240,N_19584,N_19981);
or U20241 (N_20241,N_19622,N_19892);
nor U20242 (N_20242,N_19920,N_19945);
nand U20243 (N_20243,N_19819,N_19885);
and U20244 (N_20244,N_19619,N_19724);
nor U20245 (N_20245,N_19543,N_19774);
and U20246 (N_20246,N_19992,N_19556);
or U20247 (N_20247,N_19629,N_19899);
nand U20248 (N_20248,N_19765,N_19616);
nand U20249 (N_20249,N_19511,N_19564);
nor U20250 (N_20250,N_19852,N_19670);
or U20251 (N_20251,N_19836,N_19823);
or U20252 (N_20252,N_19911,N_19744);
nor U20253 (N_20253,N_19662,N_19893);
nand U20254 (N_20254,N_19563,N_19700);
and U20255 (N_20255,N_19770,N_19776);
or U20256 (N_20256,N_19974,N_19835);
or U20257 (N_20257,N_19727,N_19672);
nand U20258 (N_20258,N_19677,N_19824);
nor U20259 (N_20259,N_19725,N_19917);
nand U20260 (N_20260,N_19756,N_19959);
nand U20261 (N_20261,N_19532,N_19510);
nand U20262 (N_20262,N_19786,N_19666);
and U20263 (N_20263,N_19833,N_19982);
nand U20264 (N_20264,N_19526,N_19893);
and U20265 (N_20265,N_19710,N_19551);
and U20266 (N_20266,N_19918,N_19550);
nand U20267 (N_20267,N_19675,N_19919);
and U20268 (N_20268,N_19865,N_19732);
or U20269 (N_20269,N_19943,N_19634);
or U20270 (N_20270,N_19644,N_19765);
nand U20271 (N_20271,N_19831,N_19973);
nand U20272 (N_20272,N_19788,N_19538);
and U20273 (N_20273,N_19994,N_19906);
and U20274 (N_20274,N_19633,N_19770);
nand U20275 (N_20275,N_19620,N_19833);
nand U20276 (N_20276,N_19500,N_19735);
nand U20277 (N_20277,N_19517,N_19933);
or U20278 (N_20278,N_19655,N_19691);
nand U20279 (N_20279,N_19970,N_19827);
nand U20280 (N_20280,N_19787,N_19720);
nor U20281 (N_20281,N_19850,N_19753);
nand U20282 (N_20282,N_19750,N_19737);
nand U20283 (N_20283,N_19849,N_19865);
and U20284 (N_20284,N_19773,N_19775);
nand U20285 (N_20285,N_19893,N_19639);
nand U20286 (N_20286,N_19501,N_19613);
nor U20287 (N_20287,N_19761,N_19856);
and U20288 (N_20288,N_19851,N_19980);
and U20289 (N_20289,N_19608,N_19693);
or U20290 (N_20290,N_19970,N_19706);
nor U20291 (N_20291,N_19888,N_19521);
or U20292 (N_20292,N_19874,N_19520);
and U20293 (N_20293,N_19610,N_19680);
nor U20294 (N_20294,N_19829,N_19788);
nor U20295 (N_20295,N_19652,N_19922);
and U20296 (N_20296,N_19670,N_19866);
nor U20297 (N_20297,N_19589,N_19531);
nor U20298 (N_20298,N_19759,N_19950);
nor U20299 (N_20299,N_19814,N_19994);
and U20300 (N_20300,N_19640,N_19679);
or U20301 (N_20301,N_19829,N_19612);
and U20302 (N_20302,N_19744,N_19933);
or U20303 (N_20303,N_19847,N_19554);
and U20304 (N_20304,N_19533,N_19726);
and U20305 (N_20305,N_19998,N_19997);
nand U20306 (N_20306,N_19880,N_19833);
nor U20307 (N_20307,N_19547,N_19731);
nor U20308 (N_20308,N_19557,N_19738);
or U20309 (N_20309,N_19636,N_19592);
or U20310 (N_20310,N_19727,N_19987);
and U20311 (N_20311,N_19534,N_19557);
or U20312 (N_20312,N_19947,N_19813);
nand U20313 (N_20313,N_19579,N_19919);
xnor U20314 (N_20314,N_19588,N_19657);
nor U20315 (N_20315,N_19882,N_19517);
or U20316 (N_20316,N_19933,N_19579);
or U20317 (N_20317,N_19936,N_19542);
nor U20318 (N_20318,N_19913,N_19683);
nor U20319 (N_20319,N_19856,N_19653);
nor U20320 (N_20320,N_19644,N_19875);
and U20321 (N_20321,N_19905,N_19647);
nand U20322 (N_20322,N_19595,N_19844);
or U20323 (N_20323,N_19654,N_19863);
and U20324 (N_20324,N_19600,N_19889);
or U20325 (N_20325,N_19511,N_19551);
and U20326 (N_20326,N_19851,N_19979);
or U20327 (N_20327,N_19930,N_19773);
or U20328 (N_20328,N_19616,N_19931);
nand U20329 (N_20329,N_19590,N_19833);
and U20330 (N_20330,N_19709,N_19684);
nand U20331 (N_20331,N_19534,N_19932);
nand U20332 (N_20332,N_19893,N_19954);
nor U20333 (N_20333,N_19995,N_19826);
nor U20334 (N_20334,N_19949,N_19634);
nand U20335 (N_20335,N_19774,N_19604);
nand U20336 (N_20336,N_19812,N_19765);
nand U20337 (N_20337,N_19761,N_19944);
or U20338 (N_20338,N_19900,N_19526);
and U20339 (N_20339,N_19597,N_19949);
nand U20340 (N_20340,N_19577,N_19927);
and U20341 (N_20341,N_19914,N_19599);
nand U20342 (N_20342,N_19815,N_19645);
nand U20343 (N_20343,N_19980,N_19603);
and U20344 (N_20344,N_19935,N_19561);
and U20345 (N_20345,N_19841,N_19672);
nand U20346 (N_20346,N_19578,N_19992);
and U20347 (N_20347,N_19898,N_19522);
nor U20348 (N_20348,N_19884,N_19964);
nand U20349 (N_20349,N_19862,N_19845);
nor U20350 (N_20350,N_19809,N_19844);
or U20351 (N_20351,N_19899,N_19817);
and U20352 (N_20352,N_19945,N_19826);
and U20353 (N_20353,N_19715,N_19934);
nand U20354 (N_20354,N_19729,N_19962);
and U20355 (N_20355,N_19604,N_19914);
nand U20356 (N_20356,N_19998,N_19857);
nor U20357 (N_20357,N_19575,N_19603);
or U20358 (N_20358,N_19683,N_19700);
nor U20359 (N_20359,N_19800,N_19608);
and U20360 (N_20360,N_19536,N_19648);
xnor U20361 (N_20361,N_19523,N_19637);
and U20362 (N_20362,N_19739,N_19798);
nor U20363 (N_20363,N_19929,N_19706);
nand U20364 (N_20364,N_19510,N_19982);
nand U20365 (N_20365,N_19750,N_19863);
xnor U20366 (N_20366,N_19671,N_19963);
nand U20367 (N_20367,N_19802,N_19751);
or U20368 (N_20368,N_19539,N_19549);
and U20369 (N_20369,N_19568,N_19977);
nand U20370 (N_20370,N_19679,N_19553);
and U20371 (N_20371,N_19742,N_19948);
nand U20372 (N_20372,N_19994,N_19609);
or U20373 (N_20373,N_19800,N_19581);
and U20374 (N_20374,N_19787,N_19754);
or U20375 (N_20375,N_19929,N_19573);
nand U20376 (N_20376,N_19930,N_19676);
and U20377 (N_20377,N_19980,N_19915);
or U20378 (N_20378,N_19750,N_19789);
nand U20379 (N_20379,N_19585,N_19663);
nand U20380 (N_20380,N_19863,N_19672);
nand U20381 (N_20381,N_19702,N_19510);
and U20382 (N_20382,N_19583,N_19652);
nor U20383 (N_20383,N_19621,N_19662);
and U20384 (N_20384,N_19934,N_19515);
and U20385 (N_20385,N_19970,N_19544);
nor U20386 (N_20386,N_19526,N_19622);
or U20387 (N_20387,N_19792,N_19773);
nor U20388 (N_20388,N_19783,N_19960);
xnor U20389 (N_20389,N_19598,N_19806);
nor U20390 (N_20390,N_19865,N_19772);
xor U20391 (N_20391,N_19704,N_19549);
and U20392 (N_20392,N_19898,N_19765);
or U20393 (N_20393,N_19567,N_19541);
or U20394 (N_20394,N_19950,N_19793);
nand U20395 (N_20395,N_19553,N_19617);
or U20396 (N_20396,N_19508,N_19869);
or U20397 (N_20397,N_19926,N_19706);
or U20398 (N_20398,N_19803,N_19752);
or U20399 (N_20399,N_19611,N_19852);
nor U20400 (N_20400,N_19759,N_19588);
nor U20401 (N_20401,N_19620,N_19559);
and U20402 (N_20402,N_19673,N_19540);
nand U20403 (N_20403,N_19651,N_19638);
nand U20404 (N_20404,N_19888,N_19527);
and U20405 (N_20405,N_19783,N_19549);
nor U20406 (N_20406,N_19724,N_19557);
and U20407 (N_20407,N_19550,N_19564);
nand U20408 (N_20408,N_19861,N_19643);
and U20409 (N_20409,N_19576,N_19956);
or U20410 (N_20410,N_19896,N_19600);
nor U20411 (N_20411,N_19973,N_19830);
and U20412 (N_20412,N_19801,N_19607);
or U20413 (N_20413,N_19897,N_19935);
or U20414 (N_20414,N_19740,N_19814);
nand U20415 (N_20415,N_19747,N_19999);
nor U20416 (N_20416,N_19860,N_19903);
nor U20417 (N_20417,N_19837,N_19563);
or U20418 (N_20418,N_19541,N_19895);
nor U20419 (N_20419,N_19741,N_19884);
or U20420 (N_20420,N_19536,N_19668);
nand U20421 (N_20421,N_19684,N_19949);
nand U20422 (N_20422,N_19801,N_19989);
or U20423 (N_20423,N_19690,N_19702);
nand U20424 (N_20424,N_19882,N_19606);
or U20425 (N_20425,N_19863,N_19980);
or U20426 (N_20426,N_19768,N_19558);
or U20427 (N_20427,N_19972,N_19815);
or U20428 (N_20428,N_19782,N_19755);
or U20429 (N_20429,N_19618,N_19834);
nor U20430 (N_20430,N_19536,N_19702);
or U20431 (N_20431,N_19545,N_19635);
or U20432 (N_20432,N_19918,N_19572);
or U20433 (N_20433,N_19688,N_19931);
nor U20434 (N_20434,N_19650,N_19796);
and U20435 (N_20435,N_19987,N_19509);
nor U20436 (N_20436,N_19885,N_19514);
nand U20437 (N_20437,N_19612,N_19837);
nor U20438 (N_20438,N_19866,N_19758);
nand U20439 (N_20439,N_19784,N_19667);
nor U20440 (N_20440,N_19690,N_19633);
nor U20441 (N_20441,N_19941,N_19947);
or U20442 (N_20442,N_19854,N_19708);
nor U20443 (N_20443,N_19638,N_19586);
and U20444 (N_20444,N_19797,N_19529);
nor U20445 (N_20445,N_19501,N_19939);
or U20446 (N_20446,N_19735,N_19638);
nand U20447 (N_20447,N_19692,N_19776);
nor U20448 (N_20448,N_19725,N_19530);
nand U20449 (N_20449,N_19780,N_19947);
xnor U20450 (N_20450,N_19521,N_19909);
or U20451 (N_20451,N_19524,N_19960);
and U20452 (N_20452,N_19667,N_19691);
or U20453 (N_20453,N_19642,N_19719);
or U20454 (N_20454,N_19705,N_19672);
or U20455 (N_20455,N_19839,N_19582);
and U20456 (N_20456,N_19767,N_19780);
or U20457 (N_20457,N_19577,N_19721);
nor U20458 (N_20458,N_19740,N_19644);
nor U20459 (N_20459,N_19677,N_19556);
or U20460 (N_20460,N_19767,N_19616);
and U20461 (N_20461,N_19761,N_19635);
or U20462 (N_20462,N_19525,N_19687);
nor U20463 (N_20463,N_19957,N_19511);
and U20464 (N_20464,N_19667,N_19858);
and U20465 (N_20465,N_19709,N_19974);
nand U20466 (N_20466,N_19653,N_19768);
and U20467 (N_20467,N_19520,N_19957);
and U20468 (N_20468,N_19816,N_19755);
and U20469 (N_20469,N_19647,N_19801);
and U20470 (N_20470,N_19947,N_19811);
and U20471 (N_20471,N_19552,N_19930);
nand U20472 (N_20472,N_19984,N_19575);
or U20473 (N_20473,N_19598,N_19888);
and U20474 (N_20474,N_19932,N_19524);
xor U20475 (N_20475,N_19636,N_19702);
and U20476 (N_20476,N_19648,N_19908);
nor U20477 (N_20477,N_19515,N_19707);
nor U20478 (N_20478,N_19590,N_19777);
and U20479 (N_20479,N_19648,N_19640);
nand U20480 (N_20480,N_19625,N_19743);
nor U20481 (N_20481,N_19533,N_19928);
nand U20482 (N_20482,N_19730,N_19824);
or U20483 (N_20483,N_19763,N_19911);
or U20484 (N_20484,N_19693,N_19914);
nor U20485 (N_20485,N_19803,N_19878);
and U20486 (N_20486,N_19814,N_19805);
nand U20487 (N_20487,N_19637,N_19589);
and U20488 (N_20488,N_19665,N_19902);
nand U20489 (N_20489,N_19568,N_19523);
and U20490 (N_20490,N_19791,N_19569);
nor U20491 (N_20491,N_19943,N_19775);
xor U20492 (N_20492,N_19803,N_19599);
and U20493 (N_20493,N_19720,N_19901);
xnor U20494 (N_20494,N_19851,N_19683);
nor U20495 (N_20495,N_19677,N_19944);
and U20496 (N_20496,N_19855,N_19535);
nand U20497 (N_20497,N_19916,N_19680);
or U20498 (N_20498,N_19509,N_19989);
nand U20499 (N_20499,N_19926,N_19762);
or U20500 (N_20500,N_20251,N_20045);
nor U20501 (N_20501,N_20041,N_20082);
nor U20502 (N_20502,N_20232,N_20153);
nor U20503 (N_20503,N_20217,N_20197);
or U20504 (N_20504,N_20346,N_20319);
nor U20505 (N_20505,N_20342,N_20241);
nand U20506 (N_20506,N_20073,N_20284);
nor U20507 (N_20507,N_20084,N_20499);
nor U20508 (N_20508,N_20252,N_20010);
nand U20509 (N_20509,N_20490,N_20332);
or U20510 (N_20510,N_20293,N_20440);
nand U20511 (N_20511,N_20442,N_20489);
and U20512 (N_20512,N_20340,N_20072);
nor U20513 (N_20513,N_20020,N_20096);
nand U20514 (N_20514,N_20427,N_20180);
or U20515 (N_20515,N_20231,N_20331);
nor U20516 (N_20516,N_20362,N_20249);
and U20517 (N_20517,N_20250,N_20453);
and U20518 (N_20518,N_20071,N_20076);
nand U20519 (N_20519,N_20289,N_20156);
nor U20520 (N_20520,N_20439,N_20060);
nor U20521 (N_20521,N_20123,N_20182);
and U20522 (N_20522,N_20325,N_20097);
nor U20523 (N_20523,N_20168,N_20318);
and U20524 (N_20524,N_20124,N_20240);
or U20525 (N_20525,N_20074,N_20094);
and U20526 (N_20526,N_20167,N_20066);
nand U20527 (N_20527,N_20134,N_20027);
and U20528 (N_20528,N_20353,N_20037);
or U20529 (N_20529,N_20000,N_20397);
or U20530 (N_20530,N_20237,N_20107);
nor U20531 (N_20531,N_20430,N_20015);
and U20532 (N_20532,N_20266,N_20159);
nand U20533 (N_20533,N_20229,N_20456);
nand U20534 (N_20534,N_20478,N_20095);
nand U20535 (N_20535,N_20259,N_20109);
or U20536 (N_20536,N_20447,N_20272);
nand U20537 (N_20537,N_20407,N_20279);
nor U20538 (N_20538,N_20363,N_20401);
nor U20539 (N_20539,N_20092,N_20434);
nor U20540 (N_20540,N_20145,N_20437);
and U20541 (N_20541,N_20222,N_20150);
nand U20542 (N_20542,N_20466,N_20303);
and U20543 (N_20543,N_20221,N_20343);
and U20544 (N_20544,N_20461,N_20006);
nand U20545 (N_20545,N_20421,N_20496);
nand U20546 (N_20546,N_20174,N_20330);
and U20547 (N_20547,N_20358,N_20425);
nand U20548 (N_20548,N_20223,N_20283);
nand U20549 (N_20549,N_20355,N_20179);
nand U20550 (N_20550,N_20133,N_20458);
nand U20551 (N_20551,N_20028,N_20274);
or U20552 (N_20552,N_20139,N_20012);
nor U20553 (N_20553,N_20151,N_20183);
and U20554 (N_20554,N_20031,N_20239);
or U20555 (N_20555,N_20386,N_20416);
or U20556 (N_20556,N_20374,N_20347);
nand U20557 (N_20557,N_20409,N_20454);
or U20558 (N_20558,N_20101,N_20307);
nor U20559 (N_20559,N_20310,N_20469);
nor U20560 (N_20560,N_20317,N_20192);
nand U20561 (N_20561,N_20057,N_20457);
or U20562 (N_20562,N_20468,N_20312);
and U20563 (N_20563,N_20455,N_20413);
or U20564 (N_20564,N_20308,N_20149);
nand U20565 (N_20565,N_20043,N_20494);
or U20566 (N_20566,N_20138,N_20282);
and U20567 (N_20567,N_20193,N_20281);
nand U20568 (N_20568,N_20077,N_20210);
or U20569 (N_20569,N_20121,N_20117);
or U20570 (N_20570,N_20388,N_20287);
nand U20571 (N_20571,N_20286,N_20370);
xnor U20572 (N_20572,N_20230,N_20474);
nand U20573 (N_20573,N_20088,N_20099);
nor U20574 (N_20574,N_20364,N_20127);
and U20575 (N_20575,N_20053,N_20348);
xor U20576 (N_20576,N_20324,N_20214);
nor U20577 (N_20577,N_20414,N_20067);
nor U20578 (N_20578,N_20435,N_20335);
and U20579 (N_20579,N_20248,N_20018);
or U20580 (N_20580,N_20079,N_20497);
or U20581 (N_20581,N_20322,N_20482);
and U20582 (N_20582,N_20298,N_20218);
xor U20583 (N_20583,N_20056,N_20061);
or U20584 (N_20584,N_20026,N_20175);
nand U20585 (N_20585,N_20338,N_20211);
nand U20586 (N_20586,N_20372,N_20431);
nor U20587 (N_20587,N_20017,N_20022);
or U20588 (N_20588,N_20140,N_20013);
and U20589 (N_20589,N_20294,N_20024);
nor U20590 (N_20590,N_20147,N_20445);
and U20591 (N_20591,N_20273,N_20007);
nor U20592 (N_20592,N_20339,N_20023);
nor U20593 (N_20593,N_20379,N_20002);
nand U20594 (N_20594,N_20393,N_20129);
nor U20595 (N_20595,N_20306,N_20199);
nand U20596 (N_20596,N_20064,N_20128);
nand U20597 (N_20597,N_20297,N_20090);
nand U20598 (N_20598,N_20087,N_20100);
or U20599 (N_20599,N_20464,N_20394);
or U20600 (N_20600,N_20450,N_20344);
nor U20601 (N_20601,N_20313,N_20033);
nor U20602 (N_20602,N_20070,N_20201);
nor U20603 (N_20603,N_20253,N_20428);
or U20604 (N_20604,N_20387,N_20368);
and U20605 (N_20605,N_20349,N_20051);
nor U20606 (N_20606,N_20004,N_20467);
nor U20607 (N_20607,N_20419,N_20327);
and U20608 (N_20608,N_20137,N_20276);
xor U20609 (N_20609,N_20102,N_20224);
nand U20610 (N_20610,N_20268,N_20191);
nor U20611 (N_20611,N_20110,N_20219);
nand U20612 (N_20612,N_20126,N_20333);
and U20613 (N_20613,N_20448,N_20105);
nor U20614 (N_20614,N_20131,N_20380);
or U20615 (N_20615,N_20366,N_20446);
and U20616 (N_20616,N_20198,N_20400);
nor U20617 (N_20617,N_20350,N_20390);
nor U20618 (N_20618,N_20356,N_20106);
or U20619 (N_20619,N_20142,N_20001);
nand U20620 (N_20620,N_20481,N_20032);
and U20621 (N_20621,N_20204,N_20256);
nand U20622 (N_20622,N_20163,N_20408);
and U20623 (N_20623,N_20058,N_20049);
or U20624 (N_20624,N_20047,N_20475);
and U20625 (N_20625,N_20209,N_20185);
nor U20626 (N_20626,N_20311,N_20227);
nor U20627 (N_20627,N_20225,N_20143);
and U20628 (N_20628,N_20320,N_20112);
nor U20629 (N_20629,N_20176,N_20396);
nand U20630 (N_20630,N_20295,N_20011);
and U20631 (N_20631,N_20405,N_20271);
and U20632 (N_20632,N_20257,N_20038);
or U20633 (N_20633,N_20173,N_20114);
or U20634 (N_20634,N_20395,N_20054);
and U20635 (N_20635,N_20152,N_20236);
nand U20636 (N_20636,N_20459,N_20476);
and U20637 (N_20637,N_20378,N_20415);
nand U20638 (N_20638,N_20160,N_20234);
nand U20639 (N_20639,N_20495,N_20177);
nor U20640 (N_20640,N_20411,N_20208);
nand U20641 (N_20641,N_20086,N_20277);
nor U20642 (N_20642,N_20423,N_20055);
and U20643 (N_20643,N_20429,N_20161);
nor U20644 (N_20644,N_20019,N_20108);
or U20645 (N_20645,N_20063,N_20089);
nor U20646 (N_20646,N_20433,N_20323);
or U20647 (N_20647,N_20369,N_20361);
nor U20648 (N_20648,N_20169,N_20166);
nor U20649 (N_20649,N_20334,N_20288);
nor U20650 (N_20650,N_20016,N_20228);
or U20651 (N_20651,N_20202,N_20402);
and U20652 (N_20652,N_20215,N_20039);
or U20653 (N_20653,N_20357,N_20203);
nand U20654 (N_20654,N_20399,N_20068);
nand U20655 (N_20655,N_20465,N_20200);
nand U20656 (N_20656,N_20485,N_20091);
or U20657 (N_20657,N_20170,N_20498);
or U20658 (N_20658,N_20492,N_20119);
and U20659 (N_20659,N_20008,N_20292);
nor U20660 (N_20660,N_20212,N_20487);
nand U20661 (N_20661,N_20162,N_20014);
or U20662 (N_20662,N_20491,N_20261);
and U20663 (N_20663,N_20462,N_20029);
xnor U20664 (N_20664,N_20085,N_20300);
xor U20665 (N_20665,N_20235,N_20329);
nor U20666 (N_20666,N_20264,N_20144);
and U20667 (N_20667,N_20280,N_20044);
nor U20668 (N_20668,N_20477,N_20354);
nor U20669 (N_20669,N_20098,N_20424);
nor U20670 (N_20670,N_20403,N_20412);
or U20671 (N_20671,N_20243,N_20392);
or U20672 (N_20672,N_20238,N_20165);
nand U20673 (N_20673,N_20410,N_20195);
or U20674 (N_20674,N_20304,N_20036);
nand U20675 (N_20675,N_20113,N_20296);
nor U20676 (N_20676,N_20463,N_20065);
and U20677 (N_20677,N_20417,N_20135);
nand U20678 (N_20678,N_20420,N_20486);
and U20679 (N_20679,N_20377,N_20194);
and U20680 (N_20680,N_20233,N_20207);
and U20681 (N_20681,N_20385,N_20383);
or U20682 (N_20682,N_20050,N_20326);
and U20683 (N_20683,N_20367,N_20484);
nor U20684 (N_20684,N_20205,N_20472);
nand U20685 (N_20685,N_20365,N_20115);
nor U20686 (N_20686,N_20125,N_20321);
and U20687 (N_20687,N_20042,N_20184);
nor U20688 (N_20688,N_20040,N_20216);
nand U20689 (N_20689,N_20375,N_20181);
nor U20690 (N_20690,N_20360,N_20245);
nand U20691 (N_20691,N_20480,N_20172);
nand U20692 (N_20692,N_20220,N_20336);
and U20693 (N_20693,N_20473,N_20267);
nand U20694 (N_20694,N_20493,N_20158);
nand U20695 (N_20695,N_20132,N_20422);
or U20696 (N_20696,N_20285,N_20406);
and U20697 (N_20697,N_20328,N_20009);
and U20698 (N_20698,N_20255,N_20382);
and U20699 (N_20699,N_20302,N_20141);
nor U20700 (N_20700,N_20451,N_20483);
nand U20701 (N_20701,N_20146,N_20337);
or U20702 (N_20702,N_20025,N_20080);
nor U20703 (N_20703,N_20265,N_20404);
nor U20704 (N_20704,N_20188,N_20301);
nand U20705 (N_20705,N_20116,N_20371);
nand U20706 (N_20706,N_20178,N_20263);
and U20707 (N_20707,N_20103,N_20242);
nand U20708 (N_20708,N_20035,N_20305);
and U20709 (N_20709,N_20470,N_20190);
or U20710 (N_20710,N_20075,N_20488);
nand U20711 (N_20711,N_20093,N_20046);
and U20712 (N_20712,N_20426,N_20246);
and U20713 (N_20713,N_20111,N_20315);
and U20714 (N_20714,N_20130,N_20436);
nor U20715 (N_20715,N_20021,N_20290);
nand U20716 (N_20716,N_20003,N_20314);
nor U20717 (N_20717,N_20244,N_20262);
and U20718 (N_20718,N_20258,N_20062);
nor U20719 (N_20719,N_20059,N_20005);
nor U20720 (N_20720,N_20275,N_20376);
or U20721 (N_20721,N_20391,N_20270);
or U20722 (N_20722,N_20048,N_20030);
xor U20723 (N_20723,N_20247,N_20345);
xnor U20724 (N_20724,N_20171,N_20254);
nor U20725 (N_20725,N_20206,N_20352);
nand U20726 (N_20726,N_20226,N_20381);
nand U20727 (N_20727,N_20081,N_20299);
or U20728 (N_20728,N_20432,N_20316);
and U20729 (N_20729,N_20452,N_20341);
and U20730 (N_20730,N_20157,N_20155);
and U20731 (N_20731,N_20154,N_20118);
and U20732 (N_20732,N_20120,N_20136);
and U20733 (N_20733,N_20479,N_20260);
nand U20734 (N_20734,N_20389,N_20034);
or U20735 (N_20735,N_20398,N_20384);
nand U20736 (N_20736,N_20291,N_20052);
or U20737 (N_20737,N_20122,N_20189);
nand U20738 (N_20738,N_20460,N_20418);
nor U20739 (N_20739,N_20187,N_20164);
nor U20740 (N_20740,N_20186,N_20443);
and U20741 (N_20741,N_20278,N_20471);
or U20742 (N_20742,N_20309,N_20083);
nor U20743 (N_20743,N_20213,N_20078);
and U20744 (N_20744,N_20449,N_20351);
nor U20745 (N_20745,N_20444,N_20148);
nand U20746 (N_20746,N_20269,N_20069);
and U20747 (N_20747,N_20196,N_20359);
or U20748 (N_20748,N_20438,N_20373);
or U20749 (N_20749,N_20104,N_20441);
nor U20750 (N_20750,N_20047,N_20431);
and U20751 (N_20751,N_20180,N_20437);
and U20752 (N_20752,N_20032,N_20249);
nand U20753 (N_20753,N_20348,N_20378);
or U20754 (N_20754,N_20450,N_20439);
nor U20755 (N_20755,N_20283,N_20435);
and U20756 (N_20756,N_20003,N_20367);
nand U20757 (N_20757,N_20240,N_20144);
or U20758 (N_20758,N_20433,N_20233);
or U20759 (N_20759,N_20186,N_20384);
xor U20760 (N_20760,N_20143,N_20461);
and U20761 (N_20761,N_20060,N_20180);
or U20762 (N_20762,N_20191,N_20474);
or U20763 (N_20763,N_20104,N_20244);
xor U20764 (N_20764,N_20132,N_20243);
or U20765 (N_20765,N_20188,N_20190);
nor U20766 (N_20766,N_20243,N_20206);
or U20767 (N_20767,N_20221,N_20140);
and U20768 (N_20768,N_20354,N_20268);
nor U20769 (N_20769,N_20151,N_20309);
or U20770 (N_20770,N_20457,N_20331);
and U20771 (N_20771,N_20465,N_20450);
and U20772 (N_20772,N_20209,N_20176);
or U20773 (N_20773,N_20429,N_20451);
nor U20774 (N_20774,N_20112,N_20188);
nand U20775 (N_20775,N_20454,N_20204);
nor U20776 (N_20776,N_20450,N_20403);
and U20777 (N_20777,N_20148,N_20495);
or U20778 (N_20778,N_20447,N_20057);
and U20779 (N_20779,N_20291,N_20452);
nand U20780 (N_20780,N_20375,N_20297);
and U20781 (N_20781,N_20096,N_20258);
nor U20782 (N_20782,N_20306,N_20002);
nor U20783 (N_20783,N_20093,N_20203);
nor U20784 (N_20784,N_20372,N_20091);
and U20785 (N_20785,N_20380,N_20088);
and U20786 (N_20786,N_20495,N_20410);
nand U20787 (N_20787,N_20101,N_20148);
or U20788 (N_20788,N_20016,N_20235);
and U20789 (N_20789,N_20026,N_20103);
or U20790 (N_20790,N_20291,N_20432);
and U20791 (N_20791,N_20075,N_20474);
nor U20792 (N_20792,N_20039,N_20064);
and U20793 (N_20793,N_20202,N_20420);
nor U20794 (N_20794,N_20259,N_20374);
nand U20795 (N_20795,N_20160,N_20452);
or U20796 (N_20796,N_20202,N_20044);
nand U20797 (N_20797,N_20012,N_20407);
nand U20798 (N_20798,N_20366,N_20181);
nand U20799 (N_20799,N_20005,N_20029);
nor U20800 (N_20800,N_20177,N_20331);
or U20801 (N_20801,N_20434,N_20070);
nand U20802 (N_20802,N_20429,N_20216);
nand U20803 (N_20803,N_20363,N_20105);
nor U20804 (N_20804,N_20142,N_20087);
nor U20805 (N_20805,N_20489,N_20481);
nor U20806 (N_20806,N_20073,N_20007);
nand U20807 (N_20807,N_20314,N_20234);
xor U20808 (N_20808,N_20369,N_20372);
or U20809 (N_20809,N_20281,N_20376);
and U20810 (N_20810,N_20351,N_20318);
and U20811 (N_20811,N_20241,N_20107);
nor U20812 (N_20812,N_20287,N_20481);
nand U20813 (N_20813,N_20296,N_20111);
and U20814 (N_20814,N_20374,N_20229);
nand U20815 (N_20815,N_20077,N_20224);
and U20816 (N_20816,N_20090,N_20182);
xor U20817 (N_20817,N_20414,N_20468);
or U20818 (N_20818,N_20013,N_20301);
or U20819 (N_20819,N_20357,N_20308);
and U20820 (N_20820,N_20429,N_20432);
and U20821 (N_20821,N_20089,N_20238);
nor U20822 (N_20822,N_20287,N_20032);
and U20823 (N_20823,N_20437,N_20330);
nand U20824 (N_20824,N_20307,N_20383);
nand U20825 (N_20825,N_20443,N_20434);
nand U20826 (N_20826,N_20247,N_20346);
or U20827 (N_20827,N_20316,N_20072);
or U20828 (N_20828,N_20498,N_20316);
nand U20829 (N_20829,N_20126,N_20145);
nand U20830 (N_20830,N_20093,N_20333);
or U20831 (N_20831,N_20236,N_20311);
nand U20832 (N_20832,N_20050,N_20340);
nor U20833 (N_20833,N_20215,N_20332);
and U20834 (N_20834,N_20419,N_20310);
or U20835 (N_20835,N_20203,N_20175);
and U20836 (N_20836,N_20448,N_20457);
and U20837 (N_20837,N_20216,N_20456);
xnor U20838 (N_20838,N_20369,N_20461);
nor U20839 (N_20839,N_20419,N_20139);
and U20840 (N_20840,N_20332,N_20227);
and U20841 (N_20841,N_20093,N_20495);
xnor U20842 (N_20842,N_20230,N_20375);
and U20843 (N_20843,N_20284,N_20317);
and U20844 (N_20844,N_20451,N_20159);
or U20845 (N_20845,N_20483,N_20433);
nor U20846 (N_20846,N_20492,N_20489);
or U20847 (N_20847,N_20060,N_20459);
nand U20848 (N_20848,N_20214,N_20198);
and U20849 (N_20849,N_20087,N_20341);
or U20850 (N_20850,N_20200,N_20159);
or U20851 (N_20851,N_20360,N_20322);
nand U20852 (N_20852,N_20238,N_20469);
nand U20853 (N_20853,N_20444,N_20267);
nand U20854 (N_20854,N_20048,N_20329);
nor U20855 (N_20855,N_20310,N_20224);
nor U20856 (N_20856,N_20159,N_20148);
nand U20857 (N_20857,N_20472,N_20180);
nand U20858 (N_20858,N_20456,N_20168);
nor U20859 (N_20859,N_20044,N_20309);
nand U20860 (N_20860,N_20049,N_20080);
nand U20861 (N_20861,N_20277,N_20245);
or U20862 (N_20862,N_20036,N_20133);
and U20863 (N_20863,N_20428,N_20082);
and U20864 (N_20864,N_20044,N_20049);
xnor U20865 (N_20865,N_20264,N_20379);
nor U20866 (N_20866,N_20470,N_20205);
nand U20867 (N_20867,N_20243,N_20482);
and U20868 (N_20868,N_20210,N_20252);
nor U20869 (N_20869,N_20238,N_20032);
nand U20870 (N_20870,N_20311,N_20408);
nand U20871 (N_20871,N_20082,N_20178);
nand U20872 (N_20872,N_20382,N_20465);
nor U20873 (N_20873,N_20089,N_20275);
nand U20874 (N_20874,N_20400,N_20158);
nand U20875 (N_20875,N_20165,N_20340);
or U20876 (N_20876,N_20439,N_20392);
nor U20877 (N_20877,N_20022,N_20143);
and U20878 (N_20878,N_20449,N_20307);
nand U20879 (N_20879,N_20175,N_20224);
and U20880 (N_20880,N_20316,N_20136);
nand U20881 (N_20881,N_20342,N_20180);
nand U20882 (N_20882,N_20376,N_20400);
or U20883 (N_20883,N_20109,N_20330);
or U20884 (N_20884,N_20415,N_20490);
and U20885 (N_20885,N_20426,N_20084);
and U20886 (N_20886,N_20030,N_20005);
nor U20887 (N_20887,N_20456,N_20160);
nor U20888 (N_20888,N_20446,N_20312);
nor U20889 (N_20889,N_20049,N_20099);
xnor U20890 (N_20890,N_20433,N_20102);
nor U20891 (N_20891,N_20326,N_20041);
or U20892 (N_20892,N_20400,N_20246);
or U20893 (N_20893,N_20405,N_20205);
nand U20894 (N_20894,N_20296,N_20367);
xor U20895 (N_20895,N_20109,N_20318);
and U20896 (N_20896,N_20252,N_20096);
nor U20897 (N_20897,N_20237,N_20317);
or U20898 (N_20898,N_20450,N_20394);
or U20899 (N_20899,N_20455,N_20223);
and U20900 (N_20900,N_20378,N_20240);
nand U20901 (N_20901,N_20109,N_20335);
or U20902 (N_20902,N_20184,N_20202);
nand U20903 (N_20903,N_20268,N_20083);
or U20904 (N_20904,N_20433,N_20220);
and U20905 (N_20905,N_20336,N_20053);
nor U20906 (N_20906,N_20138,N_20387);
nor U20907 (N_20907,N_20213,N_20313);
nor U20908 (N_20908,N_20183,N_20302);
or U20909 (N_20909,N_20120,N_20315);
nand U20910 (N_20910,N_20152,N_20279);
nand U20911 (N_20911,N_20237,N_20127);
and U20912 (N_20912,N_20475,N_20094);
nor U20913 (N_20913,N_20358,N_20315);
or U20914 (N_20914,N_20200,N_20235);
nor U20915 (N_20915,N_20404,N_20244);
and U20916 (N_20916,N_20398,N_20236);
nand U20917 (N_20917,N_20200,N_20204);
or U20918 (N_20918,N_20184,N_20334);
xor U20919 (N_20919,N_20295,N_20216);
nor U20920 (N_20920,N_20456,N_20174);
nor U20921 (N_20921,N_20293,N_20033);
or U20922 (N_20922,N_20389,N_20011);
or U20923 (N_20923,N_20333,N_20329);
nand U20924 (N_20924,N_20131,N_20183);
nand U20925 (N_20925,N_20291,N_20127);
or U20926 (N_20926,N_20491,N_20043);
nor U20927 (N_20927,N_20293,N_20015);
or U20928 (N_20928,N_20284,N_20395);
nand U20929 (N_20929,N_20281,N_20371);
nor U20930 (N_20930,N_20494,N_20382);
and U20931 (N_20931,N_20418,N_20492);
nand U20932 (N_20932,N_20416,N_20156);
or U20933 (N_20933,N_20381,N_20218);
or U20934 (N_20934,N_20320,N_20203);
and U20935 (N_20935,N_20085,N_20328);
and U20936 (N_20936,N_20161,N_20027);
nor U20937 (N_20937,N_20308,N_20458);
nand U20938 (N_20938,N_20259,N_20129);
and U20939 (N_20939,N_20304,N_20251);
or U20940 (N_20940,N_20140,N_20084);
nor U20941 (N_20941,N_20019,N_20085);
and U20942 (N_20942,N_20259,N_20336);
nand U20943 (N_20943,N_20045,N_20006);
nand U20944 (N_20944,N_20395,N_20190);
and U20945 (N_20945,N_20176,N_20030);
nand U20946 (N_20946,N_20103,N_20384);
nand U20947 (N_20947,N_20184,N_20051);
and U20948 (N_20948,N_20200,N_20484);
nand U20949 (N_20949,N_20362,N_20083);
nor U20950 (N_20950,N_20339,N_20295);
and U20951 (N_20951,N_20328,N_20298);
nand U20952 (N_20952,N_20328,N_20343);
and U20953 (N_20953,N_20203,N_20105);
or U20954 (N_20954,N_20428,N_20383);
nor U20955 (N_20955,N_20208,N_20312);
and U20956 (N_20956,N_20217,N_20371);
nor U20957 (N_20957,N_20127,N_20236);
or U20958 (N_20958,N_20115,N_20390);
nor U20959 (N_20959,N_20067,N_20433);
or U20960 (N_20960,N_20439,N_20037);
and U20961 (N_20961,N_20390,N_20107);
nand U20962 (N_20962,N_20297,N_20487);
and U20963 (N_20963,N_20074,N_20224);
nand U20964 (N_20964,N_20132,N_20021);
nand U20965 (N_20965,N_20433,N_20182);
nand U20966 (N_20966,N_20498,N_20118);
xnor U20967 (N_20967,N_20436,N_20219);
and U20968 (N_20968,N_20020,N_20157);
nor U20969 (N_20969,N_20167,N_20445);
and U20970 (N_20970,N_20481,N_20197);
nand U20971 (N_20971,N_20105,N_20137);
nand U20972 (N_20972,N_20409,N_20411);
nand U20973 (N_20973,N_20053,N_20113);
or U20974 (N_20974,N_20384,N_20123);
nor U20975 (N_20975,N_20353,N_20062);
nor U20976 (N_20976,N_20376,N_20360);
nor U20977 (N_20977,N_20309,N_20452);
nor U20978 (N_20978,N_20376,N_20459);
or U20979 (N_20979,N_20175,N_20223);
nor U20980 (N_20980,N_20196,N_20380);
and U20981 (N_20981,N_20461,N_20335);
nand U20982 (N_20982,N_20069,N_20076);
and U20983 (N_20983,N_20351,N_20026);
nor U20984 (N_20984,N_20082,N_20397);
nor U20985 (N_20985,N_20430,N_20407);
and U20986 (N_20986,N_20337,N_20437);
nor U20987 (N_20987,N_20084,N_20298);
nand U20988 (N_20988,N_20171,N_20390);
and U20989 (N_20989,N_20062,N_20418);
nor U20990 (N_20990,N_20276,N_20444);
nor U20991 (N_20991,N_20498,N_20312);
or U20992 (N_20992,N_20151,N_20272);
or U20993 (N_20993,N_20353,N_20153);
nor U20994 (N_20994,N_20334,N_20480);
or U20995 (N_20995,N_20394,N_20451);
nor U20996 (N_20996,N_20265,N_20203);
and U20997 (N_20997,N_20020,N_20299);
xor U20998 (N_20998,N_20224,N_20260);
xor U20999 (N_20999,N_20356,N_20037);
nor U21000 (N_21000,N_20559,N_20674);
nor U21001 (N_21001,N_20858,N_20751);
nand U21002 (N_21002,N_20981,N_20719);
nand U21003 (N_21003,N_20764,N_20522);
xor U21004 (N_21004,N_20814,N_20707);
nor U21005 (N_21005,N_20826,N_20575);
or U21006 (N_21006,N_20702,N_20922);
nor U21007 (N_21007,N_20528,N_20966);
nand U21008 (N_21008,N_20834,N_20668);
nand U21009 (N_21009,N_20878,N_20832);
or U21010 (N_21010,N_20830,N_20511);
nor U21011 (N_21011,N_20969,N_20554);
and U21012 (N_21012,N_20542,N_20971);
or U21013 (N_21013,N_20503,N_20925);
or U21014 (N_21014,N_20688,N_20860);
nor U21015 (N_21015,N_20510,N_20885);
nor U21016 (N_21016,N_20841,N_20909);
and U21017 (N_21017,N_20851,N_20770);
or U21018 (N_21018,N_20582,N_20653);
or U21019 (N_21019,N_20560,N_20988);
nor U21020 (N_21020,N_20984,N_20818);
nor U21021 (N_21021,N_20785,N_20899);
nor U21022 (N_21022,N_20729,N_20968);
nor U21023 (N_21023,N_20871,N_20996);
nor U21024 (N_21024,N_20580,N_20513);
nor U21025 (N_21025,N_20547,N_20853);
nor U21026 (N_21026,N_20626,N_20953);
or U21027 (N_21027,N_20935,N_20545);
and U21028 (N_21028,N_20569,N_20534);
nand U21029 (N_21029,N_20612,N_20727);
nor U21030 (N_21030,N_20952,N_20590);
and U21031 (N_21031,N_20776,N_20566);
and U21032 (N_21032,N_20556,N_20520);
or U21033 (N_21033,N_20596,N_20740);
or U21034 (N_21034,N_20624,N_20564);
and U21035 (N_21035,N_20631,N_20884);
and U21036 (N_21036,N_20954,N_20758);
nor U21037 (N_21037,N_20661,N_20804);
nor U21038 (N_21038,N_20947,N_20888);
and U21039 (N_21039,N_20930,N_20645);
or U21040 (N_21040,N_20844,N_20985);
and U21041 (N_21041,N_20722,N_20655);
nand U21042 (N_21042,N_20592,N_20839);
nor U21043 (N_21043,N_20565,N_20797);
and U21044 (N_21044,N_20618,N_20741);
or U21045 (N_21045,N_20936,N_20784);
and U21046 (N_21046,N_20763,N_20591);
or U21047 (N_21047,N_20997,N_20767);
nor U21048 (N_21048,N_20724,N_20665);
nand U21049 (N_21049,N_20583,N_20530);
nor U21050 (N_21050,N_20573,N_20505);
nor U21051 (N_21051,N_20919,N_20973);
nand U21052 (N_21052,N_20768,N_20869);
and U21053 (N_21053,N_20750,N_20684);
and U21054 (N_21054,N_20855,N_20886);
or U21055 (N_21055,N_20863,N_20803);
xnor U21056 (N_21056,N_20726,N_20551);
nor U21057 (N_21057,N_20948,N_20549);
nor U21058 (N_21058,N_20862,N_20654);
nor U21059 (N_21059,N_20731,N_20533);
nor U21060 (N_21060,N_20808,N_20584);
or U21061 (N_21061,N_20710,N_20912);
nor U21062 (N_21062,N_20623,N_20671);
and U21063 (N_21063,N_20897,N_20762);
or U21064 (N_21064,N_20649,N_20628);
nand U21065 (N_21065,N_20561,N_20896);
nand U21066 (N_21066,N_20975,N_20923);
or U21067 (N_21067,N_20926,N_20815);
xnor U21068 (N_21068,N_20721,N_20597);
nor U21069 (N_21069,N_20827,N_20526);
nand U21070 (N_21070,N_20672,N_20664);
or U21071 (N_21071,N_20536,N_20837);
nor U21072 (N_21072,N_20794,N_20715);
or U21073 (N_21073,N_20868,N_20739);
or U21074 (N_21074,N_20963,N_20516);
nor U21075 (N_21075,N_20532,N_20924);
nor U21076 (N_21076,N_20780,N_20789);
nand U21077 (N_21077,N_20994,N_20576);
or U21078 (N_21078,N_20854,N_20589);
or U21079 (N_21079,N_20941,N_20961);
nand U21080 (N_21080,N_20658,N_20543);
nand U21081 (N_21081,N_20703,N_20541);
nor U21082 (N_21082,N_20506,N_20531);
or U21083 (N_21083,N_20792,N_20680);
nor U21084 (N_21084,N_20593,N_20595);
or U21085 (N_21085,N_20605,N_20802);
and U21086 (N_21086,N_20833,N_20695);
or U21087 (N_21087,N_20856,N_20974);
or U21088 (N_21088,N_20736,N_20709);
nor U21089 (N_21089,N_20772,N_20657);
or U21090 (N_21090,N_20670,N_20544);
and U21091 (N_21091,N_20793,N_20820);
or U21092 (N_21092,N_20898,N_20989);
and U21093 (N_21093,N_20610,N_20995);
nor U21094 (N_21094,N_20900,N_20910);
nor U21095 (N_21095,N_20619,N_20681);
or U21096 (N_21096,N_20586,N_20828);
or U21097 (N_21097,N_20527,N_20810);
nor U21098 (N_21098,N_20720,N_20978);
or U21099 (N_21099,N_20791,N_20983);
and U21100 (N_21100,N_20891,N_20553);
nand U21101 (N_21101,N_20512,N_20799);
nor U21102 (N_21102,N_20976,N_20903);
and U21103 (N_21103,N_20733,N_20602);
and U21104 (N_21104,N_20894,N_20555);
and U21105 (N_21105,N_20685,N_20691);
or U21106 (N_21106,N_20625,N_20706);
nor U21107 (N_21107,N_20970,N_20660);
nor U21108 (N_21108,N_20515,N_20747);
nand U21109 (N_21109,N_20616,N_20927);
nand U21110 (N_21110,N_20678,N_20840);
or U21111 (N_21111,N_20949,N_20859);
or U21112 (N_21112,N_20849,N_20822);
nand U21113 (N_21113,N_20718,N_20982);
nand U21114 (N_21114,N_20557,N_20913);
nor U21115 (N_21115,N_20881,N_20979);
nor U21116 (N_21116,N_20906,N_20761);
nor U21117 (N_21117,N_20725,N_20964);
nor U21118 (N_21118,N_20730,N_20669);
nand U21119 (N_21119,N_20801,N_20752);
and U21120 (N_21120,N_20999,N_20940);
nor U21121 (N_21121,N_20965,N_20640);
and U21122 (N_21122,N_20972,N_20807);
nor U21123 (N_21123,N_20676,N_20836);
or U21124 (N_21124,N_20523,N_20907);
nor U21125 (N_21125,N_20921,N_20501);
and U21126 (N_21126,N_20604,N_20864);
nand U21127 (N_21127,N_20877,N_20892);
nand U21128 (N_21128,N_20829,N_20800);
or U21129 (N_21129,N_20687,N_20756);
and U21130 (N_21130,N_20621,N_20876);
or U21131 (N_21131,N_20850,N_20939);
nand U21132 (N_21132,N_20744,N_20825);
nand U21133 (N_21133,N_20987,N_20571);
and U21134 (N_21134,N_20942,N_20577);
nand U21135 (N_21135,N_20812,N_20838);
or U21136 (N_21136,N_20639,N_20537);
and U21137 (N_21137,N_20723,N_20607);
or U21138 (N_21138,N_20562,N_20614);
nand U21139 (N_21139,N_20686,N_20872);
nor U21140 (N_21140,N_20742,N_20821);
or U21141 (N_21141,N_20689,N_20809);
or U21142 (N_21142,N_20781,N_20509);
nand U21143 (N_21143,N_20622,N_20692);
or U21144 (N_21144,N_20916,N_20890);
nor U21145 (N_21145,N_20857,N_20842);
and U21146 (N_21146,N_20754,N_20880);
nand U21147 (N_21147,N_20977,N_20637);
or U21148 (N_21148,N_20956,N_20911);
or U21149 (N_21149,N_20633,N_20835);
and U21150 (N_21150,N_20986,N_20783);
nand U21151 (N_21151,N_20737,N_20502);
and U21152 (N_21152,N_20874,N_20630);
or U21153 (N_21153,N_20852,N_20749);
or U21154 (N_21154,N_20611,N_20615);
or U21155 (N_21155,N_20824,N_20711);
nand U21156 (N_21156,N_20746,N_20651);
nand U21157 (N_21157,N_20882,N_20713);
and U21158 (N_21158,N_20782,N_20777);
nor U21159 (N_21159,N_20705,N_20732);
nand U21160 (N_21160,N_20538,N_20943);
or U21161 (N_21161,N_20643,N_20717);
nand U21162 (N_21162,N_20980,N_20638);
or U21163 (N_21163,N_20682,N_20928);
nor U21164 (N_21164,N_20819,N_20908);
or U21165 (N_21165,N_20831,N_20558);
nor U21166 (N_21166,N_20748,N_20788);
and U21167 (N_21167,N_20915,N_20652);
nor U21168 (N_21168,N_20679,N_20766);
nand U21169 (N_21169,N_20959,N_20934);
nand U21170 (N_21170,N_20714,N_20945);
or U21171 (N_21171,N_20601,N_20666);
and U21172 (N_21172,N_20889,N_20938);
and U21173 (N_21173,N_20929,N_20608);
or U21174 (N_21174,N_20675,N_20518);
nand U21175 (N_21175,N_20734,N_20519);
nand U21176 (N_21176,N_20846,N_20636);
nor U21177 (N_21177,N_20873,N_20887);
nor U21178 (N_21178,N_20957,N_20587);
and U21179 (N_21179,N_20955,N_20813);
nand U21180 (N_21180,N_20958,N_20918);
nand U21181 (N_21181,N_20933,N_20775);
or U21182 (N_21182,N_20504,N_20535);
or U21183 (N_21183,N_20632,N_20698);
or U21184 (N_21184,N_20650,N_20599);
and U21185 (N_21185,N_20508,N_20529);
xnor U21186 (N_21186,N_20606,N_20779);
nor U21187 (N_21187,N_20843,N_20517);
nor U21188 (N_21188,N_20552,N_20901);
and U21189 (N_21189,N_20690,N_20743);
nor U21190 (N_21190,N_20870,N_20875);
nor U21191 (N_21191,N_20667,N_20993);
or U21192 (N_21192,N_20712,N_20704);
or U21193 (N_21193,N_20883,N_20990);
nand U21194 (N_21194,N_20594,N_20693);
or U21195 (N_21195,N_20806,N_20603);
nand U21196 (N_21196,N_20546,N_20931);
or U21197 (N_21197,N_20778,N_20944);
or U21198 (N_21198,N_20579,N_20771);
or U21199 (N_21199,N_20796,N_20951);
nor U21200 (N_21200,N_20677,N_20600);
xor U21201 (N_21201,N_20760,N_20673);
and U21202 (N_21202,N_20572,N_20735);
nor U21203 (N_21203,N_20514,N_20634);
or U21204 (N_21204,N_20795,N_20950);
and U21205 (N_21205,N_20581,N_20757);
nor U21206 (N_21206,N_20694,N_20817);
nand U21207 (N_21207,N_20644,N_20646);
and U21208 (N_21208,N_20960,N_20847);
and U21209 (N_21209,N_20627,N_20893);
or U21210 (N_21210,N_20629,N_20563);
or U21211 (N_21211,N_20728,N_20879);
or U21212 (N_21212,N_20659,N_20662);
and U21213 (N_21213,N_20902,N_20920);
or U21214 (N_21214,N_20848,N_20642);
and U21215 (N_21215,N_20816,N_20755);
and U21216 (N_21216,N_20663,N_20656);
nand U21217 (N_21217,N_20641,N_20620);
nand U21218 (N_21218,N_20905,N_20617);
nand U21219 (N_21219,N_20811,N_20647);
nor U21220 (N_21220,N_20570,N_20895);
nor U21221 (N_21221,N_20635,N_20550);
nor U21222 (N_21222,N_20500,N_20540);
xor U21223 (N_21223,N_20708,N_20525);
nor U21224 (N_21224,N_20774,N_20914);
or U21225 (N_21225,N_20798,N_20598);
nand U21226 (N_21226,N_20745,N_20701);
or U21227 (N_21227,N_20548,N_20753);
or U21228 (N_21228,N_20524,N_20917);
nand U21229 (N_21229,N_20787,N_20805);
nand U21230 (N_21230,N_20790,N_20769);
nor U21231 (N_21231,N_20609,N_20585);
and U21232 (N_21232,N_20578,N_20866);
and U21233 (N_21233,N_20946,N_20507);
and U21234 (N_21234,N_20937,N_20697);
nor U21235 (N_21235,N_20683,N_20967);
or U21236 (N_21236,N_20716,N_20567);
nand U21237 (N_21237,N_20932,N_20998);
nor U21238 (N_21238,N_20738,N_20773);
or U21239 (N_21239,N_20904,N_20867);
nor U21240 (N_21240,N_20865,N_20700);
nor U21241 (N_21241,N_20648,N_20574);
nand U21242 (N_21242,N_20696,N_20588);
nand U21243 (N_21243,N_20568,N_20613);
and U21244 (N_21244,N_20992,N_20861);
and U21245 (N_21245,N_20521,N_20786);
nor U21246 (N_21246,N_20823,N_20962);
or U21247 (N_21247,N_20991,N_20699);
or U21248 (N_21248,N_20539,N_20845);
nand U21249 (N_21249,N_20765,N_20759);
nor U21250 (N_21250,N_20808,N_20994);
or U21251 (N_21251,N_20976,N_20775);
nand U21252 (N_21252,N_20948,N_20757);
and U21253 (N_21253,N_20611,N_20729);
nor U21254 (N_21254,N_20748,N_20770);
or U21255 (N_21255,N_20558,N_20854);
nor U21256 (N_21256,N_20522,N_20915);
nand U21257 (N_21257,N_20867,N_20505);
or U21258 (N_21258,N_20775,N_20688);
and U21259 (N_21259,N_20516,N_20772);
and U21260 (N_21260,N_20889,N_20980);
or U21261 (N_21261,N_20781,N_20568);
or U21262 (N_21262,N_20834,N_20675);
or U21263 (N_21263,N_20619,N_20709);
xnor U21264 (N_21264,N_20624,N_20511);
or U21265 (N_21265,N_20678,N_20664);
nor U21266 (N_21266,N_20844,N_20704);
or U21267 (N_21267,N_20988,N_20992);
xnor U21268 (N_21268,N_20867,N_20720);
nor U21269 (N_21269,N_20632,N_20779);
or U21270 (N_21270,N_20748,N_20713);
or U21271 (N_21271,N_20588,N_20642);
xnor U21272 (N_21272,N_20613,N_20549);
and U21273 (N_21273,N_20902,N_20983);
or U21274 (N_21274,N_20514,N_20617);
nand U21275 (N_21275,N_20975,N_20831);
nor U21276 (N_21276,N_20694,N_20871);
nor U21277 (N_21277,N_20805,N_20760);
nand U21278 (N_21278,N_20598,N_20604);
nor U21279 (N_21279,N_20953,N_20644);
and U21280 (N_21280,N_20661,N_20907);
and U21281 (N_21281,N_20952,N_20616);
nor U21282 (N_21282,N_20659,N_20875);
or U21283 (N_21283,N_20863,N_20609);
or U21284 (N_21284,N_20802,N_20932);
and U21285 (N_21285,N_20538,N_20551);
nor U21286 (N_21286,N_20655,N_20663);
and U21287 (N_21287,N_20699,N_20756);
or U21288 (N_21288,N_20510,N_20622);
and U21289 (N_21289,N_20721,N_20662);
and U21290 (N_21290,N_20889,N_20577);
and U21291 (N_21291,N_20798,N_20967);
nand U21292 (N_21292,N_20914,N_20761);
or U21293 (N_21293,N_20599,N_20817);
nand U21294 (N_21294,N_20507,N_20752);
and U21295 (N_21295,N_20716,N_20864);
nand U21296 (N_21296,N_20739,N_20559);
nor U21297 (N_21297,N_20862,N_20885);
or U21298 (N_21298,N_20600,N_20810);
nor U21299 (N_21299,N_20698,N_20592);
or U21300 (N_21300,N_20984,N_20730);
nand U21301 (N_21301,N_20600,N_20789);
or U21302 (N_21302,N_20704,N_20657);
and U21303 (N_21303,N_20666,N_20551);
or U21304 (N_21304,N_20975,N_20511);
nor U21305 (N_21305,N_20716,N_20578);
and U21306 (N_21306,N_20764,N_20838);
nor U21307 (N_21307,N_20557,N_20587);
nand U21308 (N_21308,N_20607,N_20850);
nor U21309 (N_21309,N_20782,N_20681);
or U21310 (N_21310,N_20869,N_20821);
nand U21311 (N_21311,N_20554,N_20974);
or U21312 (N_21312,N_20868,N_20844);
nor U21313 (N_21313,N_20712,N_20977);
or U21314 (N_21314,N_20666,N_20685);
nor U21315 (N_21315,N_20903,N_20737);
nor U21316 (N_21316,N_20586,N_20899);
nand U21317 (N_21317,N_20987,N_20739);
nand U21318 (N_21318,N_20985,N_20720);
and U21319 (N_21319,N_20751,N_20929);
or U21320 (N_21320,N_20751,N_20568);
nand U21321 (N_21321,N_20843,N_20514);
or U21322 (N_21322,N_20955,N_20573);
or U21323 (N_21323,N_20729,N_20783);
and U21324 (N_21324,N_20501,N_20611);
or U21325 (N_21325,N_20539,N_20817);
and U21326 (N_21326,N_20666,N_20815);
and U21327 (N_21327,N_20642,N_20553);
nand U21328 (N_21328,N_20650,N_20852);
nand U21329 (N_21329,N_20657,N_20691);
or U21330 (N_21330,N_20643,N_20725);
nand U21331 (N_21331,N_20605,N_20959);
nor U21332 (N_21332,N_20587,N_20801);
nor U21333 (N_21333,N_20761,N_20850);
and U21334 (N_21334,N_20829,N_20949);
nand U21335 (N_21335,N_20785,N_20679);
or U21336 (N_21336,N_20790,N_20626);
nor U21337 (N_21337,N_20668,N_20745);
or U21338 (N_21338,N_20823,N_20767);
or U21339 (N_21339,N_20747,N_20838);
nand U21340 (N_21340,N_20762,N_20638);
nand U21341 (N_21341,N_20892,N_20644);
nand U21342 (N_21342,N_20518,N_20999);
nand U21343 (N_21343,N_20549,N_20715);
nor U21344 (N_21344,N_20801,N_20924);
nor U21345 (N_21345,N_20539,N_20629);
or U21346 (N_21346,N_20891,N_20693);
nand U21347 (N_21347,N_20931,N_20977);
or U21348 (N_21348,N_20602,N_20887);
and U21349 (N_21349,N_20816,N_20940);
nand U21350 (N_21350,N_20515,N_20988);
and U21351 (N_21351,N_20528,N_20921);
and U21352 (N_21352,N_20992,N_20941);
and U21353 (N_21353,N_20638,N_20529);
nor U21354 (N_21354,N_20558,N_20923);
and U21355 (N_21355,N_20954,N_20669);
and U21356 (N_21356,N_20956,N_20666);
nor U21357 (N_21357,N_20808,N_20587);
nand U21358 (N_21358,N_20781,N_20956);
nand U21359 (N_21359,N_20678,N_20583);
and U21360 (N_21360,N_20977,N_20867);
nand U21361 (N_21361,N_20540,N_20600);
or U21362 (N_21362,N_20978,N_20818);
and U21363 (N_21363,N_20928,N_20526);
and U21364 (N_21364,N_20733,N_20680);
nor U21365 (N_21365,N_20533,N_20621);
nor U21366 (N_21366,N_20693,N_20696);
nor U21367 (N_21367,N_20786,N_20619);
xnor U21368 (N_21368,N_20861,N_20600);
nor U21369 (N_21369,N_20722,N_20837);
xor U21370 (N_21370,N_20941,N_20910);
or U21371 (N_21371,N_20649,N_20735);
and U21372 (N_21372,N_20533,N_20959);
or U21373 (N_21373,N_20752,N_20963);
or U21374 (N_21374,N_20594,N_20678);
nor U21375 (N_21375,N_20562,N_20704);
nand U21376 (N_21376,N_20872,N_20989);
nand U21377 (N_21377,N_20936,N_20858);
nor U21378 (N_21378,N_20573,N_20555);
nor U21379 (N_21379,N_20590,N_20606);
and U21380 (N_21380,N_20808,N_20909);
and U21381 (N_21381,N_20589,N_20910);
nand U21382 (N_21382,N_20604,N_20556);
and U21383 (N_21383,N_20549,N_20995);
nand U21384 (N_21384,N_20701,N_20828);
nor U21385 (N_21385,N_20991,N_20541);
nor U21386 (N_21386,N_20893,N_20500);
and U21387 (N_21387,N_20633,N_20719);
and U21388 (N_21388,N_20797,N_20820);
or U21389 (N_21389,N_20868,N_20578);
nand U21390 (N_21390,N_20828,N_20559);
and U21391 (N_21391,N_20739,N_20794);
or U21392 (N_21392,N_20822,N_20907);
nand U21393 (N_21393,N_20579,N_20846);
nor U21394 (N_21394,N_20566,N_20835);
nand U21395 (N_21395,N_20896,N_20675);
and U21396 (N_21396,N_20851,N_20969);
nand U21397 (N_21397,N_20794,N_20796);
nor U21398 (N_21398,N_20948,N_20602);
and U21399 (N_21399,N_20679,N_20758);
nor U21400 (N_21400,N_20743,N_20526);
nor U21401 (N_21401,N_20715,N_20605);
or U21402 (N_21402,N_20553,N_20997);
nor U21403 (N_21403,N_20658,N_20747);
nor U21404 (N_21404,N_20710,N_20645);
nor U21405 (N_21405,N_20803,N_20858);
nand U21406 (N_21406,N_20551,N_20992);
and U21407 (N_21407,N_20588,N_20846);
and U21408 (N_21408,N_20565,N_20899);
nand U21409 (N_21409,N_20701,N_20906);
nand U21410 (N_21410,N_20951,N_20664);
nand U21411 (N_21411,N_20912,N_20534);
or U21412 (N_21412,N_20813,N_20632);
or U21413 (N_21413,N_20939,N_20825);
or U21414 (N_21414,N_20625,N_20983);
and U21415 (N_21415,N_20948,N_20779);
or U21416 (N_21416,N_20847,N_20922);
nand U21417 (N_21417,N_20532,N_20503);
nor U21418 (N_21418,N_20802,N_20844);
nor U21419 (N_21419,N_20559,N_20868);
and U21420 (N_21420,N_20877,N_20567);
and U21421 (N_21421,N_20614,N_20856);
nand U21422 (N_21422,N_20760,N_20533);
nand U21423 (N_21423,N_20682,N_20918);
nand U21424 (N_21424,N_20674,N_20920);
or U21425 (N_21425,N_20704,N_20963);
nor U21426 (N_21426,N_20568,N_20690);
nand U21427 (N_21427,N_20890,N_20846);
and U21428 (N_21428,N_20825,N_20595);
and U21429 (N_21429,N_20962,N_20937);
nand U21430 (N_21430,N_20569,N_20718);
nand U21431 (N_21431,N_20529,N_20651);
nor U21432 (N_21432,N_20844,N_20785);
and U21433 (N_21433,N_20713,N_20969);
and U21434 (N_21434,N_20659,N_20958);
nor U21435 (N_21435,N_20809,N_20536);
or U21436 (N_21436,N_20514,N_20869);
or U21437 (N_21437,N_20632,N_20770);
nand U21438 (N_21438,N_20829,N_20520);
xor U21439 (N_21439,N_20510,N_20822);
and U21440 (N_21440,N_20593,N_20729);
or U21441 (N_21441,N_20707,N_20769);
nor U21442 (N_21442,N_20718,N_20742);
or U21443 (N_21443,N_20910,N_20975);
and U21444 (N_21444,N_20550,N_20792);
or U21445 (N_21445,N_20755,N_20600);
or U21446 (N_21446,N_20589,N_20714);
nor U21447 (N_21447,N_20846,N_20896);
nand U21448 (N_21448,N_20652,N_20795);
or U21449 (N_21449,N_20547,N_20624);
nor U21450 (N_21450,N_20970,N_20616);
or U21451 (N_21451,N_20859,N_20734);
nand U21452 (N_21452,N_20892,N_20936);
nor U21453 (N_21453,N_20895,N_20748);
nand U21454 (N_21454,N_20818,N_20845);
or U21455 (N_21455,N_20609,N_20922);
nand U21456 (N_21456,N_20546,N_20912);
nor U21457 (N_21457,N_20843,N_20831);
and U21458 (N_21458,N_20551,N_20667);
and U21459 (N_21459,N_20532,N_20809);
nor U21460 (N_21460,N_20780,N_20792);
nor U21461 (N_21461,N_20751,N_20702);
nor U21462 (N_21462,N_20844,N_20874);
and U21463 (N_21463,N_20964,N_20506);
nand U21464 (N_21464,N_20632,N_20563);
nand U21465 (N_21465,N_20564,N_20732);
nand U21466 (N_21466,N_20637,N_20876);
or U21467 (N_21467,N_20872,N_20599);
nor U21468 (N_21468,N_20660,N_20912);
nand U21469 (N_21469,N_20656,N_20514);
nor U21470 (N_21470,N_20984,N_20856);
nor U21471 (N_21471,N_20773,N_20552);
nand U21472 (N_21472,N_20982,N_20839);
or U21473 (N_21473,N_20922,N_20570);
or U21474 (N_21474,N_20517,N_20714);
or U21475 (N_21475,N_20670,N_20705);
nand U21476 (N_21476,N_20614,N_20734);
nand U21477 (N_21477,N_20510,N_20575);
nor U21478 (N_21478,N_20937,N_20825);
nor U21479 (N_21479,N_20786,N_20528);
and U21480 (N_21480,N_20777,N_20911);
nor U21481 (N_21481,N_20602,N_20675);
or U21482 (N_21482,N_20794,N_20543);
or U21483 (N_21483,N_20767,N_20911);
and U21484 (N_21484,N_20763,N_20547);
nor U21485 (N_21485,N_20714,N_20770);
or U21486 (N_21486,N_20686,N_20821);
nor U21487 (N_21487,N_20867,N_20988);
and U21488 (N_21488,N_20686,N_20556);
or U21489 (N_21489,N_20827,N_20835);
or U21490 (N_21490,N_20512,N_20682);
and U21491 (N_21491,N_20654,N_20687);
and U21492 (N_21492,N_20636,N_20768);
nor U21493 (N_21493,N_20959,N_20713);
nor U21494 (N_21494,N_20956,N_20943);
nand U21495 (N_21495,N_20638,N_20891);
or U21496 (N_21496,N_20850,N_20721);
and U21497 (N_21497,N_20575,N_20956);
or U21498 (N_21498,N_20571,N_20644);
and U21499 (N_21499,N_20521,N_20728);
nand U21500 (N_21500,N_21053,N_21308);
or U21501 (N_21501,N_21375,N_21144);
or U21502 (N_21502,N_21159,N_21017);
or U21503 (N_21503,N_21267,N_21326);
and U21504 (N_21504,N_21285,N_21446);
or U21505 (N_21505,N_21336,N_21466);
or U21506 (N_21506,N_21158,N_21024);
or U21507 (N_21507,N_21381,N_21010);
xor U21508 (N_21508,N_21278,N_21018);
or U21509 (N_21509,N_21151,N_21030);
nand U21510 (N_21510,N_21400,N_21356);
and U21511 (N_21511,N_21404,N_21421);
or U21512 (N_21512,N_21412,N_21210);
or U21513 (N_21513,N_21273,N_21399);
nand U21514 (N_21514,N_21367,N_21318);
or U21515 (N_21515,N_21048,N_21050);
or U21516 (N_21516,N_21208,N_21320);
nor U21517 (N_21517,N_21234,N_21150);
or U21518 (N_21518,N_21259,N_21219);
nor U21519 (N_21519,N_21079,N_21137);
nand U21520 (N_21520,N_21260,N_21222);
nand U21521 (N_21521,N_21416,N_21306);
nand U21522 (N_21522,N_21346,N_21454);
xor U21523 (N_21523,N_21484,N_21450);
and U21524 (N_21524,N_21348,N_21223);
nand U21525 (N_21525,N_21052,N_21474);
nor U21526 (N_21526,N_21389,N_21483);
and U21527 (N_21527,N_21046,N_21352);
nand U21528 (N_21528,N_21269,N_21096);
and U21529 (N_21529,N_21300,N_21006);
nor U21530 (N_21530,N_21491,N_21214);
and U21531 (N_21531,N_21106,N_21410);
and U21532 (N_21532,N_21499,N_21043);
nand U21533 (N_21533,N_21255,N_21388);
nor U21534 (N_21534,N_21332,N_21155);
nor U21535 (N_21535,N_21287,N_21473);
nor U21536 (N_21536,N_21461,N_21391);
nor U21537 (N_21537,N_21495,N_21245);
nand U21538 (N_21538,N_21482,N_21098);
nor U21539 (N_21539,N_21164,N_21165);
nand U21540 (N_21540,N_21459,N_21059);
or U21541 (N_21541,N_21441,N_21369);
or U21542 (N_21542,N_21216,N_21496);
nand U21543 (N_21543,N_21221,N_21487);
and U21544 (N_21544,N_21131,N_21290);
nor U21545 (N_21545,N_21448,N_21243);
nand U21546 (N_21546,N_21019,N_21100);
nor U21547 (N_21547,N_21233,N_21022);
and U21548 (N_21548,N_21429,N_21153);
nor U21549 (N_21549,N_21277,N_21238);
or U21550 (N_21550,N_21257,N_21161);
and U21551 (N_21551,N_21136,N_21103);
and U21552 (N_21552,N_21075,N_21084);
nand U21553 (N_21553,N_21228,N_21090);
and U21554 (N_21554,N_21133,N_21088);
and U21555 (N_21555,N_21203,N_21235);
nor U21556 (N_21556,N_21177,N_21305);
or U21557 (N_21557,N_21067,N_21316);
or U21558 (N_21558,N_21392,N_21357);
nor U21559 (N_21559,N_21254,N_21353);
and U21560 (N_21560,N_21156,N_21069);
nand U21561 (N_21561,N_21071,N_21247);
or U21562 (N_21562,N_21384,N_21363);
nor U21563 (N_21563,N_21468,N_21142);
nand U21564 (N_21564,N_21185,N_21061);
and U21565 (N_21565,N_21476,N_21057);
nor U21566 (N_21566,N_21068,N_21188);
nor U21567 (N_21567,N_21029,N_21172);
nor U21568 (N_21568,N_21494,N_21250);
or U21569 (N_21569,N_21341,N_21130);
nor U21570 (N_21570,N_21288,N_21364);
nand U21571 (N_21571,N_21355,N_21311);
nor U21572 (N_21572,N_21490,N_21271);
nand U21573 (N_21573,N_21089,N_21295);
or U21574 (N_21574,N_21224,N_21117);
nor U21575 (N_21575,N_21184,N_21319);
nand U21576 (N_21576,N_21220,N_21420);
and U21577 (N_21577,N_21498,N_21325);
and U21578 (N_21578,N_21212,N_21040);
or U21579 (N_21579,N_21304,N_21148);
and U21580 (N_21580,N_21093,N_21102);
nor U21581 (N_21581,N_21372,N_21382);
or U21582 (N_21582,N_21105,N_21205);
nor U21583 (N_21583,N_21376,N_21378);
nor U21584 (N_21584,N_21012,N_21026);
nor U21585 (N_21585,N_21027,N_21160);
and U21586 (N_21586,N_21112,N_21241);
nand U21587 (N_21587,N_21343,N_21206);
or U21588 (N_21588,N_21386,N_21209);
and U21589 (N_21589,N_21011,N_21274);
or U21590 (N_21590,N_21231,N_21424);
nand U21591 (N_21591,N_21455,N_21094);
and U21592 (N_21592,N_21213,N_21331);
nand U21593 (N_21593,N_21179,N_21403);
and U21594 (N_21594,N_21362,N_21138);
nor U21595 (N_21595,N_21104,N_21072);
and U21596 (N_21596,N_21189,N_21051);
and U21597 (N_21597,N_21302,N_21080);
nor U21598 (N_21598,N_21321,N_21036);
nor U21599 (N_21599,N_21237,N_21380);
or U21600 (N_21600,N_21175,N_21147);
or U21601 (N_21601,N_21492,N_21275);
nor U21602 (N_21602,N_21281,N_21183);
or U21603 (N_21603,N_21297,N_21323);
or U21604 (N_21604,N_21240,N_21489);
nor U21605 (N_21605,N_21014,N_21481);
or U21606 (N_21606,N_21426,N_21262);
and U21607 (N_21607,N_21317,N_21201);
and U21608 (N_21608,N_21204,N_21472);
and U21609 (N_21609,N_21167,N_21191);
and U21610 (N_21610,N_21056,N_21070);
nor U21611 (N_21611,N_21101,N_21122);
and U21612 (N_21612,N_21258,N_21360);
or U21613 (N_21613,N_21091,N_21330);
and U21614 (N_21614,N_21108,N_21119);
or U21615 (N_21615,N_21293,N_21463);
or U21616 (N_21616,N_21327,N_21125);
and U21617 (N_21617,N_21286,N_21244);
nand U21618 (N_21618,N_21438,N_21015);
nand U21619 (N_21619,N_21082,N_21374);
and U21620 (N_21620,N_21251,N_21135);
xnor U21621 (N_21621,N_21408,N_21342);
nand U21622 (N_21622,N_21197,N_21301);
nand U21623 (N_21623,N_21310,N_21462);
nor U21624 (N_21624,N_21419,N_21092);
or U21625 (N_21625,N_21003,N_21460);
and U21626 (N_21626,N_21436,N_21428);
nand U21627 (N_21627,N_21291,N_21370);
nand U21628 (N_21628,N_21263,N_21371);
xor U21629 (N_21629,N_21444,N_21440);
and U21630 (N_21630,N_21478,N_21004);
or U21631 (N_21631,N_21042,N_21178);
nand U21632 (N_21632,N_21037,N_21270);
nand U21633 (N_21633,N_21198,N_21480);
and U21634 (N_21634,N_21493,N_21039);
nand U21635 (N_21635,N_21182,N_21411);
or U21636 (N_21636,N_21314,N_21236);
nor U21637 (N_21637,N_21486,N_21456);
nor U21638 (N_21638,N_21393,N_21439);
nor U21639 (N_21639,N_21129,N_21064);
nor U21640 (N_21640,N_21239,N_21433);
or U21641 (N_21641,N_21186,N_21169);
nor U21642 (N_21642,N_21414,N_21058);
or U21643 (N_21643,N_21467,N_21309);
and U21644 (N_21644,N_21207,N_21081);
nand U21645 (N_21645,N_21427,N_21335);
nand U21646 (N_21646,N_21180,N_21292);
and U21647 (N_21647,N_21111,N_21246);
nor U21648 (N_21648,N_21447,N_21171);
nand U21649 (N_21649,N_21121,N_21099);
and U21650 (N_21650,N_21422,N_21127);
and U21651 (N_21651,N_21345,N_21126);
and U21652 (N_21652,N_21115,N_21280);
or U21653 (N_21653,N_21264,N_21032);
or U21654 (N_21654,N_21021,N_21465);
nand U21655 (N_21655,N_21361,N_21008);
nor U21656 (N_21656,N_21417,N_21168);
nand U21657 (N_21657,N_21097,N_21249);
nand U21658 (N_21658,N_21116,N_21405);
and U21659 (N_21659,N_21402,N_21347);
and U21660 (N_21660,N_21095,N_21062);
nand U21661 (N_21661,N_21035,N_21470);
or U21662 (N_21662,N_21110,N_21409);
and U21663 (N_21663,N_21279,N_21329);
nand U21664 (N_21664,N_21313,N_21083);
nand U21665 (N_21665,N_21383,N_21124);
and U21666 (N_21666,N_21190,N_21398);
and U21667 (N_21667,N_21413,N_21333);
and U21668 (N_21668,N_21194,N_21049);
or U21669 (N_21669,N_21229,N_21452);
and U21670 (N_21670,N_21349,N_21034);
nor U21671 (N_21671,N_21266,N_21132);
nor U21672 (N_21672,N_21390,N_21396);
nand U21673 (N_21673,N_21366,N_21041);
or U21674 (N_21674,N_21020,N_21085);
or U21675 (N_21675,N_21000,N_21324);
or U21676 (N_21676,N_21340,N_21397);
and U21677 (N_21677,N_21256,N_21451);
and U21678 (N_21678,N_21373,N_21047);
or U21679 (N_21679,N_21261,N_21434);
nor U21680 (N_21680,N_21120,N_21031);
and U21681 (N_21681,N_21469,N_21140);
xnor U21682 (N_21682,N_21227,N_21449);
nor U21683 (N_21683,N_21038,N_21066);
nor U21684 (N_21684,N_21076,N_21453);
nor U21685 (N_21685,N_21351,N_21443);
and U21686 (N_21686,N_21272,N_21218);
nand U21687 (N_21687,N_21139,N_21149);
and U21688 (N_21688,N_21143,N_21163);
and U21689 (N_21689,N_21001,N_21128);
and U21690 (N_21690,N_21344,N_21187);
nand U21691 (N_21691,N_21337,N_21114);
nand U21692 (N_21692,N_21252,N_21118);
nor U21693 (N_21693,N_21359,N_21195);
and U21694 (N_21694,N_21028,N_21181);
and U21695 (N_21695,N_21086,N_21044);
or U21696 (N_21696,N_21387,N_21173);
and U21697 (N_21697,N_21283,N_21339);
and U21698 (N_21698,N_21312,N_21377);
nor U21699 (N_21699,N_21401,N_21230);
nand U21700 (N_21700,N_21192,N_21328);
nor U21701 (N_21701,N_21268,N_21196);
nor U21702 (N_21702,N_21475,N_21146);
and U21703 (N_21703,N_21002,N_21025);
nor U21704 (N_21704,N_21154,N_21074);
nor U21705 (N_21705,N_21479,N_21298);
or U21706 (N_21706,N_21009,N_21350);
or U21707 (N_21707,N_21430,N_21394);
nor U21708 (N_21708,N_21437,N_21007);
or U21709 (N_21709,N_21358,N_21442);
nor U21710 (N_21710,N_21226,N_21162);
nor U21711 (N_21711,N_21145,N_21307);
nand U21712 (N_21712,N_21152,N_21334);
nor U21713 (N_21713,N_21193,N_21141);
and U21714 (N_21714,N_21407,N_21087);
nand U21715 (N_21715,N_21107,N_21065);
nor U21716 (N_21716,N_21303,N_21109);
and U21717 (N_21717,N_21113,N_21418);
nand U21718 (N_21718,N_21016,N_21134);
and U21719 (N_21719,N_21299,N_21338);
and U21720 (N_21720,N_21485,N_21284);
and U21721 (N_21721,N_21242,N_21354);
or U21722 (N_21722,N_21265,N_21217);
xor U21723 (N_21723,N_21365,N_21415);
and U21724 (N_21724,N_21276,N_21176);
and U21725 (N_21725,N_21385,N_21174);
or U21726 (N_21726,N_21202,N_21060);
nor U21727 (N_21727,N_21395,N_21406);
nand U21728 (N_21728,N_21023,N_21315);
and U21729 (N_21729,N_21211,N_21055);
and U21730 (N_21730,N_21368,N_21379);
nand U21731 (N_21731,N_21458,N_21078);
or U21732 (N_21732,N_21445,N_21289);
or U21733 (N_21733,N_21253,N_21296);
nor U21734 (N_21734,N_21215,N_21033);
and U21735 (N_21735,N_21431,N_21157);
or U21736 (N_21736,N_21435,N_21005);
nand U21737 (N_21737,N_21477,N_21045);
and U21738 (N_21738,N_21488,N_21232);
or U21739 (N_21739,N_21248,N_21225);
nand U21740 (N_21740,N_21013,N_21282);
or U21741 (N_21741,N_21054,N_21423);
nor U21742 (N_21742,N_21073,N_21200);
or U21743 (N_21743,N_21077,N_21294);
and U21744 (N_21744,N_21471,N_21322);
nor U21745 (N_21745,N_21063,N_21425);
or U21746 (N_21746,N_21123,N_21457);
nor U21747 (N_21747,N_21199,N_21166);
nor U21748 (N_21748,N_21464,N_21432);
nand U21749 (N_21749,N_21497,N_21170);
and U21750 (N_21750,N_21369,N_21276);
nor U21751 (N_21751,N_21194,N_21369);
and U21752 (N_21752,N_21062,N_21068);
and U21753 (N_21753,N_21058,N_21199);
and U21754 (N_21754,N_21166,N_21198);
nand U21755 (N_21755,N_21100,N_21326);
nand U21756 (N_21756,N_21064,N_21297);
nand U21757 (N_21757,N_21104,N_21383);
and U21758 (N_21758,N_21340,N_21407);
and U21759 (N_21759,N_21227,N_21076);
nand U21760 (N_21760,N_21499,N_21209);
nand U21761 (N_21761,N_21331,N_21122);
nand U21762 (N_21762,N_21413,N_21444);
or U21763 (N_21763,N_21445,N_21416);
nand U21764 (N_21764,N_21358,N_21107);
nor U21765 (N_21765,N_21411,N_21416);
nor U21766 (N_21766,N_21356,N_21247);
nor U21767 (N_21767,N_21041,N_21082);
and U21768 (N_21768,N_21001,N_21422);
or U21769 (N_21769,N_21466,N_21398);
and U21770 (N_21770,N_21297,N_21054);
nand U21771 (N_21771,N_21221,N_21199);
nor U21772 (N_21772,N_21210,N_21428);
nand U21773 (N_21773,N_21435,N_21107);
and U21774 (N_21774,N_21145,N_21313);
and U21775 (N_21775,N_21486,N_21245);
and U21776 (N_21776,N_21358,N_21204);
nor U21777 (N_21777,N_21297,N_21087);
nand U21778 (N_21778,N_21436,N_21339);
and U21779 (N_21779,N_21492,N_21263);
nor U21780 (N_21780,N_21249,N_21071);
or U21781 (N_21781,N_21220,N_21369);
and U21782 (N_21782,N_21375,N_21148);
nor U21783 (N_21783,N_21162,N_21293);
nor U21784 (N_21784,N_21365,N_21015);
or U21785 (N_21785,N_21220,N_21007);
and U21786 (N_21786,N_21362,N_21183);
nor U21787 (N_21787,N_21248,N_21392);
or U21788 (N_21788,N_21303,N_21007);
and U21789 (N_21789,N_21334,N_21202);
and U21790 (N_21790,N_21286,N_21424);
or U21791 (N_21791,N_21452,N_21202);
xor U21792 (N_21792,N_21282,N_21488);
or U21793 (N_21793,N_21128,N_21079);
and U21794 (N_21794,N_21089,N_21458);
or U21795 (N_21795,N_21216,N_21271);
nor U21796 (N_21796,N_21348,N_21295);
or U21797 (N_21797,N_21070,N_21071);
xor U21798 (N_21798,N_21000,N_21040);
or U21799 (N_21799,N_21458,N_21421);
nand U21800 (N_21800,N_21265,N_21223);
nor U21801 (N_21801,N_21105,N_21390);
nor U21802 (N_21802,N_21214,N_21100);
nor U21803 (N_21803,N_21095,N_21423);
and U21804 (N_21804,N_21223,N_21022);
and U21805 (N_21805,N_21246,N_21297);
and U21806 (N_21806,N_21162,N_21248);
or U21807 (N_21807,N_21259,N_21474);
nor U21808 (N_21808,N_21489,N_21155);
and U21809 (N_21809,N_21499,N_21463);
nand U21810 (N_21810,N_21027,N_21221);
and U21811 (N_21811,N_21474,N_21421);
nor U21812 (N_21812,N_21343,N_21173);
nand U21813 (N_21813,N_21431,N_21042);
and U21814 (N_21814,N_21366,N_21484);
nor U21815 (N_21815,N_21400,N_21443);
or U21816 (N_21816,N_21349,N_21078);
nor U21817 (N_21817,N_21281,N_21016);
xor U21818 (N_21818,N_21055,N_21344);
nor U21819 (N_21819,N_21023,N_21382);
nor U21820 (N_21820,N_21107,N_21321);
nor U21821 (N_21821,N_21274,N_21495);
and U21822 (N_21822,N_21078,N_21439);
and U21823 (N_21823,N_21122,N_21015);
nand U21824 (N_21824,N_21447,N_21358);
and U21825 (N_21825,N_21073,N_21160);
and U21826 (N_21826,N_21416,N_21298);
or U21827 (N_21827,N_21484,N_21491);
and U21828 (N_21828,N_21332,N_21132);
nor U21829 (N_21829,N_21131,N_21370);
and U21830 (N_21830,N_21016,N_21275);
nor U21831 (N_21831,N_21402,N_21038);
and U21832 (N_21832,N_21004,N_21426);
xnor U21833 (N_21833,N_21207,N_21430);
and U21834 (N_21834,N_21231,N_21345);
nand U21835 (N_21835,N_21125,N_21183);
nand U21836 (N_21836,N_21452,N_21251);
or U21837 (N_21837,N_21312,N_21121);
or U21838 (N_21838,N_21478,N_21002);
nor U21839 (N_21839,N_21448,N_21486);
and U21840 (N_21840,N_21473,N_21378);
nor U21841 (N_21841,N_21396,N_21341);
xor U21842 (N_21842,N_21334,N_21188);
or U21843 (N_21843,N_21309,N_21448);
xor U21844 (N_21844,N_21038,N_21045);
and U21845 (N_21845,N_21256,N_21219);
and U21846 (N_21846,N_21020,N_21290);
and U21847 (N_21847,N_21162,N_21125);
or U21848 (N_21848,N_21111,N_21467);
xnor U21849 (N_21849,N_21380,N_21130);
and U21850 (N_21850,N_21453,N_21386);
nor U21851 (N_21851,N_21473,N_21409);
xnor U21852 (N_21852,N_21404,N_21040);
and U21853 (N_21853,N_21402,N_21475);
nand U21854 (N_21854,N_21367,N_21011);
xnor U21855 (N_21855,N_21100,N_21335);
or U21856 (N_21856,N_21355,N_21431);
nor U21857 (N_21857,N_21264,N_21098);
nand U21858 (N_21858,N_21439,N_21472);
nand U21859 (N_21859,N_21298,N_21146);
nor U21860 (N_21860,N_21334,N_21058);
nand U21861 (N_21861,N_21155,N_21234);
nand U21862 (N_21862,N_21202,N_21059);
nand U21863 (N_21863,N_21305,N_21394);
and U21864 (N_21864,N_21092,N_21019);
nor U21865 (N_21865,N_21423,N_21118);
and U21866 (N_21866,N_21165,N_21469);
or U21867 (N_21867,N_21091,N_21108);
and U21868 (N_21868,N_21288,N_21135);
or U21869 (N_21869,N_21423,N_21034);
xor U21870 (N_21870,N_21058,N_21123);
nand U21871 (N_21871,N_21486,N_21006);
nand U21872 (N_21872,N_21170,N_21261);
nand U21873 (N_21873,N_21474,N_21214);
nor U21874 (N_21874,N_21271,N_21064);
and U21875 (N_21875,N_21117,N_21333);
nand U21876 (N_21876,N_21050,N_21053);
or U21877 (N_21877,N_21000,N_21025);
or U21878 (N_21878,N_21335,N_21108);
nor U21879 (N_21879,N_21323,N_21383);
nand U21880 (N_21880,N_21073,N_21168);
and U21881 (N_21881,N_21209,N_21494);
nor U21882 (N_21882,N_21011,N_21160);
and U21883 (N_21883,N_21046,N_21324);
nand U21884 (N_21884,N_21151,N_21354);
or U21885 (N_21885,N_21093,N_21449);
xor U21886 (N_21886,N_21411,N_21107);
nand U21887 (N_21887,N_21271,N_21476);
and U21888 (N_21888,N_21058,N_21408);
xor U21889 (N_21889,N_21483,N_21356);
nor U21890 (N_21890,N_21171,N_21260);
nor U21891 (N_21891,N_21019,N_21378);
or U21892 (N_21892,N_21461,N_21457);
nand U21893 (N_21893,N_21417,N_21176);
nor U21894 (N_21894,N_21427,N_21029);
xor U21895 (N_21895,N_21249,N_21464);
and U21896 (N_21896,N_21083,N_21264);
and U21897 (N_21897,N_21235,N_21122);
nor U21898 (N_21898,N_21487,N_21422);
or U21899 (N_21899,N_21263,N_21106);
nand U21900 (N_21900,N_21207,N_21468);
xnor U21901 (N_21901,N_21383,N_21288);
nor U21902 (N_21902,N_21182,N_21210);
nor U21903 (N_21903,N_21321,N_21413);
and U21904 (N_21904,N_21307,N_21047);
or U21905 (N_21905,N_21297,N_21129);
and U21906 (N_21906,N_21336,N_21400);
nor U21907 (N_21907,N_21456,N_21301);
nor U21908 (N_21908,N_21309,N_21357);
nand U21909 (N_21909,N_21183,N_21181);
and U21910 (N_21910,N_21170,N_21165);
nand U21911 (N_21911,N_21079,N_21172);
nand U21912 (N_21912,N_21266,N_21046);
and U21913 (N_21913,N_21221,N_21074);
nor U21914 (N_21914,N_21443,N_21307);
nand U21915 (N_21915,N_21238,N_21470);
xnor U21916 (N_21916,N_21395,N_21276);
and U21917 (N_21917,N_21284,N_21442);
or U21918 (N_21918,N_21021,N_21396);
or U21919 (N_21919,N_21104,N_21018);
or U21920 (N_21920,N_21155,N_21404);
or U21921 (N_21921,N_21159,N_21197);
and U21922 (N_21922,N_21317,N_21320);
nor U21923 (N_21923,N_21428,N_21032);
nand U21924 (N_21924,N_21499,N_21404);
or U21925 (N_21925,N_21189,N_21136);
nor U21926 (N_21926,N_21174,N_21134);
and U21927 (N_21927,N_21174,N_21082);
nand U21928 (N_21928,N_21023,N_21001);
nor U21929 (N_21929,N_21328,N_21228);
and U21930 (N_21930,N_21152,N_21131);
or U21931 (N_21931,N_21377,N_21429);
nor U21932 (N_21932,N_21193,N_21135);
nand U21933 (N_21933,N_21089,N_21029);
nand U21934 (N_21934,N_21052,N_21448);
or U21935 (N_21935,N_21035,N_21298);
nand U21936 (N_21936,N_21023,N_21402);
and U21937 (N_21937,N_21047,N_21201);
and U21938 (N_21938,N_21403,N_21474);
nor U21939 (N_21939,N_21310,N_21033);
nand U21940 (N_21940,N_21406,N_21128);
and U21941 (N_21941,N_21008,N_21130);
or U21942 (N_21942,N_21214,N_21118);
and U21943 (N_21943,N_21192,N_21093);
nand U21944 (N_21944,N_21380,N_21486);
nand U21945 (N_21945,N_21236,N_21178);
or U21946 (N_21946,N_21108,N_21287);
nor U21947 (N_21947,N_21132,N_21447);
and U21948 (N_21948,N_21316,N_21060);
nand U21949 (N_21949,N_21242,N_21353);
xnor U21950 (N_21950,N_21305,N_21163);
or U21951 (N_21951,N_21392,N_21354);
nor U21952 (N_21952,N_21372,N_21277);
nor U21953 (N_21953,N_21217,N_21068);
and U21954 (N_21954,N_21050,N_21253);
and U21955 (N_21955,N_21343,N_21474);
and U21956 (N_21956,N_21437,N_21453);
nor U21957 (N_21957,N_21176,N_21199);
or U21958 (N_21958,N_21190,N_21338);
nor U21959 (N_21959,N_21393,N_21004);
nand U21960 (N_21960,N_21398,N_21465);
or U21961 (N_21961,N_21089,N_21231);
nand U21962 (N_21962,N_21155,N_21251);
nor U21963 (N_21963,N_21049,N_21118);
nor U21964 (N_21964,N_21123,N_21385);
and U21965 (N_21965,N_21118,N_21021);
nor U21966 (N_21966,N_21373,N_21253);
or U21967 (N_21967,N_21195,N_21128);
nand U21968 (N_21968,N_21230,N_21282);
nand U21969 (N_21969,N_21467,N_21324);
nand U21970 (N_21970,N_21247,N_21293);
nor U21971 (N_21971,N_21013,N_21422);
nand U21972 (N_21972,N_21333,N_21390);
and U21973 (N_21973,N_21203,N_21454);
and U21974 (N_21974,N_21313,N_21176);
or U21975 (N_21975,N_21259,N_21189);
or U21976 (N_21976,N_21012,N_21275);
and U21977 (N_21977,N_21223,N_21091);
nand U21978 (N_21978,N_21048,N_21088);
and U21979 (N_21979,N_21438,N_21391);
or U21980 (N_21980,N_21055,N_21250);
and U21981 (N_21981,N_21376,N_21113);
nor U21982 (N_21982,N_21213,N_21383);
or U21983 (N_21983,N_21410,N_21379);
nor U21984 (N_21984,N_21229,N_21281);
or U21985 (N_21985,N_21304,N_21078);
nor U21986 (N_21986,N_21038,N_21437);
nor U21987 (N_21987,N_21153,N_21435);
or U21988 (N_21988,N_21384,N_21071);
nand U21989 (N_21989,N_21026,N_21185);
nor U21990 (N_21990,N_21138,N_21451);
nor U21991 (N_21991,N_21241,N_21186);
or U21992 (N_21992,N_21379,N_21313);
or U21993 (N_21993,N_21143,N_21357);
or U21994 (N_21994,N_21441,N_21117);
or U21995 (N_21995,N_21067,N_21015);
and U21996 (N_21996,N_21067,N_21080);
nor U21997 (N_21997,N_21008,N_21067);
and U21998 (N_21998,N_21034,N_21370);
or U21999 (N_21999,N_21078,N_21292);
and U22000 (N_22000,N_21751,N_21592);
and U22001 (N_22001,N_21745,N_21564);
or U22002 (N_22002,N_21645,N_21691);
nand U22003 (N_22003,N_21897,N_21557);
or U22004 (N_22004,N_21898,N_21922);
or U22005 (N_22005,N_21789,N_21868);
and U22006 (N_22006,N_21579,N_21731);
xor U22007 (N_22007,N_21523,N_21967);
nand U22008 (N_22008,N_21906,N_21801);
and U22009 (N_22009,N_21627,N_21561);
nand U22010 (N_22010,N_21835,N_21762);
and U22011 (N_22011,N_21502,N_21988);
nand U22012 (N_22012,N_21573,N_21760);
and U22013 (N_22013,N_21935,N_21626);
or U22014 (N_22014,N_21952,N_21758);
nand U22015 (N_22015,N_21571,N_21820);
or U22016 (N_22016,N_21666,N_21742);
nor U22017 (N_22017,N_21697,N_21736);
nand U22018 (N_22018,N_21620,N_21668);
and U22019 (N_22019,N_21718,N_21955);
nand U22020 (N_22020,N_21830,N_21630);
nor U22021 (N_22021,N_21763,N_21601);
nor U22022 (N_22022,N_21800,N_21938);
xor U22023 (N_22023,N_21606,N_21750);
nand U22024 (N_22024,N_21546,N_21852);
and U22025 (N_22025,N_21901,N_21896);
and U22026 (N_22026,N_21554,N_21853);
and U22027 (N_22027,N_21851,N_21850);
and U22028 (N_22028,N_21644,N_21619);
and U22029 (N_22029,N_21859,N_21559);
and U22030 (N_22030,N_21844,N_21643);
nor U22031 (N_22031,N_21845,N_21791);
nand U22032 (N_22032,N_21699,N_21575);
nor U22033 (N_22033,N_21536,N_21693);
or U22034 (N_22034,N_21765,N_21858);
nand U22035 (N_22035,N_21539,N_21829);
and U22036 (N_22036,N_21827,N_21671);
nor U22037 (N_22037,N_21723,N_21681);
and U22038 (N_22038,N_21929,N_21719);
or U22039 (N_22039,N_21956,N_21819);
nor U22040 (N_22040,N_21538,N_21550);
nand U22041 (N_22041,N_21865,N_21680);
nor U22042 (N_22042,N_21921,N_21748);
nor U22043 (N_22043,N_21729,N_21872);
nand U22044 (N_22044,N_21962,N_21617);
nor U22045 (N_22045,N_21771,N_21641);
or U22046 (N_22046,N_21530,N_21517);
nor U22047 (N_22047,N_21586,N_21658);
or U22048 (N_22048,N_21522,N_21914);
nor U22049 (N_22049,N_21873,N_21806);
or U22050 (N_22050,N_21913,N_21700);
and U22051 (N_22051,N_21593,N_21945);
or U22052 (N_22052,N_21815,N_21973);
and U22053 (N_22053,N_21570,N_21611);
and U22054 (N_22054,N_21983,N_21741);
nor U22055 (N_22055,N_21552,N_21969);
nand U22056 (N_22056,N_21860,N_21650);
nand U22057 (N_22057,N_21826,N_21566);
xnor U22058 (N_22058,N_21889,N_21959);
nor U22059 (N_22059,N_21978,N_21678);
nor U22060 (N_22060,N_21995,N_21640);
nand U22061 (N_22061,N_21533,N_21932);
and U22062 (N_22062,N_21976,N_21908);
or U22063 (N_22063,N_21616,N_21847);
nand U22064 (N_22064,N_21508,N_21958);
nor U22065 (N_22065,N_21714,N_21949);
nand U22066 (N_22066,N_21796,N_21824);
or U22067 (N_22067,N_21597,N_21870);
xor U22068 (N_22068,N_21568,N_21500);
or U22069 (N_22069,N_21942,N_21934);
nand U22070 (N_22070,N_21946,N_21783);
and U22071 (N_22071,N_21940,N_21822);
nor U22072 (N_22072,N_21701,N_21948);
nand U22073 (N_22073,N_21986,N_21503);
and U22074 (N_22074,N_21738,N_21543);
nor U22075 (N_22075,N_21656,N_21866);
and U22076 (N_22076,N_21685,N_21687);
and U22077 (N_22077,N_21892,N_21980);
or U22078 (N_22078,N_21855,N_21707);
nor U22079 (N_22079,N_21911,N_21672);
nand U22080 (N_22080,N_21607,N_21977);
or U22081 (N_22081,N_21535,N_21902);
nand U22082 (N_22082,N_21909,N_21594);
nor U22083 (N_22083,N_21879,N_21628);
and U22084 (N_22084,N_21951,N_21518);
nor U22085 (N_22085,N_21505,N_21569);
and U22086 (N_22086,N_21657,N_21862);
and U22087 (N_22087,N_21524,N_21688);
nand U22088 (N_22088,N_21874,N_21917);
nand U22089 (N_22089,N_21516,N_21795);
nor U22090 (N_22090,N_21775,N_21534);
and U22091 (N_22091,N_21918,N_21884);
or U22092 (N_22092,N_21961,N_21825);
nand U22093 (N_22093,N_21904,N_21577);
and U22094 (N_22094,N_21928,N_21805);
nand U22095 (N_22095,N_21634,N_21910);
and U22096 (N_22096,N_21740,N_21793);
or U22097 (N_22097,N_21541,N_21581);
nor U22098 (N_22098,N_21567,N_21632);
or U22099 (N_22099,N_21997,N_21624);
or U22100 (N_22100,N_21991,N_21587);
and U22101 (N_22101,N_21596,N_21756);
and U22102 (N_22102,N_21814,N_21878);
xnor U22103 (N_22103,N_21583,N_21519);
or U22104 (N_22104,N_21834,N_21974);
nor U22105 (N_22105,N_21931,N_21966);
and U22106 (N_22106,N_21780,N_21778);
or U22107 (N_22107,N_21646,N_21547);
nor U22108 (N_22108,N_21836,N_21684);
or U22109 (N_22109,N_21916,N_21705);
and U22110 (N_22110,N_21711,N_21895);
and U22111 (N_22111,N_21669,N_21761);
nand U22112 (N_22112,N_21652,N_21725);
nor U22113 (N_22113,N_21580,N_21728);
and U22114 (N_22114,N_21944,N_21899);
or U22115 (N_22115,N_21506,N_21893);
and U22116 (N_22116,N_21529,N_21545);
xor U22117 (N_22117,N_21753,N_21832);
or U22118 (N_22118,N_21631,N_21989);
or U22119 (N_22119,N_21926,N_21953);
nand U22120 (N_22120,N_21735,N_21752);
or U22121 (N_22121,N_21754,N_21613);
nand U22122 (N_22122,N_21937,N_21817);
or U22123 (N_22123,N_21963,N_21578);
or U22124 (N_22124,N_21782,N_21885);
or U22125 (N_22125,N_21694,N_21662);
and U22126 (N_22126,N_21562,N_21603);
nor U22127 (N_22127,N_21722,N_21683);
nand U22128 (N_22128,N_21585,N_21553);
nand U22129 (N_22129,N_21689,N_21816);
or U22130 (N_22130,N_21621,N_21637);
nand U22131 (N_22131,N_21968,N_21837);
nand U22132 (N_22132,N_21831,N_21509);
and U22133 (N_22133,N_21883,N_21776);
nor U22134 (N_22134,N_21788,N_21739);
and U22135 (N_22135,N_21715,N_21786);
or U22136 (N_22136,N_21542,N_21664);
nor U22137 (N_22137,N_21987,N_21703);
and U22138 (N_22138,N_21724,N_21734);
or U22139 (N_22139,N_21727,N_21970);
or U22140 (N_22140,N_21591,N_21661);
and U22141 (N_22141,N_21840,N_21996);
nand U22142 (N_22142,N_21608,N_21674);
nor U22143 (N_22143,N_21686,N_21582);
nor U22144 (N_22144,N_21890,N_21981);
nand U22145 (N_22145,N_21784,N_21706);
or U22146 (N_22146,N_21954,N_21919);
nor U22147 (N_22147,N_21673,N_21900);
nor U22148 (N_22148,N_21695,N_21972);
nor U22149 (N_22149,N_21821,N_21856);
nand U22150 (N_22150,N_21807,N_21556);
nor U22151 (N_22151,N_21709,N_21894);
or U22152 (N_22152,N_21635,N_21998);
nand U22153 (N_22153,N_21623,N_21747);
or U22154 (N_22154,N_21712,N_21915);
and U22155 (N_22155,N_21609,N_21993);
and U22156 (N_22156,N_21941,N_21861);
nand U22157 (N_22157,N_21867,N_21598);
or U22158 (N_22158,N_21663,N_21651);
nand U22159 (N_22159,N_21599,N_21659);
nor U22160 (N_22160,N_21984,N_21804);
and U22161 (N_22161,N_21618,N_21720);
and U22162 (N_22162,N_21787,N_21794);
and U22163 (N_22163,N_21877,N_21511);
nor U22164 (N_22164,N_21841,N_21549);
and U22165 (N_22165,N_21649,N_21808);
nor U22166 (N_22166,N_21746,N_21614);
and U22167 (N_22167,N_21888,N_21696);
nor U22168 (N_22168,N_21513,N_21732);
nor U22169 (N_22169,N_21947,N_21797);
nor U22170 (N_22170,N_21766,N_21737);
or U22171 (N_22171,N_21558,N_21605);
nor U22172 (N_22172,N_21749,N_21743);
or U22173 (N_22173,N_21813,N_21982);
nor U22174 (N_22174,N_21653,N_21572);
or U22175 (N_22175,N_21713,N_21710);
and U22176 (N_22176,N_21773,N_21755);
or U22177 (N_22177,N_21810,N_21692);
nand U22178 (N_22178,N_21527,N_21957);
nand U22179 (N_22179,N_21768,N_21936);
and U22180 (N_22180,N_21702,N_21507);
and U22181 (N_22181,N_21759,N_21880);
nor U22182 (N_22182,N_21704,N_21504);
or U22183 (N_22183,N_21886,N_21823);
nand U22184 (N_22184,N_21544,N_21992);
or U22185 (N_22185,N_21679,N_21881);
nor U22186 (N_22186,N_21965,N_21767);
nor U22187 (N_22187,N_21876,N_21555);
nand U22188 (N_22188,N_21730,N_21802);
nor U22189 (N_22189,N_21690,N_21848);
and U22190 (N_22190,N_21799,N_21602);
and U22191 (N_22191,N_21833,N_21537);
nand U22192 (N_22192,N_21792,N_21521);
nand U22193 (N_22193,N_21924,N_21809);
and U22194 (N_22194,N_21708,N_21869);
or U22195 (N_22195,N_21975,N_21717);
and U22196 (N_22196,N_21525,N_21960);
or U22197 (N_22197,N_21846,N_21772);
nand U22198 (N_22198,N_21769,N_21595);
or U22199 (N_22199,N_21912,N_21777);
and U22200 (N_22200,N_21716,N_21584);
nand U22201 (N_22201,N_21667,N_21871);
nand U22202 (N_22202,N_21501,N_21744);
nor U22203 (N_22203,N_21994,N_21526);
and U22204 (N_22204,N_21907,N_21920);
nor U22205 (N_22205,N_21849,N_21604);
and U22206 (N_22206,N_21863,N_21629);
or U22207 (N_22207,N_21531,N_21857);
nor U22208 (N_22208,N_21574,N_21670);
and U22209 (N_22209,N_21638,N_21933);
nor U22210 (N_22210,N_21647,N_21764);
or U22211 (N_22211,N_21785,N_21864);
nor U22212 (N_22212,N_21677,N_21971);
or U22213 (N_22213,N_21639,N_21930);
or U22214 (N_22214,N_21811,N_21770);
or U22215 (N_22215,N_21903,N_21563);
or U22216 (N_22216,N_21774,N_21642);
nand U22217 (N_22217,N_21540,N_21512);
nand U22218 (N_22218,N_21633,N_21515);
nor U22219 (N_22219,N_21682,N_21950);
nand U22220 (N_22220,N_21985,N_21676);
nor U22221 (N_22221,N_21905,N_21842);
or U22222 (N_22222,N_21589,N_21979);
nand U22223 (N_22223,N_21615,N_21600);
nand U22224 (N_22224,N_21891,N_21939);
nor U22225 (N_22225,N_21576,N_21927);
nand U22226 (N_22226,N_21790,N_21565);
nor U22227 (N_22227,N_21514,N_21964);
nand U22228 (N_22228,N_21803,N_21828);
and U22229 (N_22229,N_21875,N_21551);
nor U22230 (N_22230,N_21532,N_21779);
nor U22231 (N_22231,N_21798,N_21854);
or U22232 (N_22232,N_21839,N_21610);
and U22233 (N_22233,N_21660,N_21733);
nor U22234 (N_22234,N_21812,N_21721);
and U22235 (N_22235,N_21625,N_21612);
xnor U22236 (N_22236,N_21838,N_21726);
or U22237 (N_22237,N_21675,N_21923);
nor U22238 (N_22238,N_21636,N_21528);
xnor U22239 (N_22239,N_21560,N_21843);
or U22240 (N_22240,N_21510,N_21990);
and U22241 (N_22241,N_21882,N_21665);
or U22242 (N_22242,N_21925,N_21654);
or U22243 (N_22243,N_21818,N_21999);
and U22244 (N_22244,N_21548,N_21520);
and U22245 (N_22245,N_21590,N_21757);
nor U22246 (N_22246,N_21698,N_21622);
nand U22247 (N_22247,N_21781,N_21655);
xor U22248 (N_22248,N_21648,N_21588);
and U22249 (N_22249,N_21887,N_21943);
and U22250 (N_22250,N_21576,N_21935);
or U22251 (N_22251,N_21752,N_21770);
nand U22252 (N_22252,N_21886,N_21918);
and U22253 (N_22253,N_21761,N_21520);
or U22254 (N_22254,N_21572,N_21532);
or U22255 (N_22255,N_21708,N_21718);
nor U22256 (N_22256,N_21548,N_21682);
or U22257 (N_22257,N_21740,N_21767);
nand U22258 (N_22258,N_21831,N_21693);
nor U22259 (N_22259,N_21541,N_21585);
and U22260 (N_22260,N_21773,N_21574);
nor U22261 (N_22261,N_21850,N_21609);
or U22262 (N_22262,N_21860,N_21870);
or U22263 (N_22263,N_21721,N_21817);
or U22264 (N_22264,N_21621,N_21738);
nor U22265 (N_22265,N_21575,N_21864);
xnor U22266 (N_22266,N_21842,N_21881);
nand U22267 (N_22267,N_21718,N_21799);
nor U22268 (N_22268,N_21817,N_21768);
nand U22269 (N_22269,N_21926,N_21891);
nor U22270 (N_22270,N_21807,N_21870);
or U22271 (N_22271,N_21618,N_21573);
and U22272 (N_22272,N_21605,N_21749);
nor U22273 (N_22273,N_21740,N_21833);
and U22274 (N_22274,N_21613,N_21639);
or U22275 (N_22275,N_21670,N_21891);
or U22276 (N_22276,N_21530,N_21850);
or U22277 (N_22277,N_21930,N_21694);
nand U22278 (N_22278,N_21789,N_21821);
nor U22279 (N_22279,N_21957,N_21687);
xor U22280 (N_22280,N_21762,N_21543);
and U22281 (N_22281,N_21677,N_21992);
and U22282 (N_22282,N_21794,N_21873);
nor U22283 (N_22283,N_21640,N_21737);
xor U22284 (N_22284,N_21632,N_21677);
and U22285 (N_22285,N_21621,N_21510);
nor U22286 (N_22286,N_21534,N_21942);
nand U22287 (N_22287,N_21742,N_21761);
xor U22288 (N_22288,N_21608,N_21715);
nand U22289 (N_22289,N_21621,N_21819);
nor U22290 (N_22290,N_21624,N_21756);
and U22291 (N_22291,N_21800,N_21783);
or U22292 (N_22292,N_21912,N_21833);
nor U22293 (N_22293,N_21748,N_21566);
nand U22294 (N_22294,N_21853,N_21827);
or U22295 (N_22295,N_21794,N_21811);
nor U22296 (N_22296,N_21783,N_21993);
nor U22297 (N_22297,N_21563,N_21542);
and U22298 (N_22298,N_21993,N_21936);
and U22299 (N_22299,N_21905,N_21819);
and U22300 (N_22300,N_21550,N_21778);
or U22301 (N_22301,N_21833,N_21527);
nand U22302 (N_22302,N_21588,N_21628);
nor U22303 (N_22303,N_21569,N_21748);
xnor U22304 (N_22304,N_21946,N_21924);
nor U22305 (N_22305,N_21581,N_21730);
or U22306 (N_22306,N_21560,N_21694);
or U22307 (N_22307,N_21506,N_21579);
xor U22308 (N_22308,N_21579,N_21667);
or U22309 (N_22309,N_21630,N_21548);
nor U22310 (N_22310,N_21854,N_21588);
nor U22311 (N_22311,N_21910,N_21642);
nand U22312 (N_22312,N_21926,N_21674);
or U22313 (N_22313,N_21808,N_21940);
or U22314 (N_22314,N_21521,N_21636);
nand U22315 (N_22315,N_21728,N_21602);
and U22316 (N_22316,N_21613,N_21874);
and U22317 (N_22317,N_21653,N_21910);
and U22318 (N_22318,N_21645,N_21675);
or U22319 (N_22319,N_21831,N_21589);
nand U22320 (N_22320,N_21712,N_21717);
nand U22321 (N_22321,N_21636,N_21560);
or U22322 (N_22322,N_21528,N_21875);
xnor U22323 (N_22323,N_21592,N_21663);
nor U22324 (N_22324,N_21948,N_21655);
and U22325 (N_22325,N_21533,N_21785);
and U22326 (N_22326,N_21741,N_21965);
or U22327 (N_22327,N_21842,N_21643);
and U22328 (N_22328,N_21635,N_21644);
nor U22329 (N_22329,N_21580,N_21844);
or U22330 (N_22330,N_21934,N_21781);
nand U22331 (N_22331,N_21976,N_21620);
xor U22332 (N_22332,N_21549,N_21999);
nand U22333 (N_22333,N_21669,N_21882);
and U22334 (N_22334,N_21537,N_21982);
and U22335 (N_22335,N_21911,N_21560);
or U22336 (N_22336,N_21538,N_21986);
and U22337 (N_22337,N_21920,N_21851);
nand U22338 (N_22338,N_21553,N_21825);
or U22339 (N_22339,N_21610,N_21706);
and U22340 (N_22340,N_21893,N_21508);
or U22341 (N_22341,N_21916,N_21877);
nand U22342 (N_22342,N_21831,N_21844);
or U22343 (N_22343,N_21571,N_21628);
nor U22344 (N_22344,N_21635,N_21844);
or U22345 (N_22345,N_21577,N_21803);
nand U22346 (N_22346,N_21573,N_21925);
nor U22347 (N_22347,N_21735,N_21865);
nand U22348 (N_22348,N_21854,N_21961);
nor U22349 (N_22349,N_21553,N_21865);
and U22350 (N_22350,N_21718,N_21813);
nand U22351 (N_22351,N_21870,N_21600);
and U22352 (N_22352,N_21807,N_21536);
or U22353 (N_22353,N_21719,N_21989);
or U22354 (N_22354,N_21987,N_21692);
or U22355 (N_22355,N_21796,N_21545);
xnor U22356 (N_22356,N_21555,N_21631);
and U22357 (N_22357,N_21523,N_21609);
nand U22358 (N_22358,N_21995,N_21760);
or U22359 (N_22359,N_21929,N_21845);
nand U22360 (N_22360,N_21867,N_21503);
nor U22361 (N_22361,N_21629,N_21979);
nand U22362 (N_22362,N_21578,N_21892);
or U22363 (N_22363,N_21844,N_21987);
and U22364 (N_22364,N_21885,N_21926);
nand U22365 (N_22365,N_21873,N_21749);
and U22366 (N_22366,N_21526,N_21506);
and U22367 (N_22367,N_21606,N_21773);
nor U22368 (N_22368,N_21643,N_21756);
or U22369 (N_22369,N_21567,N_21530);
or U22370 (N_22370,N_21932,N_21834);
and U22371 (N_22371,N_21523,N_21868);
nand U22372 (N_22372,N_21904,N_21952);
or U22373 (N_22373,N_21604,N_21741);
and U22374 (N_22374,N_21655,N_21627);
or U22375 (N_22375,N_21519,N_21807);
and U22376 (N_22376,N_21648,N_21860);
and U22377 (N_22377,N_21538,N_21560);
or U22378 (N_22378,N_21544,N_21754);
and U22379 (N_22379,N_21907,N_21867);
or U22380 (N_22380,N_21555,N_21883);
or U22381 (N_22381,N_21657,N_21599);
nor U22382 (N_22382,N_21536,N_21695);
nor U22383 (N_22383,N_21638,N_21507);
nand U22384 (N_22384,N_21737,N_21525);
nor U22385 (N_22385,N_21665,N_21522);
nor U22386 (N_22386,N_21562,N_21561);
or U22387 (N_22387,N_21852,N_21777);
nand U22388 (N_22388,N_21604,N_21890);
or U22389 (N_22389,N_21536,N_21664);
nor U22390 (N_22390,N_21808,N_21809);
nor U22391 (N_22391,N_21569,N_21803);
or U22392 (N_22392,N_21589,N_21676);
or U22393 (N_22393,N_21971,N_21933);
nand U22394 (N_22394,N_21937,N_21722);
and U22395 (N_22395,N_21963,N_21656);
or U22396 (N_22396,N_21886,N_21839);
and U22397 (N_22397,N_21637,N_21866);
nand U22398 (N_22398,N_21641,N_21945);
and U22399 (N_22399,N_21787,N_21651);
and U22400 (N_22400,N_21633,N_21584);
nand U22401 (N_22401,N_21676,N_21679);
or U22402 (N_22402,N_21820,N_21598);
nand U22403 (N_22403,N_21564,N_21977);
or U22404 (N_22404,N_21596,N_21906);
or U22405 (N_22405,N_21813,N_21958);
nand U22406 (N_22406,N_21877,N_21698);
and U22407 (N_22407,N_21798,N_21809);
nand U22408 (N_22408,N_21588,N_21844);
or U22409 (N_22409,N_21969,N_21842);
and U22410 (N_22410,N_21918,N_21502);
and U22411 (N_22411,N_21982,N_21547);
and U22412 (N_22412,N_21981,N_21949);
or U22413 (N_22413,N_21826,N_21635);
and U22414 (N_22414,N_21861,N_21974);
and U22415 (N_22415,N_21817,N_21500);
and U22416 (N_22416,N_21554,N_21892);
or U22417 (N_22417,N_21642,N_21753);
nand U22418 (N_22418,N_21850,N_21914);
nand U22419 (N_22419,N_21746,N_21640);
nand U22420 (N_22420,N_21585,N_21611);
and U22421 (N_22421,N_21553,N_21524);
nor U22422 (N_22422,N_21616,N_21647);
nand U22423 (N_22423,N_21765,N_21545);
and U22424 (N_22424,N_21680,N_21709);
or U22425 (N_22425,N_21754,N_21801);
and U22426 (N_22426,N_21768,N_21872);
nor U22427 (N_22427,N_21702,N_21863);
nand U22428 (N_22428,N_21671,N_21979);
and U22429 (N_22429,N_21954,N_21974);
or U22430 (N_22430,N_21501,N_21891);
nor U22431 (N_22431,N_21712,N_21841);
or U22432 (N_22432,N_21851,N_21771);
nor U22433 (N_22433,N_21682,N_21876);
nand U22434 (N_22434,N_21539,N_21652);
and U22435 (N_22435,N_21601,N_21921);
or U22436 (N_22436,N_21982,N_21779);
or U22437 (N_22437,N_21907,N_21885);
nor U22438 (N_22438,N_21651,N_21613);
or U22439 (N_22439,N_21962,N_21846);
nand U22440 (N_22440,N_21766,N_21747);
or U22441 (N_22441,N_21754,N_21558);
and U22442 (N_22442,N_21998,N_21851);
xnor U22443 (N_22443,N_21937,N_21526);
nand U22444 (N_22444,N_21845,N_21803);
nor U22445 (N_22445,N_21596,N_21770);
and U22446 (N_22446,N_21554,N_21808);
and U22447 (N_22447,N_21657,N_21578);
nand U22448 (N_22448,N_21788,N_21867);
nand U22449 (N_22449,N_21649,N_21655);
or U22450 (N_22450,N_21845,N_21706);
nor U22451 (N_22451,N_21518,N_21559);
or U22452 (N_22452,N_21991,N_21678);
or U22453 (N_22453,N_21536,N_21968);
nor U22454 (N_22454,N_21820,N_21816);
xnor U22455 (N_22455,N_21752,N_21986);
or U22456 (N_22456,N_21889,N_21819);
xor U22457 (N_22457,N_21871,N_21959);
and U22458 (N_22458,N_21518,N_21643);
or U22459 (N_22459,N_21520,N_21628);
nor U22460 (N_22460,N_21749,N_21817);
nor U22461 (N_22461,N_21756,N_21862);
or U22462 (N_22462,N_21757,N_21621);
nor U22463 (N_22463,N_21647,N_21846);
nor U22464 (N_22464,N_21546,N_21880);
nor U22465 (N_22465,N_21657,N_21856);
nand U22466 (N_22466,N_21909,N_21844);
xor U22467 (N_22467,N_21799,N_21576);
nor U22468 (N_22468,N_21698,N_21888);
nand U22469 (N_22469,N_21602,N_21761);
xor U22470 (N_22470,N_21737,N_21682);
nor U22471 (N_22471,N_21729,N_21834);
or U22472 (N_22472,N_21847,N_21647);
nor U22473 (N_22473,N_21545,N_21783);
xor U22474 (N_22474,N_21520,N_21633);
or U22475 (N_22475,N_21908,N_21914);
xnor U22476 (N_22476,N_21672,N_21989);
nand U22477 (N_22477,N_21852,N_21523);
nand U22478 (N_22478,N_21541,N_21972);
nor U22479 (N_22479,N_21766,N_21799);
and U22480 (N_22480,N_21648,N_21787);
and U22481 (N_22481,N_21535,N_21546);
nand U22482 (N_22482,N_21991,N_21912);
or U22483 (N_22483,N_21822,N_21729);
or U22484 (N_22484,N_21501,N_21681);
nor U22485 (N_22485,N_21508,N_21988);
nand U22486 (N_22486,N_21641,N_21840);
nor U22487 (N_22487,N_21708,N_21864);
or U22488 (N_22488,N_21853,N_21729);
nand U22489 (N_22489,N_21906,N_21564);
or U22490 (N_22490,N_21715,N_21989);
nor U22491 (N_22491,N_21539,N_21931);
or U22492 (N_22492,N_21700,N_21664);
nor U22493 (N_22493,N_21847,N_21774);
nand U22494 (N_22494,N_21952,N_21812);
and U22495 (N_22495,N_21792,N_21552);
or U22496 (N_22496,N_21842,N_21996);
or U22497 (N_22497,N_21613,N_21657);
nor U22498 (N_22498,N_21978,N_21562);
or U22499 (N_22499,N_21917,N_21979);
or U22500 (N_22500,N_22345,N_22217);
nor U22501 (N_22501,N_22449,N_22138);
nand U22502 (N_22502,N_22036,N_22407);
or U22503 (N_22503,N_22215,N_22146);
and U22504 (N_22504,N_22135,N_22290);
nand U22505 (N_22505,N_22056,N_22488);
nor U22506 (N_22506,N_22192,N_22332);
nor U22507 (N_22507,N_22405,N_22053);
and U22508 (N_22508,N_22214,N_22177);
xnor U22509 (N_22509,N_22253,N_22481);
or U22510 (N_22510,N_22098,N_22152);
nand U22511 (N_22511,N_22161,N_22430);
nor U22512 (N_22512,N_22327,N_22188);
nor U22513 (N_22513,N_22049,N_22221);
and U22514 (N_22514,N_22220,N_22128);
xor U22515 (N_22515,N_22232,N_22442);
xnor U22516 (N_22516,N_22140,N_22424);
or U22517 (N_22517,N_22426,N_22122);
and U22518 (N_22518,N_22074,N_22459);
or U22519 (N_22519,N_22349,N_22101);
nor U22520 (N_22520,N_22237,N_22461);
or U22521 (N_22521,N_22246,N_22040);
or U22522 (N_22522,N_22045,N_22436);
and U22523 (N_22523,N_22409,N_22181);
nand U22524 (N_22524,N_22427,N_22124);
nand U22525 (N_22525,N_22269,N_22075);
or U22526 (N_22526,N_22372,N_22418);
nand U22527 (N_22527,N_22213,N_22277);
nand U22528 (N_22528,N_22414,N_22176);
and U22529 (N_22529,N_22208,N_22266);
or U22530 (N_22530,N_22463,N_22475);
nor U22531 (N_22531,N_22298,N_22301);
or U22532 (N_22532,N_22494,N_22103);
or U22533 (N_22533,N_22441,N_22136);
nand U22534 (N_22534,N_22235,N_22199);
or U22535 (N_22535,N_22394,N_22261);
nand U22536 (N_22536,N_22273,N_22472);
nand U22537 (N_22537,N_22064,N_22158);
and U22538 (N_22538,N_22489,N_22429);
or U22539 (N_22539,N_22094,N_22398);
or U22540 (N_22540,N_22385,N_22456);
or U22541 (N_22541,N_22381,N_22236);
nand U22542 (N_22542,N_22363,N_22331);
nor U22543 (N_22543,N_22174,N_22130);
nand U22544 (N_22544,N_22412,N_22018);
and U22545 (N_22545,N_22131,N_22454);
nand U22546 (N_22546,N_22346,N_22469);
xor U22547 (N_22547,N_22184,N_22497);
nor U22548 (N_22548,N_22229,N_22143);
nor U22549 (N_22549,N_22084,N_22058);
or U22550 (N_22550,N_22115,N_22330);
xor U22551 (N_22551,N_22466,N_22343);
and U22552 (N_22552,N_22299,N_22099);
nand U22553 (N_22553,N_22303,N_22032);
or U22554 (N_22554,N_22125,N_22060);
and U22555 (N_22555,N_22357,N_22317);
nand U22556 (N_22556,N_22274,N_22382);
nand U22557 (N_22557,N_22268,N_22193);
or U22558 (N_22558,N_22389,N_22209);
and U22559 (N_22559,N_22173,N_22322);
and U22560 (N_22560,N_22249,N_22123);
nor U22561 (N_22561,N_22106,N_22300);
nor U22562 (N_22562,N_22000,N_22051);
nor U22563 (N_22563,N_22403,N_22142);
and U22564 (N_22564,N_22314,N_22117);
nor U22565 (N_22565,N_22328,N_22082);
and U22566 (N_22566,N_22026,N_22254);
and U22567 (N_22567,N_22306,N_22226);
and U22568 (N_22568,N_22499,N_22211);
or U22569 (N_22569,N_22207,N_22189);
xor U22570 (N_22570,N_22460,N_22077);
and U22571 (N_22571,N_22440,N_22020);
nor U22572 (N_22572,N_22012,N_22218);
or U22573 (N_22573,N_22336,N_22042);
nor U22574 (N_22574,N_22295,N_22275);
nand U22575 (N_22575,N_22013,N_22419);
nor U22576 (N_22576,N_22183,N_22458);
and U22577 (N_22577,N_22410,N_22470);
nand U22578 (N_22578,N_22104,N_22379);
nor U22579 (N_22579,N_22234,N_22256);
nor U22580 (N_22580,N_22196,N_22009);
nand U22581 (N_22581,N_22052,N_22384);
and U22582 (N_22582,N_22411,N_22417);
nor U22583 (N_22583,N_22027,N_22392);
and U22584 (N_22584,N_22445,N_22493);
or U22585 (N_22585,N_22329,N_22021);
or U22586 (N_22586,N_22080,N_22423);
nand U22587 (N_22587,N_22413,N_22190);
and U22588 (N_22588,N_22359,N_22244);
or U22589 (N_22589,N_22151,N_22245);
xor U22590 (N_22590,N_22311,N_22157);
and U22591 (N_22591,N_22395,N_22309);
nor U22592 (N_22592,N_22149,N_22159);
or U22593 (N_22593,N_22388,N_22095);
or U22594 (N_22594,N_22492,N_22114);
or U22595 (N_22595,N_22019,N_22421);
xnor U22596 (N_22596,N_22031,N_22210);
nor U22597 (N_22597,N_22247,N_22010);
and U22598 (N_22598,N_22008,N_22017);
or U22599 (N_22599,N_22072,N_22304);
xor U22600 (N_22600,N_22371,N_22004);
and U22601 (N_22601,N_22281,N_22396);
nand U22602 (N_22602,N_22029,N_22356);
nand U22603 (N_22603,N_22422,N_22015);
nor U22604 (N_22604,N_22258,N_22167);
nand U22605 (N_22605,N_22370,N_22353);
xnor U22606 (N_22606,N_22486,N_22374);
and U22607 (N_22607,N_22453,N_22216);
and U22608 (N_22608,N_22487,N_22178);
nand U22609 (N_22609,N_22091,N_22348);
and U22610 (N_22610,N_22230,N_22086);
nor U22611 (N_22611,N_22083,N_22380);
nor U22612 (N_22612,N_22333,N_22366);
and U22613 (N_22613,N_22404,N_22483);
and U22614 (N_22614,N_22054,N_22476);
or U22615 (N_22615,N_22068,N_22102);
or U22616 (N_22616,N_22048,N_22164);
nand U22617 (N_22617,N_22358,N_22446);
and U22618 (N_22618,N_22393,N_22090);
and U22619 (N_22619,N_22153,N_22324);
nand U22620 (N_22620,N_22365,N_22172);
nor U22621 (N_22621,N_22201,N_22386);
nand U22622 (N_22622,N_22291,N_22457);
nand U22623 (N_22623,N_22239,N_22206);
and U22624 (N_22624,N_22255,N_22127);
nor U22625 (N_22625,N_22302,N_22464);
nand U22626 (N_22626,N_22110,N_22228);
nor U22627 (N_22627,N_22399,N_22028);
nor U22628 (N_22628,N_22062,N_22066);
or U22629 (N_22629,N_22484,N_22139);
nor U22630 (N_22630,N_22313,N_22342);
or U22631 (N_22631,N_22315,N_22420);
or U22632 (N_22632,N_22197,N_22265);
and U22633 (N_22633,N_22308,N_22204);
and U22634 (N_22634,N_22170,N_22334);
nor U22635 (N_22635,N_22276,N_22039);
nor U22636 (N_22636,N_22089,N_22444);
and U22637 (N_22637,N_22169,N_22355);
nand U22638 (N_22638,N_22431,N_22495);
nor U22639 (N_22639,N_22473,N_22002);
nor U22640 (N_22640,N_22182,N_22347);
nor U22641 (N_22641,N_22383,N_22294);
nor U22642 (N_22642,N_22034,N_22326);
and U22643 (N_22643,N_22191,N_22113);
nor U22644 (N_22644,N_22227,N_22280);
nor U22645 (N_22645,N_22162,N_22271);
and U22646 (N_22646,N_22369,N_22438);
nor U22647 (N_22647,N_22225,N_22364);
and U22648 (N_22648,N_22478,N_22319);
and U22649 (N_22649,N_22378,N_22137);
nand U22650 (N_22650,N_22030,N_22490);
nor U22651 (N_22651,N_22087,N_22272);
or U22652 (N_22652,N_22033,N_22022);
or U22653 (N_22653,N_22401,N_22248);
and U22654 (N_22654,N_22377,N_22352);
nor U22655 (N_22655,N_22006,N_22450);
or U22656 (N_22656,N_22433,N_22147);
nor U22657 (N_22657,N_22491,N_22439);
or U22658 (N_22658,N_22134,N_22150);
nor U22659 (N_22659,N_22025,N_22402);
or U22660 (N_22660,N_22325,N_22014);
and U22661 (N_22661,N_22376,N_22480);
or U22662 (N_22662,N_22482,N_22195);
or U22663 (N_22663,N_22425,N_22088);
and U22664 (N_22664,N_22263,N_22289);
or U22665 (N_22665,N_22387,N_22067);
nand U22666 (N_22666,N_22479,N_22344);
nand U22667 (N_22667,N_22148,N_22055);
xor U22668 (N_22668,N_22474,N_22282);
and U22669 (N_22669,N_22452,N_22233);
or U22670 (N_22670,N_22171,N_22292);
nor U22671 (N_22671,N_22121,N_22498);
nor U22672 (N_22672,N_22316,N_22118);
or U22673 (N_22673,N_22003,N_22362);
or U22674 (N_22674,N_22360,N_22341);
nor U22675 (N_22675,N_22375,N_22085);
nand U22676 (N_22676,N_22061,N_22477);
nor U22677 (N_22677,N_22203,N_22283);
and U22678 (N_22678,N_22465,N_22415);
nand U22679 (N_22679,N_22160,N_22156);
nor U22680 (N_22680,N_22408,N_22451);
or U22681 (N_22681,N_22496,N_22050);
nor U22682 (N_22682,N_22059,N_22185);
or U22683 (N_22683,N_22321,N_22023);
and U22684 (N_22684,N_22437,N_22416);
or U22685 (N_22685,N_22043,N_22223);
and U22686 (N_22686,N_22141,N_22285);
or U22687 (N_22687,N_22129,N_22462);
or U22688 (N_22688,N_22312,N_22270);
nor U22689 (N_22689,N_22205,N_22105);
and U22690 (N_22690,N_22447,N_22071);
and U22691 (N_22691,N_22337,N_22241);
or U22692 (N_22692,N_22400,N_22264);
or U22693 (N_22693,N_22097,N_22390);
nand U22694 (N_22694,N_22350,N_22455);
nand U22695 (N_22695,N_22297,N_22373);
and U22696 (N_22696,N_22250,N_22243);
nor U22697 (N_22697,N_22468,N_22079);
nor U22698 (N_22698,N_22168,N_22198);
or U22699 (N_22699,N_22259,N_22305);
and U22700 (N_22700,N_22070,N_22320);
nor U22701 (N_22701,N_22186,N_22187);
nand U22702 (N_22702,N_22180,N_22432);
nor U22703 (N_22703,N_22163,N_22367);
xor U22704 (N_22704,N_22323,N_22011);
and U22705 (N_22705,N_22262,N_22231);
and U22706 (N_22706,N_22286,N_22267);
nand U22707 (N_22707,N_22288,N_22222);
nor U22708 (N_22708,N_22368,N_22073);
nor U22709 (N_22709,N_22252,N_22044);
nor U22710 (N_22710,N_22351,N_22038);
and U22711 (N_22711,N_22108,N_22001);
xor U22712 (N_22712,N_22251,N_22078);
or U22713 (N_22713,N_22340,N_22179);
or U22714 (N_22714,N_22240,N_22391);
nor U22715 (N_22715,N_22257,N_22278);
nor U22716 (N_22716,N_22132,N_22111);
nand U22717 (N_22717,N_22096,N_22057);
nand U22718 (N_22718,N_22016,N_22144);
or U22719 (N_22719,N_22063,N_22485);
nand U22720 (N_22720,N_22194,N_22154);
and U22721 (N_22721,N_22007,N_22145);
and U22722 (N_22722,N_22339,N_22279);
and U22723 (N_22723,N_22112,N_22041);
nor U22724 (N_22724,N_22284,N_22116);
or U22725 (N_22725,N_22126,N_22081);
and U22726 (N_22726,N_22397,N_22069);
nand U22727 (N_22727,N_22093,N_22165);
or U22728 (N_22728,N_22260,N_22107);
and U22729 (N_22729,N_22133,N_22046);
and U22730 (N_22730,N_22448,N_22076);
and U22731 (N_22731,N_22200,N_22092);
nand U22732 (N_22732,N_22219,N_22293);
and U22733 (N_22733,N_22175,N_22202);
nor U22734 (N_22734,N_22435,N_22212);
nor U22735 (N_22735,N_22119,N_22024);
nor U22736 (N_22736,N_22361,N_22307);
nand U22737 (N_22737,N_22310,N_22047);
and U22738 (N_22738,N_22005,N_22287);
and U22739 (N_22739,N_22242,N_22035);
nand U22740 (N_22740,N_22155,N_22406);
or U22741 (N_22741,N_22338,N_22109);
nor U22742 (N_22742,N_22296,N_22335);
and U22743 (N_22743,N_22467,N_22434);
or U22744 (N_22744,N_22037,N_22443);
nand U22745 (N_22745,N_22120,N_22238);
or U22746 (N_22746,N_22166,N_22471);
nor U22747 (N_22747,N_22224,N_22354);
or U22748 (N_22748,N_22065,N_22100);
nor U22749 (N_22749,N_22428,N_22318);
nor U22750 (N_22750,N_22001,N_22323);
and U22751 (N_22751,N_22047,N_22087);
and U22752 (N_22752,N_22140,N_22330);
nand U22753 (N_22753,N_22245,N_22381);
nor U22754 (N_22754,N_22027,N_22253);
and U22755 (N_22755,N_22144,N_22196);
or U22756 (N_22756,N_22100,N_22165);
nor U22757 (N_22757,N_22246,N_22100);
or U22758 (N_22758,N_22304,N_22000);
nand U22759 (N_22759,N_22210,N_22332);
and U22760 (N_22760,N_22132,N_22250);
nand U22761 (N_22761,N_22138,N_22342);
nand U22762 (N_22762,N_22078,N_22454);
and U22763 (N_22763,N_22466,N_22230);
nor U22764 (N_22764,N_22022,N_22058);
or U22765 (N_22765,N_22369,N_22251);
nor U22766 (N_22766,N_22296,N_22184);
nor U22767 (N_22767,N_22040,N_22463);
nor U22768 (N_22768,N_22493,N_22169);
nor U22769 (N_22769,N_22019,N_22111);
nand U22770 (N_22770,N_22497,N_22355);
or U22771 (N_22771,N_22418,N_22104);
nor U22772 (N_22772,N_22479,N_22044);
nand U22773 (N_22773,N_22234,N_22081);
and U22774 (N_22774,N_22279,N_22082);
or U22775 (N_22775,N_22460,N_22084);
nand U22776 (N_22776,N_22194,N_22440);
and U22777 (N_22777,N_22045,N_22029);
or U22778 (N_22778,N_22123,N_22414);
and U22779 (N_22779,N_22222,N_22421);
or U22780 (N_22780,N_22222,N_22318);
nor U22781 (N_22781,N_22050,N_22001);
or U22782 (N_22782,N_22310,N_22343);
and U22783 (N_22783,N_22191,N_22330);
or U22784 (N_22784,N_22484,N_22188);
nor U22785 (N_22785,N_22213,N_22483);
nand U22786 (N_22786,N_22471,N_22174);
nand U22787 (N_22787,N_22438,N_22400);
or U22788 (N_22788,N_22296,N_22041);
or U22789 (N_22789,N_22174,N_22246);
nand U22790 (N_22790,N_22259,N_22006);
nand U22791 (N_22791,N_22052,N_22108);
and U22792 (N_22792,N_22426,N_22078);
nand U22793 (N_22793,N_22009,N_22352);
or U22794 (N_22794,N_22390,N_22386);
nand U22795 (N_22795,N_22085,N_22314);
or U22796 (N_22796,N_22235,N_22475);
nand U22797 (N_22797,N_22474,N_22184);
nand U22798 (N_22798,N_22352,N_22209);
or U22799 (N_22799,N_22363,N_22190);
and U22800 (N_22800,N_22368,N_22484);
or U22801 (N_22801,N_22064,N_22358);
and U22802 (N_22802,N_22339,N_22381);
xnor U22803 (N_22803,N_22390,N_22473);
and U22804 (N_22804,N_22280,N_22462);
or U22805 (N_22805,N_22247,N_22331);
and U22806 (N_22806,N_22161,N_22394);
nand U22807 (N_22807,N_22277,N_22441);
and U22808 (N_22808,N_22139,N_22367);
xor U22809 (N_22809,N_22132,N_22347);
and U22810 (N_22810,N_22202,N_22467);
and U22811 (N_22811,N_22238,N_22177);
nand U22812 (N_22812,N_22065,N_22396);
nor U22813 (N_22813,N_22169,N_22363);
nand U22814 (N_22814,N_22446,N_22141);
nand U22815 (N_22815,N_22030,N_22496);
nand U22816 (N_22816,N_22330,N_22170);
and U22817 (N_22817,N_22096,N_22046);
nand U22818 (N_22818,N_22347,N_22191);
and U22819 (N_22819,N_22212,N_22194);
nor U22820 (N_22820,N_22101,N_22292);
nor U22821 (N_22821,N_22438,N_22383);
xor U22822 (N_22822,N_22310,N_22026);
nand U22823 (N_22823,N_22304,N_22135);
or U22824 (N_22824,N_22231,N_22264);
nand U22825 (N_22825,N_22403,N_22256);
nor U22826 (N_22826,N_22022,N_22299);
nand U22827 (N_22827,N_22455,N_22333);
nor U22828 (N_22828,N_22336,N_22158);
nor U22829 (N_22829,N_22378,N_22223);
or U22830 (N_22830,N_22074,N_22296);
or U22831 (N_22831,N_22126,N_22114);
nor U22832 (N_22832,N_22114,N_22280);
nor U22833 (N_22833,N_22227,N_22024);
nand U22834 (N_22834,N_22418,N_22219);
nor U22835 (N_22835,N_22295,N_22317);
or U22836 (N_22836,N_22428,N_22142);
xnor U22837 (N_22837,N_22063,N_22227);
and U22838 (N_22838,N_22384,N_22422);
nor U22839 (N_22839,N_22097,N_22488);
nand U22840 (N_22840,N_22262,N_22225);
nor U22841 (N_22841,N_22356,N_22446);
nand U22842 (N_22842,N_22150,N_22133);
nand U22843 (N_22843,N_22414,N_22348);
nor U22844 (N_22844,N_22224,N_22111);
nor U22845 (N_22845,N_22404,N_22302);
and U22846 (N_22846,N_22233,N_22378);
and U22847 (N_22847,N_22491,N_22433);
nand U22848 (N_22848,N_22101,N_22100);
and U22849 (N_22849,N_22034,N_22328);
nor U22850 (N_22850,N_22219,N_22258);
nor U22851 (N_22851,N_22334,N_22066);
or U22852 (N_22852,N_22412,N_22413);
nor U22853 (N_22853,N_22072,N_22093);
and U22854 (N_22854,N_22152,N_22423);
or U22855 (N_22855,N_22489,N_22329);
nor U22856 (N_22856,N_22181,N_22395);
nand U22857 (N_22857,N_22291,N_22164);
or U22858 (N_22858,N_22429,N_22230);
nand U22859 (N_22859,N_22106,N_22354);
and U22860 (N_22860,N_22244,N_22296);
nand U22861 (N_22861,N_22445,N_22089);
or U22862 (N_22862,N_22254,N_22219);
nor U22863 (N_22863,N_22153,N_22286);
and U22864 (N_22864,N_22184,N_22401);
or U22865 (N_22865,N_22069,N_22314);
nand U22866 (N_22866,N_22164,N_22234);
and U22867 (N_22867,N_22013,N_22350);
xnor U22868 (N_22868,N_22260,N_22423);
nand U22869 (N_22869,N_22425,N_22281);
or U22870 (N_22870,N_22033,N_22094);
or U22871 (N_22871,N_22259,N_22304);
nor U22872 (N_22872,N_22148,N_22191);
and U22873 (N_22873,N_22388,N_22346);
or U22874 (N_22874,N_22121,N_22253);
and U22875 (N_22875,N_22415,N_22369);
and U22876 (N_22876,N_22192,N_22353);
nor U22877 (N_22877,N_22201,N_22080);
or U22878 (N_22878,N_22150,N_22336);
nand U22879 (N_22879,N_22075,N_22145);
nor U22880 (N_22880,N_22030,N_22123);
and U22881 (N_22881,N_22414,N_22325);
nor U22882 (N_22882,N_22493,N_22397);
nor U22883 (N_22883,N_22288,N_22360);
and U22884 (N_22884,N_22077,N_22271);
and U22885 (N_22885,N_22047,N_22266);
nand U22886 (N_22886,N_22007,N_22050);
nor U22887 (N_22887,N_22336,N_22087);
nand U22888 (N_22888,N_22448,N_22137);
or U22889 (N_22889,N_22412,N_22217);
and U22890 (N_22890,N_22447,N_22357);
nor U22891 (N_22891,N_22101,N_22252);
and U22892 (N_22892,N_22079,N_22328);
nor U22893 (N_22893,N_22317,N_22178);
nand U22894 (N_22894,N_22442,N_22058);
or U22895 (N_22895,N_22196,N_22461);
nor U22896 (N_22896,N_22287,N_22365);
nand U22897 (N_22897,N_22452,N_22278);
nand U22898 (N_22898,N_22414,N_22106);
nand U22899 (N_22899,N_22224,N_22335);
and U22900 (N_22900,N_22216,N_22247);
nand U22901 (N_22901,N_22021,N_22347);
nor U22902 (N_22902,N_22313,N_22168);
or U22903 (N_22903,N_22085,N_22129);
xnor U22904 (N_22904,N_22195,N_22293);
or U22905 (N_22905,N_22083,N_22081);
or U22906 (N_22906,N_22091,N_22280);
or U22907 (N_22907,N_22212,N_22186);
or U22908 (N_22908,N_22482,N_22182);
nand U22909 (N_22909,N_22273,N_22026);
nor U22910 (N_22910,N_22113,N_22162);
xnor U22911 (N_22911,N_22108,N_22155);
nor U22912 (N_22912,N_22485,N_22224);
xnor U22913 (N_22913,N_22394,N_22116);
xnor U22914 (N_22914,N_22066,N_22489);
nor U22915 (N_22915,N_22495,N_22073);
and U22916 (N_22916,N_22300,N_22046);
or U22917 (N_22917,N_22481,N_22331);
and U22918 (N_22918,N_22041,N_22168);
and U22919 (N_22919,N_22402,N_22498);
nand U22920 (N_22920,N_22456,N_22292);
nor U22921 (N_22921,N_22374,N_22407);
or U22922 (N_22922,N_22434,N_22317);
or U22923 (N_22923,N_22255,N_22396);
nand U22924 (N_22924,N_22061,N_22226);
and U22925 (N_22925,N_22305,N_22103);
and U22926 (N_22926,N_22116,N_22443);
or U22927 (N_22927,N_22230,N_22395);
nor U22928 (N_22928,N_22319,N_22278);
nand U22929 (N_22929,N_22192,N_22134);
nand U22930 (N_22930,N_22027,N_22109);
nor U22931 (N_22931,N_22467,N_22438);
and U22932 (N_22932,N_22100,N_22106);
nand U22933 (N_22933,N_22021,N_22442);
and U22934 (N_22934,N_22206,N_22183);
or U22935 (N_22935,N_22209,N_22264);
or U22936 (N_22936,N_22143,N_22039);
nand U22937 (N_22937,N_22335,N_22056);
nand U22938 (N_22938,N_22062,N_22257);
nand U22939 (N_22939,N_22103,N_22481);
nand U22940 (N_22940,N_22017,N_22211);
or U22941 (N_22941,N_22435,N_22294);
nand U22942 (N_22942,N_22172,N_22262);
or U22943 (N_22943,N_22492,N_22023);
or U22944 (N_22944,N_22420,N_22453);
nand U22945 (N_22945,N_22362,N_22186);
and U22946 (N_22946,N_22330,N_22064);
and U22947 (N_22947,N_22080,N_22242);
or U22948 (N_22948,N_22277,N_22248);
or U22949 (N_22949,N_22315,N_22111);
or U22950 (N_22950,N_22342,N_22031);
and U22951 (N_22951,N_22397,N_22402);
xnor U22952 (N_22952,N_22266,N_22399);
or U22953 (N_22953,N_22472,N_22299);
xnor U22954 (N_22954,N_22251,N_22386);
nand U22955 (N_22955,N_22213,N_22092);
or U22956 (N_22956,N_22413,N_22349);
nand U22957 (N_22957,N_22456,N_22086);
or U22958 (N_22958,N_22081,N_22214);
nand U22959 (N_22959,N_22431,N_22498);
nand U22960 (N_22960,N_22156,N_22305);
nor U22961 (N_22961,N_22126,N_22157);
and U22962 (N_22962,N_22273,N_22095);
or U22963 (N_22963,N_22280,N_22021);
or U22964 (N_22964,N_22089,N_22028);
and U22965 (N_22965,N_22195,N_22085);
xnor U22966 (N_22966,N_22452,N_22226);
or U22967 (N_22967,N_22389,N_22118);
nand U22968 (N_22968,N_22165,N_22398);
nor U22969 (N_22969,N_22286,N_22308);
nor U22970 (N_22970,N_22146,N_22357);
and U22971 (N_22971,N_22393,N_22477);
and U22972 (N_22972,N_22344,N_22015);
and U22973 (N_22973,N_22254,N_22354);
nand U22974 (N_22974,N_22271,N_22299);
nor U22975 (N_22975,N_22258,N_22223);
or U22976 (N_22976,N_22295,N_22276);
nor U22977 (N_22977,N_22389,N_22372);
nand U22978 (N_22978,N_22365,N_22165);
or U22979 (N_22979,N_22417,N_22488);
nand U22980 (N_22980,N_22153,N_22437);
or U22981 (N_22981,N_22213,N_22053);
or U22982 (N_22982,N_22241,N_22472);
or U22983 (N_22983,N_22364,N_22197);
or U22984 (N_22984,N_22306,N_22164);
or U22985 (N_22985,N_22154,N_22487);
or U22986 (N_22986,N_22194,N_22023);
or U22987 (N_22987,N_22277,N_22050);
nand U22988 (N_22988,N_22056,N_22467);
nor U22989 (N_22989,N_22013,N_22331);
or U22990 (N_22990,N_22045,N_22132);
xnor U22991 (N_22991,N_22467,N_22206);
nand U22992 (N_22992,N_22234,N_22208);
and U22993 (N_22993,N_22167,N_22178);
and U22994 (N_22994,N_22135,N_22097);
nand U22995 (N_22995,N_22249,N_22426);
and U22996 (N_22996,N_22276,N_22404);
or U22997 (N_22997,N_22094,N_22186);
and U22998 (N_22998,N_22113,N_22362);
nor U22999 (N_22999,N_22383,N_22271);
nor U23000 (N_23000,N_22778,N_22770);
nor U23001 (N_23001,N_22900,N_22783);
or U23002 (N_23002,N_22595,N_22654);
nor U23003 (N_23003,N_22898,N_22531);
nor U23004 (N_23004,N_22664,N_22622);
and U23005 (N_23005,N_22751,N_22677);
or U23006 (N_23006,N_22513,N_22982);
nor U23007 (N_23007,N_22652,N_22597);
or U23008 (N_23008,N_22808,N_22838);
or U23009 (N_23009,N_22594,N_22554);
and U23010 (N_23010,N_22533,N_22601);
or U23011 (N_23011,N_22715,N_22933);
nand U23012 (N_23012,N_22888,N_22873);
nand U23013 (N_23013,N_22766,N_22916);
or U23014 (N_23014,N_22700,N_22781);
nand U23015 (N_23015,N_22951,N_22719);
or U23016 (N_23016,N_22500,N_22882);
or U23017 (N_23017,N_22532,N_22977);
and U23018 (N_23018,N_22884,N_22910);
nor U23019 (N_23019,N_22924,N_22687);
or U23020 (N_23020,N_22596,N_22765);
nor U23021 (N_23021,N_22956,N_22976);
and U23022 (N_23022,N_22787,N_22780);
nor U23023 (N_23023,N_22648,N_22929);
nor U23024 (N_23024,N_22712,N_22608);
nand U23025 (N_23025,N_22737,N_22678);
nor U23026 (N_23026,N_22840,N_22742);
or U23027 (N_23027,N_22610,N_22852);
and U23028 (N_23028,N_22602,N_22588);
nand U23029 (N_23029,N_22729,N_22774);
or U23030 (N_23030,N_22576,N_22861);
or U23031 (N_23031,N_22739,N_22673);
nor U23032 (N_23032,N_22822,N_22948);
or U23033 (N_23033,N_22716,N_22828);
nor U23034 (N_23034,N_22809,N_22943);
and U23035 (N_23035,N_22544,N_22934);
nor U23036 (N_23036,N_22877,N_22674);
nor U23037 (N_23037,N_22680,N_22965);
nor U23038 (N_23038,N_22819,N_22502);
nand U23039 (N_23039,N_22559,N_22789);
nor U23040 (N_23040,N_22607,N_22816);
and U23041 (N_23041,N_22514,N_22893);
nor U23042 (N_23042,N_22573,N_22586);
and U23043 (N_23043,N_22646,N_22551);
or U23044 (N_23044,N_22829,N_22564);
and U23045 (N_23045,N_22871,N_22713);
nor U23046 (N_23046,N_22626,N_22504);
or U23047 (N_23047,N_22591,N_22940);
or U23048 (N_23048,N_22954,N_22639);
and U23049 (N_23049,N_22864,N_22662);
and U23050 (N_23050,N_22599,N_22722);
nor U23051 (N_23051,N_22911,N_22957);
or U23052 (N_23052,N_22708,N_22892);
and U23053 (N_23053,N_22688,N_22905);
and U23054 (N_23054,N_22736,N_22914);
nor U23055 (N_23055,N_22527,N_22878);
nand U23056 (N_23056,N_22981,N_22747);
or U23057 (N_23057,N_22521,N_22985);
or U23058 (N_23058,N_22969,N_22955);
nand U23059 (N_23059,N_22696,N_22704);
nand U23060 (N_23060,N_22947,N_22690);
or U23061 (N_23061,N_22714,N_22844);
nor U23062 (N_23062,N_22579,N_22836);
nor U23063 (N_23063,N_22753,N_22612);
xor U23064 (N_23064,N_22611,N_22860);
and U23065 (N_23065,N_22849,N_22624);
nand U23066 (N_23066,N_22746,N_22897);
or U23067 (N_23067,N_22847,N_22569);
nor U23068 (N_23068,N_22663,N_22889);
nor U23069 (N_23069,N_22867,N_22725);
and U23070 (N_23070,N_22592,N_22653);
and U23071 (N_23071,N_22857,N_22813);
xnor U23072 (N_23072,N_22817,N_22640);
or U23073 (N_23073,N_22906,N_22710);
nor U23074 (N_23074,N_22647,N_22635);
or U23075 (N_23075,N_22627,N_22772);
or U23076 (N_23076,N_22741,N_22509);
and U23077 (N_23077,N_22582,N_22988);
nor U23078 (N_23078,N_22613,N_22507);
xnor U23079 (N_23079,N_22668,N_22661);
nand U23080 (N_23080,N_22767,N_22788);
and U23081 (N_23081,N_22865,N_22973);
nor U23082 (N_23082,N_22936,N_22512);
or U23083 (N_23083,N_22517,N_22935);
nor U23084 (N_23084,N_22967,N_22744);
nand U23085 (N_23085,N_22644,N_22862);
and U23086 (N_23086,N_22631,N_22705);
nor U23087 (N_23087,N_22891,N_22868);
nor U23088 (N_23088,N_22600,N_22961);
and U23089 (N_23089,N_22880,N_22615);
nor U23090 (N_23090,N_22666,N_22682);
nand U23091 (N_23091,N_22895,N_22827);
xor U23092 (N_23092,N_22960,N_22566);
nand U23093 (N_23093,N_22510,N_22524);
or U23094 (N_23094,N_22536,N_22997);
and U23095 (N_23095,N_22970,N_22885);
nor U23096 (N_23096,N_22810,N_22537);
and U23097 (N_23097,N_22749,N_22790);
or U23098 (N_23098,N_22989,N_22686);
or U23099 (N_23099,N_22676,N_22665);
nor U23100 (N_23100,N_22562,N_22720);
nor U23101 (N_23101,N_22685,N_22855);
or U23102 (N_23102,N_22724,N_22769);
or U23103 (N_23103,N_22730,N_22598);
and U23104 (N_23104,N_22773,N_22726);
or U23105 (N_23105,N_22655,N_22750);
or U23106 (N_23106,N_22565,N_22587);
or U23107 (N_23107,N_22918,N_22999);
or U23108 (N_23108,N_22980,N_22603);
and U23109 (N_23109,N_22501,N_22814);
and U23110 (N_23110,N_22856,N_22638);
nor U23111 (N_23111,N_22754,N_22614);
or U23112 (N_23112,N_22558,N_22835);
nand U23113 (N_23113,N_22959,N_22886);
nor U23114 (N_23114,N_22830,N_22826);
nand U23115 (N_23115,N_22658,N_22629);
and U23116 (N_23116,N_22863,N_22693);
or U23117 (N_23117,N_22660,N_22733);
or U23118 (N_23118,N_22557,N_22505);
and U23119 (N_23119,N_22553,N_22987);
nand U23120 (N_23120,N_22938,N_22949);
and U23121 (N_23121,N_22831,N_22552);
nand U23122 (N_23122,N_22758,N_22991);
nor U23123 (N_23123,N_22541,N_22651);
and U23124 (N_23124,N_22757,N_22921);
nand U23125 (N_23125,N_22572,N_22728);
or U23126 (N_23126,N_22815,N_22723);
nor U23127 (N_23127,N_22944,N_22529);
and U23128 (N_23128,N_22593,N_22883);
and U23129 (N_23129,N_22833,N_22811);
or U23130 (N_23130,N_22768,N_22937);
or U23131 (N_23131,N_22798,N_22584);
or U23132 (N_23132,N_22546,N_22590);
nor U23133 (N_23133,N_22968,N_22571);
and U23134 (N_23134,N_22801,N_22854);
or U23135 (N_23135,N_22657,N_22745);
nand U23136 (N_23136,N_22515,N_22667);
xnor U23137 (N_23137,N_22709,N_22915);
and U23138 (N_23138,N_22996,N_22528);
nor U23139 (N_23139,N_22649,N_22858);
nand U23140 (N_23140,N_22926,N_22998);
and U23141 (N_23141,N_22542,N_22670);
and U23142 (N_23142,N_22669,N_22843);
or U23143 (N_23143,N_22776,N_22881);
and U23144 (N_23144,N_22917,N_22605);
and U23145 (N_23145,N_22625,N_22691);
nand U23146 (N_23146,N_22630,N_22995);
and U23147 (N_23147,N_22548,N_22518);
and U23148 (N_23148,N_22894,N_22837);
or U23149 (N_23149,N_22832,N_22621);
or U23150 (N_23150,N_22699,N_22941);
or U23151 (N_23151,N_22642,N_22841);
and U23152 (N_23152,N_22805,N_22609);
or U23153 (N_23153,N_22866,N_22923);
nor U23154 (N_23154,N_22913,N_22922);
or U23155 (N_23155,N_22797,N_22577);
and U23156 (N_23156,N_22618,N_22679);
and U23157 (N_23157,N_22872,N_22526);
or U23158 (N_23158,N_22683,N_22748);
and U23159 (N_23159,N_22727,N_22784);
nand U23160 (N_23160,N_22978,N_22522);
nand U23161 (N_23161,N_22763,N_22800);
nor U23162 (N_23162,N_22964,N_22907);
nor U23163 (N_23163,N_22692,N_22650);
or U23164 (N_23164,N_22901,N_22698);
nor U23165 (N_23165,N_22792,N_22799);
nand U23166 (N_23166,N_22759,N_22636);
nand U23167 (N_23167,N_22516,N_22834);
or U23168 (N_23168,N_22549,N_22874);
and U23169 (N_23169,N_22643,N_22848);
and U23170 (N_23170,N_22920,N_22899);
and U23171 (N_23171,N_22534,N_22634);
or U23172 (N_23172,N_22623,N_22561);
or U23173 (N_23173,N_22619,N_22839);
nor U23174 (N_23174,N_22909,N_22850);
nand U23175 (N_23175,N_22823,N_22953);
or U23176 (N_23176,N_22721,N_22620);
and U23177 (N_23177,N_22804,N_22701);
and U23178 (N_23178,N_22578,N_22616);
nor U23179 (N_23179,N_22606,N_22681);
nor U23180 (N_23180,N_22545,N_22740);
nand U23181 (N_23181,N_22779,N_22580);
and U23182 (N_23182,N_22966,N_22802);
nor U23183 (N_23183,N_22743,N_22931);
and U23184 (N_23184,N_22902,N_22927);
nor U23185 (N_23185,N_22846,N_22845);
and U23186 (N_23186,N_22684,N_22503);
and U23187 (N_23187,N_22912,N_22604);
nor U23188 (N_23188,N_22971,N_22942);
xor U23189 (N_23189,N_22568,N_22793);
and U23190 (N_23190,N_22842,N_22540);
and U23191 (N_23191,N_22875,N_22930);
nor U23192 (N_23192,N_22983,N_22851);
nand U23193 (N_23193,N_22575,N_22555);
and U23194 (N_23194,N_22718,N_22585);
nand U23195 (N_23195,N_22979,N_22695);
nand U23196 (N_23196,N_22950,N_22556);
and U23197 (N_23197,N_22786,N_22795);
or U23198 (N_23198,N_22656,N_22903);
or U23199 (N_23199,N_22818,N_22617);
and U23200 (N_23200,N_22694,N_22820);
nand U23201 (N_23201,N_22511,N_22543);
nor U23202 (N_23202,N_22530,N_22589);
and U23203 (N_23203,N_22732,N_22645);
nor U23204 (N_23204,N_22946,N_22952);
or U23205 (N_23205,N_22567,N_22869);
or U23206 (N_23206,N_22932,N_22734);
or U23207 (N_23207,N_22752,N_22994);
nand U23208 (N_23208,N_22972,N_22887);
and U23209 (N_23209,N_22896,N_22570);
and U23210 (N_23210,N_22928,N_22581);
and U23211 (N_23211,N_22574,N_22538);
nor U23212 (N_23212,N_22762,N_22539);
nor U23213 (N_23213,N_22707,N_22637);
nand U23214 (N_23214,N_22519,N_22975);
or U23215 (N_23215,N_22506,N_22919);
and U23216 (N_23216,N_22756,N_22782);
or U23217 (N_23217,N_22945,N_22993);
or U23218 (N_23218,N_22702,N_22628);
and U23219 (N_23219,N_22547,N_22870);
or U23220 (N_23220,N_22785,N_22523);
and U23221 (N_23221,N_22775,N_22632);
and U23222 (N_23222,N_22633,N_22706);
and U23223 (N_23223,N_22731,N_22703);
nor U23224 (N_23224,N_22761,N_22508);
nor U23225 (N_23225,N_22825,N_22992);
or U23226 (N_23226,N_22807,N_22876);
or U23227 (N_23227,N_22520,N_22890);
and U23228 (N_23228,N_22904,N_22984);
or U23229 (N_23229,N_22908,N_22963);
or U23230 (N_23230,N_22689,N_22986);
and U23231 (N_23231,N_22939,N_22738);
xnor U23232 (N_23232,N_22717,N_22806);
nand U23233 (N_23233,N_22764,N_22794);
nor U23234 (N_23234,N_22824,N_22735);
nand U23235 (N_23235,N_22525,N_22755);
nand U23236 (N_23236,N_22879,N_22796);
and U23237 (N_23237,N_22925,N_22760);
nor U23238 (N_23238,N_22711,N_22550);
and U23239 (N_23239,N_22962,N_22563);
and U23240 (N_23240,N_22990,N_22803);
and U23241 (N_23241,N_22659,N_22697);
nand U23242 (N_23242,N_22777,N_22535);
nor U23243 (N_23243,N_22791,N_22853);
and U23244 (N_23244,N_22672,N_22560);
and U23245 (N_23245,N_22641,N_22974);
and U23246 (N_23246,N_22675,N_22671);
nor U23247 (N_23247,N_22859,N_22771);
nor U23248 (N_23248,N_22812,N_22958);
nand U23249 (N_23249,N_22821,N_22583);
nand U23250 (N_23250,N_22603,N_22540);
and U23251 (N_23251,N_22955,N_22836);
or U23252 (N_23252,N_22692,N_22962);
and U23253 (N_23253,N_22814,N_22510);
nand U23254 (N_23254,N_22629,N_22977);
xor U23255 (N_23255,N_22915,N_22828);
or U23256 (N_23256,N_22942,N_22861);
nand U23257 (N_23257,N_22510,N_22852);
nand U23258 (N_23258,N_22671,N_22993);
and U23259 (N_23259,N_22543,N_22889);
or U23260 (N_23260,N_22506,N_22826);
or U23261 (N_23261,N_22747,N_22673);
and U23262 (N_23262,N_22827,N_22866);
or U23263 (N_23263,N_22908,N_22722);
nand U23264 (N_23264,N_22909,N_22503);
or U23265 (N_23265,N_22770,N_22633);
and U23266 (N_23266,N_22535,N_22525);
and U23267 (N_23267,N_22630,N_22737);
nand U23268 (N_23268,N_22666,N_22778);
nor U23269 (N_23269,N_22881,N_22866);
nor U23270 (N_23270,N_22881,N_22992);
or U23271 (N_23271,N_22933,N_22732);
nor U23272 (N_23272,N_22761,N_22711);
nand U23273 (N_23273,N_22586,N_22617);
or U23274 (N_23274,N_22531,N_22737);
and U23275 (N_23275,N_22530,N_22958);
nor U23276 (N_23276,N_22750,N_22746);
nand U23277 (N_23277,N_22786,N_22557);
nand U23278 (N_23278,N_22851,N_22636);
nor U23279 (N_23279,N_22766,N_22674);
nor U23280 (N_23280,N_22776,N_22689);
nor U23281 (N_23281,N_22760,N_22803);
nand U23282 (N_23282,N_22677,N_22975);
nand U23283 (N_23283,N_22986,N_22993);
or U23284 (N_23284,N_22926,N_22826);
nand U23285 (N_23285,N_22783,N_22693);
and U23286 (N_23286,N_22875,N_22884);
nor U23287 (N_23287,N_22586,N_22996);
nor U23288 (N_23288,N_22504,N_22734);
nor U23289 (N_23289,N_22705,N_22860);
and U23290 (N_23290,N_22910,N_22951);
and U23291 (N_23291,N_22542,N_22736);
nor U23292 (N_23292,N_22522,N_22957);
or U23293 (N_23293,N_22930,N_22674);
nand U23294 (N_23294,N_22947,N_22541);
or U23295 (N_23295,N_22918,N_22691);
and U23296 (N_23296,N_22747,N_22849);
nand U23297 (N_23297,N_22747,N_22877);
and U23298 (N_23298,N_22700,N_22647);
nor U23299 (N_23299,N_22946,N_22696);
nor U23300 (N_23300,N_22607,N_22814);
and U23301 (N_23301,N_22927,N_22922);
nor U23302 (N_23302,N_22567,N_22528);
or U23303 (N_23303,N_22923,N_22869);
nand U23304 (N_23304,N_22816,N_22678);
nand U23305 (N_23305,N_22928,N_22507);
or U23306 (N_23306,N_22753,N_22638);
nand U23307 (N_23307,N_22549,N_22870);
or U23308 (N_23308,N_22796,N_22936);
or U23309 (N_23309,N_22997,N_22956);
nand U23310 (N_23310,N_22639,N_22703);
and U23311 (N_23311,N_22978,N_22998);
and U23312 (N_23312,N_22695,N_22580);
xnor U23313 (N_23313,N_22603,N_22889);
nor U23314 (N_23314,N_22771,N_22921);
nor U23315 (N_23315,N_22941,N_22720);
or U23316 (N_23316,N_22849,N_22912);
and U23317 (N_23317,N_22822,N_22912);
nor U23318 (N_23318,N_22586,N_22609);
nand U23319 (N_23319,N_22668,N_22819);
and U23320 (N_23320,N_22851,N_22597);
or U23321 (N_23321,N_22911,N_22907);
nand U23322 (N_23322,N_22686,N_22643);
nand U23323 (N_23323,N_22745,N_22501);
nor U23324 (N_23324,N_22793,N_22859);
and U23325 (N_23325,N_22967,N_22617);
nand U23326 (N_23326,N_22523,N_22564);
nand U23327 (N_23327,N_22805,N_22592);
nor U23328 (N_23328,N_22590,N_22793);
or U23329 (N_23329,N_22823,N_22998);
nand U23330 (N_23330,N_22626,N_22535);
nand U23331 (N_23331,N_22657,N_22937);
or U23332 (N_23332,N_22753,N_22936);
and U23333 (N_23333,N_22860,N_22578);
and U23334 (N_23334,N_22503,N_22559);
nand U23335 (N_23335,N_22578,N_22591);
xor U23336 (N_23336,N_22858,N_22684);
and U23337 (N_23337,N_22792,N_22932);
nand U23338 (N_23338,N_22859,N_22776);
nand U23339 (N_23339,N_22978,N_22719);
nand U23340 (N_23340,N_22895,N_22801);
nand U23341 (N_23341,N_22972,N_22757);
nand U23342 (N_23342,N_22578,N_22730);
nor U23343 (N_23343,N_22568,N_22800);
nor U23344 (N_23344,N_22659,N_22843);
nand U23345 (N_23345,N_22927,N_22664);
nor U23346 (N_23346,N_22618,N_22766);
and U23347 (N_23347,N_22606,N_22804);
nand U23348 (N_23348,N_22514,N_22932);
and U23349 (N_23349,N_22771,N_22540);
and U23350 (N_23350,N_22548,N_22812);
nand U23351 (N_23351,N_22570,N_22864);
and U23352 (N_23352,N_22944,N_22780);
nand U23353 (N_23353,N_22779,N_22554);
nand U23354 (N_23354,N_22557,N_22609);
or U23355 (N_23355,N_22732,N_22921);
and U23356 (N_23356,N_22958,N_22732);
and U23357 (N_23357,N_22537,N_22871);
or U23358 (N_23358,N_22682,N_22866);
or U23359 (N_23359,N_22830,N_22712);
nand U23360 (N_23360,N_22605,N_22908);
or U23361 (N_23361,N_22680,N_22868);
or U23362 (N_23362,N_22757,N_22766);
and U23363 (N_23363,N_22982,N_22646);
nor U23364 (N_23364,N_22675,N_22724);
nor U23365 (N_23365,N_22836,N_22777);
nand U23366 (N_23366,N_22506,N_22977);
and U23367 (N_23367,N_22737,N_22954);
nor U23368 (N_23368,N_22627,N_22882);
or U23369 (N_23369,N_22848,N_22987);
or U23370 (N_23370,N_22721,N_22777);
xor U23371 (N_23371,N_22573,N_22529);
nand U23372 (N_23372,N_22705,N_22515);
or U23373 (N_23373,N_22626,N_22996);
nor U23374 (N_23374,N_22506,N_22936);
or U23375 (N_23375,N_22775,N_22767);
or U23376 (N_23376,N_22947,N_22909);
nand U23377 (N_23377,N_22545,N_22648);
nand U23378 (N_23378,N_22528,N_22897);
and U23379 (N_23379,N_22528,N_22932);
and U23380 (N_23380,N_22982,N_22866);
and U23381 (N_23381,N_22619,N_22821);
or U23382 (N_23382,N_22777,N_22946);
and U23383 (N_23383,N_22777,N_22815);
nor U23384 (N_23384,N_22600,N_22682);
nor U23385 (N_23385,N_22875,N_22747);
nand U23386 (N_23386,N_22914,N_22878);
and U23387 (N_23387,N_22883,N_22537);
nor U23388 (N_23388,N_22713,N_22953);
or U23389 (N_23389,N_22707,N_22746);
nor U23390 (N_23390,N_22920,N_22615);
and U23391 (N_23391,N_22862,N_22891);
or U23392 (N_23392,N_22718,N_22964);
nor U23393 (N_23393,N_22607,N_22697);
and U23394 (N_23394,N_22628,N_22867);
or U23395 (N_23395,N_22843,N_22748);
nor U23396 (N_23396,N_22870,N_22831);
nand U23397 (N_23397,N_22731,N_22723);
and U23398 (N_23398,N_22954,N_22775);
nor U23399 (N_23399,N_22902,N_22569);
nand U23400 (N_23400,N_22566,N_22762);
nor U23401 (N_23401,N_22751,N_22691);
and U23402 (N_23402,N_22703,N_22817);
nor U23403 (N_23403,N_22951,N_22790);
nand U23404 (N_23404,N_22916,N_22696);
and U23405 (N_23405,N_22500,N_22823);
and U23406 (N_23406,N_22803,N_22984);
nor U23407 (N_23407,N_22747,N_22967);
or U23408 (N_23408,N_22966,N_22714);
or U23409 (N_23409,N_22978,N_22610);
or U23410 (N_23410,N_22680,N_22590);
nor U23411 (N_23411,N_22780,N_22595);
nand U23412 (N_23412,N_22645,N_22578);
xor U23413 (N_23413,N_22630,N_22583);
and U23414 (N_23414,N_22931,N_22590);
and U23415 (N_23415,N_22742,N_22976);
nor U23416 (N_23416,N_22781,N_22573);
nor U23417 (N_23417,N_22856,N_22504);
or U23418 (N_23418,N_22950,N_22702);
and U23419 (N_23419,N_22891,N_22813);
nand U23420 (N_23420,N_22514,N_22564);
nand U23421 (N_23421,N_22997,N_22789);
nand U23422 (N_23422,N_22595,N_22882);
or U23423 (N_23423,N_22514,N_22717);
or U23424 (N_23424,N_22946,N_22864);
nand U23425 (N_23425,N_22677,N_22888);
nand U23426 (N_23426,N_22940,N_22919);
nand U23427 (N_23427,N_22928,N_22939);
and U23428 (N_23428,N_22515,N_22563);
or U23429 (N_23429,N_22752,N_22768);
or U23430 (N_23430,N_22960,N_22759);
or U23431 (N_23431,N_22968,N_22618);
and U23432 (N_23432,N_22754,N_22571);
nor U23433 (N_23433,N_22815,N_22585);
nand U23434 (N_23434,N_22558,N_22694);
and U23435 (N_23435,N_22916,N_22940);
or U23436 (N_23436,N_22558,N_22621);
and U23437 (N_23437,N_22693,N_22679);
nand U23438 (N_23438,N_22924,N_22859);
or U23439 (N_23439,N_22771,N_22721);
or U23440 (N_23440,N_22694,N_22898);
and U23441 (N_23441,N_22569,N_22582);
and U23442 (N_23442,N_22821,N_22770);
nand U23443 (N_23443,N_22740,N_22536);
nand U23444 (N_23444,N_22866,N_22868);
nor U23445 (N_23445,N_22506,N_22770);
nor U23446 (N_23446,N_22986,N_22825);
or U23447 (N_23447,N_22519,N_22863);
xor U23448 (N_23448,N_22886,N_22678);
nor U23449 (N_23449,N_22801,N_22783);
nor U23450 (N_23450,N_22763,N_22895);
or U23451 (N_23451,N_22663,N_22804);
nand U23452 (N_23452,N_22729,N_22700);
nand U23453 (N_23453,N_22578,N_22544);
nand U23454 (N_23454,N_22693,N_22516);
and U23455 (N_23455,N_22770,N_22865);
nor U23456 (N_23456,N_22727,N_22803);
nor U23457 (N_23457,N_22795,N_22698);
nor U23458 (N_23458,N_22986,N_22923);
and U23459 (N_23459,N_22994,N_22564);
nor U23460 (N_23460,N_22826,N_22613);
nor U23461 (N_23461,N_22535,N_22772);
nand U23462 (N_23462,N_22907,N_22560);
or U23463 (N_23463,N_22587,N_22854);
or U23464 (N_23464,N_22865,N_22634);
nor U23465 (N_23465,N_22715,N_22785);
and U23466 (N_23466,N_22587,N_22828);
or U23467 (N_23467,N_22687,N_22715);
or U23468 (N_23468,N_22535,N_22739);
or U23469 (N_23469,N_22973,N_22975);
or U23470 (N_23470,N_22503,N_22880);
and U23471 (N_23471,N_22567,N_22501);
or U23472 (N_23472,N_22896,N_22712);
nand U23473 (N_23473,N_22958,N_22767);
or U23474 (N_23474,N_22953,N_22547);
nor U23475 (N_23475,N_22890,N_22771);
or U23476 (N_23476,N_22821,N_22865);
nand U23477 (N_23477,N_22762,N_22608);
and U23478 (N_23478,N_22733,N_22824);
and U23479 (N_23479,N_22915,N_22651);
nand U23480 (N_23480,N_22859,N_22768);
nand U23481 (N_23481,N_22567,N_22761);
or U23482 (N_23482,N_22610,N_22806);
or U23483 (N_23483,N_22939,N_22737);
or U23484 (N_23484,N_22879,N_22543);
nor U23485 (N_23485,N_22772,N_22943);
or U23486 (N_23486,N_22678,N_22842);
nand U23487 (N_23487,N_22989,N_22704);
nand U23488 (N_23488,N_22939,N_22936);
and U23489 (N_23489,N_22686,N_22628);
nor U23490 (N_23490,N_22671,N_22869);
and U23491 (N_23491,N_22550,N_22527);
or U23492 (N_23492,N_22799,N_22729);
or U23493 (N_23493,N_22744,N_22958);
nor U23494 (N_23494,N_22980,N_22774);
nand U23495 (N_23495,N_22862,N_22754);
and U23496 (N_23496,N_22642,N_22767);
or U23497 (N_23497,N_22656,N_22675);
or U23498 (N_23498,N_22671,N_22924);
nor U23499 (N_23499,N_22750,N_22941);
nand U23500 (N_23500,N_23058,N_23080);
nor U23501 (N_23501,N_23256,N_23332);
and U23502 (N_23502,N_23338,N_23266);
or U23503 (N_23503,N_23213,N_23091);
and U23504 (N_23504,N_23104,N_23396);
xor U23505 (N_23505,N_23054,N_23372);
nor U23506 (N_23506,N_23201,N_23002);
nor U23507 (N_23507,N_23227,N_23063);
or U23508 (N_23508,N_23430,N_23277);
and U23509 (N_23509,N_23148,N_23168);
or U23510 (N_23510,N_23440,N_23371);
nor U23511 (N_23511,N_23131,N_23146);
and U23512 (N_23512,N_23454,N_23116);
and U23513 (N_23513,N_23314,N_23283);
or U23514 (N_23514,N_23427,N_23366);
nor U23515 (N_23515,N_23084,N_23078);
nand U23516 (N_23516,N_23175,N_23388);
or U23517 (N_23517,N_23181,N_23102);
nor U23518 (N_23518,N_23018,N_23313);
and U23519 (N_23519,N_23079,N_23022);
or U23520 (N_23520,N_23111,N_23318);
nand U23521 (N_23521,N_23024,N_23470);
and U23522 (N_23522,N_23297,N_23424);
or U23523 (N_23523,N_23236,N_23442);
nand U23524 (N_23524,N_23098,N_23334);
nand U23525 (N_23525,N_23103,N_23025);
or U23526 (N_23526,N_23423,N_23289);
nor U23527 (N_23527,N_23337,N_23479);
and U23528 (N_23528,N_23205,N_23413);
or U23529 (N_23529,N_23262,N_23385);
or U23530 (N_23530,N_23398,N_23188);
or U23531 (N_23531,N_23226,N_23077);
nor U23532 (N_23532,N_23214,N_23357);
and U23533 (N_23533,N_23157,N_23496);
nand U23534 (N_23534,N_23013,N_23351);
nand U23535 (N_23535,N_23363,N_23348);
nand U23536 (N_23536,N_23315,N_23153);
and U23537 (N_23537,N_23342,N_23039);
nor U23538 (N_23538,N_23187,N_23134);
and U23539 (N_23539,N_23382,N_23114);
nor U23540 (N_23540,N_23030,N_23036);
nand U23541 (N_23541,N_23034,N_23023);
nand U23542 (N_23542,N_23020,N_23355);
nand U23543 (N_23543,N_23112,N_23478);
nand U23544 (N_23544,N_23095,N_23405);
or U23545 (N_23545,N_23070,N_23051);
or U23546 (N_23546,N_23433,N_23097);
nor U23547 (N_23547,N_23065,N_23083);
nor U23548 (N_23548,N_23199,N_23137);
and U23549 (N_23549,N_23004,N_23075);
and U23550 (N_23550,N_23124,N_23027);
or U23551 (N_23551,N_23245,N_23269);
or U23552 (N_23552,N_23295,N_23109);
nand U23553 (N_23553,N_23298,N_23432);
or U23554 (N_23554,N_23375,N_23480);
nand U23555 (N_23555,N_23100,N_23136);
and U23556 (N_23556,N_23069,N_23368);
and U23557 (N_23557,N_23411,N_23280);
nor U23558 (N_23558,N_23177,N_23281);
or U23559 (N_23559,N_23333,N_23436);
and U23560 (N_23560,N_23200,N_23272);
nor U23561 (N_23561,N_23118,N_23191);
and U23562 (N_23562,N_23317,N_23174);
or U23563 (N_23563,N_23431,N_23127);
nand U23564 (N_23564,N_23434,N_23276);
nor U23565 (N_23565,N_23308,N_23453);
or U23566 (N_23566,N_23014,N_23021);
or U23567 (N_23567,N_23015,N_23448);
nand U23568 (N_23568,N_23085,N_23158);
nand U23569 (N_23569,N_23053,N_23230);
nand U23570 (N_23570,N_23271,N_23246);
nand U23571 (N_23571,N_23299,N_23067);
nand U23572 (N_23572,N_23251,N_23301);
and U23573 (N_23573,N_23467,N_23172);
xnor U23574 (N_23574,N_23441,N_23402);
xnor U23575 (N_23575,N_23452,N_23185);
or U23576 (N_23576,N_23352,N_23090);
nor U23577 (N_23577,N_23311,N_23003);
and U23578 (N_23578,N_23224,N_23081);
nor U23579 (N_23579,N_23183,N_23225);
nor U23580 (N_23580,N_23043,N_23354);
nand U23581 (N_23581,N_23273,N_23171);
nand U23582 (N_23582,N_23082,N_23426);
and U23583 (N_23583,N_23420,N_23147);
or U23584 (N_23584,N_23094,N_23016);
nand U23585 (N_23585,N_23017,N_23229);
nor U23586 (N_23586,N_23255,N_23198);
nand U23587 (N_23587,N_23046,N_23041);
and U23588 (N_23588,N_23302,N_23037);
nor U23589 (N_23589,N_23241,N_23463);
nand U23590 (N_23590,N_23044,N_23490);
and U23591 (N_23591,N_23155,N_23005);
nor U23592 (N_23592,N_23287,N_23362);
nor U23593 (N_23593,N_23048,N_23466);
or U23594 (N_23594,N_23344,N_23202);
and U23595 (N_23595,N_23373,N_23228);
nor U23596 (N_23596,N_23026,N_23438);
and U23597 (N_23597,N_23007,N_23055);
or U23598 (N_23598,N_23247,N_23406);
or U23599 (N_23599,N_23428,N_23166);
or U23600 (N_23600,N_23123,N_23459);
nand U23601 (N_23601,N_23437,N_23403);
or U23602 (N_23602,N_23365,N_23045);
and U23603 (N_23603,N_23410,N_23071);
and U23604 (N_23604,N_23110,N_23143);
and U23605 (N_23605,N_23475,N_23282);
xor U23606 (N_23606,N_23149,N_23107);
or U23607 (N_23607,N_23326,N_23339);
or U23608 (N_23608,N_23353,N_23290);
nor U23609 (N_23609,N_23291,N_23312);
nor U23610 (N_23610,N_23439,N_23401);
nor U23611 (N_23611,N_23378,N_23167);
or U23612 (N_23612,N_23047,N_23209);
and U23613 (N_23613,N_23320,N_23232);
nor U23614 (N_23614,N_23458,N_23243);
and U23615 (N_23615,N_23456,N_23343);
nor U23616 (N_23616,N_23483,N_23336);
nor U23617 (N_23617,N_23404,N_23161);
and U23618 (N_23618,N_23092,N_23040);
or U23619 (N_23619,N_23324,N_23093);
or U23620 (N_23620,N_23208,N_23195);
or U23621 (N_23621,N_23238,N_23105);
nand U23622 (N_23622,N_23369,N_23473);
or U23623 (N_23623,N_23341,N_23468);
xnor U23624 (N_23624,N_23196,N_23407);
or U23625 (N_23625,N_23474,N_23032);
or U23626 (N_23626,N_23493,N_23293);
and U23627 (N_23627,N_23260,N_23049);
or U23628 (N_23628,N_23258,N_23261);
nand U23629 (N_23629,N_23194,N_23292);
or U23630 (N_23630,N_23010,N_23253);
nor U23631 (N_23631,N_23239,N_23395);
nor U23632 (N_23632,N_23321,N_23323);
or U23633 (N_23633,N_23384,N_23160);
and U23634 (N_23634,N_23303,N_23165);
nand U23635 (N_23635,N_23099,N_23443);
nor U23636 (N_23636,N_23215,N_23274);
nand U23637 (N_23637,N_23487,N_23150);
nand U23638 (N_23638,N_23219,N_23488);
nand U23639 (N_23639,N_23435,N_23240);
nand U23640 (N_23640,N_23176,N_23184);
nor U23641 (N_23641,N_23122,N_23064);
and U23642 (N_23642,N_23476,N_23457);
nor U23643 (N_23643,N_23374,N_23163);
and U23644 (N_23644,N_23350,N_23212);
or U23645 (N_23645,N_23254,N_23275);
nand U23646 (N_23646,N_23364,N_23267);
nand U23647 (N_23647,N_23497,N_23033);
nor U23648 (N_23648,N_23115,N_23074);
and U23649 (N_23649,N_23197,N_23327);
and U23650 (N_23650,N_23244,N_23203);
nor U23651 (N_23651,N_23133,N_23190);
or U23652 (N_23652,N_23192,N_23285);
xnor U23653 (N_23653,N_23235,N_23499);
and U23654 (N_23654,N_23050,N_23242);
and U23655 (N_23655,N_23126,N_23135);
nor U23656 (N_23656,N_23231,N_23481);
nand U23657 (N_23657,N_23062,N_23057);
xnor U23658 (N_23658,N_23393,N_23223);
and U23659 (N_23659,N_23009,N_23394);
and U23660 (N_23660,N_23408,N_23304);
and U23661 (N_23661,N_23237,N_23361);
and U23662 (N_23662,N_23417,N_23462);
nand U23663 (N_23663,N_23307,N_23495);
or U23664 (N_23664,N_23060,N_23446);
nor U23665 (N_23665,N_23390,N_23117);
nand U23666 (N_23666,N_23310,N_23469);
nand U23667 (N_23667,N_23464,N_23391);
nor U23668 (N_23668,N_23444,N_23268);
nand U23669 (N_23669,N_23300,N_23059);
nor U23670 (N_23670,N_23449,N_23011);
and U23671 (N_23671,N_23141,N_23451);
and U23672 (N_23672,N_23316,N_23106);
nor U23673 (N_23673,N_23330,N_23001);
nand U23674 (N_23674,N_23429,N_23119);
nor U23675 (N_23675,N_23249,N_23073);
nor U23676 (N_23676,N_23221,N_23207);
or U23677 (N_23677,N_23360,N_23138);
or U23678 (N_23678,N_23328,N_23486);
or U23679 (N_23679,N_23121,N_23347);
and U23680 (N_23680,N_23380,N_23415);
nand U23681 (N_23681,N_23145,N_23471);
nor U23682 (N_23682,N_23250,N_23305);
nor U23683 (N_23683,N_23220,N_23409);
nor U23684 (N_23684,N_23445,N_23399);
xnor U23685 (N_23685,N_23485,N_23216);
and U23686 (N_23686,N_23477,N_23377);
and U23687 (N_23687,N_23492,N_23180);
or U23688 (N_23688,N_23489,N_23154);
or U23689 (N_23689,N_23340,N_23113);
and U23690 (N_23690,N_23211,N_23294);
nor U23691 (N_23691,N_23329,N_23056);
nor U23692 (N_23692,N_23358,N_23455);
and U23693 (N_23693,N_23346,N_23345);
or U23694 (N_23694,N_23000,N_23173);
and U23695 (N_23695,N_23265,N_23349);
nor U23696 (N_23696,N_23164,N_23263);
nand U23697 (N_23697,N_23386,N_23381);
or U23698 (N_23698,N_23387,N_23309);
nor U23699 (N_23699,N_23139,N_23159);
nor U23700 (N_23700,N_23465,N_23052);
or U23701 (N_23701,N_23248,N_23089);
nand U23702 (N_23702,N_23233,N_23156);
xnor U23703 (N_23703,N_23096,N_23144);
nand U23704 (N_23704,N_23038,N_23484);
and U23705 (N_23705,N_23068,N_23482);
nor U23706 (N_23706,N_23331,N_23450);
nor U23707 (N_23707,N_23370,N_23425);
nor U23708 (N_23708,N_23006,N_23028);
nand U23709 (N_23709,N_23412,N_23204);
nor U23710 (N_23710,N_23008,N_23414);
nand U23711 (N_23711,N_23400,N_23072);
and U23712 (N_23712,N_23151,N_23472);
nand U23713 (N_23713,N_23418,N_23498);
and U23714 (N_23714,N_23035,N_23029);
xor U23715 (N_23715,N_23257,N_23120);
and U23716 (N_23716,N_23142,N_23367);
and U23717 (N_23717,N_23019,N_23335);
nor U23718 (N_23718,N_23288,N_23461);
nand U23719 (N_23719,N_23042,N_23132);
or U23720 (N_23720,N_23319,N_23379);
nor U23721 (N_23721,N_23088,N_23169);
or U23722 (N_23722,N_23162,N_23189);
nand U23723 (N_23723,N_23031,N_23306);
nor U23724 (N_23724,N_23128,N_23270);
nand U23725 (N_23725,N_23222,N_23125);
or U23726 (N_23726,N_23356,N_23129);
or U23727 (N_23727,N_23259,N_23076);
and U23728 (N_23728,N_23359,N_23494);
and U23729 (N_23729,N_23130,N_23422);
and U23730 (N_23730,N_23108,N_23178);
or U23731 (N_23731,N_23252,N_23086);
nor U23732 (N_23732,N_23284,N_23322);
or U23733 (N_23733,N_23389,N_23012);
or U23734 (N_23734,N_23376,N_23210);
and U23735 (N_23735,N_23325,N_23279);
and U23736 (N_23736,N_23397,N_23460);
and U23737 (N_23737,N_23286,N_23087);
and U23738 (N_23738,N_23218,N_23383);
nor U23739 (N_23739,N_23186,N_23140);
or U23740 (N_23740,N_23491,N_23179);
or U23741 (N_23741,N_23447,N_23061);
or U23742 (N_23742,N_23182,N_23193);
and U23743 (N_23743,N_23234,N_23416);
or U23744 (N_23744,N_23217,N_23101);
nor U23745 (N_23745,N_23170,N_23206);
and U23746 (N_23746,N_23419,N_23066);
and U23747 (N_23747,N_23296,N_23392);
and U23748 (N_23748,N_23421,N_23264);
or U23749 (N_23749,N_23152,N_23278);
and U23750 (N_23750,N_23313,N_23300);
or U23751 (N_23751,N_23025,N_23252);
or U23752 (N_23752,N_23351,N_23310);
and U23753 (N_23753,N_23006,N_23250);
nor U23754 (N_23754,N_23486,N_23210);
nor U23755 (N_23755,N_23339,N_23142);
nor U23756 (N_23756,N_23488,N_23492);
or U23757 (N_23757,N_23162,N_23218);
and U23758 (N_23758,N_23369,N_23301);
nand U23759 (N_23759,N_23326,N_23300);
nand U23760 (N_23760,N_23113,N_23425);
nand U23761 (N_23761,N_23498,N_23481);
nand U23762 (N_23762,N_23297,N_23470);
or U23763 (N_23763,N_23239,N_23481);
or U23764 (N_23764,N_23458,N_23068);
nor U23765 (N_23765,N_23276,N_23021);
and U23766 (N_23766,N_23222,N_23165);
and U23767 (N_23767,N_23005,N_23018);
or U23768 (N_23768,N_23279,N_23066);
and U23769 (N_23769,N_23173,N_23472);
or U23770 (N_23770,N_23143,N_23390);
and U23771 (N_23771,N_23154,N_23226);
nor U23772 (N_23772,N_23355,N_23234);
and U23773 (N_23773,N_23121,N_23496);
xor U23774 (N_23774,N_23372,N_23404);
and U23775 (N_23775,N_23387,N_23060);
nor U23776 (N_23776,N_23249,N_23305);
and U23777 (N_23777,N_23011,N_23087);
nor U23778 (N_23778,N_23271,N_23360);
nor U23779 (N_23779,N_23278,N_23177);
nor U23780 (N_23780,N_23237,N_23312);
nand U23781 (N_23781,N_23172,N_23255);
nor U23782 (N_23782,N_23193,N_23231);
or U23783 (N_23783,N_23371,N_23116);
and U23784 (N_23784,N_23303,N_23363);
or U23785 (N_23785,N_23031,N_23042);
nor U23786 (N_23786,N_23004,N_23105);
or U23787 (N_23787,N_23391,N_23050);
or U23788 (N_23788,N_23083,N_23009);
nor U23789 (N_23789,N_23436,N_23075);
nor U23790 (N_23790,N_23452,N_23233);
and U23791 (N_23791,N_23223,N_23300);
or U23792 (N_23792,N_23386,N_23091);
and U23793 (N_23793,N_23100,N_23386);
nand U23794 (N_23794,N_23478,N_23373);
and U23795 (N_23795,N_23300,N_23204);
nand U23796 (N_23796,N_23483,N_23062);
nor U23797 (N_23797,N_23171,N_23436);
and U23798 (N_23798,N_23000,N_23441);
nand U23799 (N_23799,N_23468,N_23065);
xor U23800 (N_23800,N_23188,N_23169);
nand U23801 (N_23801,N_23171,N_23023);
and U23802 (N_23802,N_23037,N_23401);
and U23803 (N_23803,N_23045,N_23382);
nand U23804 (N_23804,N_23155,N_23462);
or U23805 (N_23805,N_23170,N_23413);
and U23806 (N_23806,N_23056,N_23084);
xor U23807 (N_23807,N_23314,N_23386);
and U23808 (N_23808,N_23137,N_23424);
nor U23809 (N_23809,N_23150,N_23066);
nand U23810 (N_23810,N_23082,N_23430);
nor U23811 (N_23811,N_23176,N_23131);
nand U23812 (N_23812,N_23121,N_23182);
nor U23813 (N_23813,N_23226,N_23490);
nor U23814 (N_23814,N_23350,N_23266);
and U23815 (N_23815,N_23499,N_23026);
or U23816 (N_23816,N_23251,N_23398);
or U23817 (N_23817,N_23185,N_23475);
xor U23818 (N_23818,N_23426,N_23430);
and U23819 (N_23819,N_23381,N_23224);
xnor U23820 (N_23820,N_23404,N_23462);
nor U23821 (N_23821,N_23477,N_23140);
nor U23822 (N_23822,N_23190,N_23230);
and U23823 (N_23823,N_23076,N_23255);
or U23824 (N_23824,N_23355,N_23125);
nor U23825 (N_23825,N_23066,N_23285);
nor U23826 (N_23826,N_23470,N_23079);
or U23827 (N_23827,N_23223,N_23472);
nor U23828 (N_23828,N_23001,N_23357);
nand U23829 (N_23829,N_23188,N_23007);
and U23830 (N_23830,N_23433,N_23385);
and U23831 (N_23831,N_23180,N_23439);
or U23832 (N_23832,N_23275,N_23483);
or U23833 (N_23833,N_23382,N_23166);
nor U23834 (N_23834,N_23167,N_23371);
and U23835 (N_23835,N_23020,N_23109);
or U23836 (N_23836,N_23031,N_23311);
and U23837 (N_23837,N_23322,N_23261);
nand U23838 (N_23838,N_23137,N_23160);
or U23839 (N_23839,N_23087,N_23308);
or U23840 (N_23840,N_23052,N_23169);
nor U23841 (N_23841,N_23268,N_23109);
nor U23842 (N_23842,N_23030,N_23309);
nand U23843 (N_23843,N_23156,N_23311);
or U23844 (N_23844,N_23440,N_23355);
nor U23845 (N_23845,N_23417,N_23274);
nor U23846 (N_23846,N_23463,N_23402);
nand U23847 (N_23847,N_23023,N_23419);
nor U23848 (N_23848,N_23457,N_23233);
nor U23849 (N_23849,N_23239,N_23117);
and U23850 (N_23850,N_23019,N_23167);
or U23851 (N_23851,N_23301,N_23393);
and U23852 (N_23852,N_23100,N_23192);
nand U23853 (N_23853,N_23107,N_23157);
nand U23854 (N_23854,N_23372,N_23352);
and U23855 (N_23855,N_23277,N_23186);
or U23856 (N_23856,N_23043,N_23131);
or U23857 (N_23857,N_23392,N_23358);
nand U23858 (N_23858,N_23436,N_23180);
or U23859 (N_23859,N_23493,N_23059);
and U23860 (N_23860,N_23070,N_23166);
and U23861 (N_23861,N_23254,N_23478);
nand U23862 (N_23862,N_23131,N_23317);
nor U23863 (N_23863,N_23008,N_23206);
or U23864 (N_23864,N_23220,N_23151);
nand U23865 (N_23865,N_23388,N_23479);
nor U23866 (N_23866,N_23026,N_23298);
or U23867 (N_23867,N_23042,N_23272);
and U23868 (N_23868,N_23113,N_23284);
nand U23869 (N_23869,N_23214,N_23066);
or U23870 (N_23870,N_23037,N_23292);
and U23871 (N_23871,N_23408,N_23342);
and U23872 (N_23872,N_23364,N_23173);
nor U23873 (N_23873,N_23185,N_23372);
nor U23874 (N_23874,N_23304,N_23498);
and U23875 (N_23875,N_23377,N_23202);
and U23876 (N_23876,N_23470,N_23445);
nand U23877 (N_23877,N_23031,N_23072);
nor U23878 (N_23878,N_23227,N_23184);
nand U23879 (N_23879,N_23278,N_23222);
and U23880 (N_23880,N_23440,N_23182);
nand U23881 (N_23881,N_23122,N_23169);
and U23882 (N_23882,N_23017,N_23133);
and U23883 (N_23883,N_23143,N_23389);
and U23884 (N_23884,N_23497,N_23012);
and U23885 (N_23885,N_23375,N_23162);
or U23886 (N_23886,N_23423,N_23199);
nor U23887 (N_23887,N_23134,N_23342);
nand U23888 (N_23888,N_23178,N_23127);
nand U23889 (N_23889,N_23412,N_23237);
nand U23890 (N_23890,N_23082,N_23384);
nor U23891 (N_23891,N_23322,N_23225);
nand U23892 (N_23892,N_23201,N_23087);
nor U23893 (N_23893,N_23412,N_23481);
and U23894 (N_23894,N_23106,N_23030);
nor U23895 (N_23895,N_23292,N_23447);
nor U23896 (N_23896,N_23476,N_23315);
and U23897 (N_23897,N_23242,N_23320);
nand U23898 (N_23898,N_23266,N_23496);
and U23899 (N_23899,N_23277,N_23062);
and U23900 (N_23900,N_23451,N_23060);
nand U23901 (N_23901,N_23393,N_23164);
nor U23902 (N_23902,N_23372,N_23308);
and U23903 (N_23903,N_23241,N_23169);
nor U23904 (N_23904,N_23028,N_23163);
and U23905 (N_23905,N_23013,N_23103);
nor U23906 (N_23906,N_23363,N_23082);
nor U23907 (N_23907,N_23413,N_23491);
nand U23908 (N_23908,N_23424,N_23074);
and U23909 (N_23909,N_23059,N_23183);
nand U23910 (N_23910,N_23346,N_23054);
or U23911 (N_23911,N_23426,N_23157);
nand U23912 (N_23912,N_23374,N_23232);
nand U23913 (N_23913,N_23445,N_23353);
or U23914 (N_23914,N_23334,N_23373);
nor U23915 (N_23915,N_23354,N_23390);
nor U23916 (N_23916,N_23497,N_23442);
nand U23917 (N_23917,N_23012,N_23091);
nand U23918 (N_23918,N_23127,N_23374);
nand U23919 (N_23919,N_23066,N_23368);
xor U23920 (N_23920,N_23174,N_23291);
nand U23921 (N_23921,N_23182,N_23400);
and U23922 (N_23922,N_23271,N_23112);
nand U23923 (N_23923,N_23293,N_23442);
or U23924 (N_23924,N_23063,N_23140);
and U23925 (N_23925,N_23233,N_23087);
and U23926 (N_23926,N_23212,N_23267);
nor U23927 (N_23927,N_23337,N_23471);
nor U23928 (N_23928,N_23226,N_23199);
nand U23929 (N_23929,N_23030,N_23116);
and U23930 (N_23930,N_23481,N_23199);
nand U23931 (N_23931,N_23309,N_23278);
nand U23932 (N_23932,N_23242,N_23299);
nand U23933 (N_23933,N_23088,N_23443);
and U23934 (N_23934,N_23466,N_23496);
and U23935 (N_23935,N_23005,N_23241);
nor U23936 (N_23936,N_23128,N_23244);
and U23937 (N_23937,N_23114,N_23454);
or U23938 (N_23938,N_23323,N_23259);
nor U23939 (N_23939,N_23471,N_23404);
and U23940 (N_23940,N_23080,N_23386);
nand U23941 (N_23941,N_23468,N_23442);
nand U23942 (N_23942,N_23472,N_23443);
nor U23943 (N_23943,N_23365,N_23258);
nor U23944 (N_23944,N_23477,N_23222);
nand U23945 (N_23945,N_23175,N_23327);
or U23946 (N_23946,N_23462,N_23120);
nand U23947 (N_23947,N_23243,N_23287);
xnor U23948 (N_23948,N_23419,N_23113);
or U23949 (N_23949,N_23410,N_23143);
or U23950 (N_23950,N_23466,N_23016);
nand U23951 (N_23951,N_23186,N_23250);
or U23952 (N_23952,N_23189,N_23466);
nand U23953 (N_23953,N_23271,N_23134);
xor U23954 (N_23954,N_23256,N_23052);
nor U23955 (N_23955,N_23239,N_23186);
and U23956 (N_23956,N_23007,N_23336);
nand U23957 (N_23957,N_23293,N_23250);
nand U23958 (N_23958,N_23011,N_23367);
or U23959 (N_23959,N_23260,N_23047);
nand U23960 (N_23960,N_23416,N_23187);
and U23961 (N_23961,N_23361,N_23269);
nor U23962 (N_23962,N_23056,N_23126);
and U23963 (N_23963,N_23021,N_23437);
and U23964 (N_23964,N_23411,N_23465);
nor U23965 (N_23965,N_23462,N_23023);
and U23966 (N_23966,N_23399,N_23112);
nand U23967 (N_23967,N_23262,N_23463);
nor U23968 (N_23968,N_23201,N_23084);
nand U23969 (N_23969,N_23407,N_23496);
nand U23970 (N_23970,N_23168,N_23284);
nor U23971 (N_23971,N_23316,N_23460);
or U23972 (N_23972,N_23438,N_23214);
nor U23973 (N_23973,N_23303,N_23173);
nand U23974 (N_23974,N_23150,N_23037);
nor U23975 (N_23975,N_23232,N_23097);
or U23976 (N_23976,N_23057,N_23002);
nor U23977 (N_23977,N_23241,N_23302);
or U23978 (N_23978,N_23000,N_23464);
nor U23979 (N_23979,N_23135,N_23143);
nor U23980 (N_23980,N_23308,N_23309);
nand U23981 (N_23981,N_23186,N_23075);
and U23982 (N_23982,N_23060,N_23495);
or U23983 (N_23983,N_23345,N_23061);
or U23984 (N_23984,N_23018,N_23461);
nand U23985 (N_23985,N_23295,N_23389);
nor U23986 (N_23986,N_23192,N_23478);
or U23987 (N_23987,N_23353,N_23109);
nor U23988 (N_23988,N_23287,N_23253);
nor U23989 (N_23989,N_23397,N_23226);
or U23990 (N_23990,N_23389,N_23034);
or U23991 (N_23991,N_23285,N_23293);
nor U23992 (N_23992,N_23339,N_23330);
and U23993 (N_23993,N_23406,N_23204);
or U23994 (N_23994,N_23229,N_23065);
nand U23995 (N_23995,N_23402,N_23358);
nor U23996 (N_23996,N_23067,N_23211);
nand U23997 (N_23997,N_23332,N_23477);
and U23998 (N_23998,N_23250,N_23221);
nand U23999 (N_23999,N_23305,N_23064);
nor U24000 (N_24000,N_23602,N_23826);
nand U24001 (N_24001,N_23627,N_23673);
and U24002 (N_24002,N_23896,N_23667);
and U24003 (N_24003,N_23914,N_23768);
and U24004 (N_24004,N_23735,N_23721);
or U24005 (N_24005,N_23871,N_23639);
or U24006 (N_24006,N_23900,N_23614);
or U24007 (N_24007,N_23712,N_23903);
nor U24008 (N_24008,N_23518,N_23911);
and U24009 (N_24009,N_23631,N_23628);
or U24010 (N_24010,N_23671,N_23526);
nand U24011 (N_24011,N_23745,N_23985);
or U24012 (N_24012,N_23953,N_23623);
or U24013 (N_24013,N_23574,N_23634);
nand U24014 (N_24014,N_23845,N_23674);
nor U24015 (N_24015,N_23687,N_23913);
nand U24016 (N_24016,N_23704,N_23509);
or U24017 (N_24017,N_23626,N_23517);
nand U24018 (N_24018,N_23766,N_23759);
or U24019 (N_24019,N_23647,N_23936);
nand U24020 (N_24020,N_23863,N_23693);
or U24021 (N_24021,N_23764,N_23829);
or U24022 (N_24022,N_23749,N_23927);
or U24023 (N_24023,N_23703,N_23686);
nor U24024 (N_24024,N_23941,N_23655);
and U24025 (N_24025,N_23575,N_23661);
nand U24026 (N_24026,N_23524,N_23831);
nor U24027 (N_24027,N_23677,N_23969);
nand U24028 (N_24028,N_23888,N_23530);
nor U24029 (N_24029,N_23798,N_23547);
nor U24030 (N_24030,N_23837,N_23538);
nand U24031 (N_24031,N_23828,N_23699);
and U24032 (N_24032,N_23591,N_23556);
or U24033 (N_24033,N_23757,N_23736);
and U24034 (N_24034,N_23756,N_23600);
nand U24035 (N_24035,N_23902,N_23934);
nand U24036 (N_24036,N_23581,N_23572);
nand U24037 (N_24037,N_23617,N_23907);
nand U24038 (N_24038,N_23646,N_23862);
and U24039 (N_24039,N_23859,N_23599);
nor U24040 (N_24040,N_23963,N_23680);
nor U24041 (N_24041,N_23928,N_23970);
nor U24042 (N_24042,N_23809,N_23536);
nand U24043 (N_24043,N_23887,N_23942);
nand U24044 (N_24044,N_23998,N_23806);
and U24045 (N_24045,N_23834,N_23531);
and U24046 (N_24046,N_23874,N_23937);
or U24047 (N_24047,N_23550,N_23854);
nand U24048 (N_24048,N_23660,N_23702);
nor U24049 (N_24049,N_23891,N_23760);
or U24050 (N_24050,N_23720,N_23573);
and U24051 (N_24051,N_23543,N_23785);
and U24052 (N_24052,N_23709,N_23788);
nand U24053 (N_24053,N_23868,N_23551);
nand U24054 (N_24054,N_23801,N_23804);
or U24055 (N_24055,N_23636,N_23761);
nand U24056 (N_24056,N_23666,N_23719);
nand U24057 (N_24057,N_23637,N_23935);
or U24058 (N_24058,N_23598,N_23765);
nand U24059 (N_24059,N_23877,N_23504);
nor U24060 (N_24060,N_23762,N_23521);
nand U24061 (N_24061,N_23644,N_23813);
nand U24062 (N_24062,N_23869,N_23919);
nor U24063 (N_24063,N_23925,N_23522);
or U24064 (N_24064,N_23682,N_23571);
and U24065 (N_24065,N_23511,N_23713);
nor U24066 (N_24066,N_23563,N_23872);
xnor U24067 (N_24067,N_23830,N_23974);
or U24068 (N_24068,N_23558,N_23858);
nand U24069 (N_24069,N_23643,N_23613);
and U24070 (N_24070,N_23947,N_23839);
nor U24071 (N_24071,N_23747,N_23725);
or U24072 (N_24072,N_23577,N_23595);
and U24073 (N_24073,N_23640,N_23554);
or U24074 (N_24074,N_23909,N_23821);
or U24075 (N_24075,N_23840,N_23786);
nor U24076 (N_24076,N_23885,N_23586);
or U24077 (N_24077,N_23933,N_23773);
nor U24078 (N_24078,N_23593,N_23729);
and U24079 (N_24079,N_23592,N_23990);
nand U24080 (N_24080,N_23908,N_23691);
nor U24081 (N_24081,N_23606,N_23544);
or U24082 (N_24082,N_23578,N_23734);
nor U24083 (N_24083,N_23717,N_23791);
nor U24084 (N_24084,N_23622,N_23695);
and U24085 (N_24085,N_23815,N_23846);
or U24086 (N_24086,N_23780,N_23929);
and U24087 (N_24087,N_23860,N_23658);
nand U24088 (N_24088,N_23923,N_23535);
and U24089 (N_24089,N_23672,N_23523);
nor U24090 (N_24090,N_23799,N_23857);
or U24091 (N_24091,N_23515,N_23650);
or U24092 (N_24092,N_23656,N_23901);
xnor U24093 (N_24093,N_23549,N_23904);
and U24094 (N_24094,N_23657,N_23777);
nor U24095 (N_24095,N_23552,N_23968);
or U24096 (N_24096,N_23880,N_23890);
or U24097 (N_24097,N_23979,N_23948);
and U24098 (N_24098,N_23999,N_23564);
or U24099 (N_24099,N_23983,N_23769);
nor U24100 (N_24100,N_23584,N_23800);
or U24101 (N_24101,N_23632,N_23678);
nand U24102 (N_24102,N_23906,N_23668);
and U24103 (N_24103,N_23988,N_23844);
nor U24104 (N_24104,N_23641,N_23692);
and U24105 (N_24105,N_23866,N_23938);
nor U24106 (N_24106,N_23607,N_23560);
and U24107 (N_24107,N_23881,N_23783);
nand U24108 (N_24108,N_23710,N_23957);
xnor U24109 (N_24109,N_23951,N_23533);
nor U24110 (N_24110,N_23565,N_23782);
or U24111 (N_24111,N_23542,N_23812);
and U24112 (N_24112,N_23618,N_23705);
nor U24113 (N_24113,N_23994,N_23807);
nor U24114 (N_24114,N_23555,N_23779);
and U24115 (N_24115,N_23642,N_23527);
nand U24116 (N_24116,N_23916,N_23730);
nand U24117 (N_24117,N_23976,N_23816);
nand U24118 (N_24118,N_23700,N_23774);
or U24119 (N_24119,N_23784,N_23898);
or U24120 (N_24120,N_23507,N_23696);
or U24121 (N_24121,N_23895,N_23981);
nand U24122 (N_24122,N_23582,N_23852);
nor U24123 (N_24123,N_23993,N_23975);
or U24124 (N_24124,N_23763,N_23824);
nor U24125 (N_24125,N_23711,N_23621);
nor U24126 (N_24126,N_23733,N_23758);
nor U24127 (N_24127,N_23503,N_23810);
nor U24128 (N_24128,N_23741,N_23893);
or U24129 (N_24129,N_23648,N_23659);
or U24130 (N_24130,N_23865,N_23723);
and U24131 (N_24131,N_23594,N_23748);
and U24132 (N_24132,N_23679,N_23792);
nor U24133 (N_24133,N_23688,N_23817);
nand U24134 (N_24134,N_23850,N_23662);
or U24135 (N_24135,N_23588,N_23752);
or U24136 (N_24136,N_23669,N_23513);
or U24137 (N_24137,N_23931,N_23620);
and U24138 (N_24138,N_23864,N_23922);
and U24139 (N_24139,N_23960,N_23570);
nand U24140 (N_24140,N_23825,N_23567);
xnor U24141 (N_24141,N_23612,N_23924);
nand U24142 (N_24142,N_23851,N_23728);
and U24143 (N_24143,N_23961,N_23778);
xor U24144 (N_24144,N_23568,N_23794);
or U24145 (N_24145,N_23566,N_23849);
nor U24146 (N_24146,N_23502,N_23601);
or U24147 (N_24147,N_23793,N_23892);
nand U24148 (N_24148,N_23967,N_23982);
nor U24149 (N_24149,N_23616,N_23579);
nor U24150 (N_24150,N_23950,N_23795);
and U24151 (N_24151,N_23973,N_23589);
and U24152 (N_24152,N_23675,N_23528);
nand U24153 (N_24153,N_23753,N_23683);
nor U24154 (N_24154,N_23625,N_23603);
or U24155 (N_24155,N_23585,N_23915);
nand U24156 (N_24156,N_23819,N_23894);
nor U24157 (N_24157,N_23516,N_23797);
or U24158 (N_24158,N_23539,N_23501);
and U24159 (N_24159,N_23645,N_23611);
nor U24160 (N_24160,N_23532,N_23520);
or U24161 (N_24161,N_23724,N_23912);
nor U24162 (N_24162,N_23548,N_23883);
or U24163 (N_24163,N_23989,N_23980);
nor U24164 (N_24164,N_23789,N_23510);
and U24165 (N_24165,N_23944,N_23583);
nand U24166 (N_24166,N_23553,N_23559);
nor U24167 (N_24167,N_23820,N_23867);
nand U24168 (N_24168,N_23776,N_23932);
nand U24169 (N_24169,N_23619,N_23802);
nor U24170 (N_24170,N_23708,N_23580);
nand U24171 (N_24171,N_23525,N_23746);
nand U24172 (N_24172,N_23590,N_23847);
or U24173 (N_24173,N_23707,N_23805);
nor U24174 (N_24174,N_23905,N_23882);
and U24175 (N_24175,N_23995,N_23855);
nand U24176 (N_24176,N_23978,N_23838);
and U24177 (N_24177,N_23561,N_23926);
nand U24178 (N_24178,N_23664,N_23609);
or U24179 (N_24179,N_23884,N_23832);
nand U24180 (N_24180,N_23715,N_23822);
nor U24181 (N_24181,N_23727,N_23731);
nor U24182 (N_24182,N_23596,N_23889);
nand U24183 (N_24183,N_23615,N_23737);
and U24184 (N_24184,N_23545,N_23843);
nor U24185 (N_24185,N_23971,N_23635);
or U24186 (N_24186,N_23959,N_23608);
nor U24187 (N_24187,N_23861,N_23952);
nand U24188 (N_24188,N_23918,N_23835);
nand U24189 (N_24189,N_23811,N_23716);
nand U24190 (N_24190,N_23755,N_23964);
or U24191 (N_24191,N_23949,N_23630);
nor U24192 (N_24192,N_23886,N_23649);
nand U24193 (N_24193,N_23958,N_23651);
and U24194 (N_24194,N_23722,N_23638);
or U24195 (N_24195,N_23701,N_23943);
nor U24196 (N_24196,N_23917,N_23920);
and U24197 (N_24197,N_23663,N_23508);
nor U24198 (N_24198,N_23576,N_23781);
and U24199 (N_24199,N_23853,N_23939);
and U24200 (N_24200,N_23505,N_23875);
nor U24201 (N_24201,N_23754,N_23827);
nor U24202 (N_24202,N_23541,N_23836);
nor U24203 (N_24203,N_23899,N_23787);
nand U24204 (N_24204,N_23624,N_23685);
and U24205 (N_24205,N_23738,N_23997);
and U24206 (N_24206,N_23940,N_23587);
and U24207 (N_24207,N_23681,N_23966);
nand U24208 (N_24208,N_23629,N_23945);
nor U24209 (N_24209,N_23767,N_23742);
xnor U24210 (N_24210,N_23954,N_23546);
and U24211 (N_24211,N_23714,N_23808);
or U24212 (N_24212,N_23910,N_23654);
nor U24213 (N_24213,N_23814,N_23823);
nand U24214 (N_24214,N_23876,N_23604);
xor U24215 (N_24215,N_23514,N_23506);
and U24216 (N_24216,N_23842,N_23751);
nor U24217 (N_24217,N_23698,N_23684);
nand U24218 (N_24218,N_23740,N_23965);
and U24219 (N_24219,N_23534,N_23856);
nand U24220 (N_24220,N_23605,N_23739);
and U24221 (N_24221,N_23987,N_23743);
nand U24222 (N_24222,N_23977,N_23803);
and U24223 (N_24223,N_23930,N_23512);
and U24224 (N_24224,N_23956,N_23770);
or U24225 (N_24225,N_23706,N_23848);
and U24226 (N_24226,N_23921,N_23972);
nor U24227 (N_24227,N_23992,N_23796);
nand U24228 (N_24228,N_23962,N_23726);
nor U24229 (N_24229,N_23744,N_23519);
xnor U24230 (N_24230,N_23653,N_23897);
or U24231 (N_24231,N_23878,N_23772);
and U24232 (N_24232,N_23557,N_23690);
or U24233 (N_24233,N_23597,N_23500);
nor U24234 (N_24234,N_23529,N_23562);
nor U24235 (N_24235,N_23841,N_23955);
xor U24236 (N_24236,N_23873,N_23689);
nor U24237 (N_24237,N_23610,N_23652);
or U24238 (N_24238,N_23870,N_23718);
nor U24239 (N_24239,N_23569,N_23991);
nand U24240 (N_24240,N_23984,N_23833);
or U24241 (N_24241,N_23771,N_23537);
or U24242 (N_24242,N_23676,N_23732);
and U24243 (N_24243,N_23818,N_23670);
or U24244 (N_24244,N_23996,N_23775);
nand U24245 (N_24245,N_23879,N_23750);
or U24246 (N_24246,N_23694,N_23790);
nand U24247 (N_24247,N_23697,N_23986);
or U24248 (N_24248,N_23633,N_23540);
nor U24249 (N_24249,N_23665,N_23946);
nor U24250 (N_24250,N_23650,N_23839);
nand U24251 (N_24251,N_23844,N_23766);
or U24252 (N_24252,N_23543,N_23964);
and U24253 (N_24253,N_23740,N_23511);
nand U24254 (N_24254,N_23955,N_23770);
and U24255 (N_24255,N_23915,N_23608);
or U24256 (N_24256,N_23583,N_23907);
nand U24257 (N_24257,N_23974,N_23576);
or U24258 (N_24258,N_23902,N_23662);
and U24259 (N_24259,N_23937,N_23694);
nand U24260 (N_24260,N_23521,N_23608);
nand U24261 (N_24261,N_23542,N_23885);
and U24262 (N_24262,N_23819,N_23672);
and U24263 (N_24263,N_23649,N_23830);
and U24264 (N_24264,N_23712,N_23650);
and U24265 (N_24265,N_23832,N_23726);
xor U24266 (N_24266,N_23768,N_23968);
nor U24267 (N_24267,N_23595,N_23862);
or U24268 (N_24268,N_23584,N_23764);
nand U24269 (N_24269,N_23656,N_23728);
nand U24270 (N_24270,N_23808,N_23969);
nand U24271 (N_24271,N_23855,N_23709);
nand U24272 (N_24272,N_23905,N_23984);
nand U24273 (N_24273,N_23684,N_23843);
or U24274 (N_24274,N_23833,N_23847);
nor U24275 (N_24275,N_23674,N_23614);
and U24276 (N_24276,N_23505,N_23723);
and U24277 (N_24277,N_23760,N_23644);
or U24278 (N_24278,N_23743,N_23733);
nor U24279 (N_24279,N_23797,N_23699);
nand U24280 (N_24280,N_23524,N_23813);
or U24281 (N_24281,N_23917,N_23580);
xnor U24282 (N_24282,N_23550,N_23536);
nand U24283 (N_24283,N_23668,N_23642);
nand U24284 (N_24284,N_23630,N_23925);
or U24285 (N_24285,N_23685,N_23759);
nand U24286 (N_24286,N_23837,N_23537);
or U24287 (N_24287,N_23570,N_23732);
or U24288 (N_24288,N_23594,N_23981);
or U24289 (N_24289,N_23908,N_23984);
nand U24290 (N_24290,N_23507,N_23551);
or U24291 (N_24291,N_23612,N_23555);
or U24292 (N_24292,N_23948,N_23823);
and U24293 (N_24293,N_23864,N_23896);
or U24294 (N_24294,N_23821,N_23617);
and U24295 (N_24295,N_23707,N_23886);
and U24296 (N_24296,N_23749,N_23551);
and U24297 (N_24297,N_23795,N_23995);
and U24298 (N_24298,N_23736,N_23949);
and U24299 (N_24299,N_23976,N_23993);
nor U24300 (N_24300,N_23647,N_23721);
nor U24301 (N_24301,N_23889,N_23543);
nor U24302 (N_24302,N_23595,N_23791);
xnor U24303 (N_24303,N_23552,N_23681);
nor U24304 (N_24304,N_23730,N_23786);
nor U24305 (N_24305,N_23545,N_23965);
nand U24306 (N_24306,N_23797,N_23850);
or U24307 (N_24307,N_23990,N_23930);
nand U24308 (N_24308,N_23569,N_23555);
nor U24309 (N_24309,N_23938,N_23730);
nand U24310 (N_24310,N_23850,N_23949);
or U24311 (N_24311,N_23633,N_23707);
or U24312 (N_24312,N_23929,N_23893);
nor U24313 (N_24313,N_23924,N_23792);
nand U24314 (N_24314,N_23589,N_23825);
and U24315 (N_24315,N_23976,N_23920);
or U24316 (N_24316,N_23679,N_23540);
nor U24317 (N_24317,N_23685,N_23533);
nor U24318 (N_24318,N_23535,N_23534);
or U24319 (N_24319,N_23629,N_23695);
or U24320 (N_24320,N_23587,N_23827);
or U24321 (N_24321,N_23723,N_23645);
nor U24322 (N_24322,N_23648,N_23884);
or U24323 (N_24323,N_23954,N_23814);
nor U24324 (N_24324,N_23894,N_23601);
and U24325 (N_24325,N_23943,N_23637);
or U24326 (N_24326,N_23733,N_23814);
nor U24327 (N_24327,N_23874,N_23686);
or U24328 (N_24328,N_23714,N_23811);
and U24329 (N_24329,N_23573,N_23515);
nor U24330 (N_24330,N_23718,N_23519);
nor U24331 (N_24331,N_23897,N_23786);
and U24332 (N_24332,N_23889,N_23660);
nor U24333 (N_24333,N_23965,N_23672);
nand U24334 (N_24334,N_23695,N_23780);
and U24335 (N_24335,N_23724,N_23627);
nor U24336 (N_24336,N_23964,N_23967);
and U24337 (N_24337,N_23706,N_23698);
nor U24338 (N_24338,N_23941,N_23598);
or U24339 (N_24339,N_23526,N_23777);
or U24340 (N_24340,N_23567,N_23723);
nand U24341 (N_24341,N_23810,N_23935);
nor U24342 (N_24342,N_23628,N_23734);
nor U24343 (N_24343,N_23742,N_23932);
or U24344 (N_24344,N_23917,N_23517);
or U24345 (N_24345,N_23530,N_23861);
nor U24346 (N_24346,N_23983,N_23976);
or U24347 (N_24347,N_23843,N_23681);
or U24348 (N_24348,N_23712,N_23911);
nor U24349 (N_24349,N_23734,N_23651);
nand U24350 (N_24350,N_23545,N_23562);
and U24351 (N_24351,N_23988,N_23691);
and U24352 (N_24352,N_23837,N_23687);
and U24353 (N_24353,N_23760,N_23590);
nand U24354 (N_24354,N_23645,N_23789);
or U24355 (N_24355,N_23955,N_23934);
nand U24356 (N_24356,N_23761,N_23983);
nor U24357 (N_24357,N_23564,N_23739);
nand U24358 (N_24358,N_23578,N_23577);
and U24359 (N_24359,N_23940,N_23905);
xnor U24360 (N_24360,N_23805,N_23827);
nand U24361 (N_24361,N_23807,N_23674);
and U24362 (N_24362,N_23973,N_23595);
or U24363 (N_24363,N_23779,N_23537);
nor U24364 (N_24364,N_23526,N_23507);
or U24365 (N_24365,N_23606,N_23581);
and U24366 (N_24366,N_23659,N_23762);
nand U24367 (N_24367,N_23710,N_23788);
nor U24368 (N_24368,N_23746,N_23959);
xor U24369 (N_24369,N_23529,N_23655);
nor U24370 (N_24370,N_23986,N_23629);
nor U24371 (N_24371,N_23948,N_23949);
xor U24372 (N_24372,N_23556,N_23906);
or U24373 (N_24373,N_23916,N_23975);
nor U24374 (N_24374,N_23843,N_23677);
and U24375 (N_24375,N_23763,N_23954);
or U24376 (N_24376,N_23886,N_23686);
nand U24377 (N_24377,N_23891,N_23716);
or U24378 (N_24378,N_23975,N_23502);
or U24379 (N_24379,N_23520,N_23717);
and U24380 (N_24380,N_23669,N_23633);
nand U24381 (N_24381,N_23611,N_23661);
and U24382 (N_24382,N_23708,N_23570);
nand U24383 (N_24383,N_23998,N_23667);
nand U24384 (N_24384,N_23724,N_23915);
nand U24385 (N_24385,N_23866,N_23927);
and U24386 (N_24386,N_23794,N_23944);
and U24387 (N_24387,N_23655,N_23956);
nand U24388 (N_24388,N_23946,N_23628);
and U24389 (N_24389,N_23836,N_23902);
nor U24390 (N_24390,N_23820,N_23845);
nor U24391 (N_24391,N_23511,N_23558);
or U24392 (N_24392,N_23757,N_23713);
and U24393 (N_24393,N_23684,N_23658);
nand U24394 (N_24394,N_23617,N_23832);
nand U24395 (N_24395,N_23606,N_23914);
or U24396 (N_24396,N_23966,N_23888);
nor U24397 (N_24397,N_23764,N_23681);
nor U24398 (N_24398,N_23614,N_23719);
or U24399 (N_24399,N_23834,N_23912);
nor U24400 (N_24400,N_23852,N_23682);
or U24401 (N_24401,N_23849,N_23538);
or U24402 (N_24402,N_23582,N_23527);
or U24403 (N_24403,N_23808,N_23598);
nor U24404 (N_24404,N_23962,N_23838);
and U24405 (N_24405,N_23998,N_23960);
and U24406 (N_24406,N_23647,N_23545);
nand U24407 (N_24407,N_23930,N_23878);
nor U24408 (N_24408,N_23788,N_23643);
or U24409 (N_24409,N_23762,N_23574);
xor U24410 (N_24410,N_23824,N_23885);
nor U24411 (N_24411,N_23754,N_23562);
or U24412 (N_24412,N_23745,N_23955);
nand U24413 (N_24413,N_23723,N_23695);
or U24414 (N_24414,N_23899,N_23924);
or U24415 (N_24415,N_23823,N_23749);
nand U24416 (N_24416,N_23760,N_23985);
or U24417 (N_24417,N_23846,N_23530);
and U24418 (N_24418,N_23598,N_23811);
and U24419 (N_24419,N_23857,N_23655);
nand U24420 (N_24420,N_23913,N_23659);
and U24421 (N_24421,N_23537,N_23745);
or U24422 (N_24422,N_23628,N_23792);
and U24423 (N_24423,N_23982,N_23708);
nand U24424 (N_24424,N_23525,N_23950);
and U24425 (N_24425,N_23937,N_23738);
or U24426 (N_24426,N_23971,N_23861);
and U24427 (N_24427,N_23810,N_23870);
or U24428 (N_24428,N_23512,N_23924);
nand U24429 (N_24429,N_23692,N_23576);
nand U24430 (N_24430,N_23691,N_23540);
and U24431 (N_24431,N_23708,N_23807);
nand U24432 (N_24432,N_23668,N_23863);
and U24433 (N_24433,N_23751,N_23726);
nor U24434 (N_24434,N_23518,N_23548);
and U24435 (N_24435,N_23579,N_23676);
nor U24436 (N_24436,N_23938,N_23869);
nor U24437 (N_24437,N_23770,N_23682);
or U24438 (N_24438,N_23927,N_23579);
nor U24439 (N_24439,N_23529,N_23975);
or U24440 (N_24440,N_23522,N_23515);
nor U24441 (N_24441,N_23612,N_23967);
or U24442 (N_24442,N_23867,N_23978);
or U24443 (N_24443,N_23527,N_23672);
or U24444 (N_24444,N_23869,N_23911);
and U24445 (N_24445,N_23708,N_23646);
and U24446 (N_24446,N_23722,N_23813);
nor U24447 (N_24447,N_23925,N_23512);
or U24448 (N_24448,N_23961,N_23618);
nor U24449 (N_24449,N_23998,N_23678);
nand U24450 (N_24450,N_23765,N_23586);
and U24451 (N_24451,N_23817,N_23756);
nand U24452 (N_24452,N_23577,N_23894);
nor U24453 (N_24453,N_23657,N_23941);
and U24454 (N_24454,N_23783,N_23599);
nand U24455 (N_24455,N_23999,N_23507);
nor U24456 (N_24456,N_23739,N_23789);
nor U24457 (N_24457,N_23807,N_23860);
and U24458 (N_24458,N_23985,N_23843);
nor U24459 (N_24459,N_23736,N_23734);
nand U24460 (N_24460,N_23582,N_23719);
and U24461 (N_24461,N_23954,N_23865);
or U24462 (N_24462,N_23811,N_23699);
nor U24463 (N_24463,N_23568,N_23516);
or U24464 (N_24464,N_23727,N_23635);
and U24465 (N_24465,N_23960,N_23984);
nor U24466 (N_24466,N_23838,N_23732);
and U24467 (N_24467,N_23630,N_23640);
nand U24468 (N_24468,N_23682,N_23561);
nand U24469 (N_24469,N_23566,N_23819);
nand U24470 (N_24470,N_23686,N_23631);
nor U24471 (N_24471,N_23546,N_23718);
or U24472 (N_24472,N_23883,N_23968);
or U24473 (N_24473,N_23673,N_23993);
nor U24474 (N_24474,N_23649,N_23710);
and U24475 (N_24475,N_23602,N_23909);
nor U24476 (N_24476,N_23812,N_23562);
and U24477 (N_24477,N_23741,N_23573);
and U24478 (N_24478,N_23819,N_23791);
and U24479 (N_24479,N_23962,N_23749);
or U24480 (N_24480,N_23792,N_23980);
or U24481 (N_24481,N_23854,N_23742);
nor U24482 (N_24482,N_23518,N_23641);
and U24483 (N_24483,N_23581,N_23840);
nor U24484 (N_24484,N_23814,N_23660);
nand U24485 (N_24485,N_23531,N_23921);
and U24486 (N_24486,N_23531,N_23591);
nor U24487 (N_24487,N_23562,N_23811);
nor U24488 (N_24488,N_23786,N_23520);
nor U24489 (N_24489,N_23909,N_23708);
nand U24490 (N_24490,N_23769,N_23806);
or U24491 (N_24491,N_23767,N_23529);
or U24492 (N_24492,N_23817,N_23617);
nand U24493 (N_24493,N_23944,N_23588);
and U24494 (N_24494,N_23873,N_23708);
or U24495 (N_24495,N_23989,N_23960);
or U24496 (N_24496,N_23673,N_23867);
and U24497 (N_24497,N_23647,N_23856);
or U24498 (N_24498,N_23864,N_23925);
or U24499 (N_24499,N_23871,N_23710);
and U24500 (N_24500,N_24034,N_24076);
and U24501 (N_24501,N_24455,N_24144);
nand U24502 (N_24502,N_24122,N_24003);
nand U24503 (N_24503,N_24305,N_24470);
nor U24504 (N_24504,N_24150,N_24341);
or U24505 (N_24505,N_24307,N_24242);
nand U24506 (N_24506,N_24327,N_24213);
nor U24507 (N_24507,N_24033,N_24132);
nand U24508 (N_24508,N_24488,N_24202);
nor U24509 (N_24509,N_24416,N_24088);
and U24510 (N_24510,N_24343,N_24494);
nor U24511 (N_24511,N_24192,N_24393);
and U24512 (N_24512,N_24115,N_24475);
nor U24513 (N_24513,N_24171,N_24431);
or U24514 (N_24514,N_24415,N_24174);
nor U24515 (N_24515,N_24352,N_24075);
nor U24516 (N_24516,N_24160,N_24430);
or U24517 (N_24517,N_24273,N_24138);
xor U24518 (N_24518,N_24404,N_24186);
and U24519 (N_24519,N_24070,N_24308);
nor U24520 (N_24520,N_24460,N_24120);
or U24521 (N_24521,N_24275,N_24451);
nor U24522 (N_24522,N_24492,N_24162);
and U24523 (N_24523,N_24255,N_24353);
nor U24524 (N_24524,N_24148,N_24423);
or U24525 (N_24525,N_24454,N_24293);
or U24526 (N_24526,N_24356,N_24177);
nor U24527 (N_24527,N_24153,N_24019);
and U24528 (N_24528,N_24263,N_24024);
nor U24529 (N_24529,N_24229,N_24128);
nor U24530 (N_24530,N_24463,N_24068);
nand U24531 (N_24531,N_24052,N_24355);
nor U24532 (N_24532,N_24438,N_24061);
or U24533 (N_24533,N_24173,N_24237);
nor U24534 (N_24534,N_24127,N_24303);
and U24535 (N_24535,N_24238,N_24010);
and U24536 (N_24536,N_24047,N_24483);
and U24537 (N_24537,N_24106,N_24367);
or U24538 (N_24538,N_24007,N_24105);
nor U24539 (N_24539,N_24103,N_24471);
or U24540 (N_24540,N_24429,N_24169);
nand U24541 (N_24541,N_24296,N_24259);
xnor U24542 (N_24542,N_24087,N_24370);
or U24543 (N_24543,N_24118,N_24388);
and U24544 (N_24544,N_24385,N_24006);
nor U24545 (N_24545,N_24252,N_24264);
or U24546 (N_24546,N_24421,N_24476);
nor U24547 (N_24547,N_24321,N_24448);
nor U24548 (N_24548,N_24486,N_24278);
nor U24549 (N_24549,N_24383,N_24403);
or U24550 (N_24550,N_24204,N_24466);
nand U24551 (N_24551,N_24225,N_24465);
and U24552 (N_24552,N_24210,N_24413);
nand U24553 (N_24553,N_24155,N_24247);
nor U24554 (N_24554,N_24348,N_24437);
xor U24555 (N_24555,N_24073,N_24357);
nor U24556 (N_24556,N_24094,N_24479);
nor U24557 (N_24557,N_24095,N_24468);
nor U24558 (N_24558,N_24239,N_24085);
nor U24559 (N_24559,N_24497,N_24331);
nand U24560 (N_24560,N_24060,N_24482);
nor U24561 (N_24561,N_24198,N_24317);
and U24562 (N_24562,N_24057,N_24224);
and U24563 (N_24563,N_24441,N_24013);
or U24564 (N_24564,N_24285,N_24271);
nand U24565 (N_24565,N_24270,N_24178);
and U24566 (N_24566,N_24435,N_24261);
nand U24567 (N_24567,N_24372,N_24071);
or U24568 (N_24568,N_24334,N_24008);
nand U24569 (N_24569,N_24077,N_24040);
nand U24570 (N_24570,N_24063,N_24102);
or U24571 (N_24571,N_24265,N_24333);
xnor U24572 (N_24572,N_24112,N_24350);
and U24573 (N_24573,N_24297,N_24434);
or U24574 (N_24574,N_24228,N_24473);
nand U24575 (N_24575,N_24236,N_24302);
and U24576 (N_24576,N_24039,N_24119);
or U24577 (N_24577,N_24351,N_24014);
or U24578 (N_24578,N_24396,N_24280);
nand U24579 (N_24579,N_24272,N_24397);
and U24580 (N_24580,N_24424,N_24044);
or U24581 (N_24581,N_24243,N_24191);
nand U24582 (N_24582,N_24180,N_24098);
and U24583 (N_24583,N_24484,N_24257);
nor U24584 (N_24584,N_24166,N_24041);
nor U24585 (N_24585,N_24433,N_24309);
or U24586 (N_24586,N_24377,N_24245);
and U24587 (N_24587,N_24306,N_24189);
nor U24588 (N_24588,N_24391,N_24046);
or U24589 (N_24589,N_24190,N_24485);
nor U24590 (N_24590,N_24235,N_24375);
or U24591 (N_24591,N_24336,N_24124);
or U24592 (N_24592,N_24004,N_24140);
nand U24593 (N_24593,N_24250,N_24017);
or U24594 (N_24594,N_24290,N_24200);
and U24595 (N_24595,N_24029,N_24478);
or U24596 (N_24596,N_24090,N_24097);
and U24597 (N_24597,N_24364,N_24053);
nor U24598 (N_24598,N_24496,N_24420);
nand U24599 (N_24599,N_24168,N_24137);
nand U24600 (N_24600,N_24117,N_24025);
and U24601 (N_24601,N_24481,N_24414);
and U24602 (N_24602,N_24172,N_24092);
nor U24603 (N_24603,N_24146,N_24023);
nor U24604 (N_24604,N_24498,N_24165);
nor U24605 (N_24605,N_24042,N_24163);
nand U24606 (N_24606,N_24027,N_24459);
and U24607 (N_24607,N_24330,N_24050);
nor U24608 (N_24608,N_24176,N_24221);
nor U24609 (N_24609,N_24069,N_24011);
nand U24610 (N_24610,N_24326,N_24319);
nand U24611 (N_24611,N_24386,N_24442);
nand U24612 (N_24612,N_24474,N_24449);
and U24613 (N_24613,N_24452,N_24142);
nand U24614 (N_24614,N_24426,N_24337);
and U24615 (N_24615,N_24267,N_24164);
and U24616 (N_24616,N_24232,N_24215);
nor U24617 (N_24617,N_24458,N_24456);
xor U24618 (N_24618,N_24226,N_24318);
or U24619 (N_24619,N_24446,N_24408);
or U24620 (N_24620,N_24086,N_24187);
or U24621 (N_24621,N_24009,N_24159);
nor U24622 (N_24622,N_24109,N_24358);
nand U24623 (N_24623,N_24406,N_24480);
and U24624 (N_24624,N_24051,N_24453);
nor U24625 (N_24625,N_24443,N_24398);
nor U24626 (N_24626,N_24447,N_24314);
or U24627 (N_24627,N_24123,N_24182);
nand U24628 (N_24628,N_24373,N_24412);
and U24629 (N_24629,N_24419,N_24002);
or U24630 (N_24630,N_24129,N_24108);
or U24631 (N_24631,N_24049,N_24199);
nand U24632 (N_24632,N_24493,N_24323);
or U24633 (N_24633,N_24101,N_24445);
nand U24634 (N_24634,N_24130,N_24329);
or U24635 (N_24635,N_24405,N_24012);
nand U24636 (N_24636,N_24205,N_24266);
nor U24637 (N_24637,N_24036,N_24400);
nor U24638 (N_24638,N_24249,N_24444);
nor U24639 (N_24639,N_24432,N_24145);
or U24640 (N_24640,N_24183,N_24325);
or U24641 (N_24641,N_24167,N_24499);
and U24642 (N_24642,N_24407,N_24080);
and U24643 (N_24643,N_24234,N_24489);
nor U24644 (N_24644,N_24354,N_24207);
nor U24645 (N_24645,N_24346,N_24395);
or U24646 (N_24646,N_24113,N_24490);
nor U24647 (N_24647,N_24378,N_24147);
nand U24648 (N_24648,N_24399,N_24201);
nand U24649 (N_24649,N_24316,N_24371);
and U24650 (N_24650,N_24360,N_24276);
nand U24651 (N_24651,N_24313,N_24181);
or U24652 (N_24652,N_24427,N_24298);
nand U24653 (N_24653,N_24462,N_24216);
xor U24654 (N_24654,N_24366,N_24384);
nor U24655 (N_24655,N_24469,N_24170);
or U24656 (N_24656,N_24335,N_24206);
or U24657 (N_24657,N_24365,N_24072);
or U24658 (N_24658,N_24096,N_24032);
nand U24659 (N_24659,N_24258,N_24197);
and U24660 (N_24660,N_24212,N_24328);
or U24661 (N_24661,N_24422,N_24038);
and U24662 (N_24662,N_24196,N_24126);
nand U24663 (N_24663,N_24211,N_24300);
nor U24664 (N_24664,N_24035,N_24078);
nor U24665 (N_24665,N_24043,N_24031);
or U24666 (N_24666,N_24136,N_24209);
nand U24667 (N_24667,N_24055,N_24253);
and U24668 (N_24668,N_24368,N_24288);
nor U24669 (N_24669,N_24230,N_24054);
or U24670 (N_24670,N_24287,N_24062);
and U24671 (N_24671,N_24390,N_24310);
nor U24672 (N_24672,N_24295,N_24436);
or U24673 (N_24673,N_24067,N_24157);
nor U24674 (N_24674,N_24428,N_24125);
and U24675 (N_24675,N_24079,N_24376);
nand U24676 (N_24676,N_24477,N_24457);
nand U24677 (N_24677,N_24135,N_24081);
or U24678 (N_24678,N_24282,N_24141);
and U24679 (N_24679,N_24440,N_24450);
or U24680 (N_24680,N_24299,N_24217);
xnor U24681 (N_24681,N_24220,N_24185);
nand U24682 (N_24682,N_24254,N_24099);
nand U24683 (N_24683,N_24277,N_24315);
and U24684 (N_24684,N_24131,N_24417);
nor U24685 (N_24685,N_24401,N_24248);
and U24686 (N_24686,N_24089,N_24340);
and U24687 (N_24687,N_24048,N_24411);
nand U24688 (N_24688,N_24016,N_24304);
nand U24689 (N_24689,N_24005,N_24015);
nor U24690 (N_24690,N_24139,N_24495);
and U24691 (N_24691,N_24219,N_24322);
nor U24692 (N_24692,N_24161,N_24241);
and U24693 (N_24693,N_24110,N_24188);
and U24694 (N_24694,N_24262,N_24208);
nor U24695 (N_24695,N_24114,N_24392);
nor U24696 (N_24696,N_24214,N_24065);
nand U24697 (N_24697,N_24093,N_24320);
nand U24698 (N_24698,N_24233,N_24175);
and U24699 (N_24699,N_24133,N_24107);
and U24700 (N_24700,N_24342,N_24149);
and U24701 (N_24701,N_24256,N_24195);
nor U24702 (N_24702,N_24301,N_24154);
nor U24703 (N_24703,N_24037,N_24410);
and U24704 (N_24704,N_24179,N_24020);
nor U24705 (N_24705,N_24382,N_24283);
or U24706 (N_24706,N_24425,N_24134);
nor U24707 (N_24707,N_24152,N_24379);
or U24708 (N_24708,N_24461,N_24058);
nor U24709 (N_24709,N_24289,N_24418);
nand U24710 (N_24710,N_24292,N_24363);
and U24711 (N_24711,N_24374,N_24156);
nand U24712 (N_24712,N_24018,N_24472);
and U24713 (N_24713,N_24231,N_24359);
nand U24714 (N_24714,N_24116,N_24194);
and U24715 (N_24715,N_24269,N_24028);
nor U24716 (N_24716,N_24193,N_24022);
nand U24717 (N_24717,N_24332,N_24362);
and U24718 (N_24718,N_24361,N_24240);
nand U24719 (N_24719,N_24074,N_24151);
or U24720 (N_24720,N_24246,N_24203);
and U24721 (N_24721,N_24000,N_24222);
or U24722 (N_24722,N_24030,N_24311);
and U24723 (N_24723,N_24338,N_24344);
nor U24724 (N_24724,N_24439,N_24100);
or U24725 (N_24725,N_24026,N_24082);
and U24726 (N_24726,N_24059,N_24227);
or U24727 (N_24727,N_24158,N_24111);
and U24728 (N_24728,N_24464,N_24066);
nand U24729 (N_24729,N_24244,N_24218);
and U24730 (N_24730,N_24084,N_24387);
and U24731 (N_24731,N_24021,N_24381);
nand U24732 (N_24732,N_24487,N_24324);
nor U24733 (N_24733,N_24001,N_24260);
nor U24734 (N_24734,N_24345,N_24121);
nand U24735 (N_24735,N_24251,N_24312);
nor U24736 (N_24736,N_24223,N_24064);
and U24737 (N_24737,N_24286,N_24291);
nand U24738 (N_24738,N_24409,N_24268);
nor U24739 (N_24739,N_24104,N_24394);
nand U24740 (N_24740,N_24339,N_24091);
and U24741 (N_24741,N_24402,N_24184);
nor U24742 (N_24742,N_24380,N_24279);
nand U24743 (N_24743,N_24143,N_24274);
or U24744 (N_24744,N_24349,N_24083);
nand U24745 (N_24745,N_24389,N_24369);
nor U24746 (N_24746,N_24281,N_24491);
or U24747 (N_24747,N_24056,N_24284);
nand U24748 (N_24748,N_24347,N_24045);
and U24749 (N_24749,N_24294,N_24467);
and U24750 (N_24750,N_24317,N_24334);
nand U24751 (N_24751,N_24394,N_24156);
nand U24752 (N_24752,N_24113,N_24425);
nand U24753 (N_24753,N_24193,N_24004);
or U24754 (N_24754,N_24176,N_24435);
or U24755 (N_24755,N_24413,N_24199);
or U24756 (N_24756,N_24187,N_24278);
nor U24757 (N_24757,N_24021,N_24468);
nand U24758 (N_24758,N_24054,N_24370);
nand U24759 (N_24759,N_24314,N_24421);
and U24760 (N_24760,N_24011,N_24482);
or U24761 (N_24761,N_24126,N_24118);
and U24762 (N_24762,N_24357,N_24306);
and U24763 (N_24763,N_24491,N_24477);
and U24764 (N_24764,N_24333,N_24017);
and U24765 (N_24765,N_24316,N_24383);
nand U24766 (N_24766,N_24314,N_24038);
and U24767 (N_24767,N_24388,N_24407);
or U24768 (N_24768,N_24246,N_24250);
nand U24769 (N_24769,N_24260,N_24451);
nor U24770 (N_24770,N_24213,N_24136);
or U24771 (N_24771,N_24184,N_24112);
nor U24772 (N_24772,N_24114,N_24249);
or U24773 (N_24773,N_24159,N_24129);
or U24774 (N_24774,N_24123,N_24487);
nor U24775 (N_24775,N_24155,N_24488);
or U24776 (N_24776,N_24245,N_24439);
or U24777 (N_24777,N_24198,N_24158);
nor U24778 (N_24778,N_24241,N_24404);
nor U24779 (N_24779,N_24041,N_24338);
or U24780 (N_24780,N_24432,N_24320);
or U24781 (N_24781,N_24074,N_24315);
nand U24782 (N_24782,N_24485,N_24423);
nor U24783 (N_24783,N_24461,N_24128);
or U24784 (N_24784,N_24435,N_24420);
nand U24785 (N_24785,N_24024,N_24181);
nand U24786 (N_24786,N_24415,N_24051);
or U24787 (N_24787,N_24013,N_24050);
and U24788 (N_24788,N_24422,N_24387);
and U24789 (N_24789,N_24364,N_24159);
and U24790 (N_24790,N_24497,N_24490);
nand U24791 (N_24791,N_24037,N_24383);
and U24792 (N_24792,N_24056,N_24383);
nand U24793 (N_24793,N_24334,N_24381);
nand U24794 (N_24794,N_24300,N_24397);
and U24795 (N_24795,N_24493,N_24425);
nor U24796 (N_24796,N_24029,N_24250);
or U24797 (N_24797,N_24147,N_24197);
and U24798 (N_24798,N_24329,N_24322);
nand U24799 (N_24799,N_24310,N_24088);
nor U24800 (N_24800,N_24230,N_24486);
or U24801 (N_24801,N_24078,N_24137);
and U24802 (N_24802,N_24310,N_24452);
and U24803 (N_24803,N_24370,N_24234);
and U24804 (N_24804,N_24005,N_24498);
nor U24805 (N_24805,N_24414,N_24064);
or U24806 (N_24806,N_24051,N_24039);
or U24807 (N_24807,N_24165,N_24195);
or U24808 (N_24808,N_24316,N_24244);
nor U24809 (N_24809,N_24159,N_24392);
and U24810 (N_24810,N_24281,N_24440);
and U24811 (N_24811,N_24188,N_24377);
and U24812 (N_24812,N_24117,N_24014);
or U24813 (N_24813,N_24153,N_24211);
and U24814 (N_24814,N_24459,N_24204);
or U24815 (N_24815,N_24252,N_24026);
nand U24816 (N_24816,N_24494,N_24469);
nand U24817 (N_24817,N_24060,N_24046);
nand U24818 (N_24818,N_24253,N_24002);
and U24819 (N_24819,N_24372,N_24201);
nor U24820 (N_24820,N_24316,N_24320);
and U24821 (N_24821,N_24110,N_24139);
nor U24822 (N_24822,N_24014,N_24126);
xnor U24823 (N_24823,N_24482,N_24371);
or U24824 (N_24824,N_24481,N_24108);
and U24825 (N_24825,N_24284,N_24459);
nand U24826 (N_24826,N_24383,N_24412);
or U24827 (N_24827,N_24463,N_24387);
nand U24828 (N_24828,N_24012,N_24416);
nor U24829 (N_24829,N_24248,N_24396);
nand U24830 (N_24830,N_24410,N_24360);
and U24831 (N_24831,N_24367,N_24400);
nand U24832 (N_24832,N_24282,N_24460);
and U24833 (N_24833,N_24169,N_24351);
or U24834 (N_24834,N_24169,N_24037);
nor U24835 (N_24835,N_24171,N_24474);
and U24836 (N_24836,N_24385,N_24041);
nor U24837 (N_24837,N_24142,N_24145);
nand U24838 (N_24838,N_24159,N_24311);
nor U24839 (N_24839,N_24351,N_24440);
and U24840 (N_24840,N_24200,N_24199);
nor U24841 (N_24841,N_24387,N_24313);
nand U24842 (N_24842,N_24026,N_24000);
or U24843 (N_24843,N_24039,N_24288);
and U24844 (N_24844,N_24107,N_24101);
nand U24845 (N_24845,N_24331,N_24414);
and U24846 (N_24846,N_24011,N_24351);
or U24847 (N_24847,N_24464,N_24263);
nor U24848 (N_24848,N_24432,N_24465);
and U24849 (N_24849,N_24134,N_24088);
or U24850 (N_24850,N_24165,N_24392);
nand U24851 (N_24851,N_24128,N_24426);
and U24852 (N_24852,N_24457,N_24078);
or U24853 (N_24853,N_24443,N_24274);
nor U24854 (N_24854,N_24055,N_24206);
nand U24855 (N_24855,N_24035,N_24042);
and U24856 (N_24856,N_24074,N_24405);
or U24857 (N_24857,N_24491,N_24159);
nor U24858 (N_24858,N_24310,N_24143);
nor U24859 (N_24859,N_24117,N_24345);
and U24860 (N_24860,N_24451,N_24174);
or U24861 (N_24861,N_24050,N_24207);
or U24862 (N_24862,N_24205,N_24268);
nor U24863 (N_24863,N_24372,N_24466);
nand U24864 (N_24864,N_24072,N_24246);
and U24865 (N_24865,N_24448,N_24020);
or U24866 (N_24866,N_24279,N_24033);
and U24867 (N_24867,N_24097,N_24107);
or U24868 (N_24868,N_24208,N_24153);
or U24869 (N_24869,N_24252,N_24393);
or U24870 (N_24870,N_24150,N_24489);
nor U24871 (N_24871,N_24367,N_24489);
and U24872 (N_24872,N_24394,N_24307);
and U24873 (N_24873,N_24117,N_24334);
or U24874 (N_24874,N_24174,N_24180);
and U24875 (N_24875,N_24124,N_24430);
or U24876 (N_24876,N_24047,N_24388);
and U24877 (N_24877,N_24308,N_24010);
nand U24878 (N_24878,N_24133,N_24367);
nor U24879 (N_24879,N_24000,N_24051);
and U24880 (N_24880,N_24182,N_24460);
and U24881 (N_24881,N_24241,N_24395);
or U24882 (N_24882,N_24398,N_24342);
nand U24883 (N_24883,N_24243,N_24164);
and U24884 (N_24884,N_24389,N_24446);
and U24885 (N_24885,N_24162,N_24343);
and U24886 (N_24886,N_24135,N_24420);
or U24887 (N_24887,N_24286,N_24130);
nand U24888 (N_24888,N_24096,N_24199);
nor U24889 (N_24889,N_24000,N_24329);
xor U24890 (N_24890,N_24140,N_24183);
nand U24891 (N_24891,N_24493,N_24278);
or U24892 (N_24892,N_24225,N_24384);
or U24893 (N_24893,N_24232,N_24025);
and U24894 (N_24894,N_24361,N_24185);
nor U24895 (N_24895,N_24356,N_24400);
nand U24896 (N_24896,N_24324,N_24222);
nand U24897 (N_24897,N_24081,N_24317);
nor U24898 (N_24898,N_24069,N_24099);
and U24899 (N_24899,N_24123,N_24013);
nor U24900 (N_24900,N_24325,N_24003);
nor U24901 (N_24901,N_24210,N_24105);
xnor U24902 (N_24902,N_24023,N_24402);
nand U24903 (N_24903,N_24156,N_24160);
and U24904 (N_24904,N_24181,N_24266);
nand U24905 (N_24905,N_24093,N_24230);
nand U24906 (N_24906,N_24033,N_24203);
nand U24907 (N_24907,N_24112,N_24093);
nor U24908 (N_24908,N_24156,N_24215);
or U24909 (N_24909,N_24077,N_24422);
and U24910 (N_24910,N_24404,N_24461);
or U24911 (N_24911,N_24445,N_24292);
or U24912 (N_24912,N_24214,N_24361);
nand U24913 (N_24913,N_24319,N_24386);
or U24914 (N_24914,N_24461,N_24436);
and U24915 (N_24915,N_24230,N_24265);
nor U24916 (N_24916,N_24273,N_24407);
and U24917 (N_24917,N_24299,N_24019);
nand U24918 (N_24918,N_24084,N_24407);
xor U24919 (N_24919,N_24195,N_24242);
or U24920 (N_24920,N_24129,N_24474);
nand U24921 (N_24921,N_24268,N_24273);
and U24922 (N_24922,N_24181,N_24162);
or U24923 (N_24923,N_24175,N_24196);
nand U24924 (N_24924,N_24084,N_24456);
or U24925 (N_24925,N_24113,N_24106);
nand U24926 (N_24926,N_24469,N_24267);
or U24927 (N_24927,N_24265,N_24070);
and U24928 (N_24928,N_24247,N_24216);
or U24929 (N_24929,N_24126,N_24069);
or U24930 (N_24930,N_24497,N_24244);
nand U24931 (N_24931,N_24003,N_24225);
xnor U24932 (N_24932,N_24428,N_24456);
or U24933 (N_24933,N_24166,N_24401);
or U24934 (N_24934,N_24087,N_24052);
or U24935 (N_24935,N_24236,N_24463);
nor U24936 (N_24936,N_24195,N_24331);
nor U24937 (N_24937,N_24270,N_24076);
nor U24938 (N_24938,N_24430,N_24306);
and U24939 (N_24939,N_24210,N_24494);
or U24940 (N_24940,N_24190,N_24243);
nand U24941 (N_24941,N_24039,N_24456);
nand U24942 (N_24942,N_24074,N_24456);
nor U24943 (N_24943,N_24025,N_24113);
and U24944 (N_24944,N_24230,N_24212);
nor U24945 (N_24945,N_24148,N_24386);
nand U24946 (N_24946,N_24446,N_24047);
nand U24947 (N_24947,N_24186,N_24104);
or U24948 (N_24948,N_24348,N_24325);
nand U24949 (N_24949,N_24468,N_24224);
and U24950 (N_24950,N_24150,N_24400);
nand U24951 (N_24951,N_24432,N_24365);
and U24952 (N_24952,N_24270,N_24454);
and U24953 (N_24953,N_24018,N_24471);
nand U24954 (N_24954,N_24426,N_24273);
and U24955 (N_24955,N_24017,N_24490);
and U24956 (N_24956,N_24301,N_24458);
nor U24957 (N_24957,N_24125,N_24030);
or U24958 (N_24958,N_24394,N_24433);
or U24959 (N_24959,N_24273,N_24035);
nor U24960 (N_24960,N_24245,N_24100);
or U24961 (N_24961,N_24379,N_24287);
nand U24962 (N_24962,N_24298,N_24112);
nand U24963 (N_24963,N_24274,N_24309);
or U24964 (N_24964,N_24133,N_24388);
and U24965 (N_24965,N_24431,N_24425);
and U24966 (N_24966,N_24485,N_24021);
nor U24967 (N_24967,N_24025,N_24204);
nand U24968 (N_24968,N_24190,N_24156);
nor U24969 (N_24969,N_24315,N_24127);
and U24970 (N_24970,N_24182,N_24424);
or U24971 (N_24971,N_24035,N_24151);
and U24972 (N_24972,N_24210,N_24244);
and U24973 (N_24973,N_24287,N_24110);
or U24974 (N_24974,N_24080,N_24076);
nand U24975 (N_24975,N_24104,N_24365);
nor U24976 (N_24976,N_24467,N_24130);
or U24977 (N_24977,N_24160,N_24322);
nor U24978 (N_24978,N_24006,N_24308);
nor U24979 (N_24979,N_24356,N_24302);
and U24980 (N_24980,N_24072,N_24061);
and U24981 (N_24981,N_24047,N_24216);
or U24982 (N_24982,N_24121,N_24487);
and U24983 (N_24983,N_24084,N_24154);
or U24984 (N_24984,N_24086,N_24028);
nor U24985 (N_24985,N_24194,N_24323);
nand U24986 (N_24986,N_24219,N_24477);
nand U24987 (N_24987,N_24113,N_24336);
and U24988 (N_24988,N_24223,N_24017);
and U24989 (N_24989,N_24178,N_24461);
and U24990 (N_24990,N_24266,N_24310);
nor U24991 (N_24991,N_24274,N_24313);
xor U24992 (N_24992,N_24161,N_24040);
nor U24993 (N_24993,N_24147,N_24388);
or U24994 (N_24994,N_24335,N_24312);
nor U24995 (N_24995,N_24323,N_24482);
nor U24996 (N_24996,N_24217,N_24430);
nor U24997 (N_24997,N_24028,N_24262);
or U24998 (N_24998,N_24363,N_24368);
or U24999 (N_24999,N_24377,N_24046);
and UO_0 (O_0,N_24639,N_24941);
and UO_1 (O_1,N_24661,N_24899);
and UO_2 (O_2,N_24576,N_24850);
nand UO_3 (O_3,N_24706,N_24811);
nor UO_4 (O_4,N_24780,N_24744);
nand UO_5 (O_5,N_24813,N_24632);
and UO_6 (O_6,N_24678,N_24845);
and UO_7 (O_7,N_24594,N_24664);
nor UO_8 (O_8,N_24865,N_24978);
nand UO_9 (O_9,N_24560,N_24863);
or UO_10 (O_10,N_24585,N_24812);
nand UO_11 (O_11,N_24539,N_24603);
or UO_12 (O_12,N_24665,N_24527);
and UO_13 (O_13,N_24663,N_24529);
or UO_14 (O_14,N_24534,N_24970);
nand UO_15 (O_15,N_24691,N_24769);
nor UO_16 (O_16,N_24823,N_24902);
nand UO_17 (O_17,N_24596,N_24655);
nand UO_18 (O_18,N_24828,N_24920);
xor UO_19 (O_19,N_24720,N_24541);
or UO_20 (O_20,N_24502,N_24825);
or UO_21 (O_21,N_24647,N_24916);
or UO_22 (O_22,N_24934,N_24972);
or UO_23 (O_23,N_24894,N_24606);
nor UO_24 (O_24,N_24855,N_24508);
or UO_25 (O_25,N_24656,N_24579);
and UO_26 (O_26,N_24710,N_24771);
and UO_27 (O_27,N_24993,N_24670);
nand UO_28 (O_28,N_24878,N_24806);
nor UO_29 (O_29,N_24905,N_24924);
and UO_30 (O_30,N_24518,N_24952);
or UO_31 (O_31,N_24948,N_24524);
nand UO_32 (O_32,N_24915,N_24753);
nor UO_33 (O_33,N_24563,N_24776);
xor UO_34 (O_34,N_24758,N_24757);
or UO_35 (O_35,N_24741,N_24740);
and UO_36 (O_36,N_24985,N_24748);
nand UO_37 (O_37,N_24767,N_24848);
or UO_38 (O_38,N_24736,N_24774);
nor UO_39 (O_39,N_24766,N_24835);
or UO_40 (O_40,N_24604,N_24669);
nand UO_41 (O_41,N_24797,N_24584);
and UO_42 (O_42,N_24913,N_24533);
nor UO_43 (O_43,N_24885,N_24673);
or UO_44 (O_44,N_24857,N_24788);
and UO_45 (O_45,N_24738,N_24933);
and UO_46 (O_46,N_24625,N_24799);
and UO_47 (O_47,N_24749,N_24872);
xor UO_48 (O_48,N_24544,N_24961);
and UO_49 (O_49,N_24900,N_24616);
and UO_50 (O_50,N_24944,N_24973);
or UO_51 (O_51,N_24681,N_24930);
and UO_52 (O_52,N_24809,N_24937);
nor UO_53 (O_53,N_24784,N_24590);
and UO_54 (O_54,N_24568,N_24836);
nor UO_55 (O_55,N_24965,N_24550);
nor UO_56 (O_56,N_24507,N_24969);
nand UO_57 (O_57,N_24931,N_24554);
and UO_58 (O_58,N_24573,N_24692);
nor UO_59 (O_59,N_24715,N_24860);
nand UO_60 (O_60,N_24653,N_24723);
or UO_61 (O_61,N_24868,N_24676);
or UO_62 (O_62,N_24503,N_24896);
and UO_63 (O_63,N_24789,N_24743);
nand UO_64 (O_64,N_24979,N_24994);
or UO_65 (O_65,N_24629,N_24892);
nor UO_66 (O_66,N_24650,N_24727);
and UO_67 (O_67,N_24525,N_24912);
and UO_68 (O_68,N_24824,N_24699);
and UO_69 (O_69,N_24830,N_24976);
nand UO_70 (O_70,N_24871,N_24515);
or UO_71 (O_71,N_24737,N_24947);
nor UO_72 (O_72,N_24612,N_24731);
nand UO_73 (O_73,N_24513,N_24595);
nand UO_74 (O_74,N_24646,N_24707);
or UO_75 (O_75,N_24999,N_24523);
xnor UO_76 (O_76,N_24802,N_24853);
and UO_77 (O_77,N_24735,N_24597);
nor UO_78 (O_78,N_24903,N_24538);
and UO_79 (O_79,N_24672,N_24684);
nor UO_80 (O_80,N_24582,N_24764);
and UO_81 (O_81,N_24713,N_24546);
nor UO_82 (O_82,N_24837,N_24621);
nand UO_83 (O_83,N_24732,N_24839);
or UO_84 (O_84,N_24578,N_24927);
and UO_85 (O_85,N_24514,N_24510);
and UO_86 (O_86,N_24781,N_24638);
or UO_87 (O_87,N_24609,N_24593);
and UO_88 (O_88,N_24718,N_24875);
and UO_89 (O_89,N_24570,N_24599);
nor UO_90 (O_90,N_24636,N_24858);
or UO_91 (O_91,N_24614,N_24779);
nor UO_92 (O_92,N_24635,N_24750);
or UO_93 (O_93,N_24964,N_24679);
nand UO_94 (O_94,N_24891,N_24730);
nor UO_95 (O_95,N_24719,N_24667);
and UO_96 (O_96,N_24698,N_24628);
and UO_97 (O_97,N_24959,N_24620);
and UO_98 (O_98,N_24690,N_24775);
nor UO_99 (O_99,N_24697,N_24591);
xor UO_100 (O_100,N_24721,N_24652);
and UO_101 (O_101,N_24637,N_24537);
nand UO_102 (O_102,N_24831,N_24856);
or UO_103 (O_103,N_24666,N_24880);
nor UO_104 (O_104,N_24752,N_24548);
xnor UO_105 (O_105,N_24911,N_24587);
nand UO_106 (O_106,N_24556,N_24904);
and UO_107 (O_107,N_24887,N_24986);
or UO_108 (O_108,N_24511,N_24791);
or UO_109 (O_109,N_24956,N_24765);
nand UO_110 (O_110,N_24704,N_24962);
nand UO_111 (O_111,N_24984,N_24685);
or UO_112 (O_112,N_24649,N_24996);
xor UO_113 (O_113,N_24818,N_24693);
and UO_114 (O_114,N_24569,N_24982);
nor UO_115 (O_115,N_24938,N_24861);
nand UO_116 (O_116,N_24795,N_24528);
xor UO_117 (O_117,N_24794,N_24711);
nand UO_118 (O_118,N_24722,N_24819);
nor UO_119 (O_119,N_24910,N_24501);
nand UO_120 (O_120,N_24867,N_24909);
or UO_121 (O_121,N_24581,N_24668);
or UO_122 (O_122,N_24605,N_24989);
and UO_123 (O_123,N_24561,N_24852);
and UO_124 (O_124,N_24883,N_24553);
or UO_125 (O_125,N_24772,N_24520);
nand UO_126 (O_126,N_24907,N_24709);
nor UO_127 (O_127,N_24662,N_24798);
and UO_128 (O_128,N_24928,N_24807);
or UO_129 (O_129,N_24506,N_24901);
or UO_130 (O_130,N_24869,N_24897);
or UO_131 (O_131,N_24747,N_24572);
and UO_132 (O_132,N_24943,N_24851);
or UO_133 (O_133,N_24549,N_24695);
nand UO_134 (O_134,N_24751,N_24888);
or UO_135 (O_135,N_24622,N_24542);
nand UO_136 (O_136,N_24843,N_24577);
or UO_137 (O_137,N_24882,N_24800);
nand UO_138 (O_138,N_24700,N_24574);
or UO_139 (O_139,N_24714,N_24516);
and UO_140 (O_140,N_24626,N_24786);
nand UO_141 (O_141,N_24796,N_24547);
nand UO_142 (O_142,N_24884,N_24602);
and UO_143 (O_143,N_24558,N_24566);
nand UO_144 (O_144,N_24827,N_24623);
or UO_145 (O_145,N_24583,N_24870);
nor UO_146 (O_146,N_24658,N_24589);
or UO_147 (O_147,N_24949,N_24675);
nor UO_148 (O_148,N_24618,N_24815);
nand UO_149 (O_149,N_24512,N_24531);
nor UO_150 (O_150,N_24821,N_24725);
nand UO_151 (O_151,N_24842,N_24696);
nand UO_152 (O_152,N_24500,N_24555);
and UO_153 (O_153,N_24768,N_24906);
nand UO_154 (O_154,N_24532,N_24671);
nor UO_155 (O_155,N_24761,N_24729);
nor UO_156 (O_156,N_24847,N_24785);
nand UO_157 (O_157,N_24833,N_24873);
and UO_158 (O_158,N_24925,N_24914);
or UO_159 (O_159,N_24565,N_24659);
and UO_160 (O_160,N_24688,N_24987);
nor UO_161 (O_161,N_24728,N_24567);
nor UO_162 (O_162,N_24686,N_24677);
and UO_163 (O_163,N_24945,N_24955);
nand UO_164 (O_164,N_24586,N_24619);
xnor UO_165 (O_165,N_24866,N_24966);
or UO_166 (O_166,N_24981,N_24881);
and UO_167 (O_167,N_24963,N_24936);
or UO_168 (O_168,N_24859,N_24998);
or UO_169 (O_169,N_24643,N_24535);
nor UO_170 (O_170,N_24759,N_24680);
nor UO_171 (O_171,N_24810,N_24645);
nand UO_172 (O_172,N_24983,N_24615);
nor UO_173 (O_173,N_24841,N_24804);
or UO_174 (O_174,N_24971,N_24642);
or UO_175 (O_175,N_24694,N_24726);
nor UO_176 (O_176,N_24958,N_24530);
or UO_177 (O_177,N_24814,N_24705);
and UO_178 (O_178,N_24564,N_24504);
and UO_179 (O_179,N_24517,N_24876);
and UO_180 (O_180,N_24702,N_24838);
nor UO_181 (O_181,N_24908,N_24820);
or UO_182 (O_182,N_24509,N_24886);
or UO_183 (O_183,N_24559,N_24588);
nor UO_184 (O_184,N_24742,N_24703);
and UO_185 (O_185,N_24874,N_24519);
nand UO_186 (O_186,N_24640,N_24522);
nand UO_187 (O_187,N_24600,N_24935);
nor UO_188 (O_188,N_24536,N_24792);
and UO_189 (O_189,N_24946,N_24557);
nor UO_190 (O_190,N_24968,N_24932);
and UO_191 (O_191,N_24763,N_24617);
or UO_192 (O_192,N_24951,N_24540);
nand UO_193 (O_193,N_24980,N_24808);
and UO_194 (O_194,N_24890,N_24601);
or UO_195 (O_195,N_24580,N_24954);
nand UO_196 (O_196,N_24803,N_24687);
nand UO_197 (O_197,N_24683,N_24790);
and UO_198 (O_198,N_24975,N_24816);
and UO_199 (O_199,N_24734,N_24648);
nor UO_200 (O_200,N_24716,N_24995);
nand UO_201 (O_201,N_24926,N_24846);
and UO_202 (O_202,N_24592,N_24849);
nand UO_203 (O_203,N_24657,N_24611);
or UO_204 (O_204,N_24641,N_24608);
nand UO_205 (O_205,N_24551,N_24754);
nor UO_206 (O_206,N_24817,N_24895);
nand UO_207 (O_207,N_24575,N_24942);
nor UO_208 (O_208,N_24893,N_24552);
xor UO_209 (O_209,N_24739,N_24950);
nor UO_210 (O_210,N_24562,N_24777);
or UO_211 (O_211,N_24701,N_24783);
nand UO_212 (O_212,N_24505,N_24967);
and UO_213 (O_213,N_24834,N_24929);
xnor UO_214 (O_214,N_24793,N_24898);
and UO_215 (O_215,N_24543,N_24613);
and UO_216 (O_216,N_24829,N_24630);
nand UO_217 (O_217,N_24918,N_24877);
and UO_218 (O_218,N_24939,N_24922);
nand UO_219 (O_219,N_24545,N_24660);
and UO_220 (O_220,N_24977,N_24762);
or UO_221 (O_221,N_24805,N_24988);
nor UO_222 (O_222,N_24974,N_24844);
xor UO_223 (O_223,N_24770,N_24755);
nor UO_224 (O_224,N_24627,N_24674);
and UO_225 (O_225,N_24746,N_24864);
or UO_226 (O_226,N_24862,N_24708);
and UO_227 (O_227,N_24745,N_24801);
nand UO_228 (O_228,N_24826,N_24526);
nor UO_229 (O_229,N_24610,N_24733);
or UO_230 (O_230,N_24953,N_24756);
nor UO_231 (O_231,N_24940,N_24689);
nor UO_232 (O_232,N_24923,N_24919);
and UO_233 (O_233,N_24957,N_24598);
nand UO_234 (O_234,N_24992,N_24854);
and UO_235 (O_235,N_24634,N_24879);
nand UO_236 (O_236,N_24921,N_24997);
nand UO_237 (O_237,N_24960,N_24521);
nand UO_238 (O_238,N_24631,N_24840);
nor UO_239 (O_239,N_24760,N_24787);
nor UO_240 (O_240,N_24991,N_24778);
nand UO_241 (O_241,N_24607,N_24990);
and UO_242 (O_242,N_24682,N_24782);
and UO_243 (O_243,N_24654,N_24624);
nor UO_244 (O_244,N_24651,N_24889);
xnor UO_245 (O_245,N_24633,N_24724);
and UO_246 (O_246,N_24712,N_24773);
and UO_247 (O_247,N_24917,N_24571);
nor UO_248 (O_248,N_24832,N_24717);
nand UO_249 (O_249,N_24822,N_24644);
nor UO_250 (O_250,N_24691,N_24540);
nand UO_251 (O_251,N_24728,N_24835);
nor UO_252 (O_252,N_24903,N_24672);
nor UO_253 (O_253,N_24698,N_24925);
or UO_254 (O_254,N_24806,N_24695);
and UO_255 (O_255,N_24561,N_24728);
and UO_256 (O_256,N_24694,N_24584);
nor UO_257 (O_257,N_24704,N_24854);
nand UO_258 (O_258,N_24905,N_24968);
or UO_259 (O_259,N_24962,N_24860);
nand UO_260 (O_260,N_24555,N_24714);
nor UO_261 (O_261,N_24887,N_24699);
or UO_262 (O_262,N_24630,N_24642);
or UO_263 (O_263,N_24638,N_24530);
and UO_264 (O_264,N_24686,N_24766);
and UO_265 (O_265,N_24893,N_24737);
nand UO_266 (O_266,N_24704,N_24769);
nand UO_267 (O_267,N_24811,N_24748);
nor UO_268 (O_268,N_24806,N_24665);
or UO_269 (O_269,N_24867,N_24619);
nand UO_270 (O_270,N_24633,N_24630);
and UO_271 (O_271,N_24573,N_24925);
or UO_272 (O_272,N_24960,N_24566);
nor UO_273 (O_273,N_24586,N_24686);
and UO_274 (O_274,N_24693,N_24788);
nor UO_275 (O_275,N_24682,N_24638);
and UO_276 (O_276,N_24679,N_24798);
and UO_277 (O_277,N_24508,N_24843);
nor UO_278 (O_278,N_24682,N_24967);
and UO_279 (O_279,N_24959,N_24702);
nor UO_280 (O_280,N_24614,N_24749);
nand UO_281 (O_281,N_24888,N_24873);
or UO_282 (O_282,N_24645,N_24823);
nor UO_283 (O_283,N_24804,N_24611);
and UO_284 (O_284,N_24949,N_24665);
or UO_285 (O_285,N_24761,N_24959);
nand UO_286 (O_286,N_24556,N_24861);
or UO_287 (O_287,N_24698,N_24854);
nor UO_288 (O_288,N_24584,N_24860);
and UO_289 (O_289,N_24545,N_24600);
nor UO_290 (O_290,N_24615,N_24668);
nor UO_291 (O_291,N_24683,N_24842);
nor UO_292 (O_292,N_24527,N_24587);
nand UO_293 (O_293,N_24621,N_24568);
nor UO_294 (O_294,N_24655,N_24809);
nor UO_295 (O_295,N_24957,N_24569);
or UO_296 (O_296,N_24930,N_24646);
or UO_297 (O_297,N_24760,N_24729);
and UO_298 (O_298,N_24787,N_24588);
or UO_299 (O_299,N_24681,N_24707);
nand UO_300 (O_300,N_24776,N_24614);
nor UO_301 (O_301,N_24792,N_24949);
and UO_302 (O_302,N_24890,N_24604);
and UO_303 (O_303,N_24644,N_24951);
or UO_304 (O_304,N_24845,N_24811);
nand UO_305 (O_305,N_24639,N_24677);
nor UO_306 (O_306,N_24932,N_24953);
nand UO_307 (O_307,N_24837,N_24873);
nor UO_308 (O_308,N_24756,N_24512);
nand UO_309 (O_309,N_24871,N_24521);
or UO_310 (O_310,N_24955,N_24565);
and UO_311 (O_311,N_24609,N_24527);
and UO_312 (O_312,N_24502,N_24756);
nor UO_313 (O_313,N_24518,N_24586);
nand UO_314 (O_314,N_24919,N_24757);
and UO_315 (O_315,N_24531,N_24836);
or UO_316 (O_316,N_24977,N_24549);
nand UO_317 (O_317,N_24971,N_24596);
nand UO_318 (O_318,N_24887,N_24984);
nor UO_319 (O_319,N_24514,N_24573);
nor UO_320 (O_320,N_24558,N_24761);
or UO_321 (O_321,N_24718,N_24844);
nand UO_322 (O_322,N_24799,N_24800);
nor UO_323 (O_323,N_24565,N_24779);
nor UO_324 (O_324,N_24845,N_24667);
or UO_325 (O_325,N_24525,N_24782);
and UO_326 (O_326,N_24771,N_24685);
and UO_327 (O_327,N_24866,N_24775);
nor UO_328 (O_328,N_24880,N_24803);
nand UO_329 (O_329,N_24746,N_24953);
xor UO_330 (O_330,N_24717,N_24570);
nand UO_331 (O_331,N_24938,N_24673);
nor UO_332 (O_332,N_24793,N_24665);
or UO_333 (O_333,N_24678,N_24706);
and UO_334 (O_334,N_24727,N_24975);
nand UO_335 (O_335,N_24890,N_24822);
nand UO_336 (O_336,N_24614,N_24546);
nand UO_337 (O_337,N_24838,N_24529);
xnor UO_338 (O_338,N_24793,N_24767);
and UO_339 (O_339,N_24827,N_24932);
nand UO_340 (O_340,N_24830,N_24805);
nand UO_341 (O_341,N_24933,N_24864);
xnor UO_342 (O_342,N_24606,N_24576);
or UO_343 (O_343,N_24815,N_24969);
nand UO_344 (O_344,N_24939,N_24797);
or UO_345 (O_345,N_24576,N_24814);
nor UO_346 (O_346,N_24532,N_24926);
or UO_347 (O_347,N_24938,N_24684);
nor UO_348 (O_348,N_24749,N_24744);
or UO_349 (O_349,N_24641,N_24639);
nor UO_350 (O_350,N_24809,N_24548);
nand UO_351 (O_351,N_24856,N_24605);
nand UO_352 (O_352,N_24707,N_24960);
and UO_353 (O_353,N_24829,N_24698);
or UO_354 (O_354,N_24796,N_24990);
and UO_355 (O_355,N_24606,N_24580);
nand UO_356 (O_356,N_24978,N_24670);
nor UO_357 (O_357,N_24519,N_24745);
nand UO_358 (O_358,N_24577,N_24694);
and UO_359 (O_359,N_24789,N_24864);
nor UO_360 (O_360,N_24565,N_24596);
and UO_361 (O_361,N_24968,N_24520);
and UO_362 (O_362,N_24675,N_24565);
or UO_363 (O_363,N_24957,N_24891);
or UO_364 (O_364,N_24591,N_24534);
or UO_365 (O_365,N_24564,N_24596);
nand UO_366 (O_366,N_24717,N_24658);
and UO_367 (O_367,N_24775,N_24559);
nand UO_368 (O_368,N_24671,N_24691);
nand UO_369 (O_369,N_24995,N_24684);
nor UO_370 (O_370,N_24564,N_24841);
or UO_371 (O_371,N_24604,N_24621);
xnor UO_372 (O_372,N_24682,N_24712);
nand UO_373 (O_373,N_24589,N_24978);
and UO_374 (O_374,N_24578,N_24651);
nor UO_375 (O_375,N_24969,N_24661);
nand UO_376 (O_376,N_24970,N_24869);
or UO_377 (O_377,N_24760,N_24579);
nand UO_378 (O_378,N_24886,N_24994);
nand UO_379 (O_379,N_24854,N_24840);
or UO_380 (O_380,N_24937,N_24995);
and UO_381 (O_381,N_24684,N_24993);
and UO_382 (O_382,N_24652,N_24638);
and UO_383 (O_383,N_24982,N_24577);
xnor UO_384 (O_384,N_24515,N_24606);
nand UO_385 (O_385,N_24821,N_24670);
and UO_386 (O_386,N_24930,N_24878);
nand UO_387 (O_387,N_24838,N_24709);
nand UO_388 (O_388,N_24564,N_24587);
nor UO_389 (O_389,N_24876,N_24973);
and UO_390 (O_390,N_24874,N_24574);
and UO_391 (O_391,N_24712,N_24968);
and UO_392 (O_392,N_24735,N_24659);
or UO_393 (O_393,N_24810,N_24942);
nand UO_394 (O_394,N_24598,N_24938);
nor UO_395 (O_395,N_24909,N_24966);
or UO_396 (O_396,N_24959,N_24974);
or UO_397 (O_397,N_24639,N_24891);
and UO_398 (O_398,N_24522,N_24502);
and UO_399 (O_399,N_24567,N_24526);
or UO_400 (O_400,N_24905,N_24854);
or UO_401 (O_401,N_24518,N_24993);
or UO_402 (O_402,N_24948,N_24687);
or UO_403 (O_403,N_24592,N_24574);
nand UO_404 (O_404,N_24524,N_24633);
nand UO_405 (O_405,N_24545,N_24523);
or UO_406 (O_406,N_24828,N_24710);
and UO_407 (O_407,N_24551,N_24830);
and UO_408 (O_408,N_24595,N_24565);
or UO_409 (O_409,N_24706,N_24968);
nor UO_410 (O_410,N_24618,N_24779);
nand UO_411 (O_411,N_24552,N_24667);
and UO_412 (O_412,N_24699,N_24752);
or UO_413 (O_413,N_24768,N_24738);
and UO_414 (O_414,N_24680,N_24832);
nand UO_415 (O_415,N_24510,N_24535);
nor UO_416 (O_416,N_24570,N_24665);
and UO_417 (O_417,N_24602,N_24890);
or UO_418 (O_418,N_24656,N_24756);
nand UO_419 (O_419,N_24844,N_24831);
nor UO_420 (O_420,N_24638,N_24754);
and UO_421 (O_421,N_24747,N_24675);
nand UO_422 (O_422,N_24654,N_24863);
or UO_423 (O_423,N_24566,N_24589);
and UO_424 (O_424,N_24561,N_24597);
nor UO_425 (O_425,N_24553,N_24955);
or UO_426 (O_426,N_24855,N_24787);
xnor UO_427 (O_427,N_24664,N_24515);
or UO_428 (O_428,N_24534,N_24985);
nand UO_429 (O_429,N_24894,N_24922);
or UO_430 (O_430,N_24932,N_24808);
nand UO_431 (O_431,N_24843,N_24854);
or UO_432 (O_432,N_24665,N_24759);
and UO_433 (O_433,N_24717,N_24579);
and UO_434 (O_434,N_24894,N_24975);
nor UO_435 (O_435,N_24708,N_24509);
or UO_436 (O_436,N_24920,N_24534);
and UO_437 (O_437,N_24679,N_24614);
nor UO_438 (O_438,N_24710,N_24885);
and UO_439 (O_439,N_24708,N_24641);
and UO_440 (O_440,N_24598,N_24567);
and UO_441 (O_441,N_24600,N_24523);
nand UO_442 (O_442,N_24549,N_24991);
nand UO_443 (O_443,N_24652,N_24935);
nand UO_444 (O_444,N_24669,N_24879);
nand UO_445 (O_445,N_24840,N_24536);
nor UO_446 (O_446,N_24984,N_24860);
or UO_447 (O_447,N_24854,N_24601);
or UO_448 (O_448,N_24681,N_24876);
nand UO_449 (O_449,N_24776,N_24882);
and UO_450 (O_450,N_24932,N_24798);
nor UO_451 (O_451,N_24838,N_24858);
or UO_452 (O_452,N_24894,N_24586);
and UO_453 (O_453,N_24849,N_24577);
nor UO_454 (O_454,N_24886,N_24750);
nand UO_455 (O_455,N_24633,N_24664);
nand UO_456 (O_456,N_24747,N_24512);
and UO_457 (O_457,N_24903,N_24604);
nand UO_458 (O_458,N_24558,N_24950);
and UO_459 (O_459,N_24597,N_24820);
and UO_460 (O_460,N_24724,N_24569);
or UO_461 (O_461,N_24614,N_24750);
and UO_462 (O_462,N_24729,N_24707);
xor UO_463 (O_463,N_24563,N_24887);
and UO_464 (O_464,N_24919,N_24783);
or UO_465 (O_465,N_24673,N_24700);
and UO_466 (O_466,N_24600,N_24993);
nand UO_467 (O_467,N_24790,N_24903);
nor UO_468 (O_468,N_24761,N_24933);
nand UO_469 (O_469,N_24750,N_24522);
nor UO_470 (O_470,N_24751,N_24740);
or UO_471 (O_471,N_24645,N_24875);
nor UO_472 (O_472,N_24851,N_24960);
nand UO_473 (O_473,N_24687,N_24515);
or UO_474 (O_474,N_24810,N_24641);
and UO_475 (O_475,N_24523,N_24743);
nor UO_476 (O_476,N_24644,N_24806);
xor UO_477 (O_477,N_24941,N_24850);
nand UO_478 (O_478,N_24650,N_24949);
or UO_479 (O_479,N_24878,N_24768);
and UO_480 (O_480,N_24536,N_24957);
nor UO_481 (O_481,N_24936,N_24779);
nand UO_482 (O_482,N_24555,N_24532);
nor UO_483 (O_483,N_24832,N_24877);
and UO_484 (O_484,N_24645,N_24766);
and UO_485 (O_485,N_24726,N_24538);
nor UO_486 (O_486,N_24720,N_24711);
nand UO_487 (O_487,N_24810,N_24998);
nor UO_488 (O_488,N_24776,N_24749);
nor UO_489 (O_489,N_24619,N_24898);
and UO_490 (O_490,N_24824,N_24818);
and UO_491 (O_491,N_24582,N_24817);
nand UO_492 (O_492,N_24560,N_24930);
or UO_493 (O_493,N_24695,N_24658);
nand UO_494 (O_494,N_24779,N_24822);
xor UO_495 (O_495,N_24803,N_24526);
and UO_496 (O_496,N_24588,N_24861);
and UO_497 (O_497,N_24577,N_24819);
or UO_498 (O_498,N_24736,N_24809);
or UO_499 (O_499,N_24665,N_24639);
nand UO_500 (O_500,N_24526,N_24534);
and UO_501 (O_501,N_24513,N_24900);
and UO_502 (O_502,N_24780,N_24666);
nor UO_503 (O_503,N_24673,N_24764);
or UO_504 (O_504,N_24827,N_24547);
and UO_505 (O_505,N_24612,N_24516);
nand UO_506 (O_506,N_24623,N_24961);
nand UO_507 (O_507,N_24516,N_24888);
and UO_508 (O_508,N_24860,N_24847);
or UO_509 (O_509,N_24978,N_24931);
nand UO_510 (O_510,N_24823,N_24810);
nand UO_511 (O_511,N_24783,N_24538);
nand UO_512 (O_512,N_24683,N_24512);
nand UO_513 (O_513,N_24529,N_24856);
and UO_514 (O_514,N_24855,N_24780);
or UO_515 (O_515,N_24863,N_24504);
or UO_516 (O_516,N_24905,N_24565);
nor UO_517 (O_517,N_24617,N_24967);
and UO_518 (O_518,N_24924,N_24925);
nor UO_519 (O_519,N_24703,N_24787);
nor UO_520 (O_520,N_24620,N_24517);
or UO_521 (O_521,N_24979,N_24592);
nand UO_522 (O_522,N_24559,N_24792);
nor UO_523 (O_523,N_24826,N_24938);
nor UO_524 (O_524,N_24967,N_24975);
and UO_525 (O_525,N_24513,N_24956);
xor UO_526 (O_526,N_24762,N_24982);
and UO_527 (O_527,N_24509,N_24855);
nand UO_528 (O_528,N_24656,N_24503);
nor UO_529 (O_529,N_24639,N_24834);
and UO_530 (O_530,N_24740,N_24924);
nor UO_531 (O_531,N_24802,N_24993);
and UO_532 (O_532,N_24514,N_24689);
and UO_533 (O_533,N_24915,N_24884);
nand UO_534 (O_534,N_24621,N_24505);
and UO_535 (O_535,N_24999,N_24818);
nand UO_536 (O_536,N_24526,N_24703);
nor UO_537 (O_537,N_24853,N_24690);
or UO_538 (O_538,N_24907,N_24578);
nand UO_539 (O_539,N_24856,N_24645);
nand UO_540 (O_540,N_24591,N_24663);
and UO_541 (O_541,N_24698,N_24852);
nor UO_542 (O_542,N_24807,N_24677);
xnor UO_543 (O_543,N_24751,N_24959);
and UO_544 (O_544,N_24844,N_24841);
and UO_545 (O_545,N_24981,N_24994);
or UO_546 (O_546,N_24533,N_24928);
nand UO_547 (O_547,N_24807,N_24714);
nand UO_548 (O_548,N_24823,N_24957);
and UO_549 (O_549,N_24944,N_24873);
and UO_550 (O_550,N_24669,N_24863);
or UO_551 (O_551,N_24641,N_24764);
and UO_552 (O_552,N_24703,N_24894);
nor UO_553 (O_553,N_24620,N_24809);
and UO_554 (O_554,N_24682,N_24736);
nand UO_555 (O_555,N_24659,N_24644);
and UO_556 (O_556,N_24953,N_24794);
nor UO_557 (O_557,N_24770,N_24704);
nand UO_558 (O_558,N_24665,N_24733);
and UO_559 (O_559,N_24581,N_24721);
and UO_560 (O_560,N_24736,N_24561);
xnor UO_561 (O_561,N_24992,N_24526);
nor UO_562 (O_562,N_24707,N_24755);
nand UO_563 (O_563,N_24699,N_24971);
nand UO_564 (O_564,N_24733,N_24644);
or UO_565 (O_565,N_24901,N_24691);
or UO_566 (O_566,N_24831,N_24757);
and UO_567 (O_567,N_24547,N_24667);
nor UO_568 (O_568,N_24606,N_24523);
nor UO_569 (O_569,N_24746,N_24564);
or UO_570 (O_570,N_24523,N_24929);
nor UO_571 (O_571,N_24786,N_24956);
and UO_572 (O_572,N_24503,N_24618);
nand UO_573 (O_573,N_24946,N_24980);
or UO_574 (O_574,N_24970,N_24991);
nor UO_575 (O_575,N_24998,N_24754);
nand UO_576 (O_576,N_24645,N_24881);
and UO_577 (O_577,N_24582,N_24948);
nor UO_578 (O_578,N_24672,N_24731);
or UO_579 (O_579,N_24810,N_24931);
or UO_580 (O_580,N_24662,N_24818);
or UO_581 (O_581,N_24932,N_24673);
nor UO_582 (O_582,N_24746,N_24974);
or UO_583 (O_583,N_24886,N_24583);
nor UO_584 (O_584,N_24657,N_24616);
nand UO_585 (O_585,N_24509,N_24640);
and UO_586 (O_586,N_24614,N_24838);
nand UO_587 (O_587,N_24911,N_24823);
nor UO_588 (O_588,N_24817,N_24803);
nor UO_589 (O_589,N_24816,N_24518);
and UO_590 (O_590,N_24680,N_24730);
or UO_591 (O_591,N_24634,N_24657);
nand UO_592 (O_592,N_24903,N_24876);
nor UO_593 (O_593,N_24734,N_24777);
or UO_594 (O_594,N_24524,N_24506);
nand UO_595 (O_595,N_24728,N_24815);
nor UO_596 (O_596,N_24503,N_24668);
nand UO_597 (O_597,N_24754,N_24927);
and UO_598 (O_598,N_24765,N_24879);
xnor UO_599 (O_599,N_24857,N_24827);
nor UO_600 (O_600,N_24574,N_24798);
or UO_601 (O_601,N_24934,N_24864);
or UO_602 (O_602,N_24821,N_24956);
and UO_603 (O_603,N_24608,N_24903);
nor UO_604 (O_604,N_24691,N_24660);
or UO_605 (O_605,N_24828,N_24815);
xnor UO_606 (O_606,N_24762,N_24684);
nor UO_607 (O_607,N_24915,N_24744);
or UO_608 (O_608,N_24817,N_24833);
nor UO_609 (O_609,N_24600,N_24750);
and UO_610 (O_610,N_24752,N_24879);
nor UO_611 (O_611,N_24909,N_24802);
nor UO_612 (O_612,N_24626,N_24952);
xor UO_613 (O_613,N_24668,N_24689);
nand UO_614 (O_614,N_24979,N_24580);
and UO_615 (O_615,N_24867,N_24826);
or UO_616 (O_616,N_24795,N_24853);
nor UO_617 (O_617,N_24634,N_24503);
nand UO_618 (O_618,N_24773,N_24909);
and UO_619 (O_619,N_24600,N_24977);
nor UO_620 (O_620,N_24665,N_24621);
and UO_621 (O_621,N_24795,N_24559);
or UO_622 (O_622,N_24633,N_24831);
and UO_623 (O_623,N_24647,N_24638);
nand UO_624 (O_624,N_24981,N_24887);
and UO_625 (O_625,N_24894,N_24882);
nor UO_626 (O_626,N_24583,N_24758);
nor UO_627 (O_627,N_24905,N_24986);
nor UO_628 (O_628,N_24924,N_24522);
nor UO_629 (O_629,N_24764,N_24856);
and UO_630 (O_630,N_24660,N_24700);
nor UO_631 (O_631,N_24668,N_24561);
nand UO_632 (O_632,N_24587,N_24608);
and UO_633 (O_633,N_24700,N_24565);
and UO_634 (O_634,N_24532,N_24596);
nor UO_635 (O_635,N_24970,N_24585);
and UO_636 (O_636,N_24516,N_24611);
or UO_637 (O_637,N_24968,N_24975);
nor UO_638 (O_638,N_24587,N_24960);
and UO_639 (O_639,N_24542,N_24982);
and UO_640 (O_640,N_24579,N_24775);
and UO_641 (O_641,N_24557,N_24539);
nand UO_642 (O_642,N_24528,N_24972);
nor UO_643 (O_643,N_24623,N_24851);
or UO_644 (O_644,N_24967,N_24981);
or UO_645 (O_645,N_24913,N_24664);
nand UO_646 (O_646,N_24682,N_24985);
nor UO_647 (O_647,N_24917,N_24516);
and UO_648 (O_648,N_24981,N_24612);
nand UO_649 (O_649,N_24635,N_24975);
nor UO_650 (O_650,N_24874,N_24662);
nand UO_651 (O_651,N_24556,N_24575);
or UO_652 (O_652,N_24841,N_24629);
or UO_653 (O_653,N_24624,N_24532);
or UO_654 (O_654,N_24638,N_24833);
and UO_655 (O_655,N_24684,N_24749);
nor UO_656 (O_656,N_24612,N_24569);
nor UO_657 (O_657,N_24988,N_24886);
and UO_658 (O_658,N_24714,N_24901);
and UO_659 (O_659,N_24984,N_24795);
nand UO_660 (O_660,N_24742,N_24862);
nor UO_661 (O_661,N_24556,N_24996);
or UO_662 (O_662,N_24538,N_24682);
nor UO_663 (O_663,N_24881,N_24736);
nor UO_664 (O_664,N_24539,N_24660);
and UO_665 (O_665,N_24572,N_24540);
nor UO_666 (O_666,N_24536,N_24889);
nand UO_667 (O_667,N_24634,N_24932);
nor UO_668 (O_668,N_24953,N_24951);
nor UO_669 (O_669,N_24796,N_24804);
nor UO_670 (O_670,N_24943,N_24560);
and UO_671 (O_671,N_24528,N_24695);
nand UO_672 (O_672,N_24880,N_24812);
and UO_673 (O_673,N_24685,N_24781);
and UO_674 (O_674,N_24539,N_24930);
nand UO_675 (O_675,N_24827,N_24899);
and UO_676 (O_676,N_24961,N_24957);
nor UO_677 (O_677,N_24728,N_24931);
and UO_678 (O_678,N_24562,N_24665);
or UO_679 (O_679,N_24522,N_24827);
and UO_680 (O_680,N_24655,N_24974);
or UO_681 (O_681,N_24853,N_24706);
or UO_682 (O_682,N_24715,N_24616);
xor UO_683 (O_683,N_24795,N_24673);
nor UO_684 (O_684,N_24838,N_24741);
or UO_685 (O_685,N_24753,N_24868);
and UO_686 (O_686,N_24920,N_24807);
or UO_687 (O_687,N_24860,N_24711);
nand UO_688 (O_688,N_24763,N_24918);
nor UO_689 (O_689,N_24855,N_24752);
nor UO_690 (O_690,N_24539,N_24589);
or UO_691 (O_691,N_24698,N_24524);
and UO_692 (O_692,N_24626,N_24888);
xor UO_693 (O_693,N_24965,N_24747);
and UO_694 (O_694,N_24679,N_24632);
and UO_695 (O_695,N_24768,N_24954);
and UO_696 (O_696,N_24918,N_24759);
nand UO_697 (O_697,N_24761,N_24774);
and UO_698 (O_698,N_24605,N_24674);
or UO_699 (O_699,N_24807,N_24893);
xor UO_700 (O_700,N_24937,N_24501);
nand UO_701 (O_701,N_24794,N_24887);
nand UO_702 (O_702,N_24925,N_24817);
nand UO_703 (O_703,N_24675,N_24959);
and UO_704 (O_704,N_24846,N_24589);
and UO_705 (O_705,N_24944,N_24701);
nor UO_706 (O_706,N_24508,N_24701);
nor UO_707 (O_707,N_24576,N_24932);
or UO_708 (O_708,N_24891,N_24975);
and UO_709 (O_709,N_24986,N_24602);
or UO_710 (O_710,N_24928,N_24511);
or UO_711 (O_711,N_24592,N_24841);
nor UO_712 (O_712,N_24969,N_24500);
or UO_713 (O_713,N_24752,N_24620);
nor UO_714 (O_714,N_24835,N_24614);
nor UO_715 (O_715,N_24749,N_24791);
or UO_716 (O_716,N_24763,N_24541);
and UO_717 (O_717,N_24892,N_24644);
or UO_718 (O_718,N_24511,N_24866);
nand UO_719 (O_719,N_24916,N_24855);
nand UO_720 (O_720,N_24695,N_24566);
and UO_721 (O_721,N_24815,N_24885);
and UO_722 (O_722,N_24933,N_24842);
and UO_723 (O_723,N_24852,N_24927);
nor UO_724 (O_724,N_24705,N_24855);
nor UO_725 (O_725,N_24554,N_24934);
or UO_726 (O_726,N_24615,N_24940);
nor UO_727 (O_727,N_24895,N_24776);
or UO_728 (O_728,N_24657,N_24676);
and UO_729 (O_729,N_24721,N_24783);
nor UO_730 (O_730,N_24860,N_24739);
or UO_731 (O_731,N_24811,N_24870);
nand UO_732 (O_732,N_24713,N_24831);
or UO_733 (O_733,N_24790,N_24754);
and UO_734 (O_734,N_24635,N_24862);
nand UO_735 (O_735,N_24738,N_24629);
or UO_736 (O_736,N_24755,N_24574);
nor UO_737 (O_737,N_24508,N_24979);
nand UO_738 (O_738,N_24550,N_24920);
nor UO_739 (O_739,N_24890,N_24913);
nor UO_740 (O_740,N_24546,N_24813);
nand UO_741 (O_741,N_24842,N_24554);
nand UO_742 (O_742,N_24573,N_24963);
nand UO_743 (O_743,N_24715,N_24787);
or UO_744 (O_744,N_24659,N_24877);
nor UO_745 (O_745,N_24817,N_24711);
nor UO_746 (O_746,N_24606,N_24922);
nor UO_747 (O_747,N_24787,N_24660);
nor UO_748 (O_748,N_24920,N_24612);
nor UO_749 (O_749,N_24996,N_24576);
or UO_750 (O_750,N_24649,N_24829);
nor UO_751 (O_751,N_24713,N_24900);
nand UO_752 (O_752,N_24556,N_24821);
and UO_753 (O_753,N_24685,N_24947);
or UO_754 (O_754,N_24948,N_24696);
nand UO_755 (O_755,N_24779,N_24530);
nand UO_756 (O_756,N_24608,N_24859);
nand UO_757 (O_757,N_24884,N_24743);
or UO_758 (O_758,N_24808,N_24834);
nor UO_759 (O_759,N_24690,N_24912);
or UO_760 (O_760,N_24921,N_24814);
nor UO_761 (O_761,N_24719,N_24548);
or UO_762 (O_762,N_24585,N_24704);
and UO_763 (O_763,N_24899,N_24612);
or UO_764 (O_764,N_24763,N_24869);
nor UO_765 (O_765,N_24665,N_24525);
and UO_766 (O_766,N_24789,N_24610);
or UO_767 (O_767,N_24643,N_24688);
or UO_768 (O_768,N_24886,N_24730);
nand UO_769 (O_769,N_24744,N_24828);
nor UO_770 (O_770,N_24745,N_24821);
nand UO_771 (O_771,N_24503,N_24664);
nor UO_772 (O_772,N_24812,N_24988);
or UO_773 (O_773,N_24636,N_24778);
and UO_774 (O_774,N_24685,N_24843);
nor UO_775 (O_775,N_24529,N_24748);
or UO_776 (O_776,N_24645,N_24928);
nand UO_777 (O_777,N_24930,N_24588);
nor UO_778 (O_778,N_24824,N_24523);
nand UO_779 (O_779,N_24914,N_24802);
nor UO_780 (O_780,N_24598,N_24818);
and UO_781 (O_781,N_24549,N_24917);
and UO_782 (O_782,N_24685,N_24964);
nand UO_783 (O_783,N_24986,N_24680);
nor UO_784 (O_784,N_24514,N_24670);
and UO_785 (O_785,N_24971,N_24541);
nor UO_786 (O_786,N_24573,N_24777);
nand UO_787 (O_787,N_24939,N_24640);
nand UO_788 (O_788,N_24524,N_24511);
and UO_789 (O_789,N_24890,N_24765);
or UO_790 (O_790,N_24724,N_24558);
nand UO_791 (O_791,N_24744,N_24665);
and UO_792 (O_792,N_24742,N_24944);
and UO_793 (O_793,N_24681,N_24795);
nand UO_794 (O_794,N_24684,N_24887);
nand UO_795 (O_795,N_24518,N_24633);
nand UO_796 (O_796,N_24860,N_24756);
nor UO_797 (O_797,N_24596,N_24862);
nand UO_798 (O_798,N_24865,N_24985);
or UO_799 (O_799,N_24915,N_24689);
and UO_800 (O_800,N_24528,N_24961);
or UO_801 (O_801,N_24937,N_24663);
and UO_802 (O_802,N_24913,N_24673);
or UO_803 (O_803,N_24908,N_24860);
or UO_804 (O_804,N_24829,N_24787);
or UO_805 (O_805,N_24805,N_24856);
nor UO_806 (O_806,N_24633,N_24667);
or UO_807 (O_807,N_24946,N_24683);
or UO_808 (O_808,N_24574,N_24856);
nand UO_809 (O_809,N_24693,N_24782);
nor UO_810 (O_810,N_24617,N_24781);
nor UO_811 (O_811,N_24572,N_24966);
and UO_812 (O_812,N_24517,N_24502);
nor UO_813 (O_813,N_24741,N_24788);
and UO_814 (O_814,N_24911,N_24728);
nand UO_815 (O_815,N_24804,N_24771);
nor UO_816 (O_816,N_24913,N_24757);
and UO_817 (O_817,N_24521,N_24660);
nand UO_818 (O_818,N_24610,N_24952);
nor UO_819 (O_819,N_24874,N_24843);
or UO_820 (O_820,N_24557,N_24591);
nor UO_821 (O_821,N_24962,N_24597);
nor UO_822 (O_822,N_24974,N_24920);
nand UO_823 (O_823,N_24724,N_24521);
or UO_824 (O_824,N_24817,N_24851);
nand UO_825 (O_825,N_24548,N_24677);
or UO_826 (O_826,N_24980,N_24700);
xor UO_827 (O_827,N_24951,N_24880);
nor UO_828 (O_828,N_24662,N_24594);
nor UO_829 (O_829,N_24997,N_24601);
nand UO_830 (O_830,N_24554,N_24726);
nand UO_831 (O_831,N_24779,N_24797);
nor UO_832 (O_832,N_24599,N_24583);
and UO_833 (O_833,N_24644,N_24564);
or UO_834 (O_834,N_24827,N_24699);
and UO_835 (O_835,N_24884,N_24881);
or UO_836 (O_836,N_24549,N_24773);
and UO_837 (O_837,N_24964,N_24672);
nand UO_838 (O_838,N_24702,N_24524);
nand UO_839 (O_839,N_24899,N_24680);
nand UO_840 (O_840,N_24910,N_24782);
and UO_841 (O_841,N_24517,N_24947);
nand UO_842 (O_842,N_24561,N_24711);
nand UO_843 (O_843,N_24729,N_24943);
nand UO_844 (O_844,N_24501,N_24655);
or UO_845 (O_845,N_24979,N_24600);
and UO_846 (O_846,N_24629,N_24513);
nor UO_847 (O_847,N_24847,N_24774);
nand UO_848 (O_848,N_24704,N_24859);
nor UO_849 (O_849,N_24995,N_24981);
nand UO_850 (O_850,N_24746,N_24535);
nand UO_851 (O_851,N_24809,N_24645);
and UO_852 (O_852,N_24993,N_24726);
nand UO_853 (O_853,N_24502,N_24664);
nor UO_854 (O_854,N_24906,N_24598);
nand UO_855 (O_855,N_24525,N_24843);
and UO_856 (O_856,N_24957,N_24612);
and UO_857 (O_857,N_24894,N_24906);
xor UO_858 (O_858,N_24550,N_24942);
nand UO_859 (O_859,N_24690,N_24966);
nor UO_860 (O_860,N_24509,N_24931);
nand UO_861 (O_861,N_24536,N_24972);
or UO_862 (O_862,N_24713,N_24743);
nor UO_863 (O_863,N_24782,N_24628);
nor UO_864 (O_864,N_24550,N_24943);
nor UO_865 (O_865,N_24807,N_24711);
xor UO_866 (O_866,N_24730,N_24845);
and UO_867 (O_867,N_24699,N_24560);
nand UO_868 (O_868,N_24537,N_24718);
nand UO_869 (O_869,N_24531,N_24671);
and UO_870 (O_870,N_24856,N_24504);
and UO_871 (O_871,N_24703,N_24939);
nor UO_872 (O_872,N_24937,N_24983);
and UO_873 (O_873,N_24799,N_24594);
or UO_874 (O_874,N_24821,N_24864);
nor UO_875 (O_875,N_24935,N_24721);
or UO_876 (O_876,N_24762,N_24842);
nand UO_877 (O_877,N_24807,N_24922);
xnor UO_878 (O_878,N_24654,N_24701);
nand UO_879 (O_879,N_24737,N_24621);
nand UO_880 (O_880,N_24617,N_24639);
nand UO_881 (O_881,N_24947,N_24525);
and UO_882 (O_882,N_24819,N_24988);
nor UO_883 (O_883,N_24559,N_24779);
nand UO_884 (O_884,N_24825,N_24863);
and UO_885 (O_885,N_24771,N_24848);
and UO_886 (O_886,N_24704,N_24551);
and UO_887 (O_887,N_24902,N_24636);
and UO_888 (O_888,N_24560,N_24594);
nand UO_889 (O_889,N_24652,N_24956);
nand UO_890 (O_890,N_24570,N_24550);
nor UO_891 (O_891,N_24771,N_24638);
or UO_892 (O_892,N_24991,N_24888);
nor UO_893 (O_893,N_24863,N_24543);
nand UO_894 (O_894,N_24684,N_24641);
xnor UO_895 (O_895,N_24926,N_24922);
or UO_896 (O_896,N_24552,N_24835);
nor UO_897 (O_897,N_24878,N_24870);
nand UO_898 (O_898,N_24884,N_24634);
and UO_899 (O_899,N_24637,N_24855);
nor UO_900 (O_900,N_24756,N_24791);
nor UO_901 (O_901,N_24941,N_24596);
xnor UO_902 (O_902,N_24516,N_24615);
or UO_903 (O_903,N_24983,N_24611);
nand UO_904 (O_904,N_24966,N_24581);
nor UO_905 (O_905,N_24708,N_24992);
or UO_906 (O_906,N_24779,N_24844);
nand UO_907 (O_907,N_24928,N_24744);
nor UO_908 (O_908,N_24775,N_24915);
nor UO_909 (O_909,N_24516,N_24788);
nor UO_910 (O_910,N_24623,N_24574);
and UO_911 (O_911,N_24510,N_24615);
or UO_912 (O_912,N_24541,N_24981);
nand UO_913 (O_913,N_24631,N_24638);
nor UO_914 (O_914,N_24726,N_24873);
nand UO_915 (O_915,N_24522,N_24873);
nor UO_916 (O_916,N_24731,N_24590);
or UO_917 (O_917,N_24913,N_24619);
nor UO_918 (O_918,N_24535,N_24972);
and UO_919 (O_919,N_24952,N_24779);
nand UO_920 (O_920,N_24830,N_24766);
xnor UO_921 (O_921,N_24811,N_24911);
nor UO_922 (O_922,N_24844,N_24759);
and UO_923 (O_923,N_24967,N_24829);
and UO_924 (O_924,N_24770,N_24507);
nand UO_925 (O_925,N_24836,N_24734);
and UO_926 (O_926,N_24600,N_24923);
nor UO_927 (O_927,N_24507,N_24713);
or UO_928 (O_928,N_24970,N_24898);
nand UO_929 (O_929,N_24689,N_24727);
nand UO_930 (O_930,N_24590,N_24738);
or UO_931 (O_931,N_24707,N_24718);
and UO_932 (O_932,N_24601,N_24909);
and UO_933 (O_933,N_24671,N_24771);
and UO_934 (O_934,N_24715,N_24567);
nor UO_935 (O_935,N_24544,N_24854);
or UO_936 (O_936,N_24828,N_24915);
nor UO_937 (O_937,N_24824,N_24694);
or UO_938 (O_938,N_24778,N_24718);
nor UO_939 (O_939,N_24796,N_24634);
nand UO_940 (O_940,N_24923,N_24926);
or UO_941 (O_941,N_24676,N_24691);
and UO_942 (O_942,N_24804,N_24553);
and UO_943 (O_943,N_24548,N_24763);
nor UO_944 (O_944,N_24554,N_24626);
nor UO_945 (O_945,N_24848,N_24895);
or UO_946 (O_946,N_24798,N_24770);
or UO_947 (O_947,N_24582,N_24911);
nand UO_948 (O_948,N_24923,N_24835);
and UO_949 (O_949,N_24699,N_24595);
and UO_950 (O_950,N_24592,N_24619);
nor UO_951 (O_951,N_24514,N_24712);
nand UO_952 (O_952,N_24526,N_24790);
and UO_953 (O_953,N_24884,N_24720);
or UO_954 (O_954,N_24844,N_24503);
and UO_955 (O_955,N_24928,N_24865);
and UO_956 (O_956,N_24869,N_24939);
nor UO_957 (O_957,N_24857,N_24534);
nor UO_958 (O_958,N_24711,N_24651);
and UO_959 (O_959,N_24553,N_24999);
nor UO_960 (O_960,N_24523,N_24595);
and UO_961 (O_961,N_24960,N_24712);
or UO_962 (O_962,N_24547,N_24720);
and UO_963 (O_963,N_24875,N_24793);
nand UO_964 (O_964,N_24876,N_24844);
and UO_965 (O_965,N_24969,N_24991);
nor UO_966 (O_966,N_24625,N_24612);
nand UO_967 (O_967,N_24740,N_24730);
or UO_968 (O_968,N_24566,N_24722);
or UO_969 (O_969,N_24556,N_24873);
nor UO_970 (O_970,N_24718,N_24650);
nand UO_971 (O_971,N_24681,N_24887);
or UO_972 (O_972,N_24990,N_24735);
and UO_973 (O_973,N_24551,N_24974);
nand UO_974 (O_974,N_24768,N_24681);
nand UO_975 (O_975,N_24655,N_24594);
nand UO_976 (O_976,N_24819,N_24545);
or UO_977 (O_977,N_24546,N_24763);
nand UO_978 (O_978,N_24946,N_24906);
nand UO_979 (O_979,N_24779,N_24683);
or UO_980 (O_980,N_24989,N_24874);
or UO_981 (O_981,N_24652,N_24770);
and UO_982 (O_982,N_24732,N_24530);
nand UO_983 (O_983,N_24725,N_24650);
nand UO_984 (O_984,N_24821,N_24613);
nand UO_985 (O_985,N_24891,N_24950);
or UO_986 (O_986,N_24891,N_24837);
and UO_987 (O_987,N_24728,N_24566);
or UO_988 (O_988,N_24519,N_24956);
and UO_989 (O_989,N_24807,N_24510);
or UO_990 (O_990,N_24533,N_24552);
nor UO_991 (O_991,N_24874,N_24576);
or UO_992 (O_992,N_24913,N_24579);
and UO_993 (O_993,N_24748,N_24685);
nor UO_994 (O_994,N_24571,N_24875);
nand UO_995 (O_995,N_24867,N_24964);
nand UO_996 (O_996,N_24745,N_24629);
or UO_997 (O_997,N_24562,N_24898);
nor UO_998 (O_998,N_24757,N_24590);
nor UO_999 (O_999,N_24548,N_24748);
and UO_1000 (O_1000,N_24867,N_24532);
and UO_1001 (O_1001,N_24559,N_24613);
nor UO_1002 (O_1002,N_24664,N_24889);
and UO_1003 (O_1003,N_24522,N_24811);
or UO_1004 (O_1004,N_24840,N_24761);
or UO_1005 (O_1005,N_24900,N_24777);
nand UO_1006 (O_1006,N_24736,N_24982);
or UO_1007 (O_1007,N_24682,N_24981);
or UO_1008 (O_1008,N_24985,N_24753);
and UO_1009 (O_1009,N_24748,N_24690);
nand UO_1010 (O_1010,N_24597,N_24664);
nor UO_1011 (O_1011,N_24536,N_24867);
and UO_1012 (O_1012,N_24756,N_24956);
xnor UO_1013 (O_1013,N_24777,N_24986);
nor UO_1014 (O_1014,N_24503,N_24769);
nand UO_1015 (O_1015,N_24753,N_24623);
and UO_1016 (O_1016,N_24552,N_24693);
and UO_1017 (O_1017,N_24615,N_24629);
and UO_1018 (O_1018,N_24694,N_24541);
or UO_1019 (O_1019,N_24766,N_24924);
and UO_1020 (O_1020,N_24541,N_24531);
or UO_1021 (O_1021,N_24967,N_24907);
nand UO_1022 (O_1022,N_24960,N_24875);
and UO_1023 (O_1023,N_24794,N_24594);
and UO_1024 (O_1024,N_24989,N_24960);
nand UO_1025 (O_1025,N_24894,N_24573);
and UO_1026 (O_1026,N_24668,N_24585);
nor UO_1027 (O_1027,N_24769,N_24676);
or UO_1028 (O_1028,N_24721,N_24782);
nand UO_1029 (O_1029,N_24729,N_24921);
nand UO_1030 (O_1030,N_24991,N_24583);
or UO_1031 (O_1031,N_24856,N_24678);
and UO_1032 (O_1032,N_24894,N_24992);
nand UO_1033 (O_1033,N_24800,N_24648);
or UO_1034 (O_1034,N_24808,N_24866);
and UO_1035 (O_1035,N_24557,N_24948);
nor UO_1036 (O_1036,N_24662,N_24681);
and UO_1037 (O_1037,N_24971,N_24899);
and UO_1038 (O_1038,N_24506,N_24610);
and UO_1039 (O_1039,N_24837,N_24648);
and UO_1040 (O_1040,N_24980,N_24976);
nor UO_1041 (O_1041,N_24860,N_24633);
nand UO_1042 (O_1042,N_24934,N_24720);
and UO_1043 (O_1043,N_24771,N_24549);
nor UO_1044 (O_1044,N_24610,N_24685);
nand UO_1045 (O_1045,N_24776,N_24964);
or UO_1046 (O_1046,N_24659,N_24831);
or UO_1047 (O_1047,N_24960,N_24905);
nand UO_1048 (O_1048,N_24536,N_24504);
and UO_1049 (O_1049,N_24957,N_24750);
or UO_1050 (O_1050,N_24601,N_24689);
or UO_1051 (O_1051,N_24946,N_24565);
and UO_1052 (O_1052,N_24745,N_24747);
nand UO_1053 (O_1053,N_24537,N_24528);
and UO_1054 (O_1054,N_24942,N_24699);
nand UO_1055 (O_1055,N_24711,N_24750);
nor UO_1056 (O_1056,N_24560,N_24933);
or UO_1057 (O_1057,N_24661,N_24553);
nand UO_1058 (O_1058,N_24742,N_24922);
or UO_1059 (O_1059,N_24837,N_24602);
nand UO_1060 (O_1060,N_24823,N_24580);
or UO_1061 (O_1061,N_24837,N_24791);
nor UO_1062 (O_1062,N_24737,N_24834);
nor UO_1063 (O_1063,N_24809,N_24725);
and UO_1064 (O_1064,N_24976,N_24841);
nor UO_1065 (O_1065,N_24911,N_24619);
and UO_1066 (O_1066,N_24909,N_24914);
and UO_1067 (O_1067,N_24850,N_24806);
nand UO_1068 (O_1068,N_24904,N_24567);
or UO_1069 (O_1069,N_24585,N_24887);
or UO_1070 (O_1070,N_24532,N_24775);
or UO_1071 (O_1071,N_24717,N_24942);
and UO_1072 (O_1072,N_24927,N_24876);
nor UO_1073 (O_1073,N_24908,N_24681);
xnor UO_1074 (O_1074,N_24619,N_24593);
and UO_1075 (O_1075,N_24548,N_24904);
nand UO_1076 (O_1076,N_24604,N_24649);
nand UO_1077 (O_1077,N_24544,N_24614);
and UO_1078 (O_1078,N_24789,N_24747);
and UO_1079 (O_1079,N_24652,N_24823);
nand UO_1080 (O_1080,N_24877,N_24560);
nor UO_1081 (O_1081,N_24639,N_24829);
and UO_1082 (O_1082,N_24787,N_24850);
or UO_1083 (O_1083,N_24617,N_24715);
and UO_1084 (O_1084,N_24919,N_24681);
nor UO_1085 (O_1085,N_24706,N_24540);
or UO_1086 (O_1086,N_24627,N_24897);
and UO_1087 (O_1087,N_24593,N_24683);
and UO_1088 (O_1088,N_24958,N_24544);
or UO_1089 (O_1089,N_24880,N_24791);
xor UO_1090 (O_1090,N_24618,N_24755);
or UO_1091 (O_1091,N_24568,N_24824);
nor UO_1092 (O_1092,N_24714,N_24744);
nor UO_1093 (O_1093,N_24553,N_24823);
and UO_1094 (O_1094,N_24954,N_24500);
or UO_1095 (O_1095,N_24794,N_24811);
nor UO_1096 (O_1096,N_24802,N_24868);
nor UO_1097 (O_1097,N_24842,N_24536);
nand UO_1098 (O_1098,N_24944,N_24622);
and UO_1099 (O_1099,N_24541,N_24738);
nand UO_1100 (O_1100,N_24956,N_24834);
or UO_1101 (O_1101,N_24941,N_24691);
nand UO_1102 (O_1102,N_24891,N_24650);
and UO_1103 (O_1103,N_24687,N_24856);
and UO_1104 (O_1104,N_24710,N_24875);
or UO_1105 (O_1105,N_24875,N_24787);
nor UO_1106 (O_1106,N_24837,N_24991);
or UO_1107 (O_1107,N_24678,N_24646);
nor UO_1108 (O_1108,N_24871,N_24667);
or UO_1109 (O_1109,N_24784,N_24589);
nand UO_1110 (O_1110,N_24724,N_24784);
nor UO_1111 (O_1111,N_24882,N_24593);
or UO_1112 (O_1112,N_24933,N_24759);
nand UO_1113 (O_1113,N_24924,N_24786);
or UO_1114 (O_1114,N_24534,N_24969);
and UO_1115 (O_1115,N_24921,N_24843);
nor UO_1116 (O_1116,N_24868,N_24765);
or UO_1117 (O_1117,N_24705,N_24669);
or UO_1118 (O_1118,N_24561,N_24696);
nor UO_1119 (O_1119,N_24591,N_24660);
nand UO_1120 (O_1120,N_24713,N_24585);
nor UO_1121 (O_1121,N_24508,N_24977);
or UO_1122 (O_1122,N_24521,N_24705);
or UO_1123 (O_1123,N_24767,N_24715);
or UO_1124 (O_1124,N_24518,N_24638);
nor UO_1125 (O_1125,N_24971,N_24553);
nand UO_1126 (O_1126,N_24613,N_24691);
and UO_1127 (O_1127,N_24555,N_24611);
and UO_1128 (O_1128,N_24540,N_24689);
nor UO_1129 (O_1129,N_24504,N_24897);
or UO_1130 (O_1130,N_24737,N_24630);
nand UO_1131 (O_1131,N_24518,N_24719);
nand UO_1132 (O_1132,N_24815,N_24529);
nor UO_1133 (O_1133,N_24554,N_24540);
or UO_1134 (O_1134,N_24891,N_24936);
and UO_1135 (O_1135,N_24766,N_24811);
nor UO_1136 (O_1136,N_24954,N_24788);
or UO_1137 (O_1137,N_24873,N_24757);
nor UO_1138 (O_1138,N_24756,N_24926);
and UO_1139 (O_1139,N_24841,N_24689);
and UO_1140 (O_1140,N_24802,N_24826);
or UO_1141 (O_1141,N_24526,N_24537);
or UO_1142 (O_1142,N_24568,N_24982);
or UO_1143 (O_1143,N_24881,N_24870);
nand UO_1144 (O_1144,N_24523,N_24544);
nor UO_1145 (O_1145,N_24566,N_24878);
nor UO_1146 (O_1146,N_24670,N_24590);
nor UO_1147 (O_1147,N_24879,N_24866);
nor UO_1148 (O_1148,N_24939,N_24583);
nand UO_1149 (O_1149,N_24930,N_24830);
and UO_1150 (O_1150,N_24938,N_24605);
and UO_1151 (O_1151,N_24585,N_24752);
nor UO_1152 (O_1152,N_24910,N_24904);
nand UO_1153 (O_1153,N_24917,N_24723);
nand UO_1154 (O_1154,N_24598,N_24776);
and UO_1155 (O_1155,N_24532,N_24700);
and UO_1156 (O_1156,N_24655,N_24862);
and UO_1157 (O_1157,N_24756,N_24792);
and UO_1158 (O_1158,N_24664,N_24649);
or UO_1159 (O_1159,N_24878,N_24927);
and UO_1160 (O_1160,N_24641,N_24605);
nand UO_1161 (O_1161,N_24744,N_24522);
nand UO_1162 (O_1162,N_24572,N_24643);
or UO_1163 (O_1163,N_24956,N_24905);
nand UO_1164 (O_1164,N_24587,N_24854);
or UO_1165 (O_1165,N_24962,N_24742);
and UO_1166 (O_1166,N_24983,N_24924);
or UO_1167 (O_1167,N_24680,N_24807);
or UO_1168 (O_1168,N_24680,N_24585);
nor UO_1169 (O_1169,N_24994,N_24859);
nor UO_1170 (O_1170,N_24879,N_24766);
nor UO_1171 (O_1171,N_24776,N_24968);
nor UO_1172 (O_1172,N_24899,N_24834);
and UO_1173 (O_1173,N_24847,N_24881);
nand UO_1174 (O_1174,N_24590,N_24500);
xnor UO_1175 (O_1175,N_24877,N_24587);
and UO_1176 (O_1176,N_24756,N_24897);
nor UO_1177 (O_1177,N_24751,N_24589);
nand UO_1178 (O_1178,N_24524,N_24995);
nand UO_1179 (O_1179,N_24914,N_24886);
nor UO_1180 (O_1180,N_24687,N_24510);
and UO_1181 (O_1181,N_24712,N_24793);
nand UO_1182 (O_1182,N_24808,N_24858);
xor UO_1183 (O_1183,N_24711,N_24545);
nand UO_1184 (O_1184,N_24935,N_24608);
nand UO_1185 (O_1185,N_24807,N_24985);
nor UO_1186 (O_1186,N_24763,N_24718);
nor UO_1187 (O_1187,N_24858,N_24700);
or UO_1188 (O_1188,N_24772,N_24513);
nor UO_1189 (O_1189,N_24750,N_24807);
nand UO_1190 (O_1190,N_24932,N_24852);
and UO_1191 (O_1191,N_24909,N_24722);
nor UO_1192 (O_1192,N_24786,N_24593);
or UO_1193 (O_1193,N_24864,N_24543);
or UO_1194 (O_1194,N_24584,N_24901);
nor UO_1195 (O_1195,N_24738,N_24514);
nand UO_1196 (O_1196,N_24639,N_24584);
nand UO_1197 (O_1197,N_24642,N_24605);
and UO_1198 (O_1198,N_24697,N_24755);
nand UO_1199 (O_1199,N_24504,N_24701);
or UO_1200 (O_1200,N_24726,N_24579);
nor UO_1201 (O_1201,N_24575,N_24553);
nor UO_1202 (O_1202,N_24558,N_24854);
nor UO_1203 (O_1203,N_24707,N_24658);
nor UO_1204 (O_1204,N_24721,N_24694);
or UO_1205 (O_1205,N_24840,N_24974);
nand UO_1206 (O_1206,N_24878,N_24699);
nand UO_1207 (O_1207,N_24997,N_24734);
nand UO_1208 (O_1208,N_24744,N_24814);
or UO_1209 (O_1209,N_24592,N_24578);
and UO_1210 (O_1210,N_24701,N_24580);
nand UO_1211 (O_1211,N_24672,N_24639);
nand UO_1212 (O_1212,N_24584,N_24667);
nand UO_1213 (O_1213,N_24864,N_24622);
and UO_1214 (O_1214,N_24622,N_24875);
nor UO_1215 (O_1215,N_24921,N_24930);
nor UO_1216 (O_1216,N_24660,N_24574);
nor UO_1217 (O_1217,N_24717,N_24962);
and UO_1218 (O_1218,N_24761,N_24854);
nand UO_1219 (O_1219,N_24814,N_24687);
and UO_1220 (O_1220,N_24970,N_24988);
and UO_1221 (O_1221,N_24857,N_24950);
and UO_1222 (O_1222,N_24654,N_24911);
nand UO_1223 (O_1223,N_24512,N_24850);
or UO_1224 (O_1224,N_24744,N_24610);
or UO_1225 (O_1225,N_24716,N_24664);
and UO_1226 (O_1226,N_24788,N_24686);
nor UO_1227 (O_1227,N_24961,N_24720);
nand UO_1228 (O_1228,N_24820,N_24843);
nor UO_1229 (O_1229,N_24966,N_24596);
nand UO_1230 (O_1230,N_24977,N_24667);
and UO_1231 (O_1231,N_24526,N_24752);
nand UO_1232 (O_1232,N_24803,N_24724);
and UO_1233 (O_1233,N_24913,N_24637);
and UO_1234 (O_1234,N_24588,N_24813);
or UO_1235 (O_1235,N_24565,N_24537);
and UO_1236 (O_1236,N_24922,N_24528);
nand UO_1237 (O_1237,N_24886,N_24552);
nor UO_1238 (O_1238,N_24592,N_24813);
nand UO_1239 (O_1239,N_24974,N_24946);
and UO_1240 (O_1240,N_24504,N_24819);
or UO_1241 (O_1241,N_24920,N_24605);
or UO_1242 (O_1242,N_24564,N_24641);
or UO_1243 (O_1243,N_24623,N_24935);
or UO_1244 (O_1244,N_24559,N_24743);
nor UO_1245 (O_1245,N_24567,N_24752);
or UO_1246 (O_1246,N_24752,N_24661);
nor UO_1247 (O_1247,N_24760,N_24599);
and UO_1248 (O_1248,N_24572,N_24758);
xnor UO_1249 (O_1249,N_24590,N_24675);
xor UO_1250 (O_1250,N_24791,N_24964);
nor UO_1251 (O_1251,N_24602,N_24615);
nand UO_1252 (O_1252,N_24935,N_24977);
or UO_1253 (O_1253,N_24893,N_24993);
nor UO_1254 (O_1254,N_24888,N_24910);
nand UO_1255 (O_1255,N_24913,N_24922);
or UO_1256 (O_1256,N_24968,N_24980);
and UO_1257 (O_1257,N_24689,N_24605);
nor UO_1258 (O_1258,N_24589,N_24511);
nor UO_1259 (O_1259,N_24720,N_24565);
nor UO_1260 (O_1260,N_24807,N_24702);
and UO_1261 (O_1261,N_24796,N_24734);
nor UO_1262 (O_1262,N_24506,N_24879);
or UO_1263 (O_1263,N_24801,N_24710);
xor UO_1264 (O_1264,N_24998,N_24966);
nor UO_1265 (O_1265,N_24779,N_24640);
and UO_1266 (O_1266,N_24552,N_24959);
or UO_1267 (O_1267,N_24817,N_24700);
and UO_1268 (O_1268,N_24564,N_24790);
and UO_1269 (O_1269,N_24577,N_24899);
nor UO_1270 (O_1270,N_24942,N_24785);
and UO_1271 (O_1271,N_24766,N_24699);
and UO_1272 (O_1272,N_24666,N_24517);
nand UO_1273 (O_1273,N_24594,N_24752);
and UO_1274 (O_1274,N_24830,N_24576);
nor UO_1275 (O_1275,N_24625,N_24724);
xnor UO_1276 (O_1276,N_24785,N_24932);
nand UO_1277 (O_1277,N_24934,N_24909);
xnor UO_1278 (O_1278,N_24634,N_24561);
or UO_1279 (O_1279,N_24635,N_24782);
nand UO_1280 (O_1280,N_24618,N_24652);
and UO_1281 (O_1281,N_24689,N_24939);
nand UO_1282 (O_1282,N_24539,N_24752);
or UO_1283 (O_1283,N_24669,N_24903);
nor UO_1284 (O_1284,N_24813,N_24616);
nand UO_1285 (O_1285,N_24748,N_24939);
nand UO_1286 (O_1286,N_24892,N_24526);
and UO_1287 (O_1287,N_24966,N_24772);
nor UO_1288 (O_1288,N_24605,N_24655);
nand UO_1289 (O_1289,N_24651,N_24769);
or UO_1290 (O_1290,N_24792,N_24913);
nand UO_1291 (O_1291,N_24571,N_24792);
nor UO_1292 (O_1292,N_24761,N_24514);
nor UO_1293 (O_1293,N_24700,N_24605);
nor UO_1294 (O_1294,N_24670,N_24766);
nand UO_1295 (O_1295,N_24778,N_24867);
and UO_1296 (O_1296,N_24967,N_24697);
or UO_1297 (O_1297,N_24686,N_24826);
or UO_1298 (O_1298,N_24566,N_24546);
and UO_1299 (O_1299,N_24773,N_24652);
nand UO_1300 (O_1300,N_24863,N_24541);
and UO_1301 (O_1301,N_24899,N_24737);
nand UO_1302 (O_1302,N_24859,N_24534);
nand UO_1303 (O_1303,N_24515,N_24585);
or UO_1304 (O_1304,N_24890,N_24843);
nor UO_1305 (O_1305,N_24670,N_24802);
or UO_1306 (O_1306,N_24714,N_24916);
or UO_1307 (O_1307,N_24857,N_24606);
nand UO_1308 (O_1308,N_24687,N_24951);
xor UO_1309 (O_1309,N_24891,N_24850);
nor UO_1310 (O_1310,N_24514,N_24995);
and UO_1311 (O_1311,N_24980,N_24909);
or UO_1312 (O_1312,N_24978,N_24568);
nand UO_1313 (O_1313,N_24842,N_24594);
nor UO_1314 (O_1314,N_24681,N_24927);
and UO_1315 (O_1315,N_24759,N_24972);
and UO_1316 (O_1316,N_24650,N_24793);
nand UO_1317 (O_1317,N_24840,N_24961);
or UO_1318 (O_1318,N_24527,N_24706);
and UO_1319 (O_1319,N_24605,N_24709);
nand UO_1320 (O_1320,N_24683,N_24582);
and UO_1321 (O_1321,N_24994,N_24782);
and UO_1322 (O_1322,N_24662,N_24861);
nand UO_1323 (O_1323,N_24916,N_24940);
nand UO_1324 (O_1324,N_24930,N_24712);
nand UO_1325 (O_1325,N_24559,N_24508);
nor UO_1326 (O_1326,N_24845,N_24945);
and UO_1327 (O_1327,N_24876,N_24641);
nor UO_1328 (O_1328,N_24790,N_24981);
nand UO_1329 (O_1329,N_24820,N_24644);
and UO_1330 (O_1330,N_24858,N_24975);
or UO_1331 (O_1331,N_24633,N_24971);
nand UO_1332 (O_1332,N_24834,N_24994);
or UO_1333 (O_1333,N_24960,N_24912);
or UO_1334 (O_1334,N_24840,N_24940);
nand UO_1335 (O_1335,N_24916,N_24577);
or UO_1336 (O_1336,N_24595,N_24613);
nand UO_1337 (O_1337,N_24539,N_24768);
nand UO_1338 (O_1338,N_24558,N_24797);
nor UO_1339 (O_1339,N_24877,N_24985);
or UO_1340 (O_1340,N_24556,N_24898);
or UO_1341 (O_1341,N_24798,N_24643);
or UO_1342 (O_1342,N_24803,N_24615);
nor UO_1343 (O_1343,N_24967,N_24509);
or UO_1344 (O_1344,N_24554,N_24530);
or UO_1345 (O_1345,N_24766,N_24712);
and UO_1346 (O_1346,N_24888,N_24947);
xnor UO_1347 (O_1347,N_24831,N_24995);
nand UO_1348 (O_1348,N_24656,N_24657);
nand UO_1349 (O_1349,N_24722,N_24677);
or UO_1350 (O_1350,N_24920,N_24754);
and UO_1351 (O_1351,N_24811,N_24894);
nand UO_1352 (O_1352,N_24737,N_24948);
nor UO_1353 (O_1353,N_24550,N_24682);
and UO_1354 (O_1354,N_24873,N_24568);
nor UO_1355 (O_1355,N_24790,N_24996);
or UO_1356 (O_1356,N_24943,N_24524);
and UO_1357 (O_1357,N_24954,N_24522);
nand UO_1358 (O_1358,N_24597,N_24628);
or UO_1359 (O_1359,N_24680,N_24904);
nor UO_1360 (O_1360,N_24502,N_24537);
nor UO_1361 (O_1361,N_24597,N_24932);
or UO_1362 (O_1362,N_24937,N_24560);
or UO_1363 (O_1363,N_24516,N_24534);
and UO_1364 (O_1364,N_24514,N_24678);
or UO_1365 (O_1365,N_24798,N_24835);
nand UO_1366 (O_1366,N_24513,N_24798);
and UO_1367 (O_1367,N_24908,N_24839);
nand UO_1368 (O_1368,N_24567,N_24524);
or UO_1369 (O_1369,N_24619,N_24850);
or UO_1370 (O_1370,N_24953,N_24505);
or UO_1371 (O_1371,N_24921,N_24705);
nor UO_1372 (O_1372,N_24698,N_24754);
nor UO_1373 (O_1373,N_24813,N_24512);
and UO_1374 (O_1374,N_24720,N_24833);
nand UO_1375 (O_1375,N_24920,N_24525);
nor UO_1376 (O_1376,N_24960,N_24501);
or UO_1377 (O_1377,N_24715,N_24605);
and UO_1378 (O_1378,N_24740,N_24659);
nand UO_1379 (O_1379,N_24670,N_24721);
nor UO_1380 (O_1380,N_24684,N_24797);
nand UO_1381 (O_1381,N_24510,N_24812);
and UO_1382 (O_1382,N_24629,N_24690);
or UO_1383 (O_1383,N_24715,N_24735);
or UO_1384 (O_1384,N_24790,N_24972);
nand UO_1385 (O_1385,N_24609,N_24767);
or UO_1386 (O_1386,N_24714,N_24920);
nor UO_1387 (O_1387,N_24845,N_24938);
nor UO_1388 (O_1388,N_24597,N_24609);
nor UO_1389 (O_1389,N_24558,N_24676);
or UO_1390 (O_1390,N_24972,N_24531);
xor UO_1391 (O_1391,N_24778,N_24517);
nand UO_1392 (O_1392,N_24707,N_24923);
xnor UO_1393 (O_1393,N_24657,N_24859);
and UO_1394 (O_1394,N_24756,N_24883);
nor UO_1395 (O_1395,N_24770,N_24781);
nor UO_1396 (O_1396,N_24995,N_24822);
and UO_1397 (O_1397,N_24758,N_24934);
or UO_1398 (O_1398,N_24640,N_24637);
nand UO_1399 (O_1399,N_24645,N_24790);
or UO_1400 (O_1400,N_24705,N_24677);
nand UO_1401 (O_1401,N_24502,N_24928);
nor UO_1402 (O_1402,N_24720,N_24540);
and UO_1403 (O_1403,N_24825,N_24996);
and UO_1404 (O_1404,N_24830,N_24682);
nand UO_1405 (O_1405,N_24654,N_24527);
and UO_1406 (O_1406,N_24608,N_24796);
nor UO_1407 (O_1407,N_24921,N_24818);
nor UO_1408 (O_1408,N_24671,N_24791);
nor UO_1409 (O_1409,N_24620,N_24918);
or UO_1410 (O_1410,N_24971,N_24846);
or UO_1411 (O_1411,N_24527,N_24730);
nand UO_1412 (O_1412,N_24713,N_24669);
nor UO_1413 (O_1413,N_24645,N_24680);
or UO_1414 (O_1414,N_24807,N_24570);
or UO_1415 (O_1415,N_24619,N_24556);
nor UO_1416 (O_1416,N_24626,N_24980);
nor UO_1417 (O_1417,N_24551,N_24770);
or UO_1418 (O_1418,N_24649,N_24755);
or UO_1419 (O_1419,N_24677,N_24539);
or UO_1420 (O_1420,N_24544,N_24701);
and UO_1421 (O_1421,N_24650,N_24647);
nand UO_1422 (O_1422,N_24760,N_24961);
nor UO_1423 (O_1423,N_24669,N_24567);
nand UO_1424 (O_1424,N_24707,N_24838);
nor UO_1425 (O_1425,N_24600,N_24873);
or UO_1426 (O_1426,N_24953,N_24627);
or UO_1427 (O_1427,N_24805,N_24878);
or UO_1428 (O_1428,N_24984,N_24666);
and UO_1429 (O_1429,N_24780,N_24900);
and UO_1430 (O_1430,N_24910,N_24975);
or UO_1431 (O_1431,N_24783,N_24979);
and UO_1432 (O_1432,N_24563,N_24866);
nand UO_1433 (O_1433,N_24746,N_24657);
or UO_1434 (O_1434,N_24524,N_24703);
or UO_1435 (O_1435,N_24580,N_24523);
nor UO_1436 (O_1436,N_24522,N_24980);
or UO_1437 (O_1437,N_24767,N_24783);
nor UO_1438 (O_1438,N_24530,N_24759);
or UO_1439 (O_1439,N_24601,N_24856);
and UO_1440 (O_1440,N_24653,N_24583);
nor UO_1441 (O_1441,N_24721,N_24960);
xor UO_1442 (O_1442,N_24955,N_24887);
nor UO_1443 (O_1443,N_24754,N_24519);
nand UO_1444 (O_1444,N_24567,N_24742);
or UO_1445 (O_1445,N_24614,N_24908);
xnor UO_1446 (O_1446,N_24730,N_24782);
nand UO_1447 (O_1447,N_24700,N_24646);
nor UO_1448 (O_1448,N_24898,N_24912);
nor UO_1449 (O_1449,N_24729,N_24738);
and UO_1450 (O_1450,N_24974,N_24684);
nor UO_1451 (O_1451,N_24961,N_24740);
or UO_1452 (O_1452,N_24648,N_24515);
nor UO_1453 (O_1453,N_24744,N_24858);
and UO_1454 (O_1454,N_24641,N_24994);
nand UO_1455 (O_1455,N_24729,N_24867);
and UO_1456 (O_1456,N_24825,N_24632);
nor UO_1457 (O_1457,N_24660,N_24934);
and UO_1458 (O_1458,N_24543,N_24859);
or UO_1459 (O_1459,N_24877,N_24564);
and UO_1460 (O_1460,N_24535,N_24662);
nor UO_1461 (O_1461,N_24821,N_24852);
and UO_1462 (O_1462,N_24937,N_24741);
nand UO_1463 (O_1463,N_24654,N_24667);
or UO_1464 (O_1464,N_24598,N_24973);
and UO_1465 (O_1465,N_24626,N_24985);
and UO_1466 (O_1466,N_24928,N_24916);
and UO_1467 (O_1467,N_24573,N_24524);
nand UO_1468 (O_1468,N_24543,N_24797);
or UO_1469 (O_1469,N_24574,N_24720);
or UO_1470 (O_1470,N_24649,N_24744);
nor UO_1471 (O_1471,N_24901,N_24616);
or UO_1472 (O_1472,N_24746,N_24528);
or UO_1473 (O_1473,N_24981,N_24858);
or UO_1474 (O_1474,N_24530,N_24905);
or UO_1475 (O_1475,N_24604,N_24632);
and UO_1476 (O_1476,N_24778,N_24898);
nand UO_1477 (O_1477,N_24668,N_24576);
xnor UO_1478 (O_1478,N_24958,N_24547);
nor UO_1479 (O_1479,N_24788,N_24671);
and UO_1480 (O_1480,N_24874,N_24918);
nor UO_1481 (O_1481,N_24573,N_24620);
and UO_1482 (O_1482,N_24872,N_24972);
nor UO_1483 (O_1483,N_24692,N_24878);
and UO_1484 (O_1484,N_24891,N_24537);
xnor UO_1485 (O_1485,N_24996,N_24791);
and UO_1486 (O_1486,N_24773,N_24733);
nand UO_1487 (O_1487,N_24564,N_24721);
or UO_1488 (O_1488,N_24589,N_24726);
or UO_1489 (O_1489,N_24616,N_24927);
nor UO_1490 (O_1490,N_24788,N_24539);
or UO_1491 (O_1491,N_24599,N_24572);
and UO_1492 (O_1492,N_24983,N_24865);
or UO_1493 (O_1493,N_24945,N_24503);
and UO_1494 (O_1494,N_24584,N_24936);
nor UO_1495 (O_1495,N_24758,N_24941);
or UO_1496 (O_1496,N_24852,N_24586);
nor UO_1497 (O_1497,N_24918,N_24757);
nor UO_1498 (O_1498,N_24924,N_24515);
nor UO_1499 (O_1499,N_24802,N_24710);
or UO_1500 (O_1500,N_24624,N_24630);
nor UO_1501 (O_1501,N_24827,N_24849);
and UO_1502 (O_1502,N_24647,N_24875);
and UO_1503 (O_1503,N_24663,N_24788);
xor UO_1504 (O_1504,N_24754,N_24993);
and UO_1505 (O_1505,N_24529,N_24794);
and UO_1506 (O_1506,N_24618,N_24928);
nand UO_1507 (O_1507,N_24506,N_24822);
and UO_1508 (O_1508,N_24966,N_24513);
nor UO_1509 (O_1509,N_24806,N_24586);
nor UO_1510 (O_1510,N_24809,N_24687);
nand UO_1511 (O_1511,N_24923,N_24582);
nor UO_1512 (O_1512,N_24654,N_24852);
or UO_1513 (O_1513,N_24625,N_24793);
nor UO_1514 (O_1514,N_24924,N_24991);
nor UO_1515 (O_1515,N_24530,N_24598);
or UO_1516 (O_1516,N_24926,N_24653);
and UO_1517 (O_1517,N_24672,N_24664);
or UO_1518 (O_1518,N_24657,N_24932);
and UO_1519 (O_1519,N_24720,N_24849);
or UO_1520 (O_1520,N_24591,N_24988);
or UO_1521 (O_1521,N_24992,N_24846);
and UO_1522 (O_1522,N_24551,N_24632);
xor UO_1523 (O_1523,N_24697,N_24618);
nor UO_1524 (O_1524,N_24502,N_24526);
nor UO_1525 (O_1525,N_24500,N_24636);
nor UO_1526 (O_1526,N_24841,N_24657);
and UO_1527 (O_1527,N_24582,N_24824);
and UO_1528 (O_1528,N_24503,N_24747);
and UO_1529 (O_1529,N_24805,N_24645);
nand UO_1530 (O_1530,N_24987,N_24757);
and UO_1531 (O_1531,N_24572,N_24944);
or UO_1532 (O_1532,N_24770,N_24595);
and UO_1533 (O_1533,N_24990,N_24742);
nand UO_1534 (O_1534,N_24608,N_24831);
nor UO_1535 (O_1535,N_24543,N_24512);
nand UO_1536 (O_1536,N_24762,N_24534);
and UO_1537 (O_1537,N_24965,N_24791);
or UO_1538 (O_1538,N_24716,N_24541);
nand UO_1539 (O_1539,N_24768,N_24877);
nor UO_1540 (O_1540,N_24607,N_24940);
or UO_1541 (O_1541,N_24815,N_24895);
nand UO_1542 (O_1542,N_24723,N_24668);
or UO_1543 (O_1543,N_24546,N_24875);
or UO_1544 (O_1544,N_24629,N_24808);
nand UO_1545 (O_1545,N_24759,N_24763);
or UO_1546 (O_1546,N_24853,N_24916);
nor UO_1547 (O_1547,N_24895,N_24878);
and UO_1548 (O_1548,N_24928,N_24969);
or UO_1549 (O_1549,N_24956,N_24919);
nor UO_1550 (O_1550,N_24624,N_24824);
and UO_1551 (O_1551,N_24786,N_24718);
nor UO_1552 (O_1552,N_24806,N_24612);
or UO_1553 (O_1553,N_24739,N_24592);
nand UO_1554 (O_1554,N_24869,N_24908);
or UO_1555 (O_1555,N_24881,N_24903);
and UO_1556 (O_1556,N_24900,N_24618);
nor UO_1557 (O_1557,N_24991,N_24608);
and UO_1558 (O_1558,N_24888,N_24532);
and UO_1559 (O_1559,N_24842,N_24893);
and UO_1560 (O_1560,N_24686,N_24815);
nor UO_1561 (O_1561,N_24938,N_24534);
xnor UO_1562 (O_1562,N_24608,N_24504);
or UO_1563 (O_1563,N_24641,N_24589);
or UO_1564 (O_1564,N_24561,N_24667);
or UO_1565 (O_1565,N_24523,N_24978);
nand UO_1566 (O_1566,N_24588,N_24789);
and UO_1567 (O_1567,N_24705,N_24564);
and UO_1568 (O_1568,N_24817,N_24673);
nand UO_1569 (O_1569,N_24885,N_24735);
or UO_1570 (O_1570,N_24829,N_24744);
nand UO_1571 (O_1571,N_24873,N_24543);
and UO_1572 (O_1572,N_24847,N_24770);
nor UO_1573 (O_1573,N_24733,N_24826);
and UO_1574 (O_1574,N_24769,N_24682);
nand UO_1575 (O_1575,N_24897,N_24997);
or UO_1576 (O_1576,N_24779,N_24727);
nand UO_1577 (O_1577,N_24617,N_24935);
and UO_1578 (O_1578,N_24798,N_24839);
and UO_1579 (O_1579,N_24576,N_24997);
nand UO_1580 (O_1580,N_24525,N_24612);
nor UO_1581 (O_1581,N_24717,N_24651);
nand UO_1582 (O_1582,N_24556,N_24997);
nand UO_1583 (O_1583,N_24640,N_24786);
or UO_1584 (O_1584,N_24923,N_24678);
nand UO_1585 (O_1585,N_24573,N_24897);
nor UO_1586 (O_1586,N_24798,N_24621);
nand UO_1587 (O_1587,N_24713,N_24834);
nand UO_1588 (O_1588,N_24539,N_24708);
or UO_1589 (O_1589,N_24746,N_24761);
and UO_1590 (O_1590,N_24617,N_24859);
nor UO_1591 (O_1591,N_24728,N_24811);
nor UO_1592 (O_1592,N_24910,N_24878);
xnor UO_1593 (O_1593,N_24615,N_24600);
and UO_1594 (O_1594,N_24571,N_24666);
nand UO_1595 (O_1595,N_24570,N_24689);
nor UO_1596 (O_1596,N_24788,N_24547);
and UO_1597 (O_1597,N_24764,N_24734);
or UO_1598 (O_1598,N_24966,N_24704);
and UO_1599 (O_1599,N_24790,N_24634);
nor UO_1600 (O_1600,N_24658,N_24726);
or UO_1601 (O_1601,N_24576,N_24519);
nand UO_1602 (O_1602,N_24970,N_24762);
nand UO_1603 (O_1603,N_24640,N_24714);
nor UO_1604 (O_1604,N_24953,N_24921);
nor UO_1605 (O_1605,N_24572,N_24897);
nand UO_1606 (O_1606,N_24524,N_24517);
or UO_1607 (O_1607,N_24614,N_24842);
nand UO_1608 (O_1608,N_24953,N_24570);
nand UO_1609 (O_1609,N_24742,N_24623);
nand UO_1610 (O_1610,N_24769,N_24814);
and UO_1611 (O_1611,N_24920,N_24640);
or UO_1612 (O_1612,N_24812,N_24551);
or UO_1613 (O_1613,N_24527,N_24669);
or UO_1614 (O_1614,N_24549,N_24700);
nor UO_1615 (O_1615,N_24922,N_24514);
and UO_1616 (O_1616,N_24874,N_24866);
or UO_1617 (O_1617,N_24871,N_24698);
or UO_1618 (O_1618,N_24945,N_24693);
nand UO_1619 (O_1619,N_24830,N_24850);
nor UO_1620 (O_1620,N_24542,N_24767);
nor UO_1621 (O_1621,N_24565,N_24938);
or UO_1622 (O_1622,N_24595,N_24637);
or UO_1623 (O_1623,N_24625,N_24544);
and UO_1624 (O_1624,N_24939,N_24942);
and UO_1625 (O_1625,N_24884,N_24792);
nor UO_1626 (O_1626,N_24538,N_24535);
nand UO_1627 (O_1627,N_24905,N_24768);
nand UO_1628 (O_1628,N_24987,N_24780);
or UO_1629 (O_1629,N_24595,N_24782);
nand UO_1630 (O_1630,N_24773,N_24974);
nor UO_1631 (O_1631,N_24836,N_24547);
and UO_1632 (O_1632,N_24584,N_24713);
and UO_1633 (O_1633,N_24805,N_24631);
or UO_1634 (O_1634,N_24634,N_24919);
nand UO_1635 (O_1635,N_24962,N_24871);
xor UO_1636 (O_1636,N_24787,N_24686);
or UO_1637 (O_1637,N_24711,N_24956);
or UO_1638 (O_1638,N_24830,N_24690);
or UO_1639 (O_1639,N_24698,N_24822);
nand UO_1640 (O_1640,N_24567,N_24698);
and UO_1641 (O_1641,N_24582,N_24862);
or UO_1642 (O_1642,N_24744,N_24654);
nand UO_1643 (O_1643,N_24612,N_24956);
nor UO_1644 (O_1644,N_24543,N_24955);
or UO_1645 (O_1645,N_24865,N_24555);
nor UO_1646 (O_1646,N_24826,N_24514);
nor UO_1647 (O_1647,N_24978,N_24971);
xnor UO_1648 (O_1648,N_24849,N_24515);
nand UO_1649 (O_1649,N_24694,N_24995);
or UO_1650 (O_1650,N_24856,N_24618);
and UO_1651 (O_1651,N_24705,N_24754);
or UO_1652 (O_1652,N_24955,N_24597);
and UO_1653 (O_1653,N_24671,N_24837);
and UO_1654 (O_1654,N_24880,N_24672);
or UO_1655 (O_1655,N_24803,N_24550);
nand UO_1656 (O_1656,N_24708,N_24847);
or UO_1657 (O_1657,N_24988,N_24595);
nor UO_1658 (O_1658,N_24511,N_24947);
or UO_1659 (O_1659,N_24971,N_24852);
or UO_1660 (O_1660,N_24991,N_24544);
nor UO_1661 (O_1661,N_24766,N_24983);
nand UO_1662 (O_1662,N_24853,N_24516);
or UO_1663 (O_1663,N_24542,N_24781);
nand UO_1664 (O_1664,N_24580,N_24997);
nor UO_1665 (O_1665,N_24622,N_24871);
and UO_1666 (O_1666,N_24708,N_24536);
and UO_1667 (O_1667,N_24965,N_24802);
or UO_1668 (O_1668,N_24638,N_24822);
or UO_1669 (O_1669,N_24918,N_24981);
nor UO_1670 (O_1670,N_24932,N_24669);
or UO_1671 (O_1671,N_24703,N_24944);
or UO_1672 (O_1672,N_24879,N_24594);
or UO_1673 (O_1673,N_24953,N_24863);
or UO_1674 (O_1674,N_24657,N_24991);
nor UO_1675 (O_1675,N_24950,N_24712);
xor UO_1676 (O_1676,N_24552,N_24600);
and UO_1677 (O_1677,N_24722,N_24647);
or UO_1678 (O_1678,N_24746,N_24943);
or UO_1679 (O_1679,N_24839,N_24975);
nand UO_1680 (O_1680,N_24721,N_24716);
nand UO_1681 (O_1681,N_24529,N_24501);
and UO_1682 (O_1682,N_24635,N_24849);
nand UO_1683 (O_1683,N_24938,N_24516);
or UO_1684 (O_1684,N_24668,N_24968);
or UO_1685 (O_1685,N_24855,N_24599);
or UO_1686 (O_1686,N_24825,N_24923);
or UO_1687 (O_1687,N_24549,N_24669);
and UO_1688 (O_1688,N_24956,N_24883);
or UO_1689 (O_1689,N_24974,N_24912);
or UO_1690 (O_1690,N_24735,N_24619);
or UO_1691 (O_1691,N_24688,N_24550);
or UO_1692 (O_1692,N_24556,N_24635);
nand UO_1693 (O_1693,N_24553,N_24810);
or UO_1694 (O_1694,N_24780,N_24787);
or UO_1695 (O_1695,N_24893,N_24814);
and UO_1696 (O_1696,N_24729,N_24561);
nand UO_1697 (O_1697,N_24787,N_24566);
or UO_1698 (O_1698,N_24766,N_24959);
or UO_1699 (O_1699,N_24987,N_24999);
or UO_1700 (O_1700,N_24782,N_24966);
and UO_1701 (O_1701,N_24628,N_24911);
nand UO_1702 (O_1702,N_24869,N_24800);
nand UO_1703 (O_1703,N_24570,N_24964);
and UO_1704 (O_1704,N_24963,N_24947);
nand UO_1705 (O_1705,N_24563,N_24943);
and UO_1706 (O_1706,N_24760,N_24827);
nand UO_1707 (O_1707,N_24942,N_24641);
or UO_1708 (O_1708,N_24751,N_24585);
and UO_1709 (O_1709,N_24761,N_24767);
nor UO_1710 (O_1710,N_24755,N_24818);
nor UO_1711 (O_1711,N_24634,N_24864);
nor UO_1712 (O_1712,N_24730,N_24726);
and UO_1713 (O_1713,N_24617,N_24716);
nor UO_1714 (O_1714,N_24888,N_24924);
nor UO_1715 (O_1715,N_24659,N_24709);
and UO_1716 (O_1716,N_24879,N_24806);
and UO_1717 (O_1717,N_24903,N_24784);
and UO_1718 (O_1718,N_24787,N_24960);
nand UO_1719 (O_1719,N_24513,N_24824);
nand UO_1720 (O_1720,N_24991,N_24853);
or UO_1721 (O_1721,N_24776,N_24655);
nor UO_1722 (O_1722,N_24732,N_24928);
and UO_1723 (O_1723,N_24693,N_24630);
and UO_1724 (O_1724,N_24724,N_24883);
or UO_1725 (O_1725,N_24765,N_24616);
nand UO_1726 (O_1726,N_24552,N_24851);
nor UO_1727 (O_1727,N_24534,N_24946);
and UO_1728 (O_1728,N_24681,N_24829);
and UO_1729 (O_1729,N_24510,N_24513);
or UO_1730 (O_1730,N_24696,N_24712);
nand UO_1731 (O_1731,N_24749,N_24812);
nand UO_1732 (O_1732,N_24725,N_24717);
nor UO_1733 (O_1733,N_24694,N_24720);
or UO_1734 (O_1734,N_24665,N_24895);
xnor UO_1735 (O_1735,N_24657,N_24947);
nor UO_1736 (O_1736,N_24898,N_24663);
and UO_1737 (O_1737,N_24814,N_24722);
and UO_1738 (O_1738,N_24517,N_24839);
nor UO_1739 (O_1739,N_24601,N_24850);
nand UO_1740 (O_1740,N_24519,N_24562);
nor UO_1741 (O_1741,N_24569,N_24799);
and UO_1742 (O_1742,N_24869,N_24520);
and UO_1743 (O_1743,N_24672,N_24886);
and UO_1744 (O_1744,N_24860,N_24939);
and UO_1745 (O_1745,N_24820,N_24985);
and UO_1746 (O_1746,N_24643,N_24720);
and UO_1747 (O_1747,N_24593,N_24967);
nand UO_1748 (O_1748,N_24877,N_24666);
and UO_1749 (O_1749,N_24789,N_24983);
and UO_1750 (O_1750,N_24686,N_24847);
nor UO_1751 (O_1751,N_24554,N_24620);
or UO_1752 (O_1752,N_24784,N_24936);
or UO_1753 (O_1753,N_24618,N_24608);
xor UO_1754 (O_1754,N_24674,N_24879);
and UO_1755 (O_1755,N_24579,N_24970);
nor UO_1756 (O_1756,N_24511,N_24794);
or UO_1757 (O_1757,N_24768,N_24834);
and UO_1758 (O_1758,N_24990,N_24595);
nand UO_1759 (O_1759,N_24799,N_24663);
and UO_1760 (O_1760,N_24690,N_24920);
or UO_1761 (O_1761,N_24947,N_24925);
and UO_1762 (O_1762,N_24664,N_24989);
or UO_1763 (O_1763,N_24959,N_24522);
nor UO_1764 (O_1764,N_24644,N_24782);
xnor UO_1765 (O_1765,N_24672,N_24732);
nand UO_1766 (O_1766,N_24771,N_24949);
and UO_1767 (O_1767,N_24899,N_24894);
nand UO_1768 (O_1768,N_24848,N_24657);
nor UO_1769 (O_1769,N_24581,N_24643);
and UO_1770 (O_1770,N_24631,N_24593);
and UO_1771 (O_1771,N_24511,N_24897);
or UO_1772 (O_1772,N_24638,N_24977);
and UO_1773 (O_1773,N_24567,N_24796);
nand UO_1774 (O_1774,N_24524,N_24708);
or UO_1775 (O_1775,N_24611,N_24767);
or UO_1776 (O_1776,N_24713,N_24565);
nand UO_1777 (O_1777,N_24904,N_24512);
nor UO_1778 (O_1778,N_24863,N_24524);
or UO_1779 (O_1779,N_24679,N_24509);
nand UO_1780 (O_1780,N_24656,N_24987);
or UO_1781 (O_1781,N_24853,N_24953);
nand UO_1782 (O_1782,N_24516,N_24815);
or UO_1783 (O_1783,N_24654,N_24787);
and UO_1784 (O_1784,N_24805,N_24826);
nor UO_1785 (O_1785,N_24589,N_24944);
nor UO_1786 (O_1786,N_24750,N_24952);
nor UO_1787 (O_1787,N_24927,N_24565);
or UO_1788 (O_1788,N_24960,N_24858);
or UO_1789 (O_1789,N_24739,N_24514);
and UO_1790 (O_1790,N_24859,N_24983);
nor UO_1791 (O_1791,N_24520,N_24894);
and UO_1792 (O_1792,N_24854,N_24650);
nand UO_1793 (O_1793,N_24614,N_24972);
and UO_1794 (O_1794,N_24693,N_24761);
or UO_1795 (O_1795,N_24782,N_24639);
and UO_1796 (O_1796,N_24567,N_24948);
nand UO_1797 (O_1797,N_24518,N_24651);
and UO_1798 (O_1798,N_24969,N_24641);
nor UO_1799 (O_1799,N_24531,N_24666);
xor UO_1800 (O_1800,N_24544,N_24909);
nor UO_1801 (O_1801,N_24999,N_24649);
nor UO_1802 (O_1802,N_24718,N_24728);
nand UO_1803 (O_1803,N_24777,N_24603);
or UO_1804 (O_1804,N_24747,N_24837);
nand UO_1805 (O_1805,N_24602,N_24581);
xnor UO_1806 (O_1806,N_24553,N_24805);
nand UO_1807 (O_1807,N_24645,N_24703);
nor UO_1808 (O_1808,N_24543,N_24734);
nand UO_1809 (O_1809,N_24594,N_24669);
and UO_1810 (O_1810,N_24766,N_24687);
nand UO_1811 (O_1811,N_24756,N_24828);
and UO_1812 (O_1812,N_24605,N_24980);
xnor UO_1813 (O_1813,N_24880,N_24873);
and UO_1814 (O_1814,N_24709,N_24588);
or UO_1815 (O_1815,N_24817,N_24649);
or UO_1816 (O_1816,N_24650,N_24664);
nand UO_1817 (O_1817,N_24895,N_24925);
or UO_1818 (O_1818,N_24921,N_24959);
or UO_1819 (O_1819,N_24515,N_24546);
and UO_1820 (O_1820,N_24774,N_24963);
and UO_1821 (O_1821,N_24648,N_24924);
nand UO_1822 (O_1822,N_24757,N_24995);
nor UO_1823 (O_1823,N_24906,N_24832);
nor UO_1824 (O_1824,N_24936,N_24621);
and UO_1825 (O_1825,N_24912,N_24797);
nor UO_1826 (O_1826,N_24623,N_24588);
nor UO_1827 (O_1827,N_24787,N_24815);
and UO_1828 (O_1828,N_24931,N_24875);
or UO_1829 (O_1829,N_24674,N_24779);
nand UO_1830 (O_1830,N_24552,N_24977);
or UO_1831 (O_1831,N_24655,N_24693);
nor UO_1832 (O_1832,N_24907,N_24769);
nor UO_1833 (O_1833,N_24724,N_24594);
xor UO_1834 (O_1834,N_24801,N_24820);
and UO_1835 (O_1835,N_24851,N_24617);
xor UO_1836 (O_1836,N_24784,N_24712);
or UO_1837 (O_1837,N_24502,N_24643);
and UO_1838 (O_1838,N_24873,N_24575);
nor UO_1839 (O_1839,N_24742,N_24614);
and UO_1840 (O_1840,N_24722,N_24795);
nor UO_1841 (O_1841,N_24650,N_24605);
and UO_1842 (O_1842,N_24946,N_24656);
and UO_1843 (O_1843,N_24689,N_24687);
or UO_1844 (O_1844,N_24588,N_24905);
nor UO_1845 (O_1845,N_24613,N_24907);
or UO_1846 (O_1846,N_24603,N_24649);
or UO_1847 (O_1847,N_24512,N_24852);
nor UO_1848 (O_1848,N_24765,N_24717);
or UO_1849 (O_1849,N_24566,N_24606);
or UO_1850 (O_1850,N_24854,N_24882);
nand UO_1851 (O_1851,N_24929,N_24810);
nor UO_1852 (O_1852,N_24743,N_24896);
or UO_1853 (O_1853,N_24716,N_24668);
nand UO_1854 (O_1854,N_24961,N_24993);
or UO_1855 (O_1855,N_24646,N_24706);
nand UO_1856 (O_1856,N_24978,N_24781);
xnor UO_1857 (O_1857,N_24721,N_24815);
nand UO_1858 (O_1858,N_24845,N_24688);
nor UO_1859 (O_1859,N_24941,N_24749);
xor UO_1860 (O_1860,N_24896,N_24618);
or UO_1861 (O_1861,N_24724,N_24940);
nor UO_1862 (O_1862,N_24743,N_24887);
or UO_1863 (O_1863,N_24923,N_24799);
nand UO_1864 (O_1864,N_24795,N_24917);
nor UO_1865 (O_1865,N_24982,N_24520);
xor UO_1866 (O_1866,N_24910,N_24920);
nor UO_1867 (O_1867,N_24673,N_24987);
or UO_1868 (O_1868,N_24611,N_24621);
nand UO_1869 (O_1869,N_24621,N_24771);
nand UO_1870 (O_1870,N_24953,N_24787);
or UO_1871 (O_1871,N_24903,N_24752);
and UO_1872 (O_1872,N_24765,N_24840);
and UO_1873 (O_1873,N_24742,N_24916);
nor UO_1874 (O_1874,N_24911,N_24526);
and UO_1875 (O_1875,N_24778,N_24920);
and UO_1876 (O_1876,N_24999,N_24870);
nand UO_1877 (O_1877,N_24968,N_24730);
nand UO_1878 (O_1878,N_24771,N_24807);
or UO_1879 (O_1879,N_24952,N_24566);
nand UO_1880 (O_1880,N_24525,N_24606);
and UO_1881 (O_1881,N_24970,N_24763);
or UO_1882 (O_1882,N_24552,N_24777);
nand UO_1883 (O_1883,N_24994,N_24909);
nand UO_1884 (O_1884,N_24969,N_24777);
or UO_1885 (O_1885,N_24561,N_24838);
nor UO_1886 (O_1886,N_24501,N_24855);
nand UO_1887 (O_1887,N_24874,N_24506);
or UO_1888 (O_1888,N_24752,N_24978);
and UO_1889 (O_1889,N_24731,N_24980);
nor UO_1890 (O_1890,N_24666,N_24500);
nand UO_1891 (O_1891,N_24727,N_24716);
nor UO_1892 (O_1892,N_24545,N_24875);
and UO_1893 (O_1893,N_24544,N_24932);
and UO_1894 (O_1894,N_24659,N_24635);
nand UO_1895 (O_1895,N_24912,N_24889);
or UO_1896 (O_1896,N_24743,N_24712);
nor UO_1897 (O_1897,N_24880,N_24814);
or UO_1898 (O_1898,N_24611,N_24889);
nand UO_1899 (O_1899,N_24958,N_24880);
and UO_1900 (O_1900,N_24923,N_24826);
and UO_1901 (O_1901,N_24635,N_24723);
nor UO_1902 (O_1902,N_24962,N_24984);
xor UO_1903 (O_1903,N_24910,N_24744);
nor UO_1904 (O_1904,N_24569,N_24613);
or UO_1905 (O_1905,N_24517,N_24807);
or UO_1906 (O_1906,N_24940,N_24834);
and UO_1907 (O_1907,N_24722,N_24788);
and UO_1908 (O_1908,N_24519,N_24711);
nand UO_1909 (O_1909,N_24678,N_24792);
and UO_1910 (O_1910,N_24811,N_24776);
nor UO_1911 (O_1911,N_24511,N_24917);
nor UO_1912 (O_1912,N_24833,N_24784);
nand UO_1913 (O_1913,N_24519,N_24797);
and UO_1914 (O_1914,N_24529,N_24681);
or UO_1915 (O_1915,N_24753,N_24830);
xor UO_1916 (O_1916,N_24700,N_24745);
and UO_1917 (O_1917,N_24707,N_24520);
nand UO_1918 (O_1918,N_24706,N_24663);
nor UO_1919 (O_1919,N_24546,N_24790);
nand UO_1920 (O_1920,N_24715,N_24744);
xnor UO_1921 (O_1921,N_24676,N_24610);
nand UO_1922 (O_1922,N_24628,N_24791);
or UO_1923 (O_1923,N_24639,N_24843);
nand UO_1924 (O_1924,N_24506,N_24606);
nor UO_1925 (O_1925,N_24938,N_24868);
or UO_1926 (O_1926,N_24608,N_24901);
nor UO_1927 (O_1927,N_24594,N_24896);
and UO_1928 (O_1928,N_24677,N_24904);
nor UO_1929 (O_1929,N_24926,N_24764);
nand UO_1930 (O_1930,N_24633,N_24743);
nor UO_1931 (O_1931,N_24764,N_24537);
nor UO_1932 (O_1932,N_24841,N_24514);
nand UO_1933 (O_1933,N_24701,N_24935);
xnor UO_1934 (O_1934,N_24630,N_24673);
xor UO_1935 (O_1935,N_24857,N_24589);
or UO_1936 (O_1936,N_24923,N_24945);
and UO_1937 (O_1937,N_24870,N_24766);
or UO_1938 (O_1938,N_24846,N_24923);
or UO_1939 (O_1939,N_24933,N_24589);
or UO_1940 (O_1940,N_24536,N_24973);
or UO_1941 (O_1941,N_24567,N_24727);
nor UO_1942 (O_1942,N_24617,N_24760);
nor UO_1943 (O_1943,N_24568,N_24755);
nor UO_1944 (O_1944,N_24871,N_24509);
nand UO_1945 (O_1945,N_24676,N_24526);
nand UO_1946 (O_1946,N_24822,N_24660);
or UO_1947 (O_1947,N_24790,N_24605);
and UO_1948 (O_1948,N_24507,N_24705);
nor UO_1949 (O_1949,N_24787,N_24687);
or UO_1950 (O_1950,N_24501,N_24760);
nand UO_1951 (O_1951,N_24736,N_24977);
and UO_1952 (O_1952,N_24760,N_24656);
or UO_1953 (O_1953,N_24897,N_24646);
nand UO_1954 (O_1954,N_24913,N_24944);
nand UO_1955 (O_1955,N_24916,N_24938);
and UO_1956 (O_1956,N_24795,N_24813);
xnor UO_1957 (O_1957,N_24841,N_24543);
and UO_1958 (O_1958,N_24731,N_24580);
nand UO_1959 (O_1959,N_24675,N_24930);
nand UO_1960 (O_1960,N_24815,N_24736);
nand UO_1961 (O_1961,N_24930,N_24582);
nand UO_1962 (O_1962,N_24947,N_24868);
nor UO_1963 (O_1963,N_24652,N_24879);
nor UO_1964 (O_1964,N_24845,N_24892);
nor UO_1965 (O_1965,N_24873,N_24858);
nand UO_1966 (O_1966,N_24550,N_24661);
nand UO_1967 (O_1967,N_24616,N_24801);
nor UO_1968 (O_1968,N_24518,N_24891);
nand UO_1969 (O_1969,N_24865,N_24638);
or UO_1970 (O_1970,N_24864,N_24780);
nor UO_1971 (O_1971,N_24798,N_24511);
and UO_1972 (O_1972,N_24844,N_24784);
and UO_1973 (O_1973,N_24700,N_24851);
nor UO_1974 (O_1974,N_24722,N_24697);
and UO_1975 (O_1975,N_24678,N_24848);
nand UO_1976 (O_1976,N_24616,N_24891);
and UO_1977 (O_1977,N_24679,N_24819);
or UO_1978 (O_1978,N_24805,N_24709);
or UO_1979 (O_1979,N_24527,N_24700);
nand UO_1980 (O_1980,N_24919,N_24917);
and UO_1981 (O_1981,N_24800,N_24625);
nor UO_1982 (O_1982,N_24701,N_24831);
or UO_1983 (O_1983,N_24536,N_24624);
and UO_1984 (O_1984,N_24563,N_24688);
or UO_1985 (O_1985,N_24834,N_24759);
nor UO_1986 (O_1986,N_24893,N_24534);
nor UO_1987 (O_1987,N_24531,N_24611);
and UO_1988 (O_1988,N_24840,N_24598);
and UO_1989 (O_1989,N_24955,N_24990);
and UO_1990 (O_1990,N_24768,N_24747);
or UO_1991 (O_1991,N_24999,N_24532);
or UO_1992 (O_1992,N_24912,N_24859);
xnor UO_1993 (O_1993,N_24563,N_24615);
nor UO_1994 (O_1994,N_24908,N_24985);
nor UO_1995 (O_1995,N_24776,N_24607);
nand UO_1996 (O_1996,N_24708,N_24848);
nor UO_1997 (O_1997,N_24516,N_24821);
nor UO_1998 (O_1998,N_24719,N_24836);
and UO_1999 (O_1999,N_24902,N_24791);
and UO_2000 (O_2000,N_24615,N_24889);
nor UO_2001 (O_2001,N_24668,N_24814);
and UO_2002 (O_2002,N_24605,N_24646);
nand UO_2003 (O_2003,N_24980,N_24860);
and UO_2004 (O_2004,N_24792,N_24829);
and UO_2005 (O_2005,N_24709,N_24547);
nand UO_2006 (O_2006,N_24507,N_24546);
nor UO_2007 (O_2007,N_24885,N_24757);
or UO_2008 (O_2008,N_24940,N_24791);
and UO_2009 (O_2009,N_24826,N_24957);
and UO_2010 (O_2010,N_24891,N_24560);
nor UO_2011 (O_2011,N_24501,N_24932);
or UO_2012 (O_2012,N_24935,N_24968);
or UO_2013 (O_2013,N_24862,N_24766);
or UO_2014 (O_2014,N_24597,N_24724);
nor UO_2015 (O_2015,N_24558,N_24850);
or UO_2016 (O_2016,N_24631,N_24936);
nor UO_2017 (O_2017,N_24654,N_24950);
and UO_2018 (O_2018,N_24914,N_24952);
or UO_2019 (O_2019,N_24669,N_24806);
or UO_2020 (O_2020,N_24634,N_24671);
or UO_2021 (O_2021,N_24695,N_24708);
and UO_2022 (O_2022,N_24528,N_24765);
and UO_2023 (O_2023,N_24774,N_24539);
nor UO_2024 (O_2024,N_24638,N_24949);
and UO_2025 (O_2025,N_24870,N_24691);
or UO_2026 (O_2026,N_24580,N_24625);
or UO_2027 (O_2027,N_24839,N_24576);
and UO_2028 (O_2028,N_24505,N_24998);
xor UO_2029 (O_2029,N_24966,N_24606);
nor UO_2030 (O_2030,N_24668,N_24916);
nor UO_2031 (O_2031,N_24624,N_24694);
nor UO_2032 (O_2032,N_24747,N_24917);
and UO_2033 (O_2033,N_24660,N_24815);
or UO_2034 (O_2034,N_24985,N_24848);
nand UO_2035 (O_2035,N_24939,N_24657);
nand UO_2036 (O_2036,N_24678,N_24756);
nand UO_2037 (O_2037,N_24515,N_24788);
and UO_2038 (O_2038,N_24770,N_24573);
nor UO_2039 (O_2039,N_24524,N_24933);
or UO_2040 (O_2040,N_24553,N_24787);
nand UO_2041 (O_2041,N_24506,N_24623);
nand UO_2042 (O_2042,N_24515,N_24911);
nand UO_2043 (O_2043,N_24746,N_24851);
and UO_2044 (O_2044,N_24575,N_24932);
or UO_2045 (O_2045,N_24919,N_24516);
or UO_2046 (O_2046,N_24517,N_24569);
nor UO_2047 (O_2047,N_24687,N_24818);
nand UO_2048 (O_2048,N_24869,N_24654);
or UO_2049 (O_2049,N_24852,N_24825);
or UO_2050 (O_2050,N_24798,N_24829);
nand UO_2051 (O_2051,N_24992,N_24821);
nor UO_2052 (O_2052,N_24777,N_24793);
nand UO_2053 (O_2053,N_24859,N_24869);
and UO_2054 (O_2054,N_24606,N_24642);
nand UO_2055 (O_2055,N_24834,N_24584);
nor UO_2056 (O_2056,N_24810,N_24591);
and UO_2057 (O_2057,N_24597,N_24618);
or UO_2058 (O_2058,N_24519,N_24549);
nand UO_2059 (O_2059,N_24837,N_24918);
and UO_2060 (O_2060,N_24754,N_24548);
and UO_2061 (O_2061,N_24772,N_24551);
and UO_2062 (O_2062,N_24931,N_24838);
nor UO_2063 (O_2063,N_24595,N_24564);
nor UO_2064 (O_2064,N_24883,N_24613);
nor UO_2065 (O_2065,N_24557,N_24957);
or UO_2066 (O_2066,N_24636,N_24607);
and UO_2067 (O_2067,N_24687,N_24514);
or UO_2068 (O_2068,N_24579,N_24897);
nor UO_2069 (O_2069,N_24961,N_24782);
nand UO_2070 (O_2070,N_24654,N_24860);
nor UO_2071 (O_2071,N_24904,N_24570);
and UO_2072 (O_2072,N_24969,N_24748);
nor UO_2073 (O_2073,N_24555,N_24977);
and UO_2074 (O_2074,N_24612,N_24831);
or UO_2075 (O_2075,N_24879,N_24705);
and UO_2076 (O_2076,N_24847,N_24773);
or UO_2077 (O_2077,N_24823,N_24590);
and UO_2078 (O_2078,N_24838,N_24717);
and UO_2079 (O_2079,N_24983,N_24813);
nand UO_2080 (O_2080,N_24671,N_24738);
nor UO_2081 (O_2081,N_24843,N_24675);
and UO_2082 (O_2082,N_24725,N_24683);
nand UO_2083 (O_2083,N_24850,N_24575);
or UO_2084 (O_2084,N_24791,N_24959);
or UO_2085 (O_2085,N_24673,N_24562);
or UO_2086 (O_2086,N_24607,N_24852);
nor UO_2087 (O_2087,N_24735,N_24894);
nand UO_2088 (O_2088,N_24721,N_24978);
or UO_2089 (O_2089,N_24785,N_24885);
nand UO_2090 (O_2090,N_24608,N_24862);
nand UO_2091 (O_2091,N_24506,N_24636);
nor UO_2092 (O_2092,N_24669,N_24907);
and UO_2093 (O_2093,N_24578,N_24893);
or UO_2094 (O_2094,N_24707,N_24843);
and UO_2095 (O_2095,N_24839,N_24883);
nor UO_2096 (O_2096,N_24707,N_24717);
xor UO_2097 (O_2097,N_24860,N_24829);
nor UO_2098 (O_2098,N_24532,N_24699);
nand UO_2099 (O_2099,N_24740,N_24533);
and UO_2100 (O_2100,N_24980,N_24543);
nand UO_2101 (O_2101,N_24552,N_24618);
nand UO_2102 (O_2102,N_24590,N_24719);
nand UO_2103 (O_2103,N_24664,N_24619);
nor UO_2104 (O_2104,N_24633,N_24511);
or UO_2105 (O_2105,N_24663,N_24683);
and UO_2106 (O_2106,N_24798,N_24631);
and UO_2107 (O_2107,N_24596,N_24926);
nand UO_2108 (O_2108,N_24994,N_24984);
nand UO_2109 (O_2109,N_24780,N_24955);
nor UO_2110 (O_2110,N_24509,N_24986);
nand UO_2111 (O_2111,N_24884,N_24975);
and UO_2112 (O_2112,N_24648,N_24598);
nor UO_2113 (O_2113,N_24600,N_24589);
and UO_2114 (O_2114,N_24647,N_24717);
nand UO_2115 (O_2115,N_24900,N_24578);
or UO_2116 (O_2116,N_24555,N_24942);
or UO_2117 (O_2117,N_24667,N_24501);
and UO_2118 (O_2118,N_24597,N_24877);
nor UO_2119 (O_2119,N_24544,N_24610);
nor UO_2120 (O_2120,N_24977,N_24528);
nor UO_2121 (O_2121,N_24697,N_24656);
and UO_2122 (O_2122,N_24965,N_24701);
and UO_2123 (O_2123,N_24998,N_24501);
nor UO_2124 (O_2124,N_24977,N_24588);
nor UO_2125 (O_2125,N_24772,N_24516);
nand UO_2126 (O_2126,N_24768,N_24697);
and UO_2127 (O_2127,N_24551,N_24585);
or UO_2128 (O_2128,N_24841,N_24779);
nor UO_2129 (O_2129,N_24924,N_24931);
or UO_2130 (O_2130,N_24911,N_24564);
nor UO_2131 (O_2131,N_24599,N_24717);
nand UO_2132 (O_2132,N_24825,N_24593);
or UO_2133 (O_2133,N_24887,N_24970);
or UO_2134 (O_2134,N_24616,N_24687);
or UO_2135 (O_2135,N_24655,N_24688);
nand UO_2136 (O_2136,N_24739,N_24529);
or UO_2137 (O_2137,N_24884,N_24554);
nor UO_2138 (O_2138,N_24629,N_24725);
or UO_2139 (O_2139,N_24542,N_24637);
and UO_2140 (O_2140,N_24702,N_24939);
or UO_2141 (O_2141,N_24573,N_24921);
or UO_2142 (O_2142,N_24759,N_24568);
and UO_2143 (O_2143,N_24542,N_24817);
nand UO_2144 (O_2144,N_24762,N_24918);
nor UO_2145 (O_2145,N_24540,N_24903);
nand UO_2146 (O_2146,N_24597,N_24954);
nand UO_2147 (O_2147,N_24502,N_24989);
xor UO_2148 (O_2148,N_24855,N_24997);
nand UO_2149 (O_2149,N_24900,N_24577);
nor UO_2150 (O_2150,N_24575,N_24520);
or UO_2151 (O_2151,N_24883,N_24628);
and UO_2152 (O_2152,N_24947,N_24661);
nor UO_2153 (O_2153,N_24930,N_24640);
nor UO_2154 (O_2154,N_24518,N_24534);
nor UO_2155 (O_2155,N_24595,N_24608);
and UO_2156 (O_2156,N_24691,N_24693);
or UO_2157 (O_2157,N_24838,N_24598);
nor UO_2158 (O_2158,N_24633,N_24773);
or UO_2159 (O_2159,N_24750,N_24743);
or UO_2160 (O_2160,N_24943,N_24777);
and UO_2161 (O_2161,N_24975,N_24920);
nand UO_2162 (O_2162,N_24756,N_24712);
or UO_2163 (O_2163,N_24829,N_24834);
and UO_2164 (O_2164,N_24917,N_24829);
and UO_2165 (O_2165,N_24991,N_24530);
and UO_2166 (O_2166,N_24926,N_24931);
xor UO_2167 (O_2167,N_24722,N_24681);
or UO_2168 (O_2168,N_24942,N_24920);
or UO_2169 (O_2169,N_24711,N_24645);
xor UO_2170 (O_2170,N_24669,N_24744);
nor UO_2171 (O_2171,N_24957,N_24908);
nand UO_2172 (O_2172,N_24540,N_24960);
or UO_2173 (O_2173,N_24817,N_24915);
nor UO_2174 (O_2174,N_24701,N_24784);
nand UO_2175 (O_2175,N_24580,N_24548);
and UO_2176 (O_2176,N_24597,N_24846);
nand UO_2177 (O_2177,N_24899,N_24508);
and UO_2178 (O_2178,N_24818,N_24974);
or UO_2179 (O_2179,N_24881,N_24523);
nand UO_2180 (O_2180,N_24877,N_24690);
and UO_2181 (O_2181,N_24625,N_24692);
or UO_2182 (O_2182,N_24817,N_24877);
or UO_2183 (O_2183,N_24826,N_24959);
nor UO_2184 (O_2184,N_24757,N_24791);
or UO_2185 (O_2185,N_24600,N_24739);
nor UO_2186 (O_2186,N_24503,N_24842);
and UO_2187 (O_2187,N_24626,N_24775);
nand UO_2188 (O_2188,N_24979,N_24546);
nand UO_2189 (O_2189,N_24673,N_24950);
nor UO_2190 (O_2190,N_24700,N_24645);
and UO_2191 (O_2191,N_24525,N_24873);
nand UO_2192 (O_2192,N_24799,N_24551);
or UO_2193 (O_2193,N_24686,N_24884);
xnor UO_2194 (O_2194,N_24797,N_24753);
nor UO_2195 (O_2195,N_24812,N_24823);
xnor UO_2196 (O_2196,N_24861,N_24571);
nand UO_2197 (O_2197,N_24662,N_24676);
nor UO_2198 (O_2198,N_24556,N_24963);
and UO_2199 (O_2199,N_24875,N_24719);
nor UO_2200 (O_2200,N_24846,N_24751);
or UO_2201 (O_2201,N_24903,N_24982);
or UO_2202 (O_2202,N_24556,N_24600);
nand UO_2203 (O_2203,N_24880,N_24568);
or UO_2204 (O_2204,N_24910,N_24534);
nor UO_2205 (O_2205,N_24877,N_24577);
nand UO_2206 (O_2206,N_24756,N_24785);
and UO_2207 (O_2207,N_24709,N_24959);
nand UO_2208 (O_2208,N_24758,N_24976);
nand UO_2209 (O_2209,N_24957,N_24646);
and UO_2210 (O_2210,N_24715,N_24712);
and UO_2211 (O_2211,N_24553,N_24900);
or UO_2212 (O_2212,N_24613,N_24876);
nand UO_2213 (O_2213,N_24936,N_24605);
nand UO_2214 (O_2214,N_24902,N_24846);
nand UO_2215 (O_2215,N_24950,N_24964);
nor UO_2216 (O_2216,N_24822,N_24598);
nand UO_2217 (O_2217,N_24758,N_24769);
and UO_2218 (O_2218,N_24551,N_24553);
nor UO_2219 (O_2219,N_24800,N_24774);
and UO_2220 (O_2220,N_24681,N_24655);
or UO_2221 (O_2221,N_24835,N_24868);
nand UO_2222 (O_2222,N_24972,N_24601);
or UO_2223 (O_2223,N_24688,N_24540);
nand UO_2224 (O_2224,N_24735,N_24891);
and UO_2225 (O_2225,N_24739,N_24575);
nor UO_2226 (O_2226,N_24695,N_24619);
nor UO_2227 (O_2227,N_24935,N_24905);
xnor UO_2228 (O_2228,N_24672,N_24648);
and UO_2229 (O_2229,N_24860,N_24758);
nor UO_2230 (O_2230,N_24700,N_24505);
nor UO_2231 (O_2231,N_24534,N_24867);
nand UO_2232 (O_2232,N_24568,N_24813);
and UO_2233 (O_2233,N_24768,N_24596);
nor UO_2234 (O_2234,N_24568,N_24971);
nand UO_2235 (O_2235,N_24653,N_24703);
nor UO_2236 (O_2236,N_24547,N_24604);
nor UO_2237 (O_2237,N_24891,N_24907);
or UO_2238 (O_2238,N_24893,N_24614);
nand UO_2239 (O_2239,N_24715,N_24749);
nor UO_2240 (O_2240,N_24851,N_24767);
nand UO_2241 (O_2241,N_24708,N_24877);
xor UO_2242 (O_2242,N_24830,N_24732);
or UO_2243 (O_2243,N_24831,N_24739);
or UO_2244 (O_2244,N_24994,N_24982);
nand UO_2245 (O_2245,N_24548,N_24938);
or UO_2246 (O_2246,N_24803,N_24837);
xnor UO_2247 (O_2247,N_24817,N_24813);
and UO_2248 (O_2248,N_24578,N_24539);
nor UO_2249 (O_2249,N_24608,N_24905);
nor UO_2250 (O_2250,N_24850,N_24980);
nor UO_2251 (O_2251,N_24701,N_24842);
nor UO_2252 (O_2252,N_24914,N_24775);
nand UO_2253 (O_2253,N_24779,N_24556);
or UO_2254 (O_2254,N_24700,N_24802);
nand UO_2255 (O_2255,N_24654,N_24521);
nand UO_2256 (O_2256,N_24893,N_24976);
nor UO_2257 (O_2257,N_24661,N_24754);
nor UO_2258 (O_2258,N_24555,N_24933);
nand UO_2259 (O_2259,N_24987,N_24678);
or UO_2260 (O_2260,N_24521,N_24620);
nand UO_2261 (O_2261,N_24576,N_24723);
nor UO_2262 (O_2262,N_24952,N_24695);
nor UO_2263 (O_2263,N_24504,N_24519);
nand UO_2264 (O_2264,N_24788,N_24597);
and UO_2265 (O_2265,N_24795,N_24901);
and UO_2266 (O_2266,N_24675,N_24968);
nand UO_2267 (O_2267,N_24603,N_24936);
nor UO_2268 (O_2268,N_24972,N_24762);
nand UO_2269 (O_2269,N_24753,N_24976);
and UO_2270 (O_2270,N_24972,N_24917);
nand UO_2271 (O_2271,N_24872,N_24537);
nor UO_2272 (O_2272,N_24811,N_24646);
nand UO_2273 (O_2273,N_24938,N_24891);
nor UO_2274 (O_2274,N_24871,N_24628);
and UO_2275 (O_2275,N_24840,N_24635);
or UO_2276 (O_2276,N_24956,N_24803);
and UO_2277 (O_2277,N_24684,N_24939);
and UO_2278 (O_2278,N_24713,N_24907);
nor UO_2279 (O_2279,N_24609,N_24928);
nor UO_2280 (O_2280,N_24822,N_24834);
or UO_2281 (O_2281,N_24520,N_24961);
and UO_2282 (O_2282,N_24984,N_24702);
nand UO_2283 (O_2283,N_24998,N_24919);
nand UO_2284 (O_2284,N_24514,N_24547);
and UO_2285 (O_2285,N_24887,N_24696);
or UO_2286 (O_2286,N_24544,N_24607);
and UO_2287 (O_2287,N_24978,N_24636);
or UO_2288 (O_2288,N_24985,N_24613);
and UO_2289 (O_2289,N_24806,N_24837);
nor UO_2290 (O_2290,N_24915,N_24774);
or UO_2291 (O_2291,N_24879,N_24949);
nand UO_2292 (O_2292,N_24801,N_24909);
nand UO_2293 (O_2293,N_24996,N_24981);
xnor UO_2294 (O_2294,N_24838,N_24788);
nand UO_2295 (O_2295,N_24864,N_24961);
or UO_2296 (O_2296,N_24927,N_24886);
nand UO_2297 (O_2297,N_24790,N_24735);
or UO_2298 (O_2298,N_24999,N_24783);
or UO_2299 (O_2299,N_24962,N_24874);
nor UO_2300 (O_2300,N_24971,N_24649);
nand UO_2301 (O_2301,N_24907,N_24874);
and UO_2302 (O_2302,N_24864,N_24906);
and UO_2303 (O_2303,N_24500,N_24677);
nor UO_2304 (O_2304,N_24723,N_24616);
nor UO_2305 (O_2305,N_24961,N_24802);
and UO_2306 (O_2306,N_24631,N_24841);
nand UO_2307 (O_2307,N_24996,N_24528);
nand UO_2308 (O_2308,N_24698,N_24886);
or UO_2309 (O_2309,N_24621,N_24848);
or UO_2310 (O_2310,N_24846,N_24668);
nand UO_2311 (O_2311,N_24984,N_24550);
nand UO_2312 (O_2312,N_24852,N_24510);
nor UO_2313 (O_2313,N_24800,N_24934);
nor UO_2314 (O_2314,N_24931,N_24714);
nor UO_2315 (O_2315,N_24909,N_24820);
or UO_2316 (O_2316,N_24624,N_24802);
and UO_2317 (O_2317,N_24858,N_24572);
nand UO_2318 (O_2318,N_24524,N_24587);
nand UO_2319 (O_2319,N_24777,N_24816);
and UO_2320 (O_2320,N_24734,N_24676);
xor UO_2321 (O_2321,N_24712,N_24818);
or UO_2322 (O_2322,N_24805,N_24872);
nand UO_2323 (O_2323,N_24919,N_24641);
or UO_2324 (O_2324,N_24836,N_24767);
nor UO_2325 (O_2325,N_24911,N_24719);
nand UO_2326 (O_2326,N_24841,N_24961);
or UO_2327 (O_2327,N_24629,N_24554);
nor UO_2328 (O_2328,N_24948,N_24966);
and UO_2329 (O_2329,N_24912,N_24720);
and UO_2330 (O_2330,N_24698,N_24644);
nand UO_2331 (O_2331,N_24598,N_24849);
nor UO_2332 (O_2332,N_24770,N_24973);
nor UO_2333 (O_2333,N_24919,N_24861);
nand UO_2334 (O_2334,N_24628,N_24828);
or UO_2335 (O_2335,N_24759,N_24890);
xor UO_2336 (O_2336,N_24995,N_24786);
nor UO_2337 (O_2337,N_24712,N_24916);
nor UO_2338 (O_2338,N_24681,N_24991);
or UO_2339 (O_2339,N_24527,N_24982);
nor UO_2340 (O_2340,N_24861,N_24804);
or UO_2341 (O_2341,N_24715,N_24532);
xor UO_2342 (O_2342,N_24924,N_24788);
and UO_2343 (O_2343,N_24731,N_24937);
nor UO_2344 (O_2344,N_24526,N_24809);
nor UO_2345 (O_2345,N_24541,N_24645);
nor UO_2346 (O_2346,N_24875,N_24591);
or UO_2347 (O_2347,N_24915,N_24957);
nor UO_2348 (O_2348,N_24953,N_24894);
or UO_2349 (O_2349,N_24575,N_24983);
nand UO_2350 (O_2350,N_24776,N_24941);
nor UO_2351 (O_2351,N_24520,N_24873);
or UO_2352 (O_2352,N_24749,N_24506);
and UO_2353 (O_2353,N_24517,N_24692);
nor UO_2354 (O_2354,N_24868,N_24637);
nand UO_2355 (O_2355,N_24538,N_24916);
nand UO_2356 (O_2356,N_24576,N_24757);
nand UO_2357 (O_2357,N_24553,N_24592);
nand UO_2358 (O_2358,N_24511,N_24695);
or UO_2359 (O_2359,N_24851,N_24833);
nor UO_2360 (O_2360,N_24577,N_24591);
or UO_2361 (O_2361,N_24700,N_24875);
nand UO_2362 (O_2362,N_24567,N_24672);
and UO_2363 (O_2363,N_24798,N_24849);
nor UO_2364 (O_2364,N_24990,N_24555);
or UO_2365 (O_2365,N_24876,N_24960);
nor UO_2366 (O_2366,N_24622,N_24564);
and UO_2367 (O_2367,N_24590,N_24652);
nor UO_2368 (O_2368,N_24950,N_24784);
nor UO_2369 (O_2369,N_24726,N_24906);
and UO_2370 (O_2370,N_24954,N_24665);
and UO_2371 (O_2371,N_24794,N_24985);
nand UO_2372 (O_2372,N_24907,N_24668);
and UO_2373 (O_2373,N_24514,N_24929);
and UO_2374 (O_2374,N_24577,N_24642);
nor UO_2375 (O_2375,N_24660,N_24752);
nor UO_2376 (O_2376,N_24595,N_24558);
and UO_2377 (O_2377,N_24612,N_24778);
or UO_2378 (O_2378,N_24837,N_24542);
or UO_2379 (O_2379,N_24669,N_24547);
or UO_2380 (O_2380,N_24826,N_24709);
and UO_2381 (O_2381,N_24815,N_24863);
and UO_2382 (O_2382,N_24779,N_24909);
and UO_2383 (O_2383,N_24756,N_24567);
nand UO_2384 (O_2384,N_24761,N_24678);
and UO_2385 (O_2385,N_24573,N_24989);
or UO_2386 (O_2386,N_24843,N_24534);
xor UO_2387 (O_2387,N_24925,N_24644);
nor UO_2388 (O_2388,N_24540,N_24653);
nor UO_2389 (O_2389,N_24529,N_24765);
and UO_2390 (O_2390,N_24990,N_24654);
xnor UO_2391 (O_2391,N_24826,N_24639);
nor UO_2392 (O_2392,N_24805,N_24747);
nor UO_2393 (O_2393,N_24783,N_24864);
nor UO_2394 (O_2394,N_24537,N_24876);
and UO_2395 (O_2395,N_24879,N_24902);
nand UO_2396 (O_2396,N_24915,N_24945);
nor UO_2397 (O_2397,N_24724,N_24955);
nand UO_2398 (O_2398,N_24943,N_24870);
and UO_2399 (O_2399,N_24599,N_24939);
or UO_2400 (O_2400,N_24532,N_24857);
nand UO_2401 (O_2401,N_24654,N_24679);
nand UO_2402 (O_2402,N_24546,N_24839);
xor UO_2403 (O_2403,N_24714,N_24545);
nand UO_2404 (O_2404,N_24967,N_24798);
and UO_2405 (O_2405,N_24846,N_24669);
nor UO_2406 (O_2406,N_24756,N_24999);
or UO_2407 (O_2407,N_24888,N_24949);
and UO_2408 (O_2408,N_24537,N_24916);
nor UO_2409 (O_2409,N_24957,N_24535);
and UO_2410 (O_2410,N_24592,N_24608);
nand UO_2411 (O_2411,N_24625,N_24588);
and UO_2412 (O_2412,N_24619,N_24723);
or UO_2413 (O_2413,N_24540,N_24767);
or UO_2414 (O_2414,N_24550,N_24949);
nand UO_2415 (O_2415,N_24816,N_24806);
or UO_2416 (O_2416,N_24546,N_24846);
nand UO_2417 (O_2417,N_24959,N_24682);
or UO_2418 (O_2418,N_24772,N_24526);
or UO_2419 (O_2419,N_24663,N_24775);
nand UO_2420 (O_2420,N_24949,N_24853);
and UO_2421 (O_2421,N_24941,N_24917);
and UO_2422 (O_2422,N_24798,N_24544);
xnor UO_2423 (O_2423,N_24780,N_24710);
or UO_2424 (O_2424,N_24966,N_24654);
nand UO_2425 (O_2425,N_24856,N_24715);
nand UO_2426 (O_2426,N_24997,N_24603);
nand UO_2427 (O_2427,N_24755,N_24721);
nand UO_2428 (O_2428,N_24566,N_24761);
nor UO_2429 (O_2429,N_24991,N_24561);
or UO_2430 (O_2430,N_24708,N_24501);
nand UO_2431 (O_2431,N_24823,N_24918);
nor UO_2432 (O_2432,N_24850,N_24785);
nand UO_2433 (O_2433,N_24685,N_24925);
or UO_2434 (O_2434,N_24622,N_24669);
nand UO_2435 (O_2435,N_24845,N_24647);
or UO_2436 (O_2436,N_24847,N_24974);
and UO_2437 (O_2437,N_24882,N_24508);
or UO_2438 (O_2438,N_24994,N_24757);
nor UO_2439 (O_2439,N_24673,N_24690);
or UO_2440 (O_2440,N_24994,N_24725);
nand UO_2441 (O_2441,N_24851,N_24676);
and UO_2442 (O_2442,N_24871,N_24541);
xnor UO_2443 (O_2443,N_24756,N_24735);
xnor UO_2444 (O_2444,N_24665,N_24561);
nand UO_2445 (O_2445,N_24951,N_24520);
and UO_2446 (O_2446,N_24929,N_24642);
nor UO_2447 (O_2447,N_24744,N_24503);
or UO_2448 (O_2448,N_24784,N_24770);
or UO_2449 (O_2449,N_24681,N_24975);
and UO_2450 (O_2450,N_24907,N_24672);
and UO_2451 (O_2451,N_24544,N_24786);
nand UO_2452 (O_2452,N_24547,N_24922);
and UO_2453 (O_2453,N_24768,N_24977);
nand UO_2454 (O_2454,N_24571,N_24893);
xor UO_2455 (O_2455,N_24586,N_24908);
or UO_2456 (O_2456,N_24672,N_24968);
nor UO_2457 (O_2457,N_24962,N_24753);
or UO_2458 (O_2458,N_24736,N_24860);
or UO_2459 (O_2459,N_24778,N_24856);
or UO_2460 (O_2460,N_24788,N_24738);
nand UO_2461 (O_2461,N_24938,N_24909);
nor UO_2462 (O_2462,N_24838,N_24821);
xor UO_2463 (O_2463,N_24866,N_24951);
nor UO_2464 (O_2464,N_24652,N_24940);
and UO_2465 (O_2465,N_24738,N_24545);
or UO_2466 (O_2466,N_24902,N_24738);
or UO_2467 (O_2467,N_24853,N_24781);
and UO_2468 (O_2468,N_24726,N_24995);
nand UO_2469 (O_2469,N_24989,N_24747);
or UO_2470 (O_2470,N_24873,N_24643);
nor UO_2471 (O_2471,N_24733,N_24871);
nor UO_2472 (O_2472,N_24638,N_24984);
or UO_2473 (O_2473,N_24933,N_24993);
nor UO_2474 (O_2474,N_24581,N_24823);
or UO_2475 (O_2475,N_24780,N_24623);
and UO_2476 (O_2476,N_24910,N_24565);
and UO_2477 (O_2477,N_24741,N_24765);
and UO_2478 (O_2478,N_24573,N_24724);
nand UO_2479 (O_2479,N_24827,N_24993);
nor UO_2480 (O_2480,N_24541,N_24948);
and UO_2481 (O_2481,N_24919,N_24642);
nand UO_2482 (O_2482,N_24660,N_24749);
nor UO_2483 (O_2483,N_24519,N_24978);
or UO_2484 (O_2484,N_24872,N_24757);
nand UO_2485 (O_2485,N_24773,N_24590);
or UO_2486 (O_2486,N_24817,N_24688);
nor UO_2487 (O_2487,N_24800,N_24666);
nor UO_2488 (O_2488,N_24916,N_24508);
nor UO_2489 (O_2489,N_24952,N_24603);
or UO_2490 (O_2490,N_24941,N_24804);
and UO_2491 (O_2491,N_24905,N_24893);
or UO_2492 (O_2492,N_24626,N_24686);
or UO_2493 (O_2493,N_24931,N_24872);
and UO_2494 (O_2494,N_24626,N_24576);
or UO_2495 (O_2495,N_24746,N_24957);
nand UO_2496 (O_2496,N_24713,N_24935);
or UO_2497 (O_2497,N_24997,N_24805);
nor UO_2498 (O_2498,N_24845,N_24690);
nor UO_2499 (O_2499,N_24817,N_24608);
nand UO_2500 (O_2500,N_24826,N_24825);
nor UO_2501 (O_2501,N_24746,N_24626);
nand UO_2502 (O_2502,N_24566,N_24860);
nand UO_2503 (O_2503,N_24782,N_24789);
and UO_2504 (O_2504,N_24701,N_24812);
or UO_2505 (O_2505,N_24613,N_24599);
and UO_2506 (O_2506,N_24633,N_24845);
and UO_2507 (O_2507,N_24567,N_24811);
and UO_2508 (O_2508,N_24698,N_24785);
or UO_2509 (O_2509,N_24507,N_24768);
nand UO_2510 (O_2510,N_24652,N_24541);
nand UO_2511 (O_2511,N_24850,N_24699);
or UO_2512 (O_2512,N_24695,N_24976);
nand UO_2513 (O_2513,N_24557,N_24604);
or UO_2514 (O_2514,N_24790,N_24920);
nor UO_2515 (O_2515,N_24898,N_24645);
nand UO_2516 (O_2516,N_24557,N_24746);
and UO_2517 (O_2517,N_24795,N_24537);
or UO_2518 (O_2518,N_24938,N_24674);
and UO_2519 (O_2519,N_24898,N_24821);
or UO_2520 (O_2520,N_24979,N_24618);
and UO_2521 (O_2521,N_24656,N_24764);
nand UO_2522 (O_2522,N_24511,N_24707);
nor UO_2523 (O_2523,N_24864,N_24786);
nand UO_2524 (O_2524,N_24557,N_24810);
and UO_2525 (O_2525,N_24733,N_24615);
nor UO_2526 (O_2526,N_24994,N_24501);
nor UO_2527 (O_2527,N_24501,N_24567);
or UO_2528 (O_2528,N_24917,N_24903);
or UO_2529 (O_2529,N_24692,N_24709);
and UO_2530 (O_2530,N_24826,N_24946);
or UO_2531 (O_2531,N_24589,N_24958);
or UO_2532 (O_2532,N_24726,N_24564);
and UO_2533 (O_2533,N_24798,N_24510);
nand UO_2534 (O_2534,N_24566,N_24601);
nor UO_2535 (O_2535,N_24841,N_24756);
xor UO_2536 (O_2536,N_24517,N_24500);
nor UO_2537 (O_2537,N_24828,N_24842);
nand UO_2538 (O_2538,N_24883,N_24543);
nand UO_2539 (O_2539,N_24941,N_24760);
nand UO_2540 (O_2540,N_24562,N_24717);
and UO_2541 (O_2541,N_24666,N_24656);
xor UO_2542 (O_2542,N_24980,N_24591);
nand UO_2543 (O_2543,N_24943,N_24505);
nor UO_2544 (O_2544,N_24819,N_24887);
nand UO_2545 (O_2545,N_24814,N_24556);
nand UO_2546 (O_2546,N_24566,N_24705);
and UO_2547 (O_2547,N_24635,N_24936);
or UO_2548 (O_2548,N_24977,N_24897);
and UO_2549 (O_2549,N_24526,N_24775);
nor UO_2550 (O_2550,N_24723,N_24671);
and UO_2551 (O_2551,N_24930,N_24595);
nand UO_2552 (O_2552,N_24758,N_24894);
or UO_2553 (O_2553,N_24818,N_24982);
or UO_2554 (O_2554,N_24939,N_24624);
nand UO_2555 (O_2555,N_24606,N_24758);
nor UO_2556 (O_2556,N_24975,N_24781);
nand UO_2557 (O_2557,N_24995,N_24850);
nand UO_2558 (O_2558,N_24841,N_24531);
nand UO_2559 (O_2559,N_24610,N_24662);
or UO_2560 (O_2560,N_24726,N_24522);
or UO_2561 (O_2561,N_24643,N_24514);
and UO_2562 (O_2562,N_24750,N_24670);
or UO_2563 (O_2563,N_24533,N_24821);
nor UO_2564 (O_2564,N_24606,N_24903);
and UO_2565 (O_2565,N_24927,N_24520);
and UO_2566 (O_2566,N_24839,N_24627);
or UO_2567 (O_2567,N_24940,N_24907);
nand UO_2568 (O_2568,N_24875,N_24717);
nand UO_2569 (O_2569,N_24887,N_24858);
or UO_2570 (O_2570,N_24964,N_24693);
nor UO_2571 (O_2571,N_24659,N_24636);
and UO_2572 (O_2572,N_24952,N_24599);
xor UO_2573 (O_2573,N_24861,N_24618);
nand UO_2574 (O_2574,N_24792,N_24626);
nand UO_2575 (O_2575,N_24578,N_24627);
nand UO_2576 (O_2576,N_24863,N_24813);
nor UO_2577 (O_2577,N_24578,N_24645);
nand UO_2578 (O_2578,N_24610,N_24563);
nor UO_2579 (O_2579,N_24927,N_24654);
nand UO_2580 (O_2580,N_24900,N_24558);
or UO_2581 (O_2581,N_24511,N_24682);
or UO_2582 (O_2582,N_24900,N_24704);
nor UO_2583 (O_2583,N_24864,N_24589);
or UO_2584 (O_2584,N_24536,N_24977);
nor UO_2585 (O_2585,N_24967,N_24816);
or UO_2586 (O_2586,N_24514,N_24642);
nand UO_2587 (O_2587,N_24979,N_24859);
and UO_2588 (O_2588,N_24855,N_24596);
or UO_2589 (O_2589,N_24697,N_24724);
nor UO_2590 (O_2590,N_24638,N_24802);
or UO_2591 (O_2591,N_24891,N_24720);
and UO_2592 (O_2592,N_24916,N_24767);
nand UO_2593 (O_2593,N_24908,N_24615);
or UO_2594 (O_2594,N_24815,N_24784);
or UO_2595 (O_2595,N_24804,N_24797);
xnor UO_2596 (O_2596,N_24624,N_24815);
nand UO_2597 (O_2597,N_24701,N_24665);
xnor UO_2598 (O_2598,N_24790,N_24706);
or UO_2599 (O_2599,N_24768,N_24824);
nor UO_2600 (O_2600,N_24971,N_24931);
or UO_2601 (O_2601,N_24566,N_24942);
and UO_2602 (O_2602,N_24749,N_24557);
nor UO_2603 (O_2603,N_24903,N_24516);
nand UO_2604 (O_2604,N_24858,N_24693);
or UO_2605 (O_2605,N_24772,N_24833);
or UO_2606 (O_2606,N_24591,N_24544);
nor UO_2607 (O_2607,N_24880,N_24993);
nand UO_2608 (O_2608,N_24716,N_24855);
nand UO_2609 (O_2609,N_24843,N_24965);
nor UO_2610 (O_2610,N_24694,N_24522);
nor UO_2611 (O_2611,N_24664,N_24903);
nor UO_2612 (O_2612,N_24906,N_24910);
nand UO_2613 (O_2613,N_24769,N_24902);
or UO_2614 (O_2614,N_24720,N_24825);
or UO_2615 (O_2615,N_24563,N_24579);
and UO_2616 (O_2616,N_24674,N_24907);
nand UO_2617 (O_2617,N_24758,N_24664);
or UO_2618 (O_2618,N_24641,N_24880);
nand UO_2619 (O_2619,N_24685,N_24597);
nor UO_2620 (O_2620,N_24772,N_24674);
nor UO_2621 (O_2621,N_24827,N_24629);
xnor UO_2622 (O_2622,N_24974,N_24976);
or UO_2623 (O_2623,N_24788,N_24616);
nor UO_2624 (O_2624,N_24920,N_24857);
and UO_2625 (O_2625,N_24546,N_24964);
and UO_2626 (O_2626,N_24821,N_24594);
or UO_2627 (O_2627,N_24991,N_24772);
or UO_2628 (O_2628,N_24798,N_24720);
nor UO_2629 (O_2629,N_24995,N_24698);
or UO_2630 (O_2630,N_24833,N_24915);
or UO_2631 (O_2631,N_24675,N_24797);
or UO_2632 (O_2632,N_24571,N_24670);
or UO_2633 (O_2633,N_24735,N_24952);
or UO_2634 (O_2634,N_24692,N_24898);
nand UO_2635 (O_2635,N_24519,N_24688);
nor UO_2636 (O_2636,N_24892,N_24507);
or UO_2637 (O_2637,N_24784,N_24676);
or UO_2638 (O_2638,N_24961,N_24788);
nor UO_2639 (O_2639,N_24528,N_24580);
nor UO_2640 (O_2640,N_24709,N_24835);
nor UO_2641 (O_2641,N_24650,N_24832);
nor UO_2642 (O_2642,N_24837,N_24779);
and UO_2643 (O_2643,N_24692,N_24675);
nor UO_2644 (O_2644,N_24576,N_24528);
and UO_2645 (O_2645,N_24733,N_24834);
and UO_2646 (O_2646,N_24783,N_24983);
nand UO_2647 (O_2647,N_24870,N_24653);
or UO_2648 (O_2648,N_24691,N_24904);
nand UO_2649 (O_2649,N_24884,N_24618);
nand UO_2650 (O_2650,N_24717,N_24502);
and UO_2651 (O_2651,N_24791,N_24784);
xnor UO_2652 (O_2652,N_24536,N_24918);
nand UO_2653 (O_2653,N_24800,N_24569);
or UO_2654 (O_2654,N_24828,N_24768);
nor UO_2655 (O_2655,N_24808,N_24827);
and UO_2656 (O_2656,N_24863,N_24957);
or UO_2657 (O_2657,N_24664,N_24877);
nand UO_2658 (O_2658,N_24718,N_24831);
or UO_2659 (O_2659,N_24678,N_24755);
and UO_2660 (O_2660,N_24601,N_24733);
xor UO_2661 (O_2661,N_24678,N_24918);
and UO_2662 (O_2662,N_24955,N_24738);
nor UO_2663 (O_2663,N_24567,N_24755);
and UO_2664 (O_2664,N_24726,N_24973);
nand UO_2665 (O_2665,N_24850,N_24705);
nand UO_2666 (O_2666,N_24560,N_24757);
nand UO_2667 (O_2667,N_24832,N_24743);
and UO_2668 (O_2668,N_24642,N_24761);
or UO_2669 (O_2669,N_24947,N_24575);
or UO_2670 (O_2670,N_24891,N_24915);
nor UO_2671 (O_2671,N_24693,N_24829);
xor UO_2672 (O_2672,N_24955,N_24567);
nand UO_2673 (O_2673,N_24659,N_24995);
nand UO_2674 (O_2674,N_24992,N_24885);
or UO_2675 (O_2675,N_24810,N_24864);
and UO_2676 (O_2676,N_24674,N_24512);
or UO_2677 (O_2677,N_24629,N_24701);
nor UO_2678 (O_2678,N_24617,N_24722);
or UO_2679 (O_2679,N_24884,N_24925);
or UO_2680 (O_2680,N_24823,N_24624);
and UO_2681 (O_2681,N_24553,N_24647);
or UO_2682 (O_2682,N_24852,N_24897);
and UO_2683 (O_2683,N_24633,N_24948);
xnor UO_2684 (O_2684,N_24997,N_24903);
xnor UO_2685 (O_2685,N_24776,N_24757);
nor UO_2686 (O_2686,N_24992,N_24621);
and UO_2687 (O_2687,N_24787,N_24781);
or UO_2688 (O_2688,N_24808,N_24817);
nor UO_2689 (O_2689,N_24576,N_24811);
and UO_2690 (O_2690,N_24742,N_24810);
nor UO_2691 (O_2691,N_24924,N_24826);
and UO_2692 (O_2692,N_24648,N_24889);
nor UO_2693 (O_2693,N_24503,N_24616);
nor UO_2694 (O_2694,N_24710,N_24540);
nor UO_2695 (O_2695,N_24576,N_24805);
xor UO_2696 (O_2696,N_24595,N_24738);
and UO_2697 (O_2697,N_24844,N_24710);
and UO_2698 (O_2698,N_24560,N_24905);
and UO_2699 (O_2699,N_24873,N_24508);
and UO_2700 (O_2700,N_24969,N_24847);
nand UO_2701 (O_2701,N_24854,N_24772);
or UO_2702 (O_2702,N_24772,N_24500);
and UO_2703 (O_2703,N_24831,N_24705);
or UO_2704 (O_2704,N_24682,N_24754);
nand UO_2705 (O_2705,N_24551,N_24515);
nand UO_2706 (O_2706,N_24796,N_24732);
nor UO_2707 (O_2707,N_24677,N_24744);
nand UO_2708 (O_2708,N_24628,N_24536);
nand UO_2709 (O_2709,N_24567,N_24898);
xor UO_2710 (O_2710,N_24734,N_24787);
or UO_2711 (O_2711,N_24746,N_24879);
nand UO_2712 (O_2712,N_24953,N_24552);
nand UO_2713 (O_2713,N_24979,N_24901);
or UO_2714 (O_2714,N_24579,N_24590);
nor UO_2715 (O_2715,N_24950,N_24786);
nand UO_2716 (O_2716,N_24787,N_24638);
nor UO_2717 (O_2717,N_24844,N_24847);
xor UO_2718 (O_2718,N_24723,N_24844);
and UO_2719 (O_2719,N_24605,N_24676);
and UO_2720 (O_2720,N_24588,N_24632);
or UO_2721 (O_2721,N_24893,N_24711);
and UO_2722 (O_2722,N_24911,N_24575);
or UO_2723 (O_2723,N_24743,N_24545);
nand UO_2724 (O_2724,N_24699,N_24647);
nand UO_2725 (O_2725,N_24600,N_24856);
or UO_2726 (O_2726,N_24811,N_24625);
nor UO_2727 (O_2727,N_24953,N_24803);
nand UO_2728 (O_2728,N_24982,N_24913);
and UO_2729 (O_2729,N_24721,N_24970);
or UO_2730 (O_2730,N_24878,N_24868);
and UO_2731 (O_2731,N_24825,N_24933);
nor UO_2732 (O_2732,N_24943,N_24508);
nand UO_2733 (O_2733,N_24973,N_24815);
and UO_2734 (O_2734,N_24735,N_24896);
nor UO_2735 (O_2735,N_24920,N_24990);
or UO_2736 (O_2736,N_24924,N_24582);
nand UO_2737 (O_2737,N_24945,N_24815);
nand UO_2738 (O_2738,N_24619,N_24582);
nand UO_2739 (O_2739,N_24543,N_24902);
nor UO_2740 (O_2740,N_24811,N_24622);
nor UO_2741 (O_2741,N_24623,N_24613);
nand UO_2742 (O_2742,N_24632,N_24987);
and UO_2743 (O_2743,N_24877,N_24588);
and UO_2744 (O_2744,N_24947,N_24738);
or UO_2745 (O_2745,N_24797,N_24784);
and UO_2746 (O_2746,N_24835,N_24979);
nand UO_2747 (O_2747,N_24918,N_24572);
and UO_2748 (O_2748,N_24851,N_24843);
nor UO_2749 (O_2749,N_24802,N_24654);
nand UO_2750 (O_2750,N_24797,N_24717);
and UO_2751 (O_2751,N_24745,N_24524);
nor UO_2752 (O_2752,N_24854,N_24660);
nand UO_2753 (O_2753,N_24994,N_24758);
or UO_2754 (O_2754,N_24946,N_24516);
nand UO_2755 (O_2755,N_24558,N_24996);
nand UO_2756 (O_2756,N_24631,N_24719);
or UO_2757 (O_2757,N_24834,N_24984);
and UO_2758 (O_2758,N_24882,N_24552);
or UO_2759 (O_2759,N_24515,N_24647);
nor UO_2760 (O_2760,N_24566,N_24936);
nand UO_2761 (O_2761,N_24992,N_24852);
and UO_2762 (O_2762,N_24643,N_24994);
or UO_2763 (O_2763,N_24568,N_24891);
nand UO_2764 (O_2764,N_24689,N_24774);
or UO_2765 (O_2765,N_24616,N_24929);
nor UO_2766 (O_2766,N_24724,N_24686);
and UO_2767 (O_2767,N_24589,N_24737);
and UO_2768 (O_2768,N_24575,N_24829);
and UO_2769 (O_2769,N_24509,N_24898);
and UO_2770 (O_2770,N_24726,N_24677);
nand UO_2771 (O_2771,N_24879,N_24608);
nand UO_2772 (O_2772,N_24966,N_24883);
nor UO_2773 (O_2773,N_24575,N_24927);
nor UO_2774 (O_2774,N_24915,N_24629);
nand UO_2775 (O_2775,N_24976,N_24560);
and UO_2776 (O_2776,N_24950,N_24981);
and UO_2777 (O_2777,N_24550,N_24784);
or UO_2778 (O_2778,N_24570,N_24501);
nand UO_2779 (O_2779,N_24967,N_24500);
nand UO_2780 (O_2780,N_24905,N_24682);
nand UO_2781 (O_2781,N_24674,N_24958);
nand UO_2782 (O_2782,N_24952,N_24942);
nand UO_2783 (O_2783,N_24985,N_24832);
or UO_2784 (O_2784,N_24908,N_24975);
or UO_2785 (O_2785,N_24981,N_24968);
and UO_2786 (O_2786,N_24648,N_24542);
nand UO_2787 (O_2787,N_24648,N_24649);
and UO_2788 (O_2788,N_24668,N_24506);
nor UO_2789 (O_2789,N_24960,N_24670);
or UO_2790 (O_2790,N_24540,N_24735);
nand UO_2791 (O_2791,N_24531,N_24712);
or UO_2792 (O_2792,N_24904,N_24536);
nand UO_2793 (O_2793,N_24539,N_24895);
or UO_2794 (O_2794,N_24628,N_24627);
or UO_2795 (O_2795,N_24778,N_24897);
and UO_2796 (O_2796,N_24539,N_24571);
and UO_2797 (O_2797,N_24888,N_24928);
and UO_2798 (O_2798,N_24580,N_24848);
and UO_2799 (O_2799,N_24580,N_24518);
nor UO_2800 (O_2800,N_24984,N_24876);
nand UO_2801 (O_2801,N_24885,N_24980);
and UO_2802 (O_2802,N_24767,N_24725);
and UO_2803 (O_2803,N_24878,N_24623);
or UO_2804 (O_2804,N_24574,N_24772);
nand UO_2805 (O_2805,N_24581,N_24707);
nand UO_2806 (O_2806,N_24993,N_24594);
or UO_2807 (O_2807,N_24886,N_24880);
nand UO_2808 (O_2808,N_24737,N_24927);
or UO_2809 (O_2809,N_24847,N_24823);
nand UO_2810 (O_2810,N_24534,N_24765);
xnor UO_2811 (O_2811,N_24699,N_24635);
and UO_2812 (O_2812,N_24746,N_24931);
nand UO_2813 (O_2813,N_24710,N_24720);
nand UO_2814 (O_2814,N_24655,N_24599);
and UO_2815 (O_2815,N_24633,N_24862);
nor UO_2816 (O_2816,N_24658,N_24863);
nor UO_2817 (O_2817,N_24975,N_24528);
and UO_2818 (O_2818,N_24964,N_24757);
nand UO_2819 (O_2819,N_24719,N_24705);
and UO_2820 (O_2820,N_24921,N_24940);
nor UO_2821 (O_2821,N_24821,N_24874);
nor UO_2822 (O_2822,N_24966,N_24512);
or UO_2823 (O_2823,N_24970,N_24862);
nand UO_2824 (O_2824,N_24925,N_24682);
or UO_2825 (O_2825,N_24961,N_24532);
or UO_2826 (O_2826,N_24581,N_24624);
or UO_2827 (O_2827,N_24619,N_24859);
and UO_2828 (O_2828,N_24977,N_24929);
nor UO_2829 (O_2829,N_24648,N_24621);
nand UO_2830 (O_2830,N_24810,N_24829);
and UO_2831 (O_2831,N_24980,N_24637);
and UO_2832 (O_2832,N_24782,N_24713);
or UO_2833 (O_2833,N_24581,N_24783);
or UO_2834 (O_2834,N_24688,N_24922);
nor UO_2835 (O_2835,N_24648,N_24962);
nor UO_2836 (O_2836,N_24923,N_24583);
nand UO_2837 (O_2837,N_24670,N_24501);
nor UO_2838 (O_2838,N_24618,N_24947);
and UO_2839 (O_2839,N_24933,N_24669);
or UO_2840 (O_2840,N_24534,N_24578);
nand UO_2841 (O_2841,N_24796,N_24662);
nand UO_2842 (O_2842,N_24515,N_24825);
or UO_2843 (O_2843,N_24956,N_24503);
nor UO_2844 (O_2844,N_24981,N_24963);
or UO_2845 (O_2845,N_24849,N_24700);
nor UO_2846 (O_2846,N_24826,N_24966);
and UO_2847 (O_2847,N_24908,N_24543);
nand UO_2848 (O_2848,N_24681,N_24724);
nand UO_2849 (O_2849,N_24761,N_24788);
nand UO_2850 (O_2850,N_24558,N_24535);
nand UO_2851 (O_2851,N_24917,N_24628);
nor UO_2852 (O_2852,N_24817,N_24616);
nand UO_2853 (O_2853,N_24831,N_24623);
nand UO_2854 (O_2854,N_24504,N_24761);
or UO_2855 (O_2855,N_24971,N_24995);
nand UO_2856 (O_2856,N_24771,N_24714);
or UO_2857 (O_2857,N_24722,N_24527);
and UO_2858 (O_2858,N_24842,N_24886);
nor UO_2859 (O_2859,N_24545,N_24602);
or UO_2860 (O_2860,N_24603,N_24809);
nand UO_2861 (O_2861,N_24586,N_24860);
nor UO_2862 (O_2862,N_24982,N_24567);
and UO_2863 (O_2863,N_24971,N_24582);
or UO_2864 (O_2864,N_24643,N_24797);
nor UO_2865 (O_2865,N_24941,N_24602);
or UO_2866 (O_2866,N_24970,N_24574);
and UO_2867 (O_2867,N_24807,N_24962);
and UO_2868 (O_2868,N_24900,N_24521);
or UO_2869 (O_2869,N_24923,N_24552);
or UO_2870 (O_2870,N_24949,N_24933);
nand UO_2871 (O_2871,N_24929,N_24560);
nand UO_2872 (O_2872,N_24859,N_24658);
nor UO_2873 (O_2873,N_24601,N_24608);
nor UO_2874 (O_2874,N_24972,N_24868);
and UO_2875 (O_2875,N_24709,N_24990);
nor UO_2876 (O_2876,N_24888,N_24913);
nand UO_2877 (O_2877,N_24589,N_24592);
nor UO_2878 (O_2878,N_24546,N_24601);
nor UO_2879 (O_2879,N_24534,N_24550);
nor UO_2880 (O_2880,N_24899,N_24587);
or UO_2881 (O_2881,N_24674,N_24537);
and UO_2882 (O_2882,N_24557,N_24896);
nand UO_2883 (O_2883,N_24712,N_24553);
and UO_2884 (O_2884,N_24555,N_24501);
nor UO_2885 (O_2885,N_24935,N_24753);
nand UO_2886 (O_2886,N_24605,N_24663);
nand UO_2887 (O_2887,N_24854,N_24903);
and UO_2888 (O_2888,N_24754,N_24780);
and UO_2889 (O_2889,N_24634,N_24673);
nand UO_2890 (O_2890,N_24789,N_24840);
nand UO_2891 (O_2891,N_24624,N_24909);
nand UO_2892 (O_2892,N_24579,N_24530);
and UO_2893 (O_2893,N_24880,N_24936);
nor UO_2894 (O_2894,N_24565,N_24623);
and UO_2895 (O_2895,N_24525,N_24614);
and UO_2896 (O_2896,N_24678,N_24624);
xnor UO_2897 (O_2897,N_24509,N_24504);
nand UO_2898 (O_2898,N_24806,N_24707);
and UO_2899 (O_2899,N_24948,N_24974);
nor UO_2900 (O_2900,N_24864,N_24526);
and UO_2901 (O_2901,N_24627,N_24913);
and UO_2902 (O_2902,N_24855,N_24831);
nor UO_2903 (O_2903,N_24509,N_24919);
nor UO_2904 (O_2904,N_24834,N_24988);
and UO_2905 (O_2905,N_24634,N_24603);
nand UO_2906 (O_2906,N_24882,N_24857);
and UO_2907 (O_2907,N_24785,N_24827);
nand UO_2908 (O_2908,N_24841,N_24616);
nand UO_2909 (O_2909,N_24586,N_24765);
or UO_2910 (O_2910,N_24621,N_24659);
xnor UO_2911 (O_2911,N_24733,N_24836);
or UO_2912 (O_2912,N_24834,N_24772);
nand UO_2913 (O_2913,N_24878,N_24852);
nor UO_2914 (O_2914,N_24512,N_24565);
nand UO_2915 (O_2915,N_24616,N_24930);
and UO_2916 (O_2916,N_24569,N_24937);
and UO_2917 (O_2917,N_24652,N_24742);
nand UO_2918 (O_2918,N_24573,N_24630);
nor UO_2919 (O_2919,N_24771,N_24558);
nand UO_2920 (O_2920,N_24944,N_24820);
nor UO_2921 (O_2921,N_24715,N_24751);
nor UO_2922 (O_2922,N_24536,N_24991);
nor UO_2923 (O_2923,N_24658,N_24565);
or UO_2924 (O_2924,N_24994,N_24862);
or UO_2925 (O_2925,N_24588,N_24811);
nand UO_2926 (O_2926,N_24627,N_24603);
or UO_2927 (O_2927,N_24860,N_24612);
and UO_2928 (O_2928,N_24945,N_24590);
or UO_2929 (O_2929,N_24517,N_24936);
nand UO_2930 (O_2930,N_24774,N_24595);
nand UO_2931 (O_2931,N_24871,N_24672);
and UO_2932 (O_2932,N_24630,N_24796);
nand UO_2933 (O_2933,N_24914,N_24864);
nand UO_2934 (O_2934,N_24563,N_24797);
or UO_2935 (O_2935,N_24550,N_24646);
nor UO_2936 (O_2936,N_24872,N_24930);
nand UO_2937 (O_2937,N_24816,N_24947);
nor UO_2938 (O_2938,N_24928,N_24761);
nand UO_2939 (O_2939,N_24688,N_24865);
nor UO_2940 (O_2940,N_24697,N_24832);
nor UO_2941 (O_2941,N_24766,N_24564);
xor UO_2942 (O_2942,N_24674,N_24731);
and UO_2943 (O_2943,N_24895,N_24842);
and UO_2944 (O_2944,N_24914,N_24778);
or UO_2945 (O_2945,N_24808,N_24743);
and UO_2946 (O_2946,N_24641,N_24548);
or UO_2947 (O_2947,N_24959,N_24922);
nor UO_2948 (O_2948,N_24549,N_24684);
or UO_2949 (O_2949,N_24905,N_24505);
or UO_2950 (O_2950,N_24778,N_24840);
and UO_2951 (O_2951,N_24799,N_24742);
nand UO_2952 (O_2952,N_24984,N_24671);
nor UO_2953 (O_2953,N_24859,N_24530);
and UO_2954 (O_2954,N_24505,N_24793);
nand UO_2955 (O_2955,N_24814,N_24504);
nand UO_2956 (O_2956,N_24816,N_24594);
or UO_2957 (O_2957,N_24900,N_24965);
nor UO_2958 (O_2958,N_24636,N_24536);
or UO_2959 (O_2959,N_24875,N_24934);
nor UO_2960 (O_2960,N_24569,N_24751);
or UO_2961 (O_2961,N_24971,N_24966);
or UO_2962 (O_2962,N_24719,N_24772);
nor UO_2963 (O_2963,N_24629,N_24647);
nor UO_2964 (O_2964,N_24537,N_24937);
and UO_2965 (O_2965,N_24644,N_24798);
or UO_2966 (O_2966,N_24929,N_24780);
nand UO_2967 (O_2967,N_24682,N_24816);
and UO_2968 (O_2968,N_24838,N_24816);
nor UO_2969 (O_2969,N_24612,N_24553);
nand UO_2970 (O_2970,N_24530,N_24694);
or UO_2971 (O_2971,N_24734,N_24844);
or UO_2972 (O_2972,N_24724,N_24930);
nand UO_2973 (O_2973,N_24592,N_24630);
or UO_2974 (O_2974,N_24751,N_24753);
xnor UO_2975 (O_2975,N_24508,N_24798);
or UO_2976 (O_2976,N_24611,N_24838);
xor UO_2977 (O_2977,N_24697,N_24904);
or UO_2978 (O_2978,N_24623,N_24660);
or UO_2979 (O_2979,N_24605,N_24648);
and UO_2980 (O_2980,N_24874,N_24703);
xor UO_2981 (O_2981,N_24689,N_24724);
xnor UO_2982 (O_2982,N_24739,N_24610);
nor UO_2983 (O_2983,N_24762,N_24987);
and UO_2984 (O_2984,N_24581,N_24708);
nand UO_2985 (O_2985,N_24806,N_24549);
nor UO_2986 (O_2986,N_24756,N_24923);
or UO_2987 (O_2987,N_24687,N_24843);
and UO_2988 (O_2988,N_24702,N_24925);
nand UO_2989 (O_2989,N_24961,N_24984);
nand UO_2990 (O_2990,N_24740,N_24921);
or UO_2991 (O_2991,N_24790,N_24806);
nor UO_2992 (O_2992,N_24744,N_24707);
nor UO_2993 (O_2993,N_24636,N_24560);
or UO_2994 (O_2994,N_24930,N_24960);
or UO_2995 (O_2995,N_24938,N_24543);
and UO_2996 (O_2996,N_24596,N_24514);
nand UO_2997 (O_2997,N_24509,N_24572);
nor UO_2998 (O_2998,N_24950,N_24606);
nor UO_2999 (O_2999,N_24690,N_24869);
endmodule