module basic_1500_15000_2000_3_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10005,N_10006,N_10007,N_10009,N_10010,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10029,N_10031,N_10032,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10054,N_10055,N_10056,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10067,N_10068,N_10070,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10081,N_10082,N_10083,N_10084,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10118,N_10119,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10149,N_10150,N_10152,N_10153,N_10154,N_10155,N_10156,N_10158,N_10159,N_10160,N_10162,N_10163,N_10165,N_10167,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10187,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10211,N_10213,N_10215,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10240,N_10242,N_10243,N_10245,N_10246,N_10247,N_10250,N_10251,N_10252,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10264,N_10266,N_10267,N_10268,N_10269,N_10270,N_10272,N_10273,N_10276,N_10277,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10292,N_10293,N_10294,N_10297,N_10298,N_10300,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10309,N_10310,N_10311,N_10313,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10341,N_10344,N_10345,N_10346,N_10348,N_10349,N_10350,N_10351,N_10352,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10376,N_10377,N_10380,N_10381,N_10382,N_10383,N_10385,N_10386,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10400,N_10401,N_10402,N_10403,N_10405,N_10406,N_10408,N_10409,N_10410,N_10412,N_10413,N_10414,N_10415,N_10417,N_10418,N_10419,N_10420,N_10422,N_10423,N_10424,N_10425,N_10426,N_10428,N_10429,N_10430,N_10431,N_10432,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10464,N_10465,N_10466,N_10468,N_10469,N_10470,N_10471,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10483,N_10484,N_10485,N_10488,N_10489,N_10490,N_10491,N_10492,N_10495,N_10496,N_10497,N_10499,N_10500,N_10501,N_10502,N_10503,N_10505,N_10506,N_10507,N_10508,N_10509,N_10511,N_10513,N_10514,N_10515,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10543,N_10544,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10558,N_10561,N_10562,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10576,N_10577,N_10579,N_10580,N_10581,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10591,N_10592,N_10593,N_10594,N_10596,N_10598,N_10600,N_10602,N_10603,N_10604,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10622,N_10623,N_10624,N_10625,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10650,N_10651,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10668,N_10670,N_10671,N_10674,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10716,N_10718,N_10719,N_10720,N_10721,N_10723,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10739,N_10740,N_10741,N_10743,N_10744,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10764,N_10765,N_10766,N_10767,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10791,N_10792,N_10794,N_10795,N_10796,N_10798,N_10799,N_10801,N_10802,N_10803,N_10804,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10825,N_10826,N_10827,N_10828,N_10829,N_10831,N_10832,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10856,N_10857,N_10858,N_10861,N_10862,N_10863,N_10864,N_10865,N_10867,N_10868,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10883,N_10885,N_10886,N_10888,N_10889,N_10890,N_10891,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10903,N_10905,N_10906,N_10907,N_10909,N_10910,N_10911,N_10912,N_10913,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10944,N_10945,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10967,N_10968,N_10969,N_10970,N_10971,N_10973,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10992,N_10993,N_10995,N_10997,N_10999,N_11000,N_11001,N_11002,N_11003,N_11005,N_11006,N_11007,N_11009,N_11010,N_11011,N_11012,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11021,N_11022,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11044,N_11047,N_11048,N_11049,N_11051,N_11052,N_11053,N_11054,N_11057,N_11059,N_11060,N_11061,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11078,N_11079,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11106,N_11107,N_11108,N_11109,N_11111,N_11112,N_11113,N_11114,N_11115,N_11117,N_11118,N_11119,N_11120,N_11122,N_11123,N_11124,N_11125,N_11126,N_11129,N_11131,N_11132,N_11133,N_11134,N_11136,N_11138,N_11139,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11159,N_11161,N_11162,N_11163,N_11164,N_11165,N_11168,N_11171,N_11172,N_11173,N_11174,N_11175,N_11177,N_11178,N_11179,N_11180,N_11181,N_11183,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11195,N_11196,N_11197,N_11199,N_11200,N_11201,N_11202,N_11203,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11213,N_11215,N_11217,N_11218,N_11219,N_11220,N_11222,N_11223,N_11224,N_11227,N_11228,N_11229,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11241,N_11242,N_11243,N_11244,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11272,N_11273,N_11274,N_11276,N_11277,N_11279,N_11280,N_11282,N_11283,N_11286,N_11287,N_11288,N_11289,N_11290,N_11292,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11305,N_11306,N_11307,N_11308,N_11309,N_11311,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11327,N_11328,N_11329,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11339,N_11340,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11359,N_11360,N_11361,N_11363,N_11364,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11385,N_11386,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11427,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11471,N_11472,N_11473,N_11474,N_11475,N_11478,N_11484,N_11485,N_11488,N_11489,N_11490,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11503,N_11504,N_11505,N_11506,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11531,N_11533,N_11534,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11550,N_11551,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11561,N_11562,N_11563,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11575,N_11576,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11586,N_11587,N_11588,N_11589,N_11590,N_11594,N_11597,N_11599,N_11600,N_11601,N_11602,N_11603,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11642,N_11643,N_11644,N_11645,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11655,N_11656,N_11657,N_11659,N_11660,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11671,N_11672,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11695,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11726,N_11727,N_11728,N_11730,N_11731,N_11732,N_11734,N_11735,N_11736,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11761,N_11762,N_11763,N_11766,N_11768,N_11769,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11783,N_11784,N_11786,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11797,N_11798,N_11799,N_11801,N_11802,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11823,N_11824,N_11826,N_11828,N_11829,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11858,N_11859,N_11860,N_11861,N_11864,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11876,N_11879,N_11880,N_11881,N_11882,N_11884,N_11885,N_11887,N_11888,N_11889,N_11891,N_11892,N_11894,N_11897,N_11899,N_11900,N_11901,N_11902,N_11903,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11934,N_11935,N_11936,N_11938,N_11939,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11948,N_11949,N_11950,N_11951,N_11952,N_11954,N_11955,N_11956,N_11957,N_11958,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11982,N_11983,N_11985,N_11986,N_11987,N_11988,N_11989,N_11991,N_11992,N_11993,N_11994,N_11995,N_11998,N_11999,N_12000,N_12001,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12032,N_12033,N_12034,N_12035,N_12036,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12051,N_12052,N_12056,N_12057,N_12058,N_12059,N_12060,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12069,N_12070,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12084,N_12085,N_12086,N_12087,N_12088,N_12090,N_12091,N_12092,N_12093,N_12095,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12107,N_12108,N_12110,N_12111,N_12112,N_12114,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12123,N_12124,N_12125,N_12127,N_12129,N_12130,N_12131,N_12132,N_12133,N_12135,N_12136,N_12137,N_12138,N_12139,N_12141,N_12142,N_12144,N_12145,N_12146,N_12148,N_12149,N_12150,N_12151,N_12152,N_12154,N_12156,N_12157,N_12158,N_12159,N_12161,N_12162,N_12163,N_12164,N_12165,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12183,N_12185,N_12186,N_12187,N_12190,N_12192,N_12193,N_12195,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12207,N_12208,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12256,N_12258,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12269,N_12272,N_12273,N_12274,N_12276,N_12278,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12293,N_12294,N_12295,N_12296,N_12297,N_12299,N_12300,N_12301,N_12305,N_12307,N_12308,N_12309,N_12310,N_12312,N_12313,N_12314,N_12316,N_12317,N_12320,N_12321,N_12322,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12340,N_12341,N_12342,N_12343,N_12344,N_12346,N_12347,N_12348,N_12349,N_12351,N_12352,N_12353,N_12354,N_12355,N_12357,N_12358,N_12359,N_12360,N_12361,N_12363,N_12364,N_12365,N_12366,N_12368,N_12370,N_12371,N_12373,N_12374,N_12376,N_12377,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12396,N_12397,N_12398,N_12399,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12418,N_12420,N_12422,N_12424,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12433,N_12434,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12446,N_12447,N_12449,N_12450,N_12451,N_12453,N_12454,N_12455,N_12456,N_12458,N_12459,N_12460,N_12463,N_12464,N_12465,N_12466,N_12467,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12483,N_12484,N_12485,N_12488,N_12489,N_12491,N_12493,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12518,N_12519,N_12520,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12530,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12539,N_12540,N_12541,N_12542,N_12543,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12552,N_12553,N_12554,N_12555,N_12556,N_12559,N_12560,N_12561,N_12562,N_12564,N_12565,N_12566,N_12567,N_12568,N_12571,N_12572,N_12574,N_12576,N_12577,N_12579,N_12580,N_12581,N_12582,N_12583,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12598,N_12599,N_12600,N_12602,N_12603,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12615,N_12616,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12632,N_12634,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12647,N_12648,N_12649,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12699,N_12700,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12716,N_12717,N_12720,N_12721,N_12722,N_12723,N_12725,N_12727,N_12729,N_12730,N_12731,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12742,N_12743,N_12744,N_12746,N_12748,N_12751,N_12752,N_12754,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12784,N_12785,N_12786,N_12787,N_12788,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12802,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12819,N_12820,N_12822,N_12823,N_12825,N_12826,N_12827,N_12829,N_12830,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12840,N_12841,N_12843,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12855,N_12856,N_12857,N_12858,N_12859,N_12861,N_12863,N_12865,N_12866,N_12868,N_12869,N_12870,N_12872,N_12873,N_12874,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12886,N_12887,N_12888,N_12892,N_12893,N_12894,N_12896,N_12897,N_12901,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12912,N_12913,N_12914,N_12915,N_12918,N_12919,N_12921,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12933,N_12934,N_12935,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12951,N_12952,N_12954,N_12955,N_12958,N_12959,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12970,N_12971,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13002,N_13003,N_13004,N_13006,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13022,N_13023,N_13025,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13034,N_13035,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13046,N_13047,N_13049,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13058,N_13060,N_13062,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13075,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13102,N_13103,N_13106,N_13108,N_13109,N_13110,N_13111,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13123,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13134,N_13135,N_13137,N_13139,N_13140,N_13141,N_13142,N_13143,N_13145,N_13147,N_13148,N_13149,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13159,N_13161,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13173,N_13174,N_13178,N_13179,N_13180,N_13181,N_13182,N_13184,N_13185,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13196,N_13197,N_13198,N_13200,N_13201,N_13202,N_13203,N_13207,N_13208,N_13210,N_13211,N_13212,N_13213,N_13214,N_13216,N_13217,N_13219,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13243,N_13244,N_13245,N_13246,N_13248,N_13249,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13269,N_13270,N_13271,N_13273,N_13274,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13289,N_13290,N_13291,N_13292,N_13294,N_13295,N_13296,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13333,N_13334,N_13335,N_13336,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13352,N_13353,N_13354,N_13355,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13364,N_13365,N_13366,N_13367,N_13370,N_13371,N_13372,N_13374,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13383,N_13384,N_13385,N_13387,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13396,N_13397,N_13398,N_13399,N_13400,N_13402,N_13403,N_13405,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13416,N_13417,N_13418,N_13419,N_13421,N_13422,N_13423,N_13424,N_13425,N_13427,N_13428,N_13429,N_13431,N_13432,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13491,N_13492,N_13493,N_13495,N_13496,N_13497,N_13498,N_13499,N_13501,N_13503,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13512,N_13513,N_13514,N_13515,N_13517,N_13519,N_13520,N_13522,N_13523,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13542,N_13543,N_13544,N_13545,N_13546,N_13548,N_13549,N_13551,N_13552,N_13554,N_13555,N_13556,N_13558,N_13559,N_13560,N_13562,N_13563,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13576,N_13577,N_13578,N_13579,N_13582,N_13584,N_13586,N_13587,N_13588,N_13589,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13600,N_13601,N_13603,N_13604,N_13606,N_13607,N_13609,N_13610,N_13611,N_13612,N_13613,N_13615,N_13616,N_13617,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13626,N_13627,N_13629,N_13630,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13639,N_13640,N_13642,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13662,N_13664,N_13665,N_13666,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13689,N_13690,N_13691,N_13692,N_13694,N_13695,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13717,N_13719,N_13720,N_13721,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13733,N_13734,N_13737,N_13739,N_13740,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13753,N_13754,N_13756,N_13757,N_13758,N_13759,N_13761,N_13763,N_13766,N_13767,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13785,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13821,N_13822,N_13823,N_13824,N_13826,N_13828,N_13829,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13843,N_13844,N_13845,N_13846,N_13847,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13866,N_13868,N_13869,N_13871,N_13872,N_13873,N_13874,N_13877,N_13878,N_13880,N_13882,N_13883,N_13884,N_13885,N_13888,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13897,N_13898,N_13900,N_13901,N_13902,N_13905,N_13906,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13926,N_13927,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13950,N_13951,N_13952,N_13953,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13974,N_13975,N_13976,N_13977,N_13979,N_13981,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13992,N_13993,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14002,N_14003,N_14005,N_14006,N_14007,N_14009,N_14011,N_14012,N_14013,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14069,N_14070,N_14071,N_14072,N_14075,N_14077,N_14078,N_14079,N_14081,N_14082,N_14083,N_14084,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14099,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14115,N_14116,N_14117,N_14118,N_14119,N_14122,N_14123,N_14124,N_14126,N_14127,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14138,N_14139,N_14141,N_14142,N_14145,N_14146,N_14147,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14166,N_14167,N_14168,N_14171,N_14172,N_14173,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14193,N_14194,N_14195,N_14196,N_14197,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14210,N_14211,N_14212,N_14213,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14235,N_14236,N_14238,N_14239,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14257,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14271,N_14272,N_14273,N_14274,N_14275,N_14277,N_14278,N_14279,N_14280,N_14281,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14291,N_14292,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14318,N_14319,N_14320,N_14321,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14344,N_14345,N_14346,N_14347,N_14348,N_14351,N_14352,N_14353,N_14354,N_14355,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14369,N_14370,N_14371,N_14373,N_14374,N_14376,N_14377,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14398,N_14400,N_14402,N_14403,N_14404,N_14405,N_14407,N_14408,N_14409,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14424,N_14425,N_14426,N_14427,N_14428,N_14430,N_14433,N_14434,N_14435,N_14437,N_14438,N_14441,N_14442,N_14444,N_14445,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14456,N_14457,N_14459,N_14460,N_14462,N_14463,N_14465,N_14466,N_14467,N_14468,N_14472,N_14473,N_14475,N_14477,N_14478,N_14480,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14500,N_14502,N_14503,N_14504,N_14505,N_14507,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14525,N_14527,N_14528,N_14530,N_14531,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14543,N_14544,N_14545,N_14546,N_14547,N_14550,N_14551,N_14552,N_14553,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14574,N_14575,N_14576,N_14578,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14603,N_14605,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14616,N_14617,N_14618,N_14619,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14628,N_14630,N_14632,N_14633,N_14634,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14645,N_14646,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14665,N_14666,N_14668,N_14670,N_14671,N_14672,N_14674,N_14677,N_14678,N_14679,N_14680,N_14681,N_14684,N_14685,N_14687,N_14690,N_14691,N_14692,N_14693,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14704,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14713,N_14714,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14744,N_14745,N_14746,N_14747,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14762,N_14763,N_14766,N_14767,N_14769,N_14770,N_14772,N_14773,N_14774,N_14776,N_14778,N_14779,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14805,N_14806,N_14807,N_14808,N_14809,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14849,N_14850,N_14851,N_14852,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14863,N_14864,N_14865,N_14866,N_14867,N_14869,N_14871,N_14873,N_14874,N_14875,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14893,N_14894,N_14895,N_14896,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14913,N_14916,N_14917,N_14918,N_14919,N_14921,N_14922,N_14923,N_14925,N_14926,N_14927,N_14928,N_14929,N_14931,N_14934,N_14935,N_14937,N_14939,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14956,N_14957,N_14958,N_14959,N_14960,N_14962,N_14963,N_14964,N_14965,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14984,N_14986,N_14987,N_14988,N_14990,N_14992,N_14994,N_14995,N_14996,N_14998,N_14999;
nor U0 (N_0,In_86,In_161);
or U1 (N_1,In_151,In_718);
nand U2 (N_2,In_1054,In_694);
nor U3 (N_3,In_294,In_1365);
and U4 (N_4,In_1288,In_911);
and U5 (N_5,In_1094,In_568);
nor U6 (N_6,In_881,In_1182);
nand U7 (N_7,In_1344,In_177);
or U8 (N_8,In_436,In_229);
or U9 (N_9,In_1474,In_1368);
nand U10 (N_10,In_1356,In_1482);
or U11 (N_11,In_100,In_345);
nand U12 (N_12,In_494,In_1120);
or U13 (N_13,In_407,In_1138);
nor U14 (N_14,In_193,In_1287);
nand U15 (N_15,In_520,In_555);
nand U16 (N_16,In_526,In_1197);
and U17 (N_17,In_828,In_806);
nor U18 (N_18,In_604,In_872);
nand U19 (N_19,In_957,In_1198);
or U20 (N_20,In_706,In_114);
nand U21 (N_21,In_1099,In_120);
and U22 (N_22,In_288,In_1095);
nor U23 (N_23,In_303,In_295);
nor U24 (N_24,In_183,In_308);
nor U25 (N_25,In_674,In_1236);
nand U26 (N_26,In_880,In_1100);
nor U27 (N_27,In_328,In_645);
nor U28 (N_28,In_472,In_932);
nor U29 (N_29,In_578,In_832);
nor U30 (N_30,In_426,In_1364);
or U31 (N_31,In_1467,In_800);
and U32 (N_32,In_204,In_589);
and U33 (N_33,In_730,In_382);
or U34 (N_34,In_637,In_688);
or U35 (N_35,In_682,In_309);
nand U36 (N_36,In_1487,In_136);
and U37 (N_37,In_1471,In_349);
nor U38 (N_38,In_524,In_1176);
or U39 (N_39,In_235,In_686);
or U40 (N_40,In_1177,In_201);
or U41 (N_41,In_1475,In_1409);
or U42 (N_42,In_456,In_1234);
nor U43 (N_43,In_703,In_1440);
nor U44 (N_44,In_447,In_843);
nor U45 (N_45,In_1181,In_398);
and U46 (N_46,In_968,In_1022);
nor U47 (N_47,In_1276,In_768);
nor U48 (N_48,In_1283,In_1111);
and U49 (N_49,In_1112,In_1348);
nand U50 (N_50,In_481,In_870);
and U51 (N_51,In_52,In_338);
nor U52 (N_52,In_1196,In_534);
nand U53 (N_53,In_653,In_434);
nor U54 (N_54,In_1476,In_504);
nor U55 (N_55,In_1019,In_944);
or U56 (N_56,In_1031,In_1088);
nor U57 (N_57,In_749,In_314);
nand U58 (N_58,In_319,In_1133);
and U59 (N_59,In_28,In_242);
or U60 (N_60,In_1404,In_173);
nor U61 (N_61,In_327,In_1334);
nor U62 (N_62,In_418,In_540);
or U63 (N_63,In_929,In_226);
and U64 (N_64,In_1491,In_529);
nand U65 (N_65,In_433,In_774);
or U66 (N_66,In_897,In_72);
or U67 (N_67,In_65,In_856);
or U68 (N_68,In_149,In_1238);
or U69 (N_69,In_602,In_1465);
or U70 (N_70,In_379,In_820);
nor U71 (N_71,In_1314,In_388);
or U72 (N_72,In_482,In_250);
nor U73 (N_73,In_1466,In_885);
and U74 (N_74,In_1479,In_1067);
nor U75 (N_75,In_404,In_683);
nand U76 (N_76,In_561,In_1258);
nor U77 (N_77,In_74,In_1492);
xnor U78 (N_78,In_1290,In_143);
nand U79 (N_79,In_935,In_884);
and U80 (N_80,In_376,In_203);
and U81 (N_81,In_1011,In_1469);
nand U82 (N_82,In_876,In_80);
and U83 (N_83,In_390,In_996);
and U84 (N_84,In_521,In_284);
nand U85 (N_85,In_842,In_646);
and U86 (N_86,In_507,In_396);
or U87 (N_87,In_1030,In_89);
or U88 (N_88,In_823,In_443);
or U89 (N_89,In_855,In_1225);
nand U90 (N_90,In_1463,In_64);
nor U91 (N_91,In_454,In_457);
and U92 (N_92,In_1201,In_248);
and U93 (N_93,In_598,In_714);
or U94 (N_94,In_680,In_67);
nor U95 (N_95,In_946,In_417);
nand U96 (N_96,In_574,In_1014);
nand U97 (N_97,In_1206,In_1435);
or U98 (N_98,In_276,In_508);
nor U99 (N_99,In_792,In_1121);
or U100 (N_100,In_191,In_1423);
and U101 (N_101,In_1333,In_1412);
or U102 (N_102,In_1468,In_422);
nand U103 (N_103,In_593,In_96);
and U104 (N_104,In_1267,In_318);
or U105 (N_105,In_187,In_355);
nor U106 (N_106,In_633,In_847);
nor U107 (N_107,In_705,In_39);
and U108 (N_108,In_1457,In_770);
or U109 (N_109,In_720,In_716);
and U110 (N_110,In_59,In_926);
nor U111 (N_111,In_986,In_208);
nor U112 (N_112,In_659,In_609);
and U113 (N_113,In_906,In_1117);
and U114 (N_114,In_211,In_1322);
and U115 (N_115,In_1498,In_1449);
and U116 (N_116,In_271,In_367);
nand U117 (N_117,In_228,In_1190);
nand U118 (N_118,In_1472,In_1363);
or U119 (N_119,In_588,In_196);
nor U120 (N_120,In_1327,In_671);
nor U121 (N_121,In_1245,In_479);
and U122 (N_122,In_945,In_1066);
or U123 (N_123,In_1152,In_1172);
nand U124 (N_124,In_162,In_179);
xor U125 (N_125,In_528,In_1044);
or U126 (N_126,In_403,In_527);
nor U127 (N_127,In_232,In_697);
or U128 (N_128,In_1354,In_1216);
nor U129 (N_129,In_1091,In_970);
and U130 (N_130,In_1053,In_788);
or U131 (N_131,In_638,In_641);
nand U132 (N_132,In_901,In_743);
nand U133 (N_133,In_342,In_863);
nor U134 (N_134,In_1174,In_937);
and U135 (N_135,In_488,In_1331);
nor U136 (N_136,In_1135,In_1320);
nor U137 (N_137,In_724,In_257);
nor U138 (N_138,In_1132,In_849);
nand U139 (N_139,In_1396,In_569);
or U140 (N_140,In_585,In_894);
or U141 (N_141,In_105,In_317);
and U142 (N_142,In_950,In_809);
nor U143 (N_143,In_621,In_1146);
nand U144 (N_144,In_635,In_1230);
and U145 (N_145,In_1231,In_841);
and U146 (N_146,In_989,In_12);
and U147 (N_147,In_158,In_925);
nor U148 (N_148,In_1256,In_928);
nor U149 (N_149,In_1086,In_664);
nand U150 (N_150,In_483,In_492);
and U151 (N_151,In_631,In_1241);
nor U152 (N_152,In_1006,In_1187);
or U153 (N_153,In_839,In_550);
nor U154 (N_154,In_184,In_1336);
nor U155 (N_155,In_565,In_969);
or U156 (N_156,In_1134,In_45);
or U157 (N_157,In_735,In_1140);
nor U158 (N_158,In_1193,In_952);
nand U159 (N_159,In_141,In_728);
nand U160 (N_160,In_44,In_1394);
nor U161 (N_161,In_1040,In_1093);
and U162 (N_162,In_684,In_537);
or U163 (N_163,In_9,In_1309);
and U164 (N_164,In_1366,In_36);
nor U165 (N_165,In_461,In_907);
nand U166 (N_166,In_816,In_708);
nand U167 (N_167,In_1441,In_1321);
nor U168 (N_168,In_796,In_1384);
nand U169 (N_169,In_1185,In_163);
or U170 (N_170,In_450,In_369);
nor U171 (N_171,In_689,In_1494);
or U172 (N_172,In_316,In_640);
nor U173 (N_173,In_661,In_1299);
nand U174 (N_174,In_261,In_372);
or U175 (N_175,In_87,In_243);
or U176 (N_176,In_803,In_181);
and U177 (N_177,In_862,In_125);
and U178 (N_178,In_1183,In_1023);
nor U179 (N_179,In_1055,In_1084);
nor U180 (N_180,In_1388,In_1462);
or U181 (N_181,In_1305,In_1013);
nand U182 (N_182,In_1431,In_32);
nor U183 (N_183,In_940,In_1060);
nor U184 (N_184,In_913,In_1085);
and U185 (N_185,In_513,In_441);
nor U186 (N_186,In_4,In_98);
or U187 (N_187,In_73,In_1009);
or U188 (N_188,In_1381,In_931);
nand U189 (N_189,In_176,In_914);
nor U190 (N_190,In_124,In_547);
and U191 (N_191,In_837,In_1272);
nand U192 (N_192,In_733,In_365);
nor U193 (N_193,In_188,In_1143);
or U194 (N_194,In_954,In_500);
nor U195 (N_195,In_10,In_1255);
and U196 (N_196,In_936,In_1282);
and U197 (N_197,In_502,In_964);
or U198 (N_198,In_1422,In_1045);
and U199 (N_199,In_610,In_974);
and U200 (N_200,In_1379,In_893);
nand U201 (N_201,In_160,In_37);
xnor U202 (N_202,In_1295,In_237);
or U203 (N_203,In_990,In_363);
nand U204 (N_204,In_938,In_551);
nor U205 (N_205,In_785,In_675);
and U206 (N_206,In_1397,In_1156);
and U207 (N_207,In_84,In_824);
nor U208 (N_208,In_1136,In_767);
nand U209 (N_209,In_423,In_625);
and U210 (N_210,In_1002,In_1455);
or U211 (N_211,In_453,In_1414);
nand U212 (N_212,In_46,In_468);
nor U213 (N_213,In_627,In_459);
and U214 (N_214,In_979,In_1316);
and U215 (N_215,In_1144,In_399);
nor U216 (N_216,In_642,In_299);
nor U217 (N_217,In_2,In_1048);
and U218 (N_218,In_1046,In_651);
nand U219 (N_219,In_538,In_321);
nand U220 (N_220,In_1239,In_1035);
and U221 (N_221,In_763,In_584);
or U222 (N_222,In_614,In_1200);
and U223 (N_223,In_385,In_209);
nand U224 (N_224,In_834,In_17);
nand U225 (N_225,In_600,In_1380);
nor U226 (N_226,In_1269,In_496);
nand U227 (N_227,In_462,In_1353);
and U228 (N_228,In_1340,In_375);
and U229 (N_229,In_1421,In_498);
nor U230 (N_230,In_1259,In_1090);
nand U231 (N_231,In_343,In_993);
and U232 (N_232,In_1049,In_1056);
and U233 (N_233,In_1367,In_207);
nor U234 (N_234,In_34,In_900);
nor U235 (N_235,In_804,In_334);
nor U236 (N_236,In_464,In_206);
and U237 (N_237,In_1137,In_685);
or U238 (N_238,In_825,In_57);
nand U239 (N_239,In_634,In_557);
nand U240 (N_240,In_1203,In_643);
and U241 (N_241,In_1127,In_811);
or U242 (N_242,In_1335,In_1392);
nand U243 (N_243,In_1262,In_185);
nor U244 (N_244,In_1456,In_465);
nand U245 (N_245,In_1107,In_1173);
and U246 (N_246,In_1101,In_1124);
or U247 (N_247,In_1395,In_238);
nor U248 (N_248,In_1432,In_1192);
and U249 (N_249,In_753,In_628);
nor U250 (N_250,In_455,In_378);
nor U251 (N_251,In_1123,In_88);
nor U252 (N_252,In_1459,In_864);
and U253 (N_253,In_425,In_467);
nor U254 (N_254,In_516,In_332);
and U255 (N_255,In_411,In_967);
nor U256 (N_256,In_233,In_963);
nand U257 (N_257,In_972,In_1378);
or U258 (N_258,In_132,In_1083);
nand U259 (N_259,In_941,In_1061);
and U260 (N_260,In_808,In_566);
nor U261 (N_261,In_994,In_1279);
and U262 (N_262,In_1338,In_1115);
or U263 (N_263,In_517,In_817);
nand U264 (N_264,In_908,In_113);
nand U265 (N_265,In_1213,In_1303);
and U266 (N_266,In_23,In_1220);
and U267 (N_267,In_1000,In_1160);
and U268 (N_268,In_424,In_1105);
nor U269 (N_269,In_1062,In_51);
nor U270 (N_270,In_1485,In_882);
nand U271 (N_271,In_1376,In_655);
nand U272 (N_272,In_110,In_1142);
and U273 (N_273,In_1175,In_707);
nor U274 (N_274,In_420,In_789);
xor U275 (N_275,In_1224,In_985);
nand U276 (N_276,In_178,In_278);
nand U277 (N_277,In_750,In_874);
and U278 (N_278,In_1477,In_539);
nand U279 (N_279,In_400,In_1261);
or U280 (N_280,In_1158,In_556);
nand U281 (N_281,In_444,In_564);
nor U282 (N_282,In_1154,In_819);
nand U283 (N_283,In_1444,In_1406);
and U284 (N_284,In_868,In_346);
and U285 (N_285,In_1163,In_542);
and U286 (N_286,In_1437,In_745);
nor U287 (N_287,In_463,In_883);
and U288 (N_288,In_890,In_1222);
nor U289 (N_289,In_771,In_1411);
or U290 (N_290,In_478,In_1429);
or U291 (N_291,In_240,In_387);
or U292 (N_292,In_1063,In_1351);
nand U293 (N_293,In_713,In_779);
or U294 (N_294,In_669,In_195);
nand U295 (N_295,In_983,In_783);
and U296 (N_296,In_497,In_76);
or U297 (N_297,In_613,In_873);
nor U298 (N_298,In_106,In_111);
nor U299 (N_299,In_171,In_180);
and U300 (N_300,In_1195,In_340);
nor U301 (N_301,In_315,In_687);
or U302 (N_302,In_272,In_780);
and U303 (N_303,In_205,In_1387);
and U304 (N_304,In_1298,In_922);
nor U305 (N_305,In_899,In_335);
or U306 (N_306,In_489,In_491);
nand U307 (N_307,In_1027,In_469);
and U308 (N_308,In_1129,In_1452);
or U309 (N_309,In_1419,In_131);
and U310 (N_310,In_71,In_446);
or U311 (N_311,In_821,In_1417);
nor U312 (N_312,In_522,In_1042);
nand U313 (N_313,In_449,In_249);
and U314 (N_314,In_1403,In_354);
nand U315 (N_315,In_215,In_943);
nand U316 (N_316,In_1148,In_154);
or U317 (N_317,In_1026,In_329);
nor U318 (N_318,In_452,In_1318);
nand U319 (N_319,In_1076,In_1390);
or U320 (N_320,In_264,In_1436);
or U321 (N_321,In_1217,In_1352);
nand U322 (N_322,In_861,In_236);
nor U323 (N_323,In_1420,In_1438);
nor U324 (N_324,In_290,In_231);
nor U325 (N_325,In_761,In_818);
or U326 (N_326,In_852,In_1024);
and U327 (N_327,In_1454,In_826);
nand U328 (N_328,In_1038,In_626);
nor U329 (N_329,In_1039,In_942);
and U330 (N_330,In_953,In_719);
and U331 (N_331,In_330,In_1497);
nand U332 (N_332,In_1005,In_402);
xor U333 (N_333,In_493,In_174);
nor U334 (N_334,In_965,In_1247);
nand U335 (N_335,In_268,In_48);
and U336 (N_336,In_230,In_1306);
and U337 (N_337,In_123,In_758);
and U338 (N_338,In_930,In_0);
and U339 (N_339,In_854,In_1179);
and U340 (N_340,In_1389,In_169);
nand U341 (N_341,In_844,In_1264);
nor U342 (N_342,In_281,In_47);
nand U343 (N_343,In_1211,In_381);
nand U344 (N_344,In_756,In_148);
or U345 (N_345,In_217,In_119);
and U346 (N_346,In_1168,In_451);
and U347 (N_347,In_891,In_448);
or U348 (N_348,In_591,In_279);
or U349 (N_349,In_535,In_976);
nor U350 (N_350,In_1427,In_1128);
or U351 (N_351,In_759,In_1405);
or U352 (N_352,In_1447,In_137);
and U353 (N_353,In_1147,In_1077);
nand U354 (N_354,In_419,In_1359);
and U355 (N_355,In_128,In_917);
nand U356 (N_356,In_1265,In_416);
nor U357 (N_357,In_1189,In_150);
nor U358 (N_358,In_904,In_1229);
or U359 (N_359,In_1029,In_992);
or U360 (N_360,In_644,In_499);
or U361 (N_361,In_1235,In_1486);
or U362 (N_362,In_269,In_867);
and U363 (N_363,In_853,In_1164);
or U364 (N_364,In_1277,In_995);
and U365 (N_365,In_1329,In_81);
nand U366 (N_366,In_1202,In_797);
or U367 (N_367,In_322,In_421);
nand U368 (N_368,In_924,In_360);
and U369 (N_369,In_1080,In_186);
or U370 (N_370,In_43,In_285);
or U371 (N_371,In_153,In_1139);
nor U372 (N_372,In_672,In_898);
and U373 (N_373,In_1153,In_1311);
nor U374 (N_374,In_582,In_1481);
or U375 (N_375,In_620,In_170);
nand U376 (N_376,In_1007,In_1313);
nor U377 (N_377,In_473,In_1273);
nor U378 (N_378,In_596,In_1237);
nor U379 (N_379,In_1416,In_1243);
or U380 (N_380,In_475,In_765);
nor U381 (N_381,In_312,In_845);
and U382 (N_382,In_220,In_251);
nand U383 (N_383,In_1339,In_1242);
xor U384 (N_384,In_648,In_7);
nand U385 (N_385,In_484,In_571);
nor U386 (N_386,In_639,In_704);
nor U387 (N_387,In_1249,In_1032);
nor U388 (N_388,In_1496,In_1286);
nand U389 (N_389,In_984,In_58);
or U390 (N_390,In_1342,In_858);
and U391 (N_391,In_1480,In_1393);
nand U392 (N_392,In_658,In_301);
nand U393 (N_393,In_21,In_344);
and U394 (N_394,In_1069,In_734);
nor U395 (N_395,In_503,In_1260);
or U396 (N_396,In_695,In_977);
or U397 (N_397,In_63,In_341);
or U398 (N_398,In_33,In_962);
nand U399 (N_399,In_544,In_259);
and U400 (N_400,In_782,In_736);
or U401 (N_401,In_752,In_1223);
and U402 (N_402,In_530,In_1453);
nand U403 (N_403,In_570,In_711);
nor U404 (N_404,In_192,In_1285);
and U405 (N_405,In_1064,In_224);
nand U406 (N_406,In_833,In_19);
and U407 (N_407,In_258,In_1271);
nand U408 (N_408,In_1119,In_1297);
nand U409 (N_409,In_53,In_275);
and U410 (N_410,In_35,In_239);
or U411 (N_411,In_717,In_1377);
nand U412 (N_412,In_1489,In_617);
nor U413 (N_413,In_835,In_933);
nand U414 (N_414,In_518,In_75);
or U415 (N_415,In_723,In_117);
or U416 (N_416,In_693,In_1155);
or U417 (N_417,In_607,In_474);
and U418 (N_418,In_1433,In_118);
nor U419 (N_419,In_748,In_94);
and U420 (N_420,In_296,In_1126);
nand U421 (N_421,In_274,In_1051);
nor U422 (N_422,In_13,In_225);
or U423 (N_423,In_715,In_26);
nand U424 (N_424,In_587,In_1349);
and U425 (N_425,In_576,In_1098);
or U426 (N_426,In_265,In_624);
or U427 (N_427,In_515,In_978);
and U428 (N_428,In_189,In_337);
nand U429 (N_429,In_99,In_1018);
nand U430 (N_430,In_681,In_1375);
and U431 (N_431,In_55,In_959);
nor U432 (N_432,In_307,In_1325);
and U433 (N_433,In_1415,In_1167);
nand U434 (N_434,In_1221,In_1004);
and U435 (N_435,In_1343,In_532);
and U436 (N_436,In_1113,In_1170);
or U437 (N_437,In_573,In_1043);
nor U438 (N_438,In_138,In_406);
and U439 (N_439,In_878,In_432);
or U440 (N_440,In_49,In_895);
nand U441 (N_441,In_1490,In_351);
or U442 (N_442,In_563,In_1207);
nand U443 (N_443,In_155,In_1226);
nor U444 (N_444,In_889,In_1450);
or U445 (N_445,In_1310,In_815);
nand U446 (N_446,In_619,In_60);
or U447 (N_447,In_1347,In_438);
nor U448 (N_448,In_401,In_487);
nand U449 (N_449,In_982,In_380);
and U450 (N_450,In_213,In_24);
nor U451 (N_451,In_435,In_152);
and U452 (N_452,In_916,In_829);
and U453 (N_453,In_168,In_612);
and U454 (N_454,In_656,In_1162);
nand U455 (N_455,In_794,In_1361);
or U456 (N_456,In_888,In_200);
nand U457 (N_457,In_297,In_300);
nor U458 (N_458,In_865,In_549);
and U459 (N_459,In_310,In_601);
nor U460 (N_460,In_781,In_877);
nand U461 (N_461,In_27,In_116);
nand U462 (N_462,In_773,In_107);
nor U463 (N_463,In_840,In_1424);
or U464 (N_464,In_280,In_790);
or U465 (N_465,In_145,In_3);
nand U466 (N_466,In_1052,In_1410);
or U467 (N_467,In_79,In_164);
or U468 (N_468,In_1104,In_729);
nor U469 (N_469,In_305,In_973);
or U470 (N_470,In_395,In_199);
or U471 (N_471,In_480,In_987);
or U472 (N_472,In_552,In_56);
or U473 (N_473,In_77,In_1149);
nor U474 (N_474,In_731,In_320);
nor U475 (N_475,In_1214,In_592);
or U476 (N_476,In_1257,In_1370);
nand U477 (N_477,In_115,In_92);
and U478 (N_478,In_392,In_1263);
nand U479 (N_479,In_636,In_146);
xnor U480 (N_480,In_1087,In_869);
and U481 (N_481,In_386,In_405);
nor U482 (N_482,In_896,In_618);
xnor U483 (N_483,In_1458,In_1114);
nand U484 (N_484,In_130,In_991);
and U485 (N_485,In_1400,In_1470);
and U486 (N_486,In_1166,In_282);
or U487 (N_487,In_1199,In_966);
or U488 (N_488,In_194,In_1184);
nor U489 (N_489,In_608,In_960);
nor U490 (N_490,In_988,In_859);
nor U491 (N_491,In_1010,In_902);
nor U492 (N_492,In_241,In_223);
or U493 (N_493,In_362,In_1021);
or U494 (N_494,In_1016,In_1326);
or U495 (N_495,In_597,In_393);
nor U496 (N_496,In_927,In_439);
or U497 (N_497,In_1425,In_415);
nor U498 (N_498,In_830,In_949);
nand U499 (N_499,In_1407,In_519);
or U500 (N_500,In_325,In_353);
or U501 (N_501,In_860,In_391);
or U502 (N_502,In_159,In_630);
nor U503 (N_503,In_554,In_622);
nor U504 (N_504,In_1280,In_795);
nand U505 (N_505,In_560,In_1399);
and U506 (N_506,In_777,In_668);
nand U507 (N_507,In_616,In_747);
nand U508 (N_508,In_887,In_1483);
and U509 (N_509,In_69,In_1369);
nand U510 (N_510,In_1266,In_252);
or U511 (N_511,In_553,In_586);
nor U512 (N_512,In_590,In_667);
and U513 (N_513,In_769,In_410);
nand U514 (N_514,In_1268,In_1209);
and U515 (N_515,In_1293,In_262);
or U516 (N_516,In_256,In_1081);
nand U517 (N_517,In_1401,In_701);
and U518 (N_518,In_1362,In_541);
or U519 (N_519,In_1328,In_665);
or U520 (N_520,In_5,In_787);
or U521 (N_521,In_1037,In_1041);
nand U522 (N_522,In_583,In_266);
nor U523 (N_523,In_1284,In_1337);
and U524 (N_524,In_31,In_791);
nor U525 (N_525,In_373,In_915);
and U526 (N_526,In_650,In_358);
or U527 (N_527,In_778,In_352);
nor U528 (N_528,In_1050,In_102);
or U529 (N_529,In_1426,In_1079);
or U530 (N_530,In_1188,In_696);
nor U531 (N_531,In_595,In_848);
nor U532 (N_532,In_798,In_214);
nand U533 (N_533,In_1072,In_397);
nor U534 (N_534,In_90,In_104);
or U535 (N_535,In_1253,In_247);
nor U536 (N_536,In_850,In_323);
or U537 (N_537,In_20,In_246);
or U538 (N_538,In_1332,In_754);
or U539 (N_539,In_919,In_1034);
nand U540 (N_540,In_384,In_581);
nand U541 (N_541,In_1047,In_918);
and U542 (N_542,In_460,In_54);
nand U543 (N_543,In_6,In_732);
or U544 (N_544,In_923,In_14);
nand U545 (N_545,In_227,In_293);
or U546 (N_546,In_903,In_1012);
nand U547 (N_547,In_776,In_741);
and U548 (N_548,In_1122,In_807);
or U549 (N_549,In_1402,In_267);
xor U550 (N_550,In_1015,In_1151);
nand U551 (N_551,In_1178,In_744);
nand U552 (N_552,In_692,In_1244);
nand U553 (N_553,In_95,In_1341);
and U554 (N_554,In_1065,In_666);
nand U555 (N_555,In_905,In_1070);
nor U556 (N_556,In_722,In_1270);
or U557 (N_557,In_244,In_377);
nor U558 (N_558,In_579,In_1307);
nor U559 (N_559,In_1460,In_1408);
nand U560 (N_560,In_1473,In_22);
nor U561 (N_561,In_934,In_93);
nor U562 (N_562,In_1275,In_629);
and U563 (N_563,In_1017,In_775);
and U564 (N_564,In_721,In_1391);
or U565 (N_565,In_287,In_466);
nor U566 (N_566,In_41,In_142);
and U567 (N_567,In_662,In_350);
or U568 (N_568,In_108,In_147);
nor U569 (N_569,In_260,In_157);
xor U570 (N_570,In_62,In_1358);
nor U571 (N_571,In_359,In_394);
nor U572 (N_572,In_1131,In_366);
nor U573 (N_573,In_1291,In_414);
nand U574 (N_574,In_331,In_812);
or U575 (N_575,In_738,In_562);
nor U576 (N_576,In_66,In_140);
and U577 (N_577,In_1312,In_611);
nand U578 (N_578,In_559,In_910);
and U579 (N_579,In_980,In_663);
nor U580 (N_580,In_997,In_202);
nor U581 (N_581,In_831,In_1157);
and U582 (N_582,In_1301,In_702);
nor U583 (N_583,In_1373,In_948);
nand U584 (N_584,In_951,In_810);
or U585 (N_585,In_975,In_78);
nand U586 (N_586,In_762,In_1246);
or U587 (N_587,In_1116,In_190);
or U588 (N_588,In_112,In_357);
and U589 (N_589,In_1110,In_766);
nand U590 (N_590,In_1109,In_29);
nor U591 (N_591,In_85,In_437);
nor U592 (N_592,In_760,In_649);
nor U593 (N_593,In_298,In_383);
nor U594 (N_594,In_1252,In_1278);
or U595 (N_595,In_1484,In_165);
nand U596 (N_596,In_892,In_427);
nand U597 (N_597,In_1145,In_103);
nor U598 (N_598,In_50,In_1317);
and U599 (N_599,In_428,In_1096);
nand U600 (N_600,In_1186,In_802);
or U601 (N_601,In_1250,In_866);
and U602 (N_602,In_1371,In_1360);
nand U603 (N_603,In_691,In_97);
or U604 (N_604,In_757,In_121);
or U605 (N_605,In_886,In_921);
or U606 (N_606,In_1150,In_699);
and U607 (N_607,In_471,In_122);
and U608 (N_608,In_509,In_109);
or U609 (N_609,In_1330,In_70);
and U610 (N_610,In_476,In_1165);
or U611 (N_611,In_1057,In_1071);
nand U612 (N_612,In_1296,In_134);
nor U613 (N_613,In_175,In_222);
nand U614 (N_614,In_16,In_712);
and U615 (N_615,In_799,In_1292);
or U616 (N_616,In_575,In_673);
nand U617 (N_617,In_389,In_430);
nor U618 (N_618,In_368,In_1345);
and U619 (N_619,In_652,In_742);
and U620 (N_620,In_255,In_727);
nor U621 (N_621,In_1082,In_739);
and U622 (N_622,In_690,In_1495);
and U623 (N_623,In_289,In_751);
nor U624 (N_624,In_1169,In_709);
nand U625 (N_625,In_514,In_1205);
or U626 (N_626,In_263,In_1171);
nor U627 (N_627,In_61,In_846);
nor U628 (N_628,In_42,In_302);
or U629 (N_629,In_1191,In_700);
nand U630 (N_630,In_955,In_786);
nor U631 (N_631,In_1219,In_495);
or U632 (N_632,In_11,In_1180);
nor U633 (N_633,In_632,In_409);
or U634 (N_634,In_139,In_38);
nand U635 (N_635,In_1036,In_166);
or U636 (N_636,In_68,In_304);
nand U637 (N_637,In_1451,In_1464);
nor U638 (N_638,In_1355,In_909);
and U639 (N_639,In_431,In_291);
nand U640 (N_640,In_1078,In_533);
and U641 (N_641,In_958,In_1254);
or U642 (N_642,In_1089,In_212);
and U643 (N_643,In_603,In_133);
nor U644 (N_644,In_1304,In_254);
nor U645 (N_645,In_580,In_408);
nor U646 (N_646,In_126,In_548);
nand U647 (N_647,In_326,In_135);
or U648 (N_648,In_726,In_678);
nor U649 (N_649,In_746,In_1102);
nand U650 (N_650,In_654,In_1434);
nor U651 (N_651,In_577,In_429);
nor U652 (N_652,In_567,In_1324);
and U653 (N_653,In_273,In_920);
xnor U654 (N_654,In_1,In_1499);
and U655 (N_655,In_851,In_283);
or U656 (N_656,In_998,In_947);
nand U657 (N_657,In_531,In_361);
and U658 (N_658,In_172,In_510);
or U659 (N_659,In_144,In_543);
nor U660 (N_660,In_1442,In_1385);
or U661 (N_661,In_1446,In_1289);
nor U662 (N_662,In_1428,In_485);
or U663 (N_663,In_710,In_572);
and U664 (N_664,In_324,In_277);
and U665 (N_665,In_525,In_871);
or U666 (N_666,In_1478,In_370);
or U667 (N_667,In_270,In_82);
nand U668 (N_668,In_311,In_606);
and U669 (N_669,In_1075,In_536);
nor U670 (N_670,In_961,In_156);
and U671 (N_671,In_971,In_599);
nand U672 (N_672,In_1319,In_364);
and U673 (N_673,In_1033,In_1103);
nor U674 (N_674,In_813,In_442);
nand U675 (N_675,In_1218,In_999);
and U676 (N_676,In_857,In_511);
nor U677 (N_677,In_615,In_1281);
or U678 (N_678,In_470,In_755);
and U679 (N_679,In_40,In_523);
nand U680 (N_680,In_1108,In_91);
xor U681 (N_681,In_1208,In_127);
and U682 (N_682,In_253,In_339);
or U683 (N_683,In_1141,In_1025);
nand U684 (N_684,In_676,In_1308);
and U685 (N_685,In_875,In_1159);
xnor U686 (N_686,In_764,In_594);
nor U687 (N_687,In_221,In_1398);
nand U688 (N_688,In_1240,In_647);
nor U689 (N_689,In_1118,In_1386);
nor U690 (N_690,In_725,In_1302);
or U691 (N_691,In_827,In_814);
and U692 (N_692,In_219,In_371);
and U693 (N_693,In_8,In_545);
or U694 (N_694,In_512,In_1001);
and U695 (N_695,In_374,In_1372);
nand U696 (N_696,In_1227,In_486);
nor U697 (N_697,In_313,In_1204);
nor U698 (N_698,In_1315,In_737);
and U699 (N_699,In_216,In_1251);
or U700 (N_700,In_336,In_1445);
and U701 (N_701,In_1073,In_1430);
nor U702 (N_702,In_1493,In_1461);
nand U703 (N_703,In_1215,In_1346);
and U704 (N_704,In_1058,In_167);
nand U705 (N_705,In_306,In_1274);
nand U706 (N_706,In_1374,In_1439);
nor U707 (N_707,In_1228,In_1357);
nor U708 (N_708,In_1350,In_1020);
and U709 (N_709,In_18,In_879);
and U710 (N_710,In_939,In_956);
or U711 (N_711,In_784,In_740);
or U712 (N_712,In_912,In_83);
nor U713 (N_713,In_679,In_660);
and U714 (N_714,In_182,In_348);
nand U715 (N_715,In_445,In_1232);
nor U716 (N_716,In_1248,In_801);
xor U717 (N_717,In_1194,In_412);
and U718 (N_718,In_698,In_670);
nand U719 (N_719,In_477,In_623);
or U720 (N_720,In_1068,In_30);
and U721 (N_721,In_1323,In_1059);
nand U722 (N_722,In_1074,In_1418);
or U723 (N_723,In_333,In_838);
nor U724 (N_724,In_1212,In_1008);
nor U725 (N_725,In_1130,In_772);
nand U726 (N_726,In_347,In_101);
and U727 (N_727,In_1106,In_677);
nand U728 (N_728,In_210,In_1092);
or U729 (N_729,In_197,In_805);
and U730 (N_730,In_1028,In_1488);
nor U731 (N_731,In_822,In_356);
nor U732 (N_732,In_234,In_657);
nand U733 (N_733,In_1233,In_501);
and U734 (N_734,In_440,In_490);
nand U735 (N_735,In_1161,In_546);
nor U736 (N_736,In_1210,In_15);
xnor U737 (N_737,In_836,In_1003);
nand U738 (N_738,In_505,In_506);
or U739 (N_739,In_1443,In_1382);
nand U740 (N_740,In_218,In_1125);
nand U741 (N_741,In_245,In_1294);
nor U742 (N_742,In_1413,In_605);
nand U743 (N_743,In_1383,In_1300);
nand U744 (N_744,In_981,In_129);
or U745 (N_745,In_286,In_458);
or U746 (N_746,In_1097,In_198);
or U747 (N_747,In_292,In_558);
or U748 (N_748,In_1448,In_793);
and U749 (N_749,In_25,In_413);
or U750 (N_750,In_1495,In_150);
nand U751 (N_751,In_672,In_1178);
or U752 (N_752,In_508,In_1018);
and U753 (N_753,In_259,In_29);
nor U754 (N_754,In_1448,In_269);
nand U755 (N_755,In_538,In_1284);
or U756 (N_756,In_809,In_1419);
and U757 (N_757,In_106,In_1202);
and U758 (N_758,In_371,In_1000);
nor U759 (N_759,In_1344,In_676);
nand U760 (N_760,In_1277,In_698);
nand U761 (N_761,In_660,In_466);
or U762 (N_762,In_1122,In_24);
nor U763 (N_763,In_299,In_480);
nand U764 (N_764,In_897,In_7);
or U765 (N_765,In_54,In_1144);
nand U766 (N_766,In_1199,In_319);
nand U767 (N_767,In_373,In_887);
or U768 (N_768,In_1371,In_803);
and U769 (N_769,In_866,In_1225);
or U770 (N_770,In_331,In_44);
nand U771 (N_771,In_1018,In_333);
nor U772 (N_772,In_1063,In_207);
or U773 (N_773,In_663,In_1409);
nor U774 (N_774,In_1444,In_1245);
nand U775 (N_775,In_210,In_1459);
xor U776 (N_776,In_239,In_977);
nor U777 (N_777,In_937,In_1002);
nor U778 (N_778,In_68,In_532);
nor U779 (N_779,In_1469,In_1490);
nor U780 (N_780,In_1391,In_1208);
nand U781 (N_781,In_518,In_174);
nand U782 (N_782,In_26,In_253);
nand U783 (N_783,In_496,In_223);
and U784 (N_784,In_518,In_297);
and U785 (N_785,In_1329,In_1074);
nor U786 (N_786,In_1096,In_1458);
and U787 (N_787,In_764,In_1093);
and U788 (N_788,In_651,In_1157);
or U789 (N_789,In_522,In_501);
nor U790 (N_790,In_260,In_121);
nand U791 (N_791,In_1329,In_1352);
nand U792 (N_792,In_18,In_1019);
and U793 (N_793,In_301,In_779);
and U794 (N_794,In_866,In_173);
nand U795 (N_795,In_1077,In_557);
and U796 (N_796,In_1025,In_172);
and U797 (N_797,In_1334,In_120);
and U798 (N_798,In_1345,In_1105);
nor U799 (N_799,In_314,In_1061);
nor U800 (N_800,In_1415,In_46);
nand U801 (N_801,In_207,In_1335);
and U802 (N_802,In_146,In_785);
nor U803 (N_803,In_1344,In_1324);
nor U804 (N_804,In_523,In_599);
or U805 (N_805,In_114,In_1419);
or U806 (N_806,In_1137,In_1375);
nand U807 (N_807,In_81,In_757);
or U808 (N_808,In_1441,In_106);
nor U809 (N_809,In_216,In_279);
or U810 (N_810,In_922,In_887);
nor U811 (N_811,In_1040,In_1478);
and U812 (N_812,In_713,In_393);
or U813 (N_813,In_223,In_431);
or U814 (N_814,In_431,In_765);
and U815 (N_815,In_70,In_370);
and U816 (N_816,In_271,In_108);
or U817 (N_817,In_1059,In_1260);
and U818 (N_818,In_844,In_505);
nand U819 (N_819,In_613,In_670);
nor U820 (N_820,In_1019,In_601);
xor U821 (N_821,In_1263,In_694);
nor U822 (N_822,In_1097,In_641);
nand U823 (N_823,In_880,In_1460);
or U824 (N_824,In_545,In_992);
nor U825 (N_825,In_715,In_458);
or U826 (N_826,In_480,In_1356);
nand U827 (N_827,In_874,In_106);
nand U828 (N_828,In_857,In_1467);
nor U829 (N_829,In_866,In_1098);
nor U830 (N_830,In_357,In_1087);
and U831 (N_831,In_798,In_1011);
nor U832 (N_832,In_271,In_1372);
and U833 (N_833,In_195,In_136);
and U834 (N_834,In_1330,In_300);
nor U835 (N_835,In_1355,In_1478);
nand U836 (N_836,In_1128,In_312);
nand U837 (N_837,In_529,In_386);
nor U838 (N_838,In_950,In_1283);
or U839 (N_839,In_678,In_238);
or U840 (N_840,In_358,In_608);
and U841 (N_841,In_1080,In_1450);
nor U842 (N_842,In_1493,In_389);
and U843 (N_843,In_1108,In_363);
nand U844 (N_844,In_111,In_572);
and U845 (N_845,In_1188,In_239);
xor U846 (N_846,In_718,In_123);
or U847 (N_847,In_1465,In_1090);
nor U848 (N_848,In_1389,In_1088);
nor U849 (N_849,In_833,In_1085);
nand U850 (N_850,In_867,In_1239);
nor U851 (N_851,In_825,In_849);
or U852 (N_852,In_787,In_932);
or U853 (N_853,In_1383,In_1449);
and U854 (N_854,In_250,In_1139);
or U855 (N_855,In_1312,In_1165);
xor U856 (N_856,In_569,In_1417);
nand U857 (N_857,In_599,In_406);
or U858 (N_858,In_738,In_1453);
nor U859 (N_859,In_1128,In_866);
or U860 (N_860,In_574,In_1419);
or U861 (N_861,In_221,In_453);
nand U862 (N_862,In_437,In_536);
nor U863 (N_863,In_996,In_1159);
nor U864 (N_864,In_24,In_192);
nand U865 (N_865,In_1065,In_1313);
nor U866 (N_866,In_1100,In_1151);
nor U867 (N_867,In_753,In_819);
nand U868 (N_868,In_1186,In_300);
nand U869 (N_869,In_1331,In_469);
nor U870 (N_870,In_122,In_742);
nand U871 (N_871,In_1168,In_1392);
or U872 (N_872,In_1170,In_1160);
or U873 (N_873,In_905,In_142);
nor U874 (N_874,In_207,In_525);
nand U875 (N_875,In_552,In_129);
nor U876 (N_876,In_948,In_593);
or U877 (N_877,In_91,In_864);
nand U878 (N_878,In_1111,In_1432);
and U879 (N_879,In_750,In_758);
nand U880 (N_880,In_13,In_304);
or U881 (N_881,In_1264,In_821);
nand U882 (N_882,In_29,In_1496);
and U883 (N_883,In_193,In_1061);
nor U884 (N_884,In_1174,In_32);
nand U885 (N_885,In_943,In_1079);
and U886 (N_886,In_685,In_1309);
or U887 (N_887,In_120,In_1358);
and U888 (N_888,In_930,In_1099);
and U889 (N_889,In_658,In_1298);
nand U890 (N_890,In_217,In_934);
nor U891 (N_891,In_1431,In_166);
nand U892 (N_892,In_813,In_543);
nand U893 (N_893,In_380,In_607);
or U894 (N_894,In_120,In_1256);
nor U895 (N_895,In_387,In_677);
nand U896 (N_896,In_651,In_1493);
nand U897 (N_897,In_993,In_980);
and U898 (N_898,In_446,In_431);
and U899 (N_899,In_266,In_105);
and U900 (N_900,In_676,In_1286);
or U901 (N_901,In_1071,In_253);
and U902 (N_902,In_746,In_32);
or U903 (N_903,In_598,In_1005);
or U904 (N_904,In_1088,In_1029);
and U905 (N_905,In_1376,In_1239);
nor U906 (N_906,In_524,In_203);
nor U907 (N_907,In_343,In_785);
nor U908 (N_908,In_319,In_851);
and U909 (N_909,In_858,In_519);
nor U910 (N_910,In_1205,In_330);
nand U911 (N_911,In_491,In_304);
nor U912 (N_912,In_784,In_978);
nand U913 (N_913,In_309,In_1013);
nand U914 (N_914,In_1461,In_1456);
nor U915 (N_915,In_939,In_1173);
and U916 (N_916,In_907,In_136);
nand U917 (N_917,In_1019,In_958);
or U918 (N_918,In_420,In_880);
and U919 (N_919,In_131,In_24);
or U920 (N_920,In_115,In_290);
nor U921 (N_921,In_1422,In_1297);
and U922 (N_922,In_1180,In_1495);
and U923 (N_923,In_794,In_386);
nand U924 (N_924,In_1388,In_368);
or U925 (N_925,In_677,In_405);
nand U926 (N_926,In_835,In_690);
nor U927 (N_927,In_63,In_1215);
or U928 (N_928,In_395,In_1299);
nor U929 (N_929,In_1461,In_72);
nand U930 (N_930,In_888,In_622);
or U931 (N_931,In_884,In_113);
and U932 (N_932,In_171,In_845);
and U933 (N_933,In_410,In_1001);
nand U934 (N_934,In_175,In_797);
and U935 (N_935,In_861,In_940);
xor U936 (N_936,In_1244,In_1358);
nor U937 (N_937,In_520,In_875);
nor U938 (N_938,In_239,In_741);
and U939 (N_939,In_188,In_39);
or U940 (N_940,In_885,In_968);
nor U941 (N_941,In_1005,In_509);
and U942 (N_942,In_241,In_522);
nor U943 (N_943,In_1315,In_420);
and U944 (N_944,In_1489,In_1435);
or U945 (N_945,In_545,In_116);
nor U946 (N_946,In_1374,In_1001);
nor U947 (N_947,In_894,In_1019);
or U948 (N_948,In_85,In_0);
and U949 (N_949,In_744,In_1041);
nor U950 (N_950,In_270,In_906);
or U951 (N_951,In_1399,In_694);
and U952 (N_952,In_1011,In_926);
and U953 (N_953,In_857,In_1117);
nand U954 (N_954,In_918,In_1433);
or U955 (N_955,In_1322,In_846);
or U956 (N_956,In_251,In_673);
nor U957 (N_957,In_856,In_607);
or U958 (N_958,In_535,In_499);
nand U959 (N_959,In_940,In_1438);
or U960 (N_960,In_1309,In_639);
nand U961 (N_961,In_250,In_994);
or U962 (N_962,In_311,In_1053);
nand U963 (N_963,In_916,In_690);
and U964 (N_964,In_1413,In_1);
nand U965 (N_965,In_1010,In_342);
nand U966 (N_966,In_194,In_1204);
nor U967 (N_967,In_845,In_564);
and U968 (N_968,In_1239,In_1257);
nor U969 (N_969,In_245,In_1355);
or U970 (N_970,In_599,In_125);
nand U971 (N_971,In_382,In_998);
nand U972 (N_972,In_603,In_422);
nor U973 (N_973,In_851,In_294);
or U974 (N_974,In_1370,In_995);
or U975 (N_975,In_721,In_339);
nand U976 (N_976,In_134,In_771);
or U977 (N_977,In_509,In_1113);
nand U978 (N_978,In_1251,In_387);
or U979 (N_979,In_515,In_669);
and U980 (N_980,In_1476,In_681);
nor U981 (N_981,In_43,In_13);
nand U982 (N_982,In_696,In_240);
or U983 (N_983,In_542,In_1199);
or U984 (N_984,In_1339,In_961);
nand U985 (N_985,In_1445,In_196);
nand U986 (N_986,In_1342,In_1129);
nor U987 (N_987,In_436,In_18);
or U988 (N_988,In_1261,In_714);
or U989 (N_989,In_498,In_888);
and U990 (N_990,In_700,In_823);
nand U991 (N_991,In_1235,In_765);
nor U992 (N_992,In_1083,In_354);
or U993 (N_993,In_140,In_1232);
or U994 (N_994,In_83,In_193);
or U995 (N_995,In_1283,In_1122);
and U996 (N_996,In_918,In_1328);
nor U997 (N_997,In_591,In_292);
nand U998 (N_998,In_339,In_204);
nand U999 (N_999,In_397,In_1036);
nor U1000 (N_1000,In_40,In_24);
nand U1001 (N_1001,In_431,In_2);
or U1002 (N_1002,In_67,In_445);
nor U1003 (N_1003,In_1132,In_324);
nor U1004 (N_1004,In_92,In_18);
nand U1005 (N_1005,In_1052,In_71);
and U1006 (N_1006,In_1110,In_36);
or U1007 (N_1007,In_505,In_635);
nand U1008 (N_1008,In_313,In_847);
xnor U1009 (N_1009,In_590,In_503);
or U1010 (N_1010,In_707,In_1462);
nor U1011 (N_1011,In_176,In_685);
nand U1012 (N_1012,In_1367,In_970);
nor U1013 (N_1013,In_130,In_400);
nand U1014 (N_1014,In_1118,In_219);
and U1015 (N_1015,In_1439,In_1038);
or U1016 (N_1016,In_882,In_348);
nand U1017 (N_1017,In_753,In_1370);
nor U1018 (N_1018,In_660,In_1067);
and U1019 (N_1019,In_645,In_76);
nand U1020 (N_1020,In_690,In_62);
nor U1021 (N_1021,In_190,In_934);
nand U1022 (N_1022,In_832,In_346);
nand U1023 (N_1023,In_1165,In_33);
and U1024 (N_1024,In_191,In_817);
or U1025 (N_1025,In_271,In_493);
nor U1026 (N_1026,In_1367,In_295);
nand U1027 (N_1027,In_729,In_1225);
nor U1028 (N_1028,In_1089,In_1142);
nor U1029 (N_1029,In_1311,In_669);
nor U1030 (N_1030,In_656,In_652);
nor U1031 (N_1031,In_1259,In_688);
and U1032 (N_1032,In_173,In_544);
or U1033 (N_1033,In_861,In_1212);
and U1034 (N_1034,In_967,In_506);
and U1035 (N_1035,In_149,In_627);
or U1036 (N_1036,In_794,In_381);
nor U1037 (N_1037,In_383,In_41);
and U1038 (N_1038,In_750,In_998);
and U1039 (N_1039,In_1350,In_1289);
nand U1040 (N_1040,In_470,In_1257);
and U1041 (N_1041,In_1461,In_881);
nor U1042 (N_1042,In_683,In_97);
nor U1043 (N_1043,In_902,In_1114);
nand U1044 (N_1044,In_234,In_113);
nor U1045 (N_1045,In_767,In_1366);
and U1046 (N_1046,In_258,In_814);
or U1047 (N_1047,In_1191,In_886);
and U1048 (N_1048,In_1124,In_1056);
or U1049 (N_1049,In_701,In_1017);
xnor U1050 (N_1050,In_877,In_1034);
nor U1051 (N_1051,In_833,In_1382);
nor U1052 (N_1052,In_83,In_237);
nand U1053 (N_1053,In_1400,In_93);
and U1054 (N_1054,In_1323,In_1458);
or U1055 (N_1055,In_1217,In_602);
or U1056 (N_1056,In_1392,In_1079);
nor U1057 (N_1057,In_1486,In_1137);
nand U1058 (N_1058,In_1428,In_1272);
nand U1059 (N_1059,In_232,In_1138);
nand U1060 (N_1060,In_533,In_594);
nand U1061 (N_1061,In_49,In_207);
and U1062 (N_1062,In_651,In_1321);
or U1063 (N_1063,In_123,In_81);
nand U1064 (N_1064,In_1440,In_1485);
or U1065 (N_1065,In_1044,In_1494);
nor U1066 (N_1066,In_369,In_797);
nor U1067 (N_1067,In_1288,In_690);
xor U1068 (N_1068,In_53,In_1364);
nor U1069 (N_1069,In_1343,In_1139);
nand U1070 (N_1070,In_1428,In_520);
and U1071 (N_1071,In_377,In_659);
and U1072 (N_1072,In_915,In_994);
xnor U1073 (N_1073,In_1449,In_141);
nand U1074 (N_1074,In_1444,In_492);
nor U1075 (N_1075,In_1455,In_1059);
and U1076 (N_1076,In_834,In_1365);
nand U1077 (N_1077,In_167,In_394);
and U1078 (N_1078,In_1139,In_629);
nor U1079 (N_1079,In_1038,In_1268);
and U1080 (N_1080,In_1223,In_150);
nor U1081 (N_1081,In_986,In_240);
nand U1082 (N_1082,In_597,In_563);
nand U1083 (N_1083,In_517,In_413);
and U1084 (N_1084,In_661,In_872);
or U1085 (N_1085,In_1182,In_406);
nand U1086 (N_1086,In_1226,In_1104);
or U1087 (N_1087,In_310,In_1034);
or U1088 (N_1088,In_1131,In_649);
nor U1089 (N_1089,In_571,In_129);
nand U1090 (N_1090,In_72,In_672);
or U1091 (N_1091,In_905,In_100);
nor U1092 (N_1092,In_921,In_1388);
nor U1093 (N_1093,In_63,In_285);
nand U1094 (N_1094,In_1377,In_224);
and U1095 (N_1095,In_115,In_1418);
or U1096 (N_1096,In_603,In_860);
and U1097 (N_1097,In_180,In_460);
nand U1098 (N_1098,In_1413,In_927);
nand U1099 (N_1099,In_1297,In_790);
nand U1100 (N_1100,In_1061,In_286);
nand U1101 (N_1101,In_997,In_1255);
and U1102 (N_1102,In_513,In_851);
nor U1103 (N_1103,In_924,In_238);
and U1104 (N_1104,In_804,In_342);
nor U1105 (N_1105,In_277,In_1006);
nand U1106 (N_1106,In_28,In_340);
or U1107 (N_1107,In_1113,In_810);
nor U1108 (N_1108,In_1205,In_1336);
and U1109 (N_1109,In_1034,In_1111);
nand U1110 (N_1110,In_1197,In_1240);
nand U1111 (N_1111,In_1478,In_135);
or U1112 (N_1112,In_110,In_841);
nor U1113 (N_1113,In_154,In_738);
nand U1114 (N_1114,In_1065,In_64);
and U1115 (N_1115,In_1224,In_29);
and U1116 (N_1116,In_1106,In_1390);
or U1117 (N_1117,In_371,In_246);
or U1118 (N_1118,In_1138,In_674);
and U1119 (N_1119,In_833,In_79);
or U1120 (N_1120,In_21,In_1081);
nor U1121 (N_1121,In_430,In_1133);
and U1122 (N_1122,In_206,In_168);
nand U1123 (N_1123,In_118,In_43);
nor U1124 (N_1124,In_805,In_544);
or U1125 (N_1125,In_573,In_651);
or U1126 (N_1126,In_1494,In_1280);
nor U1127 (N_1127,In_385,In_1431);
and U1128 (N_1128,In_436,In_1007);
and U1129 (N_1129,In_322,In_215);
nor U1130 (N_1130,In_179,In_419);
or U1131 (N_1131,In_328,In_492);
or U1132 (N_1132,In_1122,In_857);
nor U1133 (N_1133,In_277,In_1078);
xor U1134 (N_1134,In_1074,In_705);
nor U1135 (N_1135,In_1285,In_781);
nor U1136 (N_1136,In_773,In_587);
nor U1137 (N_1137,In_214,In_23);
and U1138 (N_1138,In_1125,In_557);
and U1139 (N_1139,In_1419,In_66);
nand U1140 (N_1140,In_643,In_527);
nor U1141 (N_1141,In_1020,In_65);
nor U1142 (N_1142,In_856,In_1293);
nor U1143 (N_1143,In_468,In_1256);
and U1144 (N_1144,In_477,In_1218);
and U1145 (N_1145,In_1236,In_1387);
or U1146 (N_1146,In_621,In_1447);
nand U1147 (N_1147,In_1377,In_974);
or U1148 (N_1148,In_246,In_1487);
nand U1149 (N_1149,In_547,In_893);
and U1150 (N_1150,In_943,In_417);
and U1151 (N_1151,In_475,In_37);
or U1152 (N_1152,In_1434,In_1306);
nor U1153 (N_1153,In_239,In_405);
or U1154 (N_1154,In_1363,In_369);
nor U1155 (N_1155,In_478,In_999);
or U1156 (N_1156,In_1214,In_92);
nand U1157 (N_1157,In_668,In_560);
and U1158 (N_1158,In_181,In_1302);
and U1159 (N_1159,In_47,In_593);
nor U1160 (N_1160,In_714,In_638);
and U1161 (N_1161,In_281,In_1375);
xnor U1162 (N_1162,In_791,In_1049);
or U1163 (N_1163,In_877,In_204);
or U1164 (N_1164,In_93,In_414);
nor U1165 (N_1165,In_688,In_690);
or U1166 (N_1166,In_1475,In_924);
or U1167 (N_1167,In_1056,In_41);
and U1168 (N_1168,In_266,In_1283);
nand U1169 (N_1169,In_986,In_982);
nor U1170 (N_1170,In_121,In_873);
and U1171 (N_1171,In_1440,In_1355);
nand U1172 (N_1172,In_1210,In_83);
nand U1173 (N_1173,In_510,In_1204);
nor U1174 (N_1174,In_966,In_207);
nand U1175 (N_1175,In_807,In_554);
nor U1176 (N_1176,In_1439,In_783);
nand U1177 (N_1177,In_1215,In_1364);
nand U1178 (N_1178,In_1171,In_228);
and U1179 (N_1179,In_357,In_621);
nor U1180 (N_1180,In_1136,In_78);
nor U1181 (N_1181,In_834,In_726);
or U1182 (N_1182,In_421,In_377);
xor U1183 (N_1183,In_789,In_339);
nand U1184 (N_1184,In_998,In_158);
or U1185 (N_1185,In_1306,In_1484);
and U1186 (N_1186,In_495,In_370);
nor U1187 (N_1187,In_778,In_133);
and U1188 (N_1188,In_916,In_954);
or U1189 (N_1189,In_677,In_1423);
or U1190 (N_1190,In_695,In_642);
or U1191 (N_1191,In_628,In_156);
or U1192 (N_1192,In_637,In_955);
nand U1193 (N_1193,In_978,In_1230);
nand U1194 (N_1194,In_909,In_781);
or U1195 (N_1195,In_337,In_850);
and U1196 (N_1196,In_539,In_1103);
and U1197 (N_1197,In_442,In_602);
and U1198 (N_1198,In_1103,In_945);
nor U1199 (N_1199,In_272,In_1169);
nor U1200 (N_1200,In_398,In_592);
nor U1201 (N_1201,In_1485,In_24);
or U1202 (N_1202,In_1361,In_1369);
nor U1203 (N_1203,In_1446,In_1135);
nand U1204 (N_1204,In_1291,In_1425);
nand U1205 (N_1205,In_1274,In_159);
and U1206 (N_1206,In_150,In_1496);
and U1207 (N_1207,In_84,In_107);
or U1208 (N_1208,In_1376,In_800);
nand U1209 (N_1209,In_991,In_1412);
or U1210 (N_1210,In_533,In_245);
and U1211 (N_1211,In_667,In_327);
and U1212 (N_1212,In_215,In_19);
and U1213 (N_1213,In_950,In_15);
nand U1214 (N_1214,In_225,In_967);
or U1215 (N_1215,In_514,In_516);
or U1216 (N_1216,In_723,In_791);
nand U1217 (N_1217,In_135,In_931);
xor U1218 (N_1218,In_895,In_1337);
and U1219 (N_1219,In_272,In_121);
or U1220 (N_1220,In_1498,In_1054);
or U1221 (N_1221,In_864,In_66);
or U1222 (N_1222,In_401,In_707);
nand U1223 (N_1223,In_76,In_1169);
or U1224 (N_1224,In_231,In_789);
nor U1225 (N_1225,In_59,In_1460);
nand U1226 (N_1226,In_1,In_489);
and U1227 (N_1227,In_1018,In_1392);
and U1228 (N_1228,In_1469,In_486);
or U1229 (N_1229,In_342,In_1180);
and U1230 (N_1230,In_987,In_542);
nand U1231 (N_1231,In_48,In_1176);
nor U1232 (N_1232,In_1017,In_507);
nand U1233 (N_1233,In_1305,In_1309);
nand U1234 (N_1234,In_733,In_1447);
nor U1235 (N_1235,In_745,In_1370);
nor U1236 (N_1236,In_1315,In_960);
nor U1237 (N_1237,In_380,In_870);
nand U1238 (N_1238,In_861,In_1156);
nor U1239 (N_1239,In_1401,In_1423);
nor U1240 (N_1240,In_728,In_710);
or U1241 (N_1241,In_581,In_1119);
or U1242 (N_1242,In_959,In_1428);
and U1243 (N_1243,In_726,In_441);
or U1244 (N_1244,In_1442,In_241);
nand U1245 (N_1245,In_1489,In_970);
nor U1246 (N_1246,In_249,In_721);
nor U1247 (N_1247,In_1163,In_1015);
nor U1248 (N_1248,In_588,In_239);
and U1249 (N_1249,In_1250,In_750);
and U1250 (N_1250,In_685,In_1175);
and U1251 (N_1251,In_1214,In_58);
nor U1252 (N_1252,In_607,In_166);
xnor U1253 (N_1253,In_943,In_1272);
nand U1254 (N_1254,In_857,In_1090);
or U1255 (N_1255,In_114,In_237);
nor U1256 (N_1256,In_1153,In_1177);
nand U1257 (N_1257,In_482,In_453);
nor U1258 (N_1258,In_5,In_783);
nor U1259 (N_1259,In_322,In_93);
or U1260 (N_1260,In_952,In_867);
nand U1261 (N_1261,In_1070,In_640);
xnor U1262 (N_1262,In_840,In_1210);
nand U1263 (N_1263,In_413,In_883);
and U1264 (N_1264,In_398,In_404);
or U1265 (N_1265,In_1486,In_39);
nand U1266 (N_1266,In_377,In_867);
or U1267 (N_1267,In_1315,In_1267);
or U1268 (N_1268,In_364,In_1046);
and U1269 (N_1269,In_269,In_40);
xor U1270 (N_1270,In_1012,In_747);
and U1271 (N_1271,In_93,In_1073);
nor U1272 (N_1272,In_1191,In_195);
nor U1273 (N_1273,In_400,In_575);
nand U1274 (N_1274,In_1189,In_819);
or U1275 (N_1275,In_1235,In_1258);
nand U1276 (N_1276,In_865,In_1497);
and U1277 (N_1277,In_651,In_168);
and U1278 (N_1278,In_900,In_944);
nor U1279 (N_1279,In_629,In_353);
nor U1280 (N_1280,In_999,In_1186);
nand U1281 (N_1281,In_1132,In_1217);
and U1282 (N_1282,In_974,In_964);
nor U1283 (N_1283,In_423,In_360);
nand U1284 (N_1284,In_1155,In_469);
or U1285 (N_1285,In_76,In_588);
nor U1286 (N_1286,In_8,In_218);
or U1287 (N_1287,In_142,In_876);
and U1288 (N_1288,In_302,In_282);
or U1289 (N_1289,In_1386,In_624);
and U1290 (N_1290,In_992,In_1308);
or U1291 (N_1291,In_276,In_160);
and U1292 (N_1292,In_1014,In_231);
nand U1293 (N_1293,In_449,In_65);
or U1294 (N_1294,In_1438,In_654);
nor U1295 (N_1295,In_1462,In_1302);
and U1296 (N_1296,In_1496,In_298);
and U1297 (N_1297,In_127,In_1210);
or U1298 (N_1298,In_143,In_291);
or U1299 (N_1299,In_1115,In_353);
nand U1300 (N_1300,In_590,In_993);
and U1301 (N_1301,In_1115,In_459);
nand U1302 (N_1302,In_822,In_908);
nand U1303 (N_1303,In_1369,In_111);
nor U1304 (N_1304,In_1049,In_1402);
nand U1305 (N_1305,In_603,In_476);
nand U1306 (N_1306,In_1010,In_1102);
and U1307 (N_1307,In_1351,In_160);
or U1308 (N_1308,In_731,In_715);
xnor U1309 (N_1309,In_1365,In_729);
nand U1310 (N_1310,In_643,In_1008);
nand U1311 (N_1311,In_1484,In_404);
nand U1312 (N_1312,In_798,In_491);
nand U1313 (N_1313,In_1196,In_1084);
nor U1314 (N_1314,In_183,In_1346);
or U1315 (N_1315,In_404,In_671);
or U1316 (N_1316,In_226,In_664);
or U1317 (N_1317,In_710,In_905);
and U1318 (N_1318,In_167,In_479);
nand U1319 (N_1319,In_959,In_731);
nand U1320 (N_1320,In_12,In_318);
nor U1321 (N_1321,In_191,In_632);
nor U1322 (N_1322,In_416,In_921);
or U1323 (N_1323,In_1315,In_625);
and U1324 (N_1324,In_463,In_205);
nand U1325 (N_1325,In_1179,In_261);
or U1326 (N_1326,In_712,In_1168);
and U1327 (N_1327,In_1398,In_593);
or U1328 (N_1328,In_481,In_604);
nor U1329 (N_1329,In_835,In_944);
nand U1330 (N_1330,In_983,In_31);
nor U1331 (N_1331,In_1088,In_566);
and U1332 (N_1332,In_1218,In_622);
or U1333 (N_1333,In_1070,In_844);
or U1334 (N_1334,In_281,In_1292);
nand U1335 (N_1335,In_1129,In_1369);
or U1336 (N_1336,In_1219,In_447);
nor U1337 (N_1337,In_1328,In_1403);
nor U1338 (N_1338,In_458,In_1115);
or U1339 (N_1339,In_1326,In_170);
nor U1340 (N_1340,In_1031,In_673);
nor U1341 (N_1341,In_463,In_1329);
nand U1342 (N_1342,In_1249,In_764);
or U1343 (N_1343,In_378,In_873);
nand U1344 (N_1344,In_1481,In_1458);
and U1345 (N_1345,In_1287,In_44);
and U1346 (N_1346,In_1478,In_749);
or U1347 (N_1347,In_1453,In_329);
or U1348 (N_1348,In_558,In_1186);
or U1349 (N_1349,In_350,In_712);
nand U1350 (N_1350,In_560,In_504);
nand U1351 (N_1351,In_1394,In_397);
nand U1352 (N_1352,In_1434,In_1152);
and U1353 (N_1353,In_941,In_44);
and U1354 (N_1354,In_1419,In_289);
nand U1355 (N_1355,In_928,In_729);
nor U1356 (N_1356,In_561,In_854);
or U1357 (N_1357,In_909,In_976);
nor U1358 (N_1358,In_238,In_403);
and U1359 (N_1359,In_556,In_440);
and U1360 (N_1360,In_1262,In_581);
nand U1361 (N_1361,In_1316,In_1348);
and U1362 (N_1362,In_851,In_1088);
or U1363 (N_1363,In_441,In_300);
or U1364 (N_1364,In_1412,In_1044);
nand U1365 (N_1365,In_488,In_591);
or U1366 (N_1366,In_1479,In_1253);
nor U1367 (N_1367,In_141,In_181);
nor U1368 (N_1368,In_74,In_939);
nand U1369 (N_1369,In_1443,In_711);
nand U1370 (N_1370,In_39,In_561);
nand U1371 (N_1371,In_555,In_1472);
or U1372 (N_1372,In_1147,In_501);
and U1373 (N_1373,In_534,In_190);
nor U1374 (N_1374,In_1228,In_440);
nor U1375 (N_1375,In_1274,In_921);
nor U1376 (N_1376,In_555,In_846);
and U1377 (N_1377,In_258,In_350);
nand U1378 (N_1378,In_782,In_1216);
xor U1379 (N_1379,In_478,In_983);
or U1380 (N_1380,In_610,In_172);
nand U1381 (N_1381,In_86,In_1240);
nor U1382 (N_1382,In_563,In_1311);
or U1383 (N_1383,In_210,In_574);
and U1384 (N_1384,In_33,In_619);
or U1385 (N_1385,In_202,In_1333);
nor U1386 (N_1386,In_880,In_653);
nor U1387 (N_1387,In_547,In_978);
nand U1388 (N_1388,In_336,In_851);
nand U1389 (N_1389,In_867,In_857);
or U1390 (N_1390,In_1043,In_406);
or U1391 (N_1391,In_300,In_1244);
or U1392 (N_1392,In_859,In_845);
or U1393 (N_1393,In_1236,In_1382);
nand U1394 (N_1394,In_679,In_250);
or U1395 (N_1395,In_445,In_868);
nand U1396 (N_1396,In_620,In_638);
or U1397 (N_1397,In_1004,In_392);
and U1398 (N_1398,In_990,In_644);
and U1399 (N_1399,In_133,In_1482);
nor U1400 (N_1400,In_148,In_109);
and U1401 (N_1401,In_1312,In_1095);
xor U1402 (N_1402,In_521,In_1243);
or U1403 (N_1403,In_1074,In_1107);
and U1404 (N_1404,In_640,In_48);
and U1405 (N_1405,In_1217,In_1002);
nand U1406 (N_1406,In_766,In_959);
and U1407 (N_1407,In_1491,In_1417);
and U1408 (N_1408,In_810,In_179);
nor U1409 (N_1409,In_1075,In_469);
or U1410 (N_1410,In_801,In_518);
nor U1411 (N_1411,In_262,In_158);
nand U1412 (N_1412,In_1127,In_896);
nand U1413 (N_1413,In_1352,In_870);
nor U1414 (N_1414,In_420,In_372);
or U1415 (N_1415,In_902,In_621);
or U1416 (N_1416,In_905,In_1098);
and U1417 (N_1417,In_872,In_882);
or U1418 (N_1418,In_33,In_609);
nand U1419 (N_1419,In_377,In_1381);
or U1420 (N_1420,In_61,In_963);
nor U1421 (N_1421,In_350,In_1162);
nand U1422 (N_1422,In_1177,In_1049);
nand U1423 (N_1423,In_1435,In_626);
or U1424 (N_1424,In_1441,In_514);
nand U1425 (N_1425,In_41,In_1173);
nor U1426 (N_1426,In_1451,In_75);
nand U1427 (N_1427,In_230,In_331);
nor U1428 (N_1428,In_781,In_846);
or U1429 (N_1429,In_1310,In_268);
or U1430 (N_1430,In_248,In_837);
and U1431 (N_1431,In_374,In_897);
and U1432 (N_1432,In_25,In_1173);
nor U1433 (N_1433,In_339,In_379);
and U1434 (N_1434,In_1325,In_541);
and U1435 (N_1435,In_311,In_1035);
or U1436 (N_1436,In_1183,In_1232);
or U1437 (N_1437,In_868,In_471);
nor U1438 (N_1438,In_176,In_27);
nand U1439 (N_1439,In_1164,In_77);
nand U1440 (N_1440,In_403,In_1066);
or U1441 (N_1441,In_290,In_736);
nand U1442 (N_1442,In_75,In_112);
nor U1443 (N_1443,In_363,In_75);
nor U1444 (N_1444,In_1186,In_268);
and U1445 (N_1445,In_946,In_1299);
or U1446 (N_1446,In_617,In_407);
or U1447 (N_1447,In_353,In_915);
nand U1448 (N_1448,In_216,In_405);
nand U1449 (N_1449,In_1207,In_262);
nand U1450 (N_1450,In_645,In_903);
and U1451 (N_1451,In_1106,In_314);
and U1452 (N_1452,In_1295,In_1113);
nand U1453 (N_1453,In_1346,In_898);
and U1454 (N_1454,In_289,In_529);
or U1455 (N_1455,In_685,In_455);
or U1456 (N_1456,In_1319,In_834);
nor U1457 (N_1457,In_1100,In_1078);
nand U1458 (N_1458,In_687,In_986);
nor U1459 (N_1459,In_480,In_886);
and U1460 (N_1460,In_784,In_249);
nor U1461 (N_1461,In_1127,In_864);
and U1462 (N_1462,In_1108,In_752);
or U1463 (N_1463,In_1308,In_316);
nor U1464 (N_1464,In_768,In_1379);
nand U1465 (N_1465,In_817,In_270);
nor U1466 (N_1466,In_205,In_579);
or U1467 (N_1467,In_1347,In_574);
nor U1468 (N_1468,In_369,In_792);
or U1469 (N_1469,In_654,In_726);
nand U1470 (N_1470,In_202,In_511);
nand U1471 (N_1471,In_724,In_997);
nor U1472 (N_1472,In_739,In_1100);
or U1473 (N_1473,In_1044,In_774);
nor U1474 (N_1474,In_311,In_122);
nor U1475 (N_1475,In_13,In_620);
nor U1476 (N_1476,In_554,In_446);
and U1477 (N_1477,In_1156,In_1193);
or U1478 (N_1478,In_287,In_799);
and U1479 (N_1479,In_294,In_1459);
and U1480 (N_1480,In_842,In_433);
and U1481 (N_1481,In_323,In_977);
and U1482 (N_1482,In_560,In_467);
and U1483 (N_1483,In_989,In_1129);
nor U1484 (N_1484,In_100,In_1498);
nor U1485 (N_1485,In_1086,In_581);
and U1486 (N_1486,In_280,In_589);
and U1487 (N_1487,In_1181,In_226);
nor U1488 (N_1488,In_651,In_840);
or U1489 (N_1489,In_124,In_8);
nor U1490 (N_1490,In_1444,In_1065);
and U1491 (N_1491,In_480,In_791);
and U1492 (N_1492,In_911,In_1494);
or U1493 (N_1493,In_403,In_188);
nand U1494 (N_1494,In_321,In_455);
nand U1495 (N_1495,In_1276,In_887);
and U1496 (N_1496,In_1067,In_805);
nor U1497 (N_1497,In_322,In_1494);
and U1498 (N_1498,In_1194,In_1227);
and U1499 (N_1499,In_1037,In_83);
and U1500 (N_1500,In_1418,In_1278);
and U1501 (N_1501,In_1348,In_1088);
nor U1502 (N_1502,In_94,In_177);
nor U1503 (N_1503,In_38,In_807);
nand U1504 (N_1504,In_309,In_1183);
and U1505 (N_1505,In_507,In_323);
nand U1506 (N_1506,In_846,In_1122);
and U1507 (N_1507,In_572,In_1041);
and U1508 (N_1508,In_384,In_1092);
or U1509 (N_1509,In_1261,In_1453);
nand U1510 (N_1510,In_716,In_1098);
nor U1511 (N_1511,In_627,In_1357);
nor U1512 (N_1512,In_1493,In_33);
nor U1513 (N_1513,In_93,In_185);
or U1514 (N_1514,In_1457,In_1360);
nor U1515 (N_1515,In_250,In_784);
nand U1516 (N_1516,In_456,In_835);
or U1517 (N_1517,In_879,In_587);
and U1518 (N_1518,In_1485,In_1362);
or U1519 (N_1519,In_1098,In_603);
or U1520 (N_1520,In_1004,In_1276);
nand U1521 (N_1521,In_443,In_1001);
nor U1522 (N_1522,In_539,In_776);
or U1523 (N_1523,In_1304,In_704);
and U1524 (N_1524,In_1417,In_1182);
nand U1525 (N_1525,In_1270,In_89);
nor U1526 (N_1526,In_263,In_7);
nand U1527 (N_1527,In_1215,In_1389);
nand U1528 (N_1528,In_1278,In_330);
or U1529 (N_1529,In_1288,In_258);
and U1530 (N_1530,In_207,In_1177);
nand U1531 (N_1531,In_1083,In_937);
and U1532 (N_1532,In_471,In_1238);
or U1533 (N_1533,In_696,In_1354);
or U1534 (N_1534,In_355,In_1348);
or U1535 (N_1535,In_1301,In_1061);
nor U1536 (N_1536,In_1304,In_1357);
xnor U1537 (N_1537,In_398,In_617);
or U1538 (N_1538,In_648,In_283);
nor U1539 (N_1539,In_99,In_1418);
nor U1540 (N_1540,In_1257,In_258);
nand U1541 (N_1541,In_819,In_35);
nand U1542 (N_1542,In_411,In_232);
nor U1543 (N_1543,In_651,In_380);
nor U1544 (N_1544,In_744,In_1014);
nor U1545 (N_1545,In_716,In_552);
and U1546 (N_1546,In_646,In_288);
or U1547 (N_1547,In_502,In_564);
nor U1548 (N_1548,In_375,In_282);
nand U1549 (N_1549,In_966,In_187);
and U1550 (N_1550,In_646,In_314);
or U1551 (N_1551,In_1024,In_1377);
nand U1552 (N_1552,In_879,In_606);
nand U1553 (N_1553,In_1379,In_827);
and U1554 (N_1554,In_43,In_77);
nor U1555 (N_1555,In_110,In_1082);
nand U1556 (N_1556,In_1056,In_378);
nor U1557 (N_1557,In_828,In_550);
or U1558 (N_1558,In_1314,In_1319);
nand U1559 (N_1559,In_347,In_1470);
nor U1560 (N_1560,In_979,In_1250);
nor U1561 (N_1561,In_1299,In_81);
nor U1562 (N_1562,In_250,In_543);
and U1563 (N_1563,In_296,In_887);
nor U1564 (N_1564,In_23,In_1124);
and U1565 (N_1565,In_1021,In_182);
nor U1566 (N_1566,In_84,In_623);
or U1567 (N_1567,In_1028,In_871);
nor U1568 (N_1568,In_317,In_1454);
or U1569 (N_1569,In_880,In_1200);
nand U1570 (N_1570,In_227,In_656);
and U1571 (N_1571,In_1272,In_1211);
nand U1572 (N_1572,In_925,In_1134);
nor U1573 (N_1573,In_1325,In_787);
and U1574 (N_1574,In_735,In_990);
or U1575 (N_1575,In_1386,In_323);
nor U1576 (N_1576,In_1479,In_364);
nand U1577 (N_1577,In_730,In_724);
and U1578 (N_1578,In_427,In_839);
or U1579 (N_1579,In_16,In_1204);
or U1580 (N_1580,In_910,In_754);
and U1581 (N_1581,In_357,In_628);
and U1582 (N_1582,In_479,In_32);
nand U1583 (N_1583,In_139,In_1002);
and U1584 (N_1584,In_1276,In_1320);
nand U1585 (N_1585,In_76,In_641);
and U1586 (N_1586,In_984,In_861);
nand U1587 (N_1587,In_110,In_51);
and U1588 (N_1588,In_351,In_161);
or U1589 (N_1589,In_564,In_1221);
nor U1590 (N_1590,In_269,In_898);
nand U1591 (N_1591,In_532,In_860);
nand U1592 (N_1592,In_133,In_130);
nand U1593 (N_1593,In_152,In_805);
or U1594 (N_1594,In_0,In_66);
nor U1595 (N_1595,In_1454,In_1105);
and U1596 (N_1596,In_286,In_929);
and U1597 (N_1597,In_1241,In_1042);
and U1598 (N_1598,In_1131,In_1127);
and U1599 (N_1599,In_422,In_1019);
nor U1600 (N_1600,In_233,In_1350);
nor U1601 (N_1601,In_427,In_1400);
or U1602 (N_1602,In_212,In_233);
nor U1603 (N_1603,In_1174,In_9);
nand U1604 (N_1604,In_353,In_632);
nand U1605 (N_1605,In_648,In_237);
or U1606 (N_1606,In_567,In_336);
or U1607 (N_1607,In_1254,In_1486);
nor U1608 (N_1608,In_1418,In_1376);
and U1609 (N_1609,In_425,In_19);
or U1610 (N_1610,In_0,In_769);
or U1611 (N_1611,In_36,In_1287);
and U1612 (N_1612,In_953,In_808);
nor U1613 (N_1613,In_444,In_1439);
and U1614 (N_1614,In_1311,In_411);
nand U1615 (N_1615,In_411,In_1128);
nand U1616 (N_1616,In_416,In_117);
or U1617 (N_1617,In_770,In_344);
and U1618 (N_1618,In_863,In_886);
nor U1619 (N_1619,In_301,In_350);
nand U1620 (N_1620,In_561,In_733);
or U1621 (N_1621,In_368,In_1121);
or U1622 (N_1622,In_463,In_399);
nor U1623 (N_1623,In_885,In_1093);
or U1624 (N_1624,In_1201,In_1193);
nor U1625 (N_1625,In_219,In_655);
and U1626 (N_1626,In_1145,In_609);
nor U1627 (N_1627,In_823,In_564);
nor U1628 (N_1628,In_145,In_1347);
nand U1629 (N_1629,In_497,In_1101);
nor U1630 (N_1630,In_571,In_1209);
nor U1631 (N_1631,In_92,In_859);
or U1632 (N_1632,In_918,In_1446);
or U1633 (N_1633,In_60,In_231);
or U1634 (N_1634,In_922,In_820);
nand U1635 (N_1635,In_1292,In_1085);
or U1636 (N_1636,In_584,In_800);
nand U1637 (N_1637,In_366,In_1148);
nor U1638 (N_1638,In_757,In_1432);
nor U1639 (N_1639,In_582,In_39);
nand U1640 (N_1640,In_1464,In_889);
nor U1641 (N_1641,In_1074,In_560);
nor U1642 (N_1642,In_1106,In_762);
nor U1643 (N_1643,In_430,In_214);
or U1644 (N_1644,In_1149,In_777);
nor U1645 (N_1645,In_756,In_1079);
or U1646 (N_1646,In_1220,In_842);
nand U1647 (N_1647,In_189,In_252);
nor U1648 (N_1648,In_523,In_1429);
nor U1649 (N_1649,In_1357,In_40);
and U1650 (N_1650,In_1229,In_127);
nand U1651 (N_1651,In_239,In_1404);
nor U1652 (N_1652,In_147,In_521);
nand U1653 (N_1653,In_379,In_66);
or U1654 (N_1654,In_560,In_1424);
and U1655 (N_1655,In_350,In_66);
and U1656 (N_1656,In_45,In_183);
or U1657 (N_1657,In_1252,In_1341);
and U1658 (N_1658,In_812,In_1448);
nor U1659 (N_1659,In_470,In_930);
nor U1660 (N_1660,In_153,In_1350);
and U1661 (N_1661,In_1096,In_743);
nand U1662 (N_1662,In_1119,In_1232);
or U1663 (N_1663,In_767,In_507);
nor U1664 (N_1664,In_754,In_627);
or U1665 (N_1665,In_439,In_1361);
nor U1666 (N_1666,In_874,In_661);
or U1667 (N_1667,In_68,In_1371);
nand U1668 (N_1668,In_769,In_697);
nor U1669 (N_1669,In_502,In_1134);
nor U1670 (N_1670,In_960,In_232);
nor U1671 (N_1671,In_1299,In_406);
or U1672 (N_1672,In_824,In_1417);
nand U1673 (N_1673,In_1309,In_259);
or U1674 (N_1674,In_833,In_936);
or U1675 (N_1675,In_284,In_1478);
nor U1676 (N_1676,In_604,In_751);
nand U1677 (N_1677,In_781,In_203);
and U1678 (N_1678,In_517,In_124);
and U1679 (N_1679,In_924,In_671);
nor U1680 (N_1680,In_186,In_770);
or U1681 (N_1681,In_37,In_164);
nand U1682 (N_1682,In_1116,In_973);
nor U1683 (N_1683,In_460,In_972);
nor U1684 (N_1684,In_693,In_1219);
and U1685 (N_1685,In_1443,In_743);
or U1686 (N_1686,In_389,In_1419);
or U1687 (N_1687,In_1474,In_9);
nand U1688 (N_1688,In_1216,In_535);
nor U1689 (N_1689,In_479,In_456);
nor U1690 (N_1690,In_297,In_974);
or U1691 (N_1691,In_502,In_1256);
and U1692 (N_1692,In_389,In_892);
nand U1693 (N_1693,In_580,In_460);
nor U1694 (N_1694,In_1264,In_512);
or U1695 (N_1695,In_119,In_367);
nor U1696 (N_1696,In_27,In_750);
or U1697 (N_1697,In_80,In_1474);
or U1698 (N_1698,In_1305,In_1055);
nor U1699 (N_1699,In_259,In_35);
and U1700 (N_1700,In_643,In_104);
or U1701 (N_1701,In_281,In_1177);
and U1702 (N_1702,In_741,In_1378);
nor U1703 (N_1703,In_1104,In_262);
nand U1704 (N_1704,In_22,In_818);
or U1705 (N_1705,In_1488,In_779);
nor U1706 (N_1706,In_1213,In_820);
or U1707 (N_1707,In_849,In_1064);
nand U1708 (N_1708,In_1060,In_1113);
or U1709 (N_1709,In_265,In_525);
nand U1710 (N_1710,In_319,In_626);
nor U1711 (N_1711,In_424,In_214);
nor U1712 (N_1712,In_1258,In_864);
nand U1713 (N_1713,In_818,In_530);
nor U1714 (N_1714,In_636,In_775);
nor U1715 (N_1715,In_1451,In_688);
or U1716 (N_1716,In_606,In_131);
and U1717 (N_1717,In_215,In_982);
nor U1718 (N_1718,In_1303,In_458);
nor U1719 (N_1719,In_590,In_85);
or U1720 (N_1720,In_1166,In_401);
xor U1721 (N_1721,In_365,In_1126);
xor U1722 (N_1722,In_1366,In_879);
and U1723 (N_1723,In_184,In_266);
nor U1724 (N_1724,In_913,In_1118);
or U1725 (N_1725,In_599,In_1145);
and U1726 (N_1726,In_1194,In_43);
and U1727 (N_1727,In_1383,In_1018);
or U1728 (N_1728,In_627,In_1285);
nor U1729 (N_1729,In_706,In_378);
nand U1730 (N_1730,In_426,In_1040);
and U1731 (N_1731,In_681,In_1295);
and U1732 (N_1732,In_984,In_89);
nand U1733 (N_1733,In_588,In_1393);
nand U1734 (N_1734,In_446,In_661);
and U1735 (N_1735,In_942,In_213);
nand U1736 (N_1736,In_119,In_501);
or U1737 (N_1737,In_210,In_255);
and U1738 (N_1738,In_1421,In_1075);
or U1739 (N_1739,In_683,In_998);
xnor U1740 (N_1740,In_719,In_1025);
nor U1741 (N_1741,In_233,In_706);
and U1742 (N_1742,In_1177,In_470);
or U1743 (N_1743,In_1352,In_82);
nor U1744 (N_1744,In_856,In_1160);
and U1745 (N_1745,In_1390,In_1480);
nor U1746 (N_1746,In_493,In_661);
nand U1747 (N_1747,In_78,In_332);
or U1748 (N_1748,In_1354,In_73);
nor U1749 (N_1749,In_666,In_827);
nor U1750 (N_1750,In_1213,In_143);
or U1751 (N_1751,In_486,In_814);
nor U1752 (N_1752,In_1268,In_652);
and U1753 (N_1753,In_1234,In_945);
or U1754 (N_1754,In_744,In_1393);
nand U1755 (N_1755,In_855,In_759);
nor U1756 (N_1756,In_452,In_984);
nor U1757 (N_1757,In_841,In_488);
nand U1758 (N_1758,In_724,In_48);
or U1759 (N_1759,In_1102,In_1250);
nor U1760 (N_1760,In_809,In_1095);
nor U1761 (N_1761,In_1393,In_155);
or U1762 (N_1762,In_651,In_216);
or U1763 (N_1763,In_904,In_1405);
nand U1764 (N_1764,In_624,In_105);
nand U1765 (N_1765,In_394,In_539);
nor U1766 (N_1766,In_45,In_1184);
nand U1767 (N_1767,In_441,In_333);
nor U1768 (N_1768,In_1103,In_317);
nor U1769 (N_1769,In_387,In_1224);
or U1770 (N_1770,In_526,In_1374);
and U1771 (N_1771,In_570,In_528);
and U1772 (N_1772,In_318,In_158);
and U1773 (N_1773,In_212,In_1342);
nand U1774 (N_1774,In_993,In_1288);
or U1775 (N_1775,In_609,In_814);
nand U1776 (N_1776,In_866,In_1486);
or U1777 (N_1777,In_1038,In_94);
or U1778 (N_1778,In_439,In_711);
nor U1779 (N_1779,In_1054,In_964);
nand U1780 (N_1780,In_545,In_1224);
or U1781 (N_1781,In_39,In_1379);
nor U1782 (N_1782,In_1077,In_272);
or U1783 (N_1783,In_1282,In_581);
and U1784 (N_1784,In_2,In_1111);
nand U1785 (N_1785,In_1054,In_639);
or U1786 (N_1786,In_513,In_844);
and U1787 (N_1787,In_275,In_1272);
nand U1788 (N_1788,In_269,In_324);
and U1789 (N_1789,In_739,In_1125);
or U1790 (N_1790,In_597,In_1158);
and U1791 (N_1791,In_772,In_305);
and U1792 (N_1792,In_1033,In_818);
nor U1793 (N_1793,In_1496,In_1359);
or U1794 (N_1794,In_1337,In_969);
and U1795 (N_1795,In_1092,In_44);
or U1796 (N_1796,In_412,In_894);
nand U1797 (N_1797,In_998,In_333);
and U1798 (N_1798,In_1009,In_1092);
nor U1799 (N_1799,In_1310,In_1044);
or U1800 (N_1800,In_1032,In_161);
or U1801 (N_1801,In_219,In_627);
nor U1802 (N_1802,In_848,In_863);
nor U1803 (N_1803,In_284,In_699);
or U1804 (N_1804,In_716,In_645);
nand U1805 (N_1805,In_643,In_1175);
and U1806 (N_1806,In_1427,In_181);
nor U1807 (N_1807,In_341,In_1022);
nand U1808 (N_1808,In_601,In_345);
or U1809 (N_1809,In_426,In_946);
nand U1810 (N_1810,In_1394,In_1390);
nand U1811 (N_1811,In_668,In_328);
or U1812 (N_1812,In_270,In_461);
and U1813 (N_1813,In_418,In_156);
or U1814 (N_1814,In_1107,In_716);
nand U1815 (N_1815,In_819,In_249);
or U1816 (N_1816,In_288,In_902);
nand U1817 (N_1817,In_745,In_215);
nand U1818 (N_1818,In_660,In_535);
nand U1819 (N_1819,In_1323,In_1156);
or U1820 (N_1820,In_1205,In_620);
and U1821 (N_1821,In_841,In_481);
or U1822 (N_1822,In_410,In_596);
nor U1823 (N_1823,In_359,In_179);
nor U1824 (N_1824,In_169,In_1455);
and U1825 (N_1825,In_608,In_1357);
nand U1826 (N_1826,In_58,In_956);
or U1827 (N_1827,In_1101,In_891);
nand U1828 (N_1828,In_1363,In_618);
nand U1829 (N_1829,In_885,In_963);
or U1830 (N_1830,In_80,In_255);
nand U1831 (N_1831,In_1455,In_378);
and U1832 (N_1832,In_141,In_655);
nand U1833 (N_1833,In_1195,In_1220);
and U1834 (N_1834,In_763,In_1470);
or U1835 (N_1835,In_924,In_1418);
or U1836 (N_1836,In_442,In_1069);
and U1837 (N_1837,In_1498,In_842);
and U1838 (N_1838,In_565,In_1240);
or U1839 (N_1839,In_1161,In_746);
and U1840 (N_1840,In_619,In_156);
nand U1841 (N_1841,In_1390,In_960);
and U1842 (N_1842,In_921,In_662);
nand U1843 (N_1843,In_73,In_946);
nand U1844 (N_1844,In_345,In_682);
or U1845 (N_1845,In_1412,In_1469);
nand U1846 (N_1846,In_534,In_915);
or U1847 (N_1847,In_1312,In_649);
or U1848 (N_1848,In_231,In_637);
and U1849 (N_1849,In_461,In_348);
nand U1850 (N_1850,In_1136,In_703);
nor U1851 (N_1851,In_1250,In_1392);
and U1852 (N_1852,In_926,In_617);
and U1853 (N_1853,In_770,In_751);
and U1854 (N_1854,In_261,In_279);
and U1855 (N_1855,In_1473,In_497);
and U1856 (N_1856,In_60,In_850);
nand U1857 (N_1857,In_1236,In_180);
nand U1858 (N_1858,In_592,In_191);
nand U1859 (N_1859,In_1183,In_1269);
and U1860 (N_1860,In_473,In_298);
nand U1861 (N_1861,In_1483,In_1076);
and U1862 (N_1862,In_89,In_530);
and U1863 (N_1863,In_1199,In_461);
or U1864 (N_1864,In_640,In_1323);
and U1865 (N_1865,In_1249,In_1279);
or U1866 (N_1866,In_676,In_410);
and U1867 (N_1867,In_1193,In_1336);
or U1868 (N_1868,In_119,In_1176);
or U1869 (N_1869,In_559,In_596);
nor U1870 (N_1870,In_742,In_242);
nor U1871 (N_1871,In_311,In_954);
or U1872 (N_1872,In_801,In_705);
nand U1873 (N_1873,In_532,In_915);
or U1874 (N_1874,In_1340,In_68);
nor U1875 (N_1875,In_1348,In_1496);
or U1876 (N_1876,In_774,In_307);
nor U1877 (N_1877,In_1029,In_863);
and U1878 (N_1878,In_1138,In_868);
or U1879 (N_1879,In_1495,In_8);
nor U1880 (N_1880,In_1073,In_832);
and U1881 (N_1881,In_322,In_1293);
or U1882 (N_1882,In_1139,In_1098);
nor U1883 (N_1883,In_1189,In_1092);
and U1884 (N_1884,In_531,In_492);
nand U1885 (N_1885,In_741,In_1349);
and U1886 (N_1886,In_787,In_1283);
nor U1887 (N_1887,In_1132,In_1190);
nor U1888 (N_1888,In_1116,In_147);
nor U1889 (N_1889,In_40,In_344);
or U1890 (N_1890,In_385,In_392);
and U1891 (N_1891,In_342,In_408);
and U1892 (N_1892,In_1229,In_837);
nand U1893 (N_1893,In_145,In_214);
xor U1894 (N_1894,In_337,In_57);
nor U1895 (N_1895,In_740,In_189);
or U1896 (N_1896,In_190,In_75);
nand U1897 (N_1897,In_588,In_262);
nor U1898 (N_1898,In_1373,In_721);
nand U1899 (N_1899,In_1234,In_1010);
nor U1900 (N_1900,In_195,In_1182);
or U1901 (N_1901,In_1486,In_505);
and U1902 (N_1902,In_1118,In_268);
or U1903 (N_1903,In_1450,In_594);
nand U1904 (N_1904,In_662,In_862);
nand U1905 (N_1905,In_1473,In_1471);
nor U1906 (N_1906,In_602,In_1162);
and U1907 (N_1907,In_1326,In_1406);
nor U1908 (N_1908,In_929,In_790);
nand U1909 (N_1909,In_725,In_1402);
or U1910 (N_1910,In_1099,In_450);
nand U1911 (N_1911,In_1127,In_798);
or U1912 (N_1912,In_315,In_928);
nor U1913 (N_1913,In_283,In_304);
nand U1914 (N_1914,In_566,In_1045);
or U1915 (N_1915,In_734,In_1436);
and U1916 (N_1916,In_10,In_793);
or U1917 (N_1917,In_598,In_938);
nand U1918 (N_1918,In_167,In_849);
or U1919 (N_1919,In_164,In_663);
xor U1920 (N_1920,In_1420,In_749);
and U1921 (N_1921,In_307,In_1332);
or U1922 (N_1922,In_754,In_1001);
and U1923 (N_1923,In_1064,In_992);
nand U1924 (N_1924,In_129,In_395);
nand U1925 (N_1925,In_376,In_1437);
nor U1926 (N_1926,In_903,In_486);
nor U1927 (N_1927,In_826,In_703);
nand U1928 (N_1928,In_752,In_40);
nor U1929 (N_1929,In_1187,In_1361);
or U1930 (N_1930,In_1491,In_1399);
nand U1931 (N_1931,In_163,In_921);
nor U1932 (N_1932,In_622,In_897);
nand U1933 (N_1933,In_1426,In_946);
nand U1934 (N_1934,In_1363,In_1306);
nand U1935 (N_1935,In_594,In_365);
and U1936 (N_1936,In_1323,In_540);
or U1937 (N_1937,In_909,In_1034);
nand U1938 (N_1938,In_952,In_856);
or U1939 (N_1939,In_863,In_256);
or U1940 (N_1940,In_450,In_957);
nand U1941 (N_1941,In_568,In_145);
nor U1942 (N_1942,In_76,In_1035);
nor U1943 (N_1943,In_1094,In_18);
or U1944 (N_1944,In_265,In_1374);
nor U1945 (N_1945,In_1042,In_116);
nor U1946 (N_1946,In_819,In_675);
or U1947 (N_1947,In_1493,In_357);
or U1948 (N_1948,In_906,In_11);
or U1949 (N_1949,In_624,In_577);
or U1950 (N_1950,In_1207,In_1153);
and U1951 (N_1951,In_1101,In_1032);
and U1952 (N_1952,In_301,In_414);
and U1953 (N_1953,In_801,In_1411);
nand U1954 (N_1954,In_775,In_415);
nand U1955 (N_1955,In_980,In_735);
nand U1956 (N_1956,In_361,In_1057);
or U1957 (N_1957,In_862,In_416);
nand U1958 (N_1958,In_822,In_1049);
nand U1959 (N_1959,In_1335,In_137);
nand U1960 (N_1960,In_170,In_652);
and U1961 (N_1961,In_1473,In_1334);
nand U1962 (N_1962,In_1060,In_1016);
and U1963 (N_1963,In_954,In_451);
nor U1964 (N_1964,In_662,In_737);
xnor U1965 (N_1965,In_711,In_303);
nand U1966 (N_1966,In_499,In_1348);
nand U1967 (N_1967,In_94,In_1332);
nor U1968 (N_1968,In_275,In_573);
xnor U1969 (N_1969,In_51,In_865);
nor U1970 (N_1970,In_493,In_1429);
or U1971 (N_1971,In_253,In_38);
or U1972 (N_1972,In_799,In_897);
and U1973 (N_1973,In_713,In_487);
nand U1974 (N_1974,In_720,In_1049);
nand U1975 (N_1975,In_1156,In_559);
nor U1976 (N_1976,In_881,In_748);
or U1977 (N_1977,In_115,In_985);
and U1978 (N_1978,In_1074,In_2);
nand U1979 (N_1979,In_48,In_81);
nor U1980 (N_1980,In_888,In_458);
nand U1981 (N_1981,In_845,In_1419);
and U1982 (N_1982,In_736,In_927);
and U1983 (N_1983,In_480,In_1368);
and U1984 (N_1984,In_110,In_49);
or U1985 (N_1985,In_1447,In_95);
nor U1986 (N_1986,In_967,In_777);
and U1987 (N_1987,In_1492,In_145);
or U1988 (N_1988,In_1348,In_300);
nor U1989 (N_1989,In_265,In_1424);
or U1990 (N_1990,In_314,In_653);
or U1991 (N_1991,In_1026,In_1236);
or U1992 (N_1992,In_1414,In_277);
nor U1993 (N_1993,In_173,In_943);
and U1994 (N_1994,In_467,In_793);
nand U1995 (N_1995,In_326,In_729);
xor U1996 (N_1996,In_108,In_85);
and U1997 (N_1997,In_1483,In_1126);
and U1998 (N_1998,In_1211,In_437);
nand U1999 (N_1999,In_321,In_435);
or U2000 (N_2000,In_973,In_218);
nand U2001 (N_2001,In_1359,In_52);
or U2002 (N_2002,In_92,In_206);
nand U2003 (N_2003,In_1237,In_128);
nand U2004 (N_2004,In_125,In_368);
nor U2005 (N_2005,In_1272,In_596);
or U2006 (N_2006,In_732,In_773);
and U2007 (N_2007,In_163,In_611);
and U2008 (N_2008,In_153,In_1189);
nand U2009 (N_2009,In_437,In_461);
and U2010 (N_2010,In_1421,In_560);
or U2011 (N_2011,In_965,In_1362);
and U2012 (N_2012,In_1129,In_1091);
or U2013 (N_2013,In_1457,In_202);
or U2014 (N_2014,In_1234,In_970);
xor U2015 (N_2015,In_646,In_55);
nor U2016 (N_2016,In_648,In_398);
nor U2017 (N_2017,In_1023,In_229);
nor U2018 (N_2018,In_912,In_153);
or U2019 (N_2019,In_186,In_903);
and U2020 (N_2020,In_272,In_1150);
and U2021 (N_2021,In_1381,In_23);
nor U2022 (N_2022,In_962,In_227);
and U2023 (N_2023,In_261,In_136);
nand U2024 (N_2024,In_1296,In_664);
nand U2025 (N_2025,In_430,In_1484);
nand U2026 (N_2026,In_1034,In_1153);
nand U2027 (N_2027,In_1355,In_304);
nor U2028 (N_2028,In_744,In_1170);
nand U2029 (N_2029,In_348,In_1340);
and U2030 (N_2030,In_254,In_38);
or U2031 (N_2031,In_334,In_1106);
and U2032 (N_2032,In_462,In_833);
nand U2033 (N_2033,In_1425,In_1447);
xnor U2034 (N_2034,In_1319,In_1234);
and U2035 (N_2035,In_1261,In_485);
and U2036 (N_2036,In_39,In_1424);
nand U2037 (N_2037,In_306,In_88);
or U2038 (N_2038,In_1407,In_370);
or U2039 (N_2039,In_469,In_389);
and U2040 (N_2040,In_1351,In_424);
nand U2041 (N_2041,In_1119,In_790);
or U2042 (N_2042,In_1499,In_1477);
nand U2043 (N_2043,In_1230,In_1425);
nor U2044 (N_2044,In_1025,In_1337);
and U2045 (N_2045,In_235,In_458);
nor U2046 (N_2046,In_353,In_919);
nand U2047 (N_2047,In_1256,In_1469);
nor U2048 (N_2048,In_979,In_1490);
xnor U2049 (N_2049,In_100,In_851);
and U2050 (N_2050,In_808,In_899);
nor U2051 (N_2051,In_1146,In_146);
and U2052 (N_2052,In_226,In_1434);
nor U2053 (N_2053,In_821,In_1275);
nor U2054 (N_2054,In_529,In_26);
and U2055 (N_2055,In_1075,In_1073);
and U2056 (N_2056,In_1007,In_524);
or U2057 (N_2057,In_725,In_1323);
and U2058 (N_2058,In_513,In_23);
and U2059 (N_2059,In_1240,In_1066);
or U2060 (N_2060,In_1089,In_925);
nor U2061 (N_2061,In_596,In_1216);
nand U2062 (N_2062,In_423,In_1372);
nor U2063 (N_2063,In_1290,In_196);
nor U2064 (N_2064,In_1421,In_678);
xnor U2065 (N_2065,In_1100,In_824);
and U2066 (N_2066,In_955,In_42);
and U2067 (N_2067,In_1452,In_184);
or U2068 (N_2068,In_143,In_125);
nand U2069 (N_2069,In_557,In_870);
nand U2070 (N_2070,In_661,In_1042);
or U2071 (N_2071,In_142,In_90);
or U2072 (N_2072,In_1092,In_744);
nor U2073 (N_2073,In_931,In_1474);
nand U2074 (N_2074,In_390,In_659);
nand U2075 (N_2075,In_515,In_797);
or U2076 (N_2076,In_1102,In_311);
nand U2077 (N_2077,In_823,In_1274);
and U2078 (N_2078,In_1138,In_873);
or U2079 (N_2079,In_1374,In_676);
nor U2080 (N_2080,In_517,In_724);
and U2081 (N_2081,In_716,In_1270);
nand U2082 (N_2082,In_671,In_98);
and U2083 (N_2083,In_434,In_91);
nand U2084 (N_2084,In_1294,In_790);
and U2085 (N_2085,In_464,In_654);
or U2086 (N_2086,In_672,In_192);
and U2087 (N_2087,In_932,In_499);
or U2088 (N_2088,In_1360,In_301);
and U2089 (N_2089,In_508,In_929);
and U2090 (N_2090,In_464,In_865);
nand U2091 (N_2091,In_733,In_173);
and U2092 (N_2092,In_697,In_1482);
nor U2093 (N_2093,In_142,In_405);
nor U2094 (N_2094,In_872,In_1375);
or U2095 (N_2095,In_861,In_2);
or U2096 (N_2096,In_1295,In_831);
or U2097 (N_2097,In_1402,In_461);
nand U2098 (N_2098,In_727,In_1350);
and U2099 (N_2099,In_494,In_585);
nand U2100 (N_2100,In_1499,In_1229);
and U2101 (N_2101,In_1454,In_227);
and U2102 (N_2102,In_886,In_1113);
nor U2103 (N_2103,In_1333,In_1471);
or U2104 (N_2104,In_243,In_498);
or U2105 (N_2105,In_737,In_1318);
nand U2106 (N_2106,In_578,In_1353);
or U2107 (N_2107,In_118,In_967);
nand U2108 (N_2108,In_944,In_310);
nor U2109 (N_2109,In_1441,In_1415);
nand U2110 (N_2110,In_1358,In_419);
nand U2111 (N_2111,In_90,In_292);
and U2112 (N_2112,In_33,In_53);
nand U2113 (N_2113,In_219,In_373);
or U2114 (N_2114,In_1180,In_883);
or U2115 (N_2115,In_1164,In_823);
or U2116 (N_2116,In_1096,In_1401);
nor U2117 (N_2117,In_1386,In_953);
nand U2118 (N_2118,In_34,In_1232);
or U2119 (N_2119,In_1136,In_1356);
nor U2120 (N_2120,In_667,In_989);
and U2121 (N_2121,In_916,In_317);
nor U2122 (N_2122,In_1099,In_291);
or U2123 (N_2123,In_1012,In_845);
nor U2124 (N_2124,In_1005,In_982);
nor U2125 (N_2125,In_1061,In_1371);
nor U2126 (N_2126,In_1088,In_1021);
or U2127 (N_2127,In_496,In_187);
or U2128 (N_2128,In_6,In_308);
nor U2129 (N_2129,In_1278,In_932);
and U2130 (N_2130,In_972,In_1254);
nor U2131 (N_2131,In_950,In_1177);
or U2132 (N_2132,In_1313,In_1045);
and U2133 (N_2133,In_1151,In_288);
nand U2134 (N_2134,In_488,In_146);
nand U2135 (N_2135,In_904,In_1449);
nand U2136 (N_2136,In_1026,In_300);
or U2137 (N_2137,In_965,In_767);
or U2138 (N_2138,In_691,In_614);
or U2139 (N_2139,In_664,In_589);
nand U2140 (N_2140,In_647,In_581);
xor U2141 (N_2141,In_358,In_1257);
nor U2142 (N_2142,In_738,In_956);
and U2143 (N_2143,In_660,In_1193);
nand U2144 (N_2144,In_252,In_1203);
and U2145 (N_2145,In_486,In_1308);
nand U2146 (N_2146,In_377,In_164);
nand U2147 (N_2147,In_1381,In_1177);
nand U2148 (N_2148,In_191,In_1233);
nand U2149 (N_2149,In_489,In_433);
nor U2150 (N_2150,In_155,In_749);
nand U2151 (N_2151,In_335,In_1438);
or U2152 (N_2152,In_132,In_1194);
or U2153 (N_2153,In_274,In_275);
and U2154 (N_2154,In_1369,In_196);
or U2155 (N_2155,In_901,In_596);
or U2156 (N_2156,In_397,In_947);
or U2157 (N_2157,In_294,In_473);
nand U2158 (N_2158,In_1408,In_1214);
nor U2159 (N_2159,In_894,In_1320);
nor U2160 (N_2160,In_910,In_1188);
nand U2161 (N_2161,In_40,In_1302);
or U2162 (N_2162,In_781,In_461);
nand U2163 (N_2163,In_381,In_1276);
nor U2164 (N_2164,In_1049,In_1352);
nand U2165 (N_2165,In_998,In_414);
or U2166 (N_2166,In_1357,In_690);
and U2167 (N_2167,In_148,In_578);
nor U2168 (N_2168,In_444,In_260);
or U2169 (N_2169,In_279,In_149);
nand U2170 (N_2170,In_1040,In_923);
nand U2171 (N_2171,In_1355,In_1463);
nand U2172 (N_2172,In_1403,In_1130);
and U2173 (N_2173,In_227,In_1491);
and U2174 (N_2174,In_1406,In_26);
and U2175 (N_2175,In_1027,In_849);
and U2176 (N_2176,In_564,In_89);
nor U2177 (N_2177,In_1072,In_99);
or U2178 (N_2178,In_657,In_1471);
or U2179 (N_2179,In_176,In_1097);
nor U2180 (N_2180,In_194,In_1089);
and U2181 (N_2181,In_1387,In_278);
or U2182 (N_2182,In_1039,In_49);
nand U2183 (N_2183,In_384,In_1160);
or U2184 (N_2184,In_540,In_1485);
nand U2185 (N_2185,In_220,In_551);
and U2186 (N_2186,In_375,In_177);
and U2187 (N_2187,In_512,In_308);
or U2188 (N_2188,In_1404,In_1339);
or U2189 (N_2189,In_1126,In_327);
nor U2190 (N_2190,In_1295,In_1496);
or U2191 (N_2191,In_980,In_918);
nor U2192 (N_2192,In_676,In_1212);
or U2193 (N_2193,In_490,In_579);
nand U2194 (N_2194,In_1436,In_448);
or U2195 (N_2195,In_1115,In_1494);
nand U2196 (N_2196,In_889,In_1089);
nand U2197 (N_2197,In_989,In_1148);
or U2198 (N_2198,In_76,In_338);
or U2199 (N_2199,In_880,In_740);
or U2200 (N_2200,In_113,In_964);
nand U2201 (N_2201,In_1092,In_1242);
or U2202 (N_2202,In_40,In_643);
nand U2203 (N_2203,In_1026,In_734);
and U2204 (N_2204,In_1176,In_593);
or U2205 (N_2205,In_854,In_894);
nor U2206 (N_2206,In_1188,In_301);
nand U2207 (N_2207,In_1337,In_603);
nand U2208 (N_2208,In_1355,In_424);
xnor U2209 (N_2209,In_1362,In_1240);
nor U2210 (N_2210,In_611,In_1263);
and U2211 (N_2211,In_1414,In_364);
and U2212 (N_2212,In_1190,In_682);
or U2213 (N_2213,In_167,In_888);
nor U2214 (N_2214,In_651,In_306);
nor U2215 (N_2215,In_85,In_1339);
and U2216 (N_2216,In_1169,In_164);
and U2217 (N_2217,In_536,In_516);
and U2218 (N_2218,In_723,In_232);
nand U2219 (N_2219,In_299,In_1024);
and U2220 (N_2220,In_169,In_819);
nand U2221 (N_2221,In_219,In_97);
and U2222 (N_2222,In_90,In_998);
nand U2223 (N_2223,In_810,In_97);
and U2224 (N_2224,In_56,In_433);
and U2225 (N_2225,In_1021,In_1293);
or U2226 (N_2226,In_593,In_1497);
and U2227 (N_2227,In_1084,In_824);
nor U2228 (N_2228,In_375,In_135);
nor U2229 (N_2229,In_1286,In_989);
and U2230 (N_2230,In_198,In_1209);
or U2231 (N_2231,In_1037,In_1193);
nand U2232 (N_2232,In_1373,In_337);
nand U2233 (N_2233,In_408,In_155);
nand U2234 (N_2234,In_515,In_820);
or U2235 (N_2235,In_877,In_747);
or U2236 (N_2236,In_1034,In_344);
nor U2237 (N_2237,In_1357,In_1131);
and U2238 (N_2238,In_1120,In_40);
or U2239 (N_2239,In_106,In_127);
or U2240 (N_2240,In_482,In_1037);
nor U2241 (N_2241,In_597,In_1277);
nor U2242 (N_2242,In_1425,In_577);
nand U2243 (N_2243,In_645,In_1371);
nor U2244 (N_2244,In_496,In_153);
or U2245 (N_2245,In_1455,In_1328);
nor U2246 (N_2246,In_1026,In_711);
nor U2247 (N_2247,In_213,In_95);
and U2248 (N_2248,In_109,In_665);
and U2249 (N_2249,In_743,In_25);
nand U2250 (N_2250,In_565,In_875);
or U2251 (N_2251,In_1043,In_435);
or U2252 (N_2252,In_187,In_273);
nand U2253 (N_2253,In_490,In_781);
or U2254 (N_2254,In_148,In_1420);
nor U2255 (N_2255,In_574,In_1446);
nor U2256 (N_2256,In_1114,In_1259);
or U2257 (N_2257,In_503,In_1236);
and U2258 (N_2258,In_253,In_1129);
and U2259 (N_2259,In_262,In_293);
nor U2260 (N_2260,In_1022,In_0);
or U2261 (N_2261,In_402,In_1076);
nor U2262 (N_2262,In_1322,In_27);
and U2263 (N_2263,In_516,In_762);
nor U2264 (N_2264,In_54,In_501);
nor U2265 (N_2265,In_1213,In_1495);
nor U2266 (N_2266,In_734,In_666);
or U2267 (N_2267,In_979,In_227);
nand U2268 (N_2268,In_65,In_1090);
nor U2269 (N_2269,In_1032,In_1337);
and U2270 (N_2270,In_546,In_124);
and U2271 (N_2271,In_183,In_565);
or U2272 (N_2272,In_1303,In_866);
nand U2273 (N_2273,In_830,In_680);
or U2274 (N_2274,In_753,In_1019);
nor U2275 (N_2275,In_624,In_775);
nand U2276 (N_2276,In_494,In_1392);
or U2277 (N_2277,In_527,In_232);
and U2278 (N_2278,In_483,In_1240);
or U2279 (N_2279,In_1115,In_1384);
nor U2280 (N_2280,In_545,In_1275);
and U2281 (N_2281,In_252,In_715);
and U2282 (N_2282,In_342,In_1464);
nor U2283 (N_2283,In_449,In_1253);
nor U2284 (N_2284,In_908,In_963);
and U2285 (N_2285,In_1427,In_435);
nand U2286 (N_2286,In_595,In_1465);
or U2287 (N_2287,In_132,In_363);
or U2288 (N_2288,In_218,In_984);
or U2289 (N_2289,In_177,In_1003);
nand U2290 (N_2290,In_1003,In_1032);
nor U2291 (N_2291,In_83,In_1179);
nor U2292 (N_2292,In_1057,In_572);
xor U2293 (N_2293,In_1089,In_1146);
or U2294 (N_2294,In_477,In_743);
nor U2295 (N_2295,In_1312,In_509);
and U2296 (N_2296,In_552,In_919);
or U2297 (N_2297,In_137,In_109);
or U2298 (N_2298,In_556,In_745);
and U2299 (N_2299,In_407,In_723);
and U2300 (N_2300,In_1092,In_1305);
nor U2301 (N_2301,In_746,In_117);
nor U2302 (N_2302,In_584,In_196);
and U2303 (N_2303,In_72,In_877);
nand U2304 (N_2304,In_488,In_1046);
or U2305 (N_2305,In_1191,In_1460);
or U2306 (N_2306,In_359,In_1219);
xnor U2307 (N_2307,In_1032,In_947);
nand U2308 (N_2308,In_1364,In_1218);
and U2309 (N_2309,In_392,In_532);
nand U2310 (N_2310,In_1297,In_250);
and U2311 (N_2311,In_746,In_540);
nand U2312 (N_2312,In_551,In_1443);
or U2313 (N_2313,In_725,In_1270);
nand U2314 (N_2314,In_767,In_998);
or U2315 (N_2315,In_27,In_1114);
nand U2316 (N_2316,In_695,In_498);
xnor U2317 (N_2317,In_1479,In_163);
nand U2318 (N_2318,In_404,In_199);
or U2319 (N_2319,In_76,In_189);
and U2320 (N_2320,In_399,In_277);
nand U2321 (N_2321,In_1213,In_828);
nor U2322 (N_2322,In_828,In_33);
nor U2323 (N_2323,In_1197,In_993);
nor U2324 (N_2324,In_1449,In_491);
and U2325 (N_2325,In_976,In_257);
or U2326 (N_2326,In_480,In_15);
and U2327 (N_2327,In_807,In_966);
nand U2328 (N_2328,In_507,In_1173);
or U2329 (N_2329,In_552,In_25);
nand U2330 (N_2330,In_1278,In_1092);
and U2331 (N_2331,In_942,In_904);
and U2332 (N_2332,In_45,In_664);
or U2333 (N_2333,In_352,In_1377);
nand U2334 (N_2334,In_454,In_850);
nand U2335 (N_2335,In_798,In_186);
nand U2336 (N_2336,In_1451,In_302);
and U2337 (N_2337,In_999,In_48);
nand U2338 (N_2338,In_395,In_543);
nor U2339 (N_2339,In_1082,In_1162);
and U2340 (N_2340,In_1369,In_1424);
or U2341 (N_2341,In_1334,In_669);
nand U2342 (N_2342,In_881,In_636);
xor U2343 (N_2343,In_1280,In_1110);
nand U2344 (N_2344,In_266,In_469);
nand U2345 (N_2345,In_1262,In_1465);
nor U2346 (N_2346,In_613,In_1352);
nand U2347 (N_2347,In_342,In_378);
and U2348 (N_2348,In_563,In_1347);
or U2349 (N_2349,In_877,In_713);
nor U2350 (N_2350,In_71,In_383);
nor U2351 (N_2351,In_80,In_1384);
or U2352 (N_2352,In_1308,In_640);
or U2353 (N_2353,In_280,In_883);
or U2354 (N_2354,In_1323,In_1093);
nand U2355 (N_2355,In_1234,In_1378);
or U2356 (N_2356,In_628,In_1499);
nand U2357 (N_2357,In_90,In_1131);
and U2358 (N_2358,In_871,In_385);
nor U2359 (N_2359,In_1171,In_584);
and U2360 (N_2360,In_1248,In_1107);
nor U2361 (N_2361,In_328,In_238);
nor U2362 (N_2362,In_1047,In_251);
and U2363 (N_2363,In_1261,In_1179);
or U2364 (N_2364,In_342,In_134);
nand U2365 (N_2365,In_88,In_203);
nand U2366 (N_2366,In_464,In_914);
and U2367 (N_2367,In_563,In_74);
and U2368 (N_2368,In_1395,In_315);
or U2369 (N_2369,In_430,In_93);
or U2370 (N_2370,In_1418,In_459);
nand U2371 (N_2371,In_187,In_1420);
or U2372 (N_2372,In_873,In_1432);
nand U2373 (N_2373,In_1154,In_293);
or U2374 (N_2374,In_1166,In_787);
or U2375 (N_2375,In_996,In_1445);
nand U2376 (N_2376,In_187,In_385);
nand U2377 (N_2377,In_330,In_605);
nor U2378 (N_2378,In_1201,In_1077);
nand U2379 (N_2379,In_1478,In_536);
and U2380 (N_2380,In_181,In_1392);
or U2381 (N_2381,In_620,In_525);
nor U2382 (N_2382,In_852,In_319);
or U2383 (N_2383,In_1002,In_297);
nand U2384 (N_2384,In_53,In_775);
or U2385 (N_2385,In_1082,In_5);
nor U2386 (N_2386,In_7,In_145);
nand U2387 (N_2387,In_370,In_8);
or U2388 (N_2388,In_1084,In_826);
nand U2389 (N_2389,In_529,In_250);
nand U2390 (N_2390,In_929,In_809);
xnor U2391 (N_2391,In_17,In_383);
and U2392 (N_2392,In_979,In_1113);
and U2393 (N_2393,In_384,In_599);
nor U2394 (N_2394,In_219,In_432);
or U2395 (N_2395,In_941,In_119);
xor U2396 (N_2396,In_196,In_793);
nor U2397 (N_2397,In_800,In_637);
nor U2398 (N_2398,In_527,In_1388);
nor U2399 (N_2399,In_1460,In_546);
nand U2400 (N_2400,In_22,In_388);
nor U2401 (N_2401,In_121,In_479);
or U2402 (N_2402,In_577,In_578);
or U2403 (N_2403,In_1361,In_1233);
nor U2404 (N_2404,In_954,In_448);
nor U2405 (N_2405,In_989,In_248);
nor U2406 (N_2406,In_982,In_64);
nor U2407 (N_2407,In_190,In_567);
nor U2408 (N_2408,In_427,In_308);
or U2409 (N_2409,In_168,In_1097);
nor U2410 (N_2410,In_1241,In_808);
or U2411 (N_2411,In_1320,In_391);
and U2412 (N_2412,In_1166,In_1204);
nor U2413 (N_2413,In_1053,In_689);
or U2414 (N_2414,In_758,In_468);
nor U2415 (N_2415,In_1315,In_1374);
nand U2416 (N_2416,In_465,In_521);
or U2417 (N_2417,In_767,In_832);
nand U2418 (N_2418,In_277,In_1454);
nand U2419 (N_2419,In_558,In_1315);
nor U2420 (N_2420,In_1468,In_135);
or U2421 (N_2421,In_1287,In_151);
or U2422 (N_2422,In_1150,In_773);
nand U2423 (N_2423,In_311,In_429);
or U2424 (N_2424,In_1418,In_85);
and U2425 (N_2425,In_885,In_1421);
nand U2426 (N_2426,In_1059,In_1405);
nor U2427 (N_2427,In_1413,In_660);
nor U2428 (N_2428,In_502,In_1171);
and U2429 (N_2429,In_718,In_1370);
or U2430 (N_2430,In_410,In_207);
or U2431 (N_2431,In_1193,In_1087);
nand U2432 (N_2432,In_911,In_311);
and U2433 (N_2433,In_487,In_610);
and U2434 (N_2434,In_1457,In_1136);
and U2435 (N_2435,In_1105,In_373);
nor U2436 (N_2436,In_86,In_1468);
and U2437 (N_2437,In_1470,In_4);
and U2438 (N_2438,In_921,In_1478);
nor U2439 (N_2439,In_506,In_358);
or U2440 (N_2440,In_1119,In_440);
nand U2441 (N_2441,In_1309,In_141);
nor U2442 (N_2442,In_26,In_809);
nor U2443 (N_2443,In_286,In_307);
and U2444 (N_2444,In_981,In_661);
nor U2445 (N_2445,In_1135,In_244);
nor U2446 (N_2446,In_171,In_54);
and U2447 (N_2447,In_179,In_386);
or U2448 (N_2448,In_63,In_220);
and U2449 (N_2449,In_148,In_646);
nor U2450 (N_2450,In_22,In_1000);
nor U2451 (N_2451,In_883,In_1322);
nor U2452 (N_2452,In_102,In_64);
nand U2453 (N_2453,In_139,In_36);
nand U2454 (N_2454,In_1329,In_1215);
nand U2455 (N_2455,In_1379,In_711);
nor U2456 (N_2456,In_517,In_1349);
nand U2457 (N_2457,In_507,In_1042);
nand U2458 (N_2458,In_606,In_1223);
and U2459 (N_2459,In_1365,In_1371);
nand U2460 (N_2460,In_1299,In_52);
nand U2461 (N_2461,In_1153,In_1377);
and U2462 (N_2462,In_1301,In_1366);
nor U2463 (N_2463,In_1129,In_1075);
nor U2464 (N_2464,In_1433,In_1076);
nor U2465 (N_2465,In_1221,In_1194);
and U2466 (N_2466,In_1391,In_407);
or U2467 (N_2467,In_555,In_631);
nand U2468 (N_2468,In_763,In_1072);
nor U2469 (N_2469,In_1495,In_699);
or U2470 (N_2470,In_1465,In_1383);
or U2471 (N_2471,In_1107,In_1273);
or U2472 (N_2472,In_716,In_99);
nand U2473 (N_2473,In_431,In_229);
or U2474 (N_2474,In_27,In_818);
and U2475 (N_2475,In_874,In_129);
nand U2476 (N_2476,In_788,In_1425);
or U2477 (N_2477,In_1270,In_1192);
and U2478 (N_2478,In_919,In_721);
or U2479 (N_2479,In_1168,In_1436);
and U2480 (N_2480,In_779,In_190);
nor U2481 (N_2481,In_1144,In_830);
nand U2482 (N_2482,In_102,In_1448);
or U2483 (N_2483,In_442,In_629);
nand U2484 (N_2484,In_307,In_954);
nand U2485 (N_2485,In_848,In_238);
nand U2486 (N_2486,In_502,In_267);
or U2487 (N_2487,In_477,In_705);
nor U2488 (N_2488,In_305,In_1096);
nand U2489 (N_2489,In_415,In_577);
nand U2490 (N_2490,In_1494,In_1294);
or U2491 (N_2491,In_1008,In_945);
nor U2492 (N_2492,In_663,In_154);
or U2493 (N_2493,In_399,In_838);
and U2494 (N_2494,In_732,In_591);
or U2495 (N_2495,In_435,In_1351);
nor U2496 (N_2496,In_1396,In_740);
nor U2497 (N_2497,In_911,In_271);
nor U2498 (N_2498,In_190,In_108);
or U2499 (N_2499,In_1022,In_1042);
or U2500 (N_2500,In_1082,In_679);
or U2501 (N_2501,In_773,In_952);
nor U2502 (N_2502,In_1480,In_1239);
or U2503 (N_2503,In_33,In_275);
nor U2504 (N_2504,In_1241,In_1424);
nor U2505 (N_2505,In_820,In_1225);
or U2506 (N_2506,In_1005,In_570);
or U2507 (N_2507,In_205,In_114);
and U2508 (N_2508,In_1020,In_1279);
nand U2509 (N_2509,In_145,In_684);
xor U2510 (N_2510,In_1359,In_532);
nand U2511 (N_2511,In_1393,In_781);
and U2512 (N_2512,In_382,In_835);
nor U2513 (N_2513,In_1093,In_664);
and U2514 (N_2514,In_93,In_1007);
nor U2515 (N_2515,In_757,In_753);
and U2516 (N_2516,In_895,In_453);
nand U2517 (N_2517,In_1328,In_923);
nor U2518 (N_2518,In_1020,In_150);
nand U2519 (N_2519,In_114,In_629);
and U2520 (N_2520,In_715,In_1107);
or U2521 (N_2521,In_487,In_1404);
and U2522 (N_2522,In_310,In_882);
nand U2523 (N_2523,In_551,In_1174);
nor U2524 (N_2524,In_662,In_54);
and U2525 (N_2525,In_850,In_68);
and U2526 (N_2526,In_316,In_449);
nor U2527 (N_2527,In_1227,In_768);
nor U2528 (N_2528,In_1100,In_43);
nor U2529 (N_2529,In_636,In_955);
and U2530 (N_2530,In_1250,In_77);
nand U2531 (N_2531,In_604,In_412);
and U2532 (N_2532,In_423,In_883);
or U2533 (N_2533,In_1285,In_1454);
or U2534 (N_2534,In_806,In_1175);
nand U2535 (N_2535,In_1006,In_687);
nor U2536 (N_2536,In_1112,In_387);
or U2537 (N_2537,In_664,In_645);
nor U2538 (N_2538,In_783,In_1420);
and U2539 (N_2539,In_1259,In_270);
or U2540 (N_2540,In_931,In_1405);
and U2541 (N_2541,In_764,In_1381);
nand U2542 (N_2542,In_888,In_592);
nand U2543 (N_2543,In_159,In_1333);
nand U2544 (N_2544,In_631,In_1493);
and U2545 (N_2545,In_1178,In_97);
nor U2546 (N_2546,In_1065,In_981);
nand U2547 (N_2547,In_198,In_599);
or U2548 (N_2548,In_655,In_912);
nand U2549 (N_2549,In_1323,In_1260);
nor U2550 (N_2550,In_829,In_1013);
nand U2551 (N_2551,In_1210,In_66);
nor U2552 (N_2552,In_1023,In_576);
nor U2553 (N_2553,In_1186,In_630);
or U2554 (N_2554,In_1477,In_1066);
or U2555 (N_2555,In_590,In_153);
nand U2556 (N_2556,In_507,In_714);
nor U2557 (N_2557,In_923,In_513);
or U2558 (N_2558,In_1312,In_790);
or U2559 (N_2559,In_1458,In_195);
nand U2560 (N_2560,In_1131,In_457);
nor U2561 (N_2561,In_1001,In_842);
and U2562 (N_2562,In_566,In_1113);
nor U2563 (N_2563,In_345,In_152);
or U2564 (N_2564,In_195,In_198);
nand U2565 (N_2565,In_1270,In_1017);
and U2566 (N_2566,In_1482,In_946);
and U2567 (N_2567,In_611,In_1084);
nand U2568 (N_2568,In_489,In_949);
nor U2569 (N_2569,In_534,In_228);
nand U2570 (N_2570,In_271,In_644);
and U2571 (N_2571,In_472,In_708);
or U2572 (N_2572,In_658,In_623);
or U2573 (N_2573,In_1295,In_81);
or U2574 (N_2574,In_1189,In_701);
and U2575 (N_2575,In_392,In_1421);
nand U2576 (N_2576,In_1164,In_973);
nand U2577 (N_2577,In_972,In_611);
nand U2578 (N_2578,In_431,In_1099);
nand U2579 (N_2579,In_1304,In_1395);
nand U2580 (N_2580,In_1390,In_134);
xnor U2581 (N_2581,In_600,In_907);
or U2582 (N_2582,In_545,In_945);
or U2583 (N_2583,In_556,In_362);
or U2584 (N_2584,In_372,In_510);
and U2585 (N_2585,In_911,In_122);
nor U2586 (N_2586,In_544,In_1060);
nor U2587 (N_2587,In_302,In_221);
nand U2588 (N_2588,In_980,In_965);
or U2589 (N_2589,In_1183,In_224);
nand U2590 (N_2590,In_207,In_252);
or U2591 (N_2591,In_201,In_1444);
or U2592 (N_2592,In_280,In_512);
nor U2593 (N_2593,In_46,In_1143);
or U2594 (N_2594,In_749,In_638);
nor U2595 (N_2595,In_882,In_652);
and U2596 (N_2596,In_775,In_272);
nor U2597 (N_2597,In_1297,In_303);
nor U2598 (N_2598,In_775,In_496);
nand U2599 (N_2599,In_482,In_374);
xor U2600 (N_2600,In_1373,In_1110);
nand U2601 (N_2601,In_1431,In_10);
and U2602 (N_2602,In_153,In_1469);
or U2603 (N_2603,In_586,In_104);
or U2604 (N_2604,In_580,In_1039);
and U2605 (N_2605,In_1086,In_1443);
and U2606 (N_2606,In_50,In_1238);
nor U2607 (N_2607,In_204,In_63);
and U2608 (N_2608,In_909,In_636);
and U2609 (N_2609,In_528,In_1118);
and U2610 (N_2610,In_304,In_761);
and U2611 (N_2611,In_1333,In_1222);
nand U2612 (N_2612,In_840,In_540);
nor U2613 (N_2613,In_1006,In_1410);
and U2614 (N_2614,In_1065,In_912);
and U2615 (N_2615,In_73,In_1411);
or U2616 (N_2616,In_764,In_1057);
nor U2617 (N_2617,In_682,In_1318);
nand U2618 (N_2618,In_901,In_73);
xor U2619 (N_2619,In_209,In_825);
nor U2620 (N_2620,In_436,In_932);
nand U2621 (N_2621,In_1084,In_536);
nor U2622 (N_2622,In_549,In_210);
nand U2623 (N_2623,In_341,In_519);
nand U2624 (N_2624,In_987,In_108);
or U2625 (N_2625,In_1426,In_487);
nor U2626 (N_2626,In_394,In_973);
or U2627 (N_2627,In_1405,In_1470);
nor U2628 (N_2628,In_333,In_868);
or U2629 (N_2629,In_772,In_535);
or U2630 (N_2630,In_227,In_848);
or U2631 (N_2631,In_968,In_847);
and U2632 (N_2632,In_139,In_1323);
nand U2633 (N_2633,In_644,In_1244);
or U2634 (N_2634,In_277,In_171);
nor U2635 (N_2635,In_1409,In_754);
nand U2636 (N_2636,In_1329,In_225);
nand U2637 (N_2637,In_1331,In_847);
or U2638 (N_2638,In_1163,In_198);
nor U2639 (N_2639,In_653,In_174);
and U2640 (N_2640,In_483,In_711);
nand U2641 (N_2641,In_658,In_838);
and U2642 (N_2642,In_1130,In_1035);
or U2643 (N_2643,In_1144,In_1492);
and U2644 (N_2644,In_161,In_946);
or U2645 (N_2645,In_974,In_1271);
nor U2646 (N_2646,In_1430,In_431);
or U2647 (N_2647,In_752,In_197);
and U2648 (N_2648,In_881,In_798);
nand U2649 (N_2649,In_23,In_158);
nor U2650 (N_2650,In_1010,In_279);
or U2651 (N_2651,In_885,In_1367);
nor U2652 (N_2652,In_60,In_924);
and U2653 (N_2653,In_881,In_202);
nor U2654 (N_2654,In_767,In_1269);
or U2655 (N_2655,In_1091,In_983);
nand U2656 (N_2656,In_1381,In_1001);
nand U2657 (N_2657,In_47,In_460);
nor U2658 (N_2658,In_225,In_109);
nor U2659 (N_2659,In_216,In_1168);
nor U2660 (N_2660,In_1350,In_449);
and U2661 (N_2661,In_72,In_849);
or U2662 (N_2662,In_464,In_209);
nor U2663 (N_2663,In_821,In_1122);
nand U2664 (N_2664,In_688,In_336);
and U2665 (N_2665,In_629,In_1250);
nand U2666 (N_2666,In_557,In_813);
or U2667 (N_2667,In_1086,In_674);
nor U2668 (N_2668,In_1036,In_525);
or U2669 (N_2669,In_861,In_85);
nor U2670 (N_2670,In_20,In_819);
and U2671 (N_2671,In_143,In_1051);
or U2672 (N_2672,In_1157,In_1350);
nor U2673 (N_2673,In_1304,In_1473);
nor U2674 (N_2674,In_1,In_112);
nor U2675 (N_2675,In_1097,In_816);
and U2676 (N_2676,In_225,In_14);
or U2677 (N_2677,In_295,In_18);
or U2678 (N_2678,In_1220,In_1324);
and U2679 (N_2679,In_1099,In_1290);
and U2680 (N_2680,In_899,In_1340);
and U2681 (N_2681,In_1249,In_1226);
and U2682 (N_2682,In_1449,In_1240);
nor U2683 (N_2683,In_263,In_937);
or U2684 (N_2684,In_132,In_98);
nor U2685 (N_2685,In_863,In_442);
and U2686 (N_2686,In_28,In_1057);
and U2687 (N_2687,In_4,In_956);
xnor U2688 (N_2688,In_756,In_1261);
or U2689 (N_2689,In_543,In_258);
and U2690 (N_2690,In_186,In_526);
nand U2691 (N_2691,In_148,In_1209);
and U2692 (N_2692,In_1120,In_702);
or U2693 (N_2693,In_683,In_425);
or U2694 (N_2694,In_374,In_4);
nor U2695 (N_2695,In_399,In_904);
and U2696 (N_2696,In_533,In_81);
nor U2697 (N_2697,In_109,In_293);
nand U2698 (N_2698,In_1360,In_699);
nand U2699 (N_2699,In_803,In_1403);
and U2700 (N_2700,In_719,In_1297);
and U2701 (N_2701,In_741,In_489);
nor U2702 (N_2702,In_1191,In_163);
nand U2703 (N_2703,In_295,In_610);
and U2704 (N_2704,In_186,In_532);
or U2705 (N_2705,In_967,In_793);
nor U2706 (N_2706,In_1233,In_1198);
and U2707 (N_2707,In_619,In_864);
and U2708 (N_2708,In_9,In_585);
nand U2709 (N_2709,In_295,In_341);
nor U2710 (N_2710,In_505,In_360);
and U2711 (N_2711,In_530,In_1198);
xnor U2712 (N_2712,In_164,In_1317);
nor U2713 (N_2713,In_242,In_1086);
nand U2714 (N_2714,In_254,In_542);
and U2715 (N_2715,In_57,In_204);
nand U2716 (N_2716,In_637,In_802);
nand U2717 (N_2717,In_217,In_125);
and U2718 (N_2718,In_1078,In_101);
and U2719 (N_2719,In_1482,In_306);
and U2720 (N_2720,In_767,In_1292);
nand U2721 (N_2721,In_1091,In_1263);
or U2722 (N_2722,In_215,In_439);
and U2723 (N_2723,In_433,In_27);
and U2724 (N_2724,In_343,In_691);
nand U2725 (N_2725,In_970,In_868);
and U2726 (N_2726,In_14,In_1005);
nand U2727 (N_2727,In_587,In_441);
nand U2728 (N_2728,In_156,In_739);
nor U2729 (N_2729,In_877,In_767);
or U2730 (N_2730,In_685,In_1187);
nor U2731 (N_2731,In_1295,In_946);
or U2732 (N_2732,In_39,In_1034);
nor U2733 (N_2733,In_876,In_243);
or U2734 (N_2734,In_701,In_277);
or U2735 (N_2735,In_478,In_894);
and U2736 (N_2736,In_798,In_1203);
nor U2737 (N_2737,In_1326,In_699);
nand U2738 (N_2738,In_639,In_546);
and U2739 (N_2739,In_634,In_1022);
nor U2740 (N_2740,In_559,In_431);
nand U2741 (N_2741,In_557,In_1147);
and U2742 (N_2742,In_662,In_1059);
nand U2743 (N_2743,In_696,In_521);
or U2744 (N_2744,In_752,In_700);
or U2745 (N_2745,In_1075,In_103);
nand U2746 (N_2746,In_385,In_554);
or U2747 (N_2747,In_254,In_131);
nor U2748 (N_2748,In_1448,In_1136);
and U2749 (N_2749,In_1329,In_1361);
nand U2750 (N_2750,In_1235,In_87);
nand U2751 (N_2751,In_145,In_368);
and U2752 (N_2752,In_674,In_657);
nand U2753 (N_2753,In_798,In_901);
xnor U2754 (N_2754,In_1374,In_788);
and U2755 (N_2755,In_551,In_1280);
nand U2756 (N_2756,In_962,In_945);
and U2757 (N_2757,In_1345,In_560);
nand U2758 (N_2758,In_1163,In_323);
nand U2759 (N_2759,In_450,In_513);
and U2760 (N_2760,In_1385,In_530);
nor U2761 (N_2761,In_954,In_770);
and U2762 (N_2762,In_1073,In_1484);
nor U2763 (N_2763,In_729,In_279);
nand U2764 (N_2764,In_1331,In_1142);
nand U2765 (N_2765,In_300,In_1449);
nand U2766 (N_2766,In_162,In_126);
nor U2767 (N_2767,In_194,In_981);
nand U2768 (N_2768,In_1139,In_248);
and U2769 (N_2769,In_13,In_234);
and U2770 (N_2770,In_676,In_337);
or U2771 (N_2771,In_48,In_1474);
and U2772 (N_2772,In_69,In_73);
nand U2773 (N_2773,In_899,In_745);
nor U2774 (N_2774,In_1010,In_843);
nand U2775 (N_2775,In_1075,In_1015);
and U2776 (N_2776,In_225,In_794);
nand U2777 (N_2777,In_1430,In_1026);
nor U2778 (N_2778,In_551,In_1139);
nand U2779 (N_2779,In_987,In_970);
nand U2780 (N_2780,In_325,In_1336);
or U2781 (N_2781,In_778,In_613);
and U2782 (N_2782,In_1263,In_673);
and U2783 (N_2783,In_46,In_803);
and U2784 (N_2784,In_1155,In_1166);
or U2785 (N_2785,In_513,In_1209);
nand U2786 (N_2786,In_1000,In_1200);
nor U2787 (N_2787,In_597,In_261);
and U2788 (N_2788,In_453,In_601);
and U2789 (N_2789,In_1084,In_62);
or U2790 (N_2790,In_165,In_780);
nand U2791 (N_2791,In_1175,In_877);
or U2792 (N_2792,In_1048,In_465);
and U2793 (N_2793,In_821,In_637);
or U2794 (N_2794,In_133,In_731);
or U2795 (N_2795,In_1458,In_281);
nand U2796 (N_2796,In_319,In_1184);
nor U2797 (N_2797,In_985,In_815);
nor U2798 (N_2798,In_614,In_224);
and U2799 (N_2799,In_1151,In_68);
or U2800 (N_2800,In_67,In_198);
nor U2801 (N_2801,In_140,In_1152);
and U2802 (N_2802,In_394,In_1143);
nand U2803 (N_2803,In_1432,In_616);
and U2804 (N_2804,In_971,In_1309);
and U2805 (N_2805,In_459,In_1375);
or U2806 (N_2806,In_393,In_752);
and U2807 (N_2807,In_1096,In_1433);
nand U2808 (N_2808,In_1207,In_25);
and U2809 (N_2809,In_118,In_476);
nor U2810 (N_2810,In_1374,In_243);
nor U2811 (N_2811,In_1358,In_774);
and U2812 (N_2812,In_1276,In_762);
nor U2813 (N_2813,In_1108,In_709);
nor U2814 (N_2814,In_378,In_170);
and U2815 (N_2815,In_794,In_810);
nand U2816 (N_2816,In_14,In_731);
nand U2817 (N_2817,In_779,In_1194);
nand U2818 (N_2818,In_362,In_1289);
and U2819 (N_2819,In_776,In_403);
and U2820 (N_2820,In_809,In_954);
nor U2821 (N_2821,In_416,In_1202);
nand U2822 (N_2822,In_1421,In_1297);
and U2823 (N_2823,In_277,In_510);
or U2824 (N_2824,In_193,In_637);
xor U2825 (N_2825,In_465,In_340);
or U2826 (N_2826,In_710,In_124);
or U2827 (N_2827,In_883,In_1145);
and U2828 (N_2828,In_386,In_176);
and U2829 (N_2829,In_997,In_591);
nor U2830 (N_2830,In_349,In_398);
and U2831 (N_2831,In_1303,In_1406);
nor U2832 (N_2832,In_75,In_573);
nand U2833 (N_2833,In_1014,In_699);
xnor U2834 (N_2834,In_201,In_607);
and U2835 (N_2835,In_1322,In_1416);
and U2836 (N_2836,In_516,In_307);
or U2837 (N_2837,In_1043,In_1488);
or U2838 (N_2838,In_169,In_1291);
and U2839 (N_2839,In_1175,In_463);
nor U2840 (N_2840,In_303,In_521);
xor U2841 (N_2841,In_1254,In_839);
or U2842 (N_2842,In_538,In_593);
nand U2843 (N_2843,In_1328,In_503);
nor U2844 (N_2844,In_219,In_459);
nand U2845 (N_2845,In_502,In_1254);
nor U2846 (N_2846,In_506,In_1366);
nand U2847 (N_2847,In_805,In_433);
and U2848 (N_2848,In_1140,In_1431);
or U2849 (N_2849,In_1283,In_509);
nor U2850 (N_2850,In_977,In_484);
and U2851 (N_2851,In_298,In_1394);
or U2852 (N_2852,In_1217,In_15);
or U2853 (N_2853,In_185,In_988);
or U2854 (N_2854,In_1116,In_195);
or U2855 (N_2855,In_1196,In_1053);
nor U2856 (N_2856,In_1224,In_1327);
and U2857 (N_2857,In_498,In_1007);
or U2858 (N_2858,In_971,In_640);
nand U2859 (N_2859,In_6,In_30);
nand U2860 (N_2860,In_245,In_170);
nand U2861 (N_2861,In_485,In_548);
or U2862 (N_2862,In_580,In_493);
nor U2863 (N_2863,In_1445,In_821);
nand U2864 (N_2864,In_1200,In_1453);
nand U2865 (N_2865,In_1179,In_22);
nor U2866 (N_2866,In_760,In_1077);
or U2867 (N_2867,In_54,In_427);
nand U2868 (N_2868,In_169,In_636);
nor U2869 (N_2869,In_102,In_1297);
nand U2870 (N_2870,In_932,In_103);
nand U2871 (N_2871,In_115,In_837);
nand U2872 (N_2872,In_1464,In_1053);
and U2873 (N_2873,In_1163,In_1229);
and U2874 (N_2874,In_146,In_817);
nor U2875 (N_2875,In_1498,In_1187);
and U2876 (N_2876,In_830,In_243);
nand U2877 (N_2877,In_825,In_1383);
nand U2878 (N_2878,In_335,In_370);
and U2879 (N_2879,In_391,In_970);
and U2880 (N_2880,In_1417,In_412);
or U2881 (N_2881,In_6,In_224);
nor U2882 (N_2882,In_966,In_1266);
nor U2883 (N_2883,In_400,In_834);
nand U2884 (N_2884,In_684,In_261);
and U2885 (N_2885,In_631,In_388);
xnor U2886 (N_2886,In_994,In_1109);
nor U2887 (N_2887,In_1497,In_619);
and U2888 (N_2888,In_131,In_470);
or U2889 (N_2889,In_783,In_565);
nor U2890 (N_2890,In_18,In_611);
nand U2891 (N_2891,In_216,In_109);
xnor U2892 (N_2892,In_1232,In_775);
and U2893 (N_2893,In_1077,In_1493);
nor U2894 (N_2894,In_459,In_183);
nand U2895 (N_2895,In_270,In_1189);
nand U2896 (N_2896,In_1483,In_138);
xor U2897 (N_2897,In_1254,In_1469);
or U2898 (N_2898,In_1320,In_355);
nor U2899 (N_2899,In_31,In_16);
and U2900 (N_2900,In_530,In_642);
and U2901 (N_2901,In_408,In_802);
nor U2902 (N_2902,In_549,In_919);
nand U2903 (N_2903,In_1081,In_321);
and U2904 (N_2904,In_608,In_797);
nand U2905 (N_2905,In_881,In_73);
or U2906 (N_2906,In_89,In_1467);
nor U2907 (N_2907,In_375,In_662);
nor U2908 (N_2908,In_494,In_402);
or U2909 (N_2909,In_472,In_1487);
or U2910 (N_2910,In_338,In_297);
nand U2911 (N_2911,In_1357,In_809);
and U2912 (N_2912,In_859,In_1283);
or U2913 (N_2913,In_365,In_534);
nor U2914 (N_2914,In_1368,In_732);
nor U2915 (N_2915,In_875,In_1348);
nor U2916 (N_2916,In_16,In_165);
or U2917 (N_2917,In_805,In_88);
nand U2918 (N_2918,In_803,In_585);
and U2919 (N_2919,In_669,In_1008);
or U2920 (N_2920,In_1320,In_806);
and U2921 (N_2921,In_38,In_1026);
nand U2922 (N_2922,In_1005,In_1318);
nor U2923 (N_2923,In_233,In_75);
nor U2924 (N_2924,In_1022,In_659);
and U2925 (N_2925,In_841,In_123);
and U2926 (N_2926,In_1389,In_673);
or U2927 (N_2927,In_1076,In_26);
and U2928 (N_2928,In_504,In_1312);
or U2929 (N_2929,In_272,In_1064);
xor U2930 (N_2930,In_415,In_311);
nand U2931 (N_2931,In_1256,In_640);
nor U2932 (N_2932,In_119,In_570);
nor U2933 (N_2933,In_564,In_621);
or U2934 (N_2934,In_625,In_12);
nor U2935 (N_2935,In_1013,In_1221);
nand U2936 (N_2936,In_404,In_480);
and U2937 (N_2937,In_268,In_1296);
or U2938 (N_2938,In_387,In_1069);
nand U2939 (N_2939,In_1047,In_1055);
and U2940 (N_2940,In_847,In_285);
and U2941 (N_2941,In_855,In_1078);
nor U2942 (N_2942,In_792,In_1431);
nand U2943 (N_2943,In_1438,In_1251);
nand U2944 (N_2944,In_1214,In_8);
nand U2945 (N_2945,In_1225,In_1435);
or U2946 (N_2946,In_998,In_890);
and U2947 (N_2947,In_1499,In_498);
nor U2948 (N_2948,In_1264,In_865);
nand U2949 (N_2949,In_198,In_1184);
and U2950 (N_2950,In_670,In_1211);
or U2951 (N_2951,In_1480,In_415);
and U2952 (N_2952,In_1210,In_30);
and U2953 (N_2953,In_1124,In_1165);
and U2954 (N_2954,In_787,In_697);
and U2955 (N_2955,In_465,In_864);
nor U2956 (N_2956,In_1205,In_970);
and U2957 (N_2957,In_985,In_1260);
and U2958 (N_2958,In_408,In_78);
nand U2959 (N_2959,In_1495,In_1498);
and U2960 (N_2960,In_43,In_1107);
nor U2961 (N_2961,In_1470,In_1002);
and U2962 (N_2962,In_1340,In_1073);
and U2963 (N_2963,In_724,In_1366);
or U2964 (N_2964,In_1129,In_1098);
nand U2965 (N_2965,In_1295,In_326);
nor U2966 (N_2966,In_166,In_1226);
nor U2967 (N_2967,In_1192,In_392);
nor U2968 (N_2968,In_18,In_29);
and U2969 (N_2969,In_1203,In_133);
or U2970 (N_2970,In_58,In_1314);
nand U2971 (N_2971,In_1052,In_13);
and U2972 (N_2972,In_887,In_1115);
and U2973 (N_2973,In_97,In_931);
nor U2974 (N_2974,In_667,In_1115);
nand U2975 (N_2975,In_687,In_877);
nor U2976 (N_2976,In_1457,In_760);
nor U2977 (N_2977,In_1171,In_1163);
or U2978 (N_2978,In_122,In_229);
nor U2979 (N_2979,In_862,In_480);
or U2980 (N_2980,In_1450,In_192);
or U2981 (N_2981,In_1123,In_1305);
or U2982 (N_2982,In_1090,In_1115);
or U2983 (N_2983,In_1216,In_194);
or U2984 (N_2984,In_1010,In_434);
and U2985 (N_2985,In_702,In_222);
nor U2986 (N_2986,In_703,In_375);
nand U2987 (N_2987,In_509,In_31);
and U2988 (N_2988,In_782,In_537);
or U2989 (N_2989,In_432,In_658);
nor U2990 (N_2990,In_908,In_102);
or U2991 (N_2991,In_659,In_1372);
or U2992 (N_2992,In_271,In_124);
and U2993 (N_2993,In_463,In_719);
nor U2994 (N_2994,In_1342,In_554);
and U2995 (N_2995,In_467,In_351);
and U2996 (N_2996,In_286,In_211);
nor U2997 (N_2997,In_1104,In_75);
xnor U2998 (N_2998,In_992,In_175);
and U2999 (N_2999,In_1312,In_413);
or U3000 (N_3000,In_872,In_954);
nor U3001 (N_3001,In_1169,In_471);
or U3002 (N_3002,In_1421,In_8);
nor U3003 (N_3003,In_1480,In_23);
nor U3004 (N_3004,In_786,In_223);
and U3005 (N_3005,In_883,In_756);
or U3006 (N_3006,In_135,In_505);
nand U3007 (N_3007,In_771,In_1017);
nand U3008 (N_3008,In_1182,In_887);
nor U3009 (N_3009,In_146,In_1181);
nor U3010 (N_3010,In_590,In_322);
nand U3011 (N_3011,In_936,In_1411);
and U3012 (N_3012,In_745,In_737);
and U3013 (N_3013,In_954,In_861);
nor U3014 (N_3014,In_99,In_998);
nor U3015 (N_3015,In_965,In_976);
xnor U3016 (N_3016,In_1443,In_852);
and U3017 (N_3017,In_316,In_353);
or U3018 (N_3018,In_1467,In_1468);
and U3019 (N_3019,In_423,In_821);
nor U3020 (N_3020,In_334,In_889);
nand U3021 (N_3021,In_1335,In_385);
nand U3022 (N_3022,In_576,In_1000);
or U3023 (N_3023,In_820,In_1007);
nand U3024 (N_3024,In_783,In_1460);
and U3025 (N_3025,In_1456,In_46);
and U3026 (N_3026,In_1240,In_262);
nor U3027 (N_3027,In_643,In_1115);
nand U3028 (N_3028,In_1352,In_844);
nor U3029 (N_3029,In_624,In_1035);
or U3030 (N_3030,In_1175,In_59);
or U3031 (N_3031,In_331,In_1487);
nor U3032 (N_3032,In_952,In_1090);
and U3033 (N_3033,In_390,In_97);
or U3034 (N_3034,In_617,In_742);
and U3035 (N_3035,In_764,In_612);
nor U3036 (N_3036,In_85,In_1325);
and U3037 (N_3037,In_147,In_186);
nor U3038 (N_3038,In_847,In_1372);
nand U3039 (N_3039,In_52,In_994);
and U3040 (N_3040,In_1371,In_1358);
nor U3041 (N_3041,In_606,In_217);
or U3042 (N_3042,In_1291,In_265);
and U3043 (N_3043,In_1469,In_1108);
nor U3044 (N_3044,In_1152,In_655);
nor U3045 (N_3045,In_757,In_1023);
and U3046 (N_3046,In_1290,In_716);
or U3047 (N_3047,In_341,In_466);
xnor U3048 (N_3048,In_1124,In_408);
nor U3049 (N_3049,In_1007,In_578);
nor U3050 (N_3050,In_1117,In_933);
nand U3051 (N_3051,In_1477,In_1196);
or U3052 (N_3052,In_882,In_536);
nor U3053 (N_3053,In_116,In_660);
nand U3054 (N_3054,In_1382,In_350);
nor U3055 (N_3055,In_1227,In_366);
nor U3056 (N_3056,In_463,In_881);
and U3057 (N_3057,In_543,In_1128);
or U3058 (N_3058,In_933,In_800);
or U3059 (N_3059,In_665,In_1114);
nand U3060 (N_3060,In_18,In_992);
and U3061 (N_3061,In_757,In_649);
or U3062 (N_3062,In_1384,In_713);
and U3063 (N_3063,In_1209,In_440);
or U3064 (N_3064,In_895,In_178);
and U3065 (N_3065,In_161,In_194);
nand U3066 (N_3066,In_935,In_78);
nor U3067 (N_3067,In_879,In_78);
nand U3068 (N_3068,In_366,In_556);
nor U3069 (N_3069,In_784,In_878);
or U3070 (N_3070,In_1094,In_1362);
nand U3071 (N_3071,In_679,In_1347);
nor U3072 (N_3072,In_988,In_406);
nand U3073 (N_3073,In_502,In_1125);
nand U3074 (N_3074,In_1069,In_1333);
or U3075 (N_3075,In_1277,In_817);
nand U3076 (N_3076,In_967,In_656);
nand U3077 (N_3077,In_818,In_517);
nand U3078 (N_3078,In_302,In_386);
nand U3079 (N_3079,In_647,In_980);
nor U3080 (N_3080,In_325,In_875);
and U3081 (N_3081,In_1205,In_659);
and U3082 (N_3082,In_1229,In_285);
nand U3083 (N_3083,In_1426,In_462);
and U3084 (N_3084,In_1002,In_142);
nand U3085 (N_3085,In_330,In_1165);
or U3086 (N_3086,In_1476,In_697);
nand U3087 (N_3087,In_299,In_752);
or U3088 (N_3088,In_1493,In_515);
xnor U3089 (N_3089,In_1277,In_465);
and U3090 (N_3090,In_637,In_772);
and U3091 (N_3091,In_131,In_831);
and U3092 (N_3092,In_69,In_688);
and U3093 (N_3093,In_1365,In_753);
nor U3094 (N_3094,In_1192,In_339);
nand U3095 (N_3095,In_182,In_1218);
and U3096 (N_3096,In_768,In_869);
and U3097 (N_3097,In_828,In_310);
nor U3098 (N_3098,In_1173,In_504);
nand U3099 (N_3099,In_251,In_390);
or U3100 (N_3100,In_736,In_1423);
nor U3101 (N_3101,In_891,In_1009);
and U3102 (N_3102,In_290,In_1283);
nand U3103 (N_3103,In_1283,In_575);
nor U3104 (N_3104,In_1183,In_743);
nand U3105 (N_3105,In_208,In_1491);
or U3106 (N_3106,In_1493,In_325);
nor U3107 (N_3107,In_849,In_864);
and U3108 (N_3108,In_1073,In_333);
nor U3109 (N_3109,In_193,In_492);
and U3110 (N_3110,In_1412,In_1159);
nor U3111 (N_3111,In_653,In_1491);
or U3112 (N_3112,In_1235,In_227);
and U3113 (N_3113,In_246,In_496);
nand U3114 (N_3114,In_1054,In_599);
nand U3115 (N_3115,In_1351,In_1211);
and U3116 (N_3116,In_734,In_982);
nor U3117 (N_3117,In_1241,In_1460);
nor U3118 (N_3118,In_551,In_1372);
nand U3119 (N_3119,In_44,In_1193);
nor U3120 (N_3120,In_44,In_1055);
nand U3121 (N_3121,In_428,In_603);
nor U3122 (N_3122,In_690,In_855);
nand U3123 (N_3123,In_1420,In_733);
nor U3124 (N_3124,In_500,In_867);
nand U3125 (N_3125,In_1006,In_1186);
or U3126 (N_3126,In_1286,In_652);
and U3127 (N_3127,In_1393,In_416);
or U3128 (N_3128,In_311,In_971);
or U3129 (N_3129,In_1183,In_1481);
nand U3130 (N_3130,In_182,In_1104);
nand U3131 (N_3131,In_1475,In_77);
and U3132 (N_3132,In_561,In_1228);
nor U3133 (N_3133,In_49,In_1421);
nand U3134 (N_3134,In_389,In_1361);
or U3135 (N_3135,In_82,In_1496);
nand U3136 (N_3136,In_1085,In_967);
nor U3137 (N_3137,In_362,In_1032);
nand U3138 (N_3138,In_931,In_232);
nor U3139 (N_3139,In_760,In_728);
and U3140 (N_3140,In_438,In_665);
nor U3141 (N_3141,In_1244,In_254);
nor U3142 (N_3142,In_1127,In_882);
nor U3143 (N_3143,In_772,In_1342);
or U3144 (N_3144,In_1162,In_698);
nor U3145 (N_3145,In_1015,In_421);
and U3146 (N_3146,In_405,In_296);
nand U3147 (N_3147,In_1471,In_939);
nand U3148 (N_3148,In_944,In_611);
and U3149 (N_3149,In_868,In_62);
or U3150 (N_3150,In_883,In_1125);
and U3151 (N_3151,In_1284,In_680);
nand U3152 (N_3152,In_641,In_880);
or U3153 (N_3153,In_1252,In_290);
xnor U3154 (N_3154,In_1347,In_767);
or U3155 (N_3155,In_267,In_878);
or U3156 (N_3156,In_1010,In_498);
or U3157 (N_3157,In_1285,In_1453);
nand U3158 (N_3158,In_1271,In_1188);
and U3159 (N_3159,In_551,In_604);
and U3160 (N_3160,In_1368,In_194);
nor U3161 (N_3161,In_1275,In_239);
nor U3162 (N_3162,In_106,In_979);
and U3163 (N_3163,In_680,In_578);
and U3164 (N_3164,In_1003,In_443);
and U3165 (N_3165,In_633,In_664);
and U3166 (N_3166,In_1176,In_1381);
nand U3167 (N_3167,In_262,In_1304);
and U3168 (N_3168,In_1039,In_584);
nand U3169 (N_3169,In_970,In_52);
nand U3170 (N_3170,In_1258,In_1408);
nand U3171 (N_3171,In_1256,In_512);
nand U3172 (N_3172,In_255,In_1173);
and U3173 (N_3173,In_157,In_1481);
and U3174 (N_3174,In_612,In_412);
or U3175 (N_3175,In_852,In_1203);
and U3176 (N_3176,In_429,In_569);
nor U3177 (N_3177,In_517,In_62);
nand U3178 (N_3178,In_5,In_411);
or U3179 (N_3179,In_509,In_1425);
nor U3180 (N_3180,In_806,In_366);
or U3181 (N_3181,In_1442,In_1030);
and U3182 (N_3182,In_695,In_853);
or U3183 (N_3183,In_1458,In_121);
nor U3184 (N_3184,In_344,In_515);
or U3185 (N_3185,In_591,In_715);
or U3186 (N_3186,In_85,In_1198);
and U3187 (N_3187,In_880,In_1416);
and U3188 (N_3188,In_1395,In_126);
or U3189 (N_3189,In_371,In_185);
and U3190 (N_3190,In_26,In_109);
nor U3191 (N_3191,In_596,In_1077);
or U3192 (N_3192,In_1156,In_625);
or U3193 (N_3193,In_780,In_614);
and U3194 (N_3194,In_909,In_179);
and U3195 (N_3195,In_566,In_1239);
nor U3196 (N_3196,In_1159,In_1200);
and U3197 (N_3197,In_974,In_426);
xnor U3198 (N_3198,In_258,In_675);
or U3199 (N_3199,In_1316,In_749);
and U3200 (N_3200,In_1102,In_1049);
and U3201 (N_3201,In_1405,In_620);
and U3202 (N_3202,In_379,In_1366);
nor U3203 (N_3203,In_591,In_1260);
nand U3204 (N_3204,In_455,In_710);
nor U3205 (N_3205,In_1412,In_74);
nor U3206 (N_3206,In_1459,In_759);
nand U3207 (N_3207,In_1205,In_515);
nand U3208 (N_3208,In_1377,In_139);
nor U3209 (N_3209,In_218,In_442);
or U3210 (N_3210,In_661,In_873);
and U3211 (N_3211,In_1304,In_522);
nand U3212 (N_3212,In_627,In_1300);
nor U3213 (N_3213,In_27,In_726);
or U3214 (N_3214,In_44,In_811);
and U3215 (N_3215,In_386,In_1494);
nand U3216 (N_3216,In_211,In_667);
nand U3217 (N_3217,In_540,In_1389);
or U3218 (N_3218,In_133,In_1320);
and U3219 (N_3219,In_858,In_543);
or U3220 (N_3220,In_861,In_489);
or U3221 (N_3221,In_9,In_1043);
or U3222 (N_3222,In_401,In_1219);
and U3223 (N_3223,In_201,In_325);
or U3224 (N_3224,In_1466,In_1354);
nor U3225 (N_3225,In_1237,In_102);
nor U3226 (N_3226,In_1317,In_407);
and U3227 (N_3227,In_332,In_875);
or U3228 (N_3228,In_1347,In_354);
nor U3229 (N_3229,In_1441,In_1342);
or U3230 (N_3230,In_829,In_169);
nand U3231 (N_3231,In_689,In_355);
nand U3232 (N_3232,In_695,In_413);
nor U3233 (N_3233,In_823,In_789);
nand U3234 (N_3234,In_390,In_1388);
nor U3235 (N_3235,In_177,In_264);
and U3236 (N_3236,In_796,In_343);
nor U3237 (N_3237,In_527,In_910);
or U3238 (N_3238,In_261,In_217);
xnor U3239 (N_3239,In_1437,In_86);
or U3240 (N_3240,In_1424,In_1196);
or U3241 (N_3241,In_271,In_335);
nand U3242 (N_3242,In_841,In_782);
nor U3243 (N_3243,In_985,In_1268);
and U3244 (N_3244,In_14,In_403);
nor U3245 (N_3245,In_807,In_1280);
nand U3246 (N_3246,In_524,In_467);
or U3247 (N_3247,In_295,In_697);
or U3248 (N_3248,In_831,In_705);
or U3249 (N_3249,In_431,In_244);
nand U3250 (N_3250,In_793,In_1183);
nor U3251 (N_3251,In_267,In_589);
nand U3252 (N_3252,In_824,In_788);
and U3253 (N_3253,In_1333,In_698);
and U3254 (N_3254,In_1267,In_848);
or U3255 (N_3255,In_776,In_967);
nand U3256 (N_3256,In_1274,In_244);
nor U3257 (N_3257,In_679,In_1338);
or U3258 (N_3258,In_1435,In_902);
nand U3259 (N_3259,In_1470,In_840);
or U3260 (N_3260,In_589,In_200);
and U3261 (N_3261,In_1209,In_309);
nand U3262 (N_3262,In_88,In_344);
nand U3263 (N_3263,In_625,In_888);
nor U3264 (N_3264,In_1264,In_910);
or U3265 (N_3265,In_1127,In_927);
nor U3266 (N_3266,In_1191,In_965);
nor U3267 (N_3267,In_760,In_290);
or U3268 (N_3268,In_301,In_120);
nand U3269 (N_3269,In_1383,In_576);
nor U3270 (N_3270,In_1196,In_898);
and U3271 (N_3271,In_46,In_274);
or U3272 (N_3272,In_538,In_650);
and U3273 (N_3273,In_436,In_639);
or U3274 (N_3274,In_1348,In_1225);
nand U3275 (N_3275,In_1005,In_489);
nor U3276 (N_3276,In_960,In_540);
nor U3277 (N_3277,In_1205,In_254);
and U3278 (N_3278,In_1060,In_862);
nand U3279 (N_3279,In_1424,In_1359);
nand U3280 (N_3280,In_217,In_1151);
nand U3281 (N_3281,In_317,In_319);
and U3282 (N_3282,In_303,In_158);
and U3283 (N_3283,In_1428,In_201);
or U3284 (N_3284,In_447,In_644);
and U3285 (N_3285,In_456,In_768);
nand U3286 (N_3286,In_285,In_718);
or U3287 (N_3287,In_235,In_805);
nand U3288 (N_3288,In_1442,In_715);
nor U3289 (N_3289,In_1395,In_1433);
nor U3290 (N_3290,In_779,In_55);
nor U3291 (N_3291,In_1125,In_811);
nor U3292 (N_3292,In_478,In_701);
nor U3293 (N_3293,In_1261,In_1056);
nand U3294 (N_3294,In_401,In_865);
nor U3295 (N_3295,In_594,In_202);
and U3296 (N_3296,In_823,In_691);
or U3297 (N_3297,In_423,In_1270);
nand U3298 (N_3298,In_59,In_93);
nand U3299 (N_3299,In_1488,In_478);
and U3300 (N_3300,In_1061,In_1236);
nor U3301 (N_3301,In_1435,In_667);
nor U3302 (N_3302,In_1334,In_1478);
nor U3303 (N_3303,In_479,In_1095);
nor U3304 (N_3304,In_645,In_926);
nand U3305 (N_3305,In_890,In_1155);
or U3306 (N_3306,In_1176,In_904);
nand U3307 (N_3307,In_277,In_425);
nand U3308 (N_3308,In_775,In_800);
or U3309 (N_3309,In_1268,In_73);
nor U3310 (N_3310,In_29,In_124);
nor U3311 (N_3311,In_1007,In_573);
and U3312 (N_3312,In_352,In_156);
and U3313 (N_3313,In_1357,In_1221);
nor U3314 (N_3314,In_515,In_590);
nor U3315 (N_3315,In_130,In_354);
or U3316 (N_3316,In_159,In_1196);
nor U3317 (N_3317,In_1026,In_275);
or U3318 (N_3318,In_1398,In_819);
or U3319 (N_3319,In_1332,In_567);
and U3320 (N_3320,In_734,In_1033);
nor U3321 (N_3321,In_1194,In_705);
and U3322 (N_3322,In_144,In_529);
or U3323 (N_3323,In_1455,In_382);
or U3324 (N_3324,In_160,In_881);
or U3325 (N_3325,In_741,In_537);
and U3326 (N_3326,In_1041,In_62);
and U3327 (N_3327,In_782,In_1044);
and U3328 (N_3328,In_916,In_482);
nand U3329 (N_3329,In_1248,In_52);
and U3330 (N_3330,In_945,In_1471);
nor U3331 (N_3331,In_794,In_995);
and U3332 (N_3332,In_982,In_1160);
and U3333 (N_3333,In_1403,In_417);
nand U3334 (N_3334,In_1404,In_574);
or U3335 (N_3335,In_1309,In_1055);
nand U3336 (N_3336,In_1162,In_1184);
nand U3337 (N_3337,In_874,In_16);
and U3338 (N_3338,In_90,In_175);
nor U3339 (N_3339,In_1048,In_1097);
or U3340 (N_3340,In_134,In_1428);
nand U3341 (N_3341,In_447,In_699);
or U3342 (N_3342,In_598,In_1370);
nor U3343 (N_3343,In_274,In_909);
nor U3344 (N_3344,In_253,In_152);
and U3345 (N_3345,In_895,In_1070);
nand U3346 (N_3346,In_1032,In_694);
nor U3347 (N_3347,In_1197,In_156);
nor U3348 (N_3348,In_1214,In_1373);
nand U3349 (N_3349,In_482,In_1302);
or U3350 (N_3350,In_1340,In_643);
or U3351 (N_3351,In_1471,In_1474);
and U3352 (N_3352,In_1221,In_710);
and U3353 (N_3353,In_1178,In_1225);
nor U3354 (N_3354,In_708,In_1099);
nand U3355 (N_3355,In_1100,In_687);
and U3356 (N_3356,In_75,In_213);
or U3357 (N_3357,In_558,In_94);
and U3358 (N_3358,In_259,In_904);
or U3359 (N_3359,In_468,In_966);
and U3360 (N_3360,In_496,In_84);
or U3361 (N_3361,In_1307,In_570);
nand U3362 (N_3362,In_1195,In_400);
nand U3363 (N_3363,In_627,In_425);
or U3364 (N_3364,In_1065,In_993);
or U3365 (N_3365,In_49,In_364);
nor U3366 (N_3366,In_1363,In_417);
nand U3367 (N_3367,In_265,In_1090);
nor U3368 (N_3368,In_1175,In_300);
nand U3369 (N_3369,In_555,In_578);
or U3370 (N_3370,In_805,In_526);
and U3371 (N_3371,In_584,In_730);
or U3372 (N_3372,In_379,In_975);
and U3373 (N_3373,In_1484,In_1148);
nor U3374 (N_3374,In_519,In_189);
nor U3375 (N_3375,In_264,In_1376);
or U3376 (N_3376,In_68,In_947);
and U3377 (N_3377,In_1408,In_630);
or U3378 (N_3378,In_48,In_980);
nor U3379 (N_3379,In_1376,In_235);
or U3380 (N_3380,In_321,In_1052);
and U3381 (N_3381,In_427,In_459);
nand U3382 (N_3382,In_426,In_362);
or U3383 (N_3383,In_63,In_1328);
or U3384 (N_3384,In_517,In_637);
or U3385 (N_3385,In_661,In_1100);
nand U3386 (N_3386,In_429,In_136);
or U3387 (N_3387,In_809,In_982);
or U3388 (N_3388,In_1372,In_736);
or U3389 (N_3389,In_1316,In_702);
or U3390 (N_3390,In_953,In_747);
or U3391 (N_3391,In_447,In_81);
or U3392 (N_3392,In_1310,In_754);
nand U3393 (N_3393,In_207,In_1192);
or U3394 (N_3394,In_272,In_1108);
nor U3395 (N_3395,In_1278,In_417);
nand U3396 (N_3396,In_534,In_411);
nor U3397 (N_3397,In_411,In_604);
nor U3398 (N_3398,In_680,In_230);
nor U3399 (N_3399,In_296,In_1032);
and U3400 (N_3400,In_689,In_250);
or U3401 (N_3401,In_151,In_584);
or U3402 (N_3402,In_792,In_1416);
or U3403 (N_3403,In_778,In_372);
nor U3404 (N_3404,In_886,In_27);
or U3405 (N_3405,In_1093,In_100);
nor U3406 (N_3406,In_99,In_473);
and U3407 (N_3407,In_367,In_31);
or U3408 (N_3408,In_47,In_1075);
nand U3409 (N_3409,In_665,In_445);
nand U3410 (N_3410,In_58,In_437);
and U3411 (N_3411,In_193,In_802);
and U3412 (N_3412,In_646,In_1350);
or U3413 (N_3413,In_906,In_998);
or U3414 (N_3414,In_247,In_1231);
nor U3415 (N_3415,In_1293,In_1412);
or U3416 (N_3416,In_1334,In_832);
xor U3417 (N_3417,In_334,In_188);
nand U3418 (N_3418,In_95,In_6);
nand U3419 (N_3419,In_1019,In_1328);
nand U3420 (N_3420,In_856,In_420);
nand U3421 (N_3421,In_731,In_74);
nand U3422 (N_3422,In_1043,In_1321);
and U3423 (N_3423,In_972,In_837);
and U3424 (N_3424,In_1176,In_990);
nand U3425 (N_3425,In_932,In_1241);
nor U3426 (N_3426,In_983,In_1178);
nand U3427 (N_3427,In_515,In_303);
or U3428 (N_3428,In_1012,In_195);
or U3429 (N_3429,In_131,In_799);
nand U3430 (N_3430,In_1302,In_1310);
and U3431 (N_3431,In_979,In_1448);
nor U3432 (N_3432,In_621,In_504);
nor U3433 (N_3433,In_405,In_468);
or U3434 (N_3434,In_465,In_567);
and U3435 (N_3435,In_1160,In_560);
and U3436 (N_3436,In_41,In_147);
nor U3437 (N_3437,In_894,In_347);
nand U3438 (N_3438,In_827,In_257);
and U3439 (N_3439,In_136,In_438);
nand U3440 (N_3440,In_558,In_110);
and U3441 (N_3441,In_339,In_385);
nor U3442 (N_3442,In_712,In_1307);
nand U3443 (N_3443,In_1228,In_91);
or U3444 (N_3444,In_854,In_853);
and U3445 (N_3445,In_839,In_1335);
and U3446 (N_3446,In_719,In_716);
or U3447 (N_3447,In_747,In_1108);
nand U3448 (N_3448,In_384,In_841);
or U3449 (N_3449,In_909,In_1278);
nand U3450 (N_3450,In_808,In_189);
or U3451 (N_3451,In_686,In_1349);
or U3452 (N_3452,In_780,In_1382);
or U3453 (N_3453,In_354,In_1286);
and U3454 (N_3454,In_37,In_678);
nand U3455 (N_3455,In_1363,In_1141);
and U3456 (N_3456,In_957,In_405);
nand U3457 (N_3457,In_756,In_765);
or U3458 (N_3458,In_394,In_1319);
and U3459 (N_3459,In_790,In_60);
and U3460 (N_3460,In_903,In_1094);
or U3461 (N_3461,In_856,In_754);
and U3462 (N_3462,In_178,In_941);
or U3463 (N_3463,In_1419,In_93);
nand U3464 (N_3464,In_385,In_1405);
and U3465 (N_3465,In_12,In_800);
nand U3466 (N_3466,In_590,In_1355);
and U3467 (N_3467,In_998,In_275);
nand U3468 (N_3468,In_911,In_293);
and U3469 (N_3469,In_808,In_942);
and U3470 (N_3470,In_1479,In_658);
and U3471 (N_3471,In_747,In_256);
nor U3472 (N_3472,In_581,In_1112);
and U3473 (N_3473,In_1059,In_1198);
nand U3474 (N_3474,In_464,In_1440);
nand U3475 (N_3475,In_386,In_477);
nand U3476 (N_3476,In_77,In_931);
or U3477 (N_3477,In_848,In_199);
or U3478 (N_3478,In_864,In_461);
and U3479 (N_3479,In_1165,In_870);
nand U3480 (N_3480,In_187,In_506);
nor U3481 (N_3481,In_177,In_1269);
nand U3482 (N_3482,In_143,In_1091);
nand U3483 (N_3483,In_1440,In_88);
nor U3484 (N_3484,In_1098,In_1255);
nand U3485 (N_3485,In_1291,In_438);
nor U3486 (N_3486,In_1074,In_180);
nand U3487 (N_3487,In_1200,In_130);
and U3488 (N_3488,In_518,In_636);
nor U3489 (N_3489,In_74,In_1154);
nand U3490 (N_3490,In_102,In_1077);
or U3491 (N_3491,In_761,In_1296);
and U3492 (N_3492,In_75,In_1381);
nand U3493 (N_3493,In_888,In_1375);
and U3494 (N_3494,In_269,In_682);
nor U3495 (N_3495,In_845,In_886);
or U3496 (N_3496,In_1498,In_766);
nor U3497 (N_3497,In_832,In_684);
nand U3498 (N_3498,In_830,In_702);
nand U3499 (N_3499,In_643,In_429);
nor U3500 (N_3500,In_64,In_467);
and U3501 (N_3501,In_409,In_157);
and U3502 (N_3502,In_648,In_252);
nand U3503 (N_3503,In_556,In_1467);
nand U3504 (N_3504,In_740,In_1399);
nor U3505 (N_3505,In_617,In_1225);
nand U3506 (N_3506,In_675,In_834);
and U3507 (N_3507,In_140,In_1068);
and U3508 (N_3508,In_1133,In_1437);
and U3509 (N_3509,In_933,In_952);
nand U3510 (N_3510,In_691,In_75);
nand U3511 (N_3511,In_461,In_230);
nand U3512 (N_3512,In_463,In_1426);
or U3513 (N_3513,In_874,In_1352);
nor U3514 (N_3514,In_1175,In_186);
or U3515 (N_3515,In_1372,In_278);
nand U3516 (N_3516,In_280,In_1097);
or U3517 (N_3517,In_754,In_1249);
and U3518 (N_3518,In_1079,In_7);
and U3519 (N_3519,In_892,In_1380);
nand U3520 (N_3520,In_150,In_783);
or U3521 (N_3521,In_1364,In_1399);
nand U3522 (N_3522,In_386,In_1440);
nand U3523 (N_3523,In_1209,In_380);
nand U3524 (N_3524,In_1119,In_1330);
or U3525 (N_3525,In_753,In_549);
or U3526 (N_3526,In_1150,In_1275);
and U3527 (N_3527,In_618,In_172);
or U3528 (N_3528,In_629,In_87);
and U3529 (N_3529,In_111,In_660);
and U3530 (N_3530,In_845,In_570);
nand U3531 (N_3531,In_617,In_545);
nor U3532 (N_3532,In_793,In_1262);
or U3533 (N_3533,In_1362,In_1370);
or U3534 (N_3534,In_1461,In_807);
nand U3535 (N_3535,In_1123,In_188);
nand U3536 (N_3536,In_1155,In_202);
or U3537 (N_3537,In_538,In_558);
and U3538 (N_3538,In_358,In_999);
nand U3539 (N_3539,In_47,In_308);
nor U3540 (N_3540,In_144,In_588);
or U3541 (N_3541,In_1306,In_842);
nand U3542 (N_3542,In_934,In_279);
or U3543 (N_3543,In_265,In_231);
or U3544 (N_3544,In_413,In_354);
and U3545 (N_3545,In_1099,In_321);
nand U3546 (N_3546,In_527,In_878);
nor U3547 (N_3547,In_56,In_1458);
nor U3548 (N_3548,In_577,In_1470);
nand U3549 (N_3549,In_447,In_709);
nor U3550 (N_3550,In_584,In_1155);
or U3551 (N_3551,In_1469,In_140);
and U3552 (N_3552,In_117,In_1327);
or U3553 (N_3553,In_1291,In_984);
or U3554 (N_3554,In_430,In_1354);
or U3555 (N_3555,In_156,In_512);
nor U3556 (N_3556,In_1124,In_1495);
or U3557 (N_3557,In_1426,In_958);
or U3558 (N_3558,In_1479,In_261);
nand U3559 (N_3559,In_835,In_654);
nor U3560 (N_3560,In_956,In_469);
nand U3561 (N_3561,In_216,In_785);
nor U3562 (N_3562,In_121,In_1203);
nand U3563 (N_3563,In_1199,In_1157);
nand U3564 (N_3564,In_960,In_789);
nand U3565 (N_3565,In_434,In_554);
and U3566 (N_3566,In_1377,In_913);
nor U3567 (N_3567,In_737,In_730);
or U3568 (N_3568,In_782,In_36);
nand U3569 (N_3569,In_620,In_234);
and U3570 (N_3570,In_297,In_1332);
nand U3571 (N_3571,In_860,In_1107);
nor U3572 (N_3572,In_625,In_1083);
nor U3573 (N_3573,In_1094,In_739);
or U3574 (N_3574,In_1325,In_1159);
or U3575 (N_3575,In_970,In_16);
nand U3576 (N_3576,In_1267,In_264);
nand U3577 (N_3577,In_1466,In_372);
nand U3578 (N_3578,In_673,In_704);
nand U3579 (N_3579,In_1296,In_1024);
or U3580 (N_3580,In_262,In_83);
and U3581 (N_3581,In_1432,In_1356);
nand U3582 (N_3582,In_1436,In_634);
nor U3583 (N_3583,In_861,In_1310);
nor U3584 (N_3584,In_577,In_644);
nand U3585 (N_3585,In_976,In_271);
nor U3586 (N_3586,In_96,In_947);
or U3587 (N_3587,In_1077,In_59);
and U3588 (N_3588,In_1381,In_335);
and U3589 (N_3589,In_1046,In_853);
and U3590 (N_3590,In_1074,In_413);
and U3591 (N_3591,In_866,In_906);
nand U3592 (N_3592,In_66,In_1129);
and U3593 (N_3593,In_554,In_355);
or U3594 (N_3594,In_894,In_260);
nand U3595 (N_3595,In_365,In_1279);
or U3596 (N_3596,In_747,In_912);
nand U3597 (N_3597,In_992,In_1122);
or U3598 (N_3598,In_1165,In_957);
and U3599 (N_3599,In_364,In_1382);
nand U3600 (N_3600,In_1238,In_282);
nor U3601 (N_3601,In_113,In_1377);
and U3602 (N_3602,In_574,In_212);
xor U3603 (N_3603,In_1018,In_687);
nor U3604 (N_3604,In_1183,In_723);
nand U3605 (N_3605,In_1359,In_1030);
or U3606 (N_3606,In_744,In_1366);
or U3607 (N_3607,In_83,In_349);
nor U3608 (N_3608,In_60,In_51);
nand U3609 (N_3609,In_256,In_846);
and U3610 (N_3610,In_633,In_1081);
or U3611 (N_3611,In_551,In_336);
nand U3612 (N_3612,In_843,In_1391);
or U3613 (N_3613,In_17,In_1474);
or U3614 (N_3614,In_920,In_1011);
nand U3615 (N_3615,In_1064,In_1393);
and U3616 (N_3616,In_391,In_1410);
nand U3617 (N_3617,In_682,In_1130);
and U3618 (N_3618,In_1286,In_326);
nor U3619 (N_3619,In_129,In_753);
or U3620 (N_3620,In_1277,In_1259);
or U3621 (N_3621,In_1432,In_25);
nand U3622 (N_3622,In_470,In_4);
nor U3623 (N_3623,In_432,In_977);
nor U3624 (N_3624,In_555,In_515);
or U3625 (N_3625,In_1283,In_1420);
or U3626 (N_3626,In_382,In_525);
or U3627 (N_3627,In_1054,In_258);
nor U3628 (N_3628,In_570,In_591);
nand U3629 (N_3629,In_144,In_1046);
or U3630 (N_3630,In_950,In_891);
or U3631 (N_3631,In_445,In_1270);
nor U3632 (N_3632,In_714,In_1162);
and U3633 (N_3633,In_772,In_956);
and U3634 (N_3634,In_519,In_417);
nor U3635 (N_3635,In_1200,In_573);
nand U3636 (N_3636,In_18,In_1200);
nor U3637 (N_3637,In_30,In_604);
and U3638 (N_3638,In_107,In_583);
and U3639 (N_3639,In_472,In_836);
nand U3640 (N_3640,In_605,In_1179);
nor U3641 (N_3641,In_710,In_745);
or U3642 (N_3642,In_924,In_900);
nor U3643 (N_3643,In_1441,In_1404);
and U3644 (N_3644,In_449,In_438);
nand U3645 (N_3645,In_109,In_355);
or U3646 (N_3646,In_550,In_865);
or U3647 (N_3647,In_1152,In_670);
and U3648 (N_3648,In_1408,In_1078);
nor U3649 (N_3649,In_1180,In_719);
and U3650 (N_3650,In_1270,In_914);
or U3651 (N_3651,In_1084,In_768);
and U3652 (N_3652,In_1170,In_727);
nor U3653 (N_3653,In_994,In_18);
and U3654 (N_3654,In_848,In_1123);
and U3655 (N_3655,In_354,In_1313);
nor U3656 (N_3656,In_1172,In_1412);
and U3657 (N_3657,In_1023,In_935);
nor U3658 (N_3658,In_118,In_846);
nor U3659 (N_3659,In_212,In_706);
nor U3660 (N_3660,In_757,In_161);
nand U3661 (N_3661,In_782,In_154);
nor U3662 (N_3662,In_250,In_1428);
or U3663 (N_3663,In_1229,In_252);
nand U3664 (N_3664,In_460,In_747);
and U3665 (N_3665,In_1288,In_1192);
nor U3666 (N_3666,In_242,In_1297);
xnor U3667 (N_3667,In_156,In_1258);
nand U3668 (N_3668,In_1449,In_989);
and U3669 (N_3669,In_1128,In_728);
and U3670 (N_3670,In_1415,In_1053);
nand U3671 (N_3671,In_975,In_511);
nand U3672 (N_3672,In_1139,In_143);
nor U3673 (N_3673,In_17,In_1485);
or U3674 (N_3674,In_1291,In_937);
nand U3675 (N_3675,In_305,In_653);
nor U3676 (N_3676,In_687,In_1173);
or U3677 (N_3677,In_94,In_568);
nor U3678 (N_3678,In_29,In_1301);
and U3679 (N_3679,In_743,In_1398);
xnor U3680 (N_3680,In_1184,In_1211);
or U3681 (N_3681,In_55,In_1384);
xnor U3682 (N_3682,In_164,In_1190);
or U3683 (N_3683,In_491,In_402);
and U3684 (N_3684,In_1055,In_176);
nor U3685 (N_3685,In_827,In_1281);
or U3686 (N_3686,In_565,In_38);
or U3687 (N_3687,In_1219,In_191);
nand U3688 (N_3688,In_1005,In_238);
and U3689 (N_3689,In_1195,In_523);
or U3690 (N_3690,In_1285,In_822);
nor U3691 (N_3691,In_247,In_1470);
nand U3692 (N_3692,In_39,In_312);
or U3693 (N_3693,In_1337,In_68);
or U3694 (N_3694,In_110,In_921);
and U3695 (N_3695,In_685,In_379);
and U3696 (N_3696,In_1073,In_788);
nor U3697 (N_3697,In_970,In_899);
nor U3698 (N_3698,In_33,In_613);
or U3699 (N_3699,In_1183,In_473);
or U3700 (N_3700,In_564,In_1430);
or U3701 (N_3701,In_972,In_1452);
nor U3702 (N_3702,In_927,In_1384);
or U3703 (N_3703,In_1403,In_717);
nor U3704 (N_3704,In_229,In_809);
or U3705 (N_3705,In_912,In_1443);
nand U3706 (N_3706,In_503,In_526);
and U3707 (N_3707,In_387,In_744);
nand U3708 (N_3708,In_1446,In_1210);
nand U3709 (N_3709,In_200,In_187);
and U3710 (N_3710,In_113,In_232);
nand U3711 (N_3711,In_354,In_498);
nor U3712 (N_3712,In_1386,In_764);
nor U3713 (N_3713,In_786,In_511);
nand U3714 (N_3714,In_467,In_1142);
or U3715 (N_3715,In_1047,In_808);
nand U3716 (N_3716,In_185,In_209);
nand U3717 (N_3717,In_648,In_643);
nand U3718 (N_3718,In_1444,In_273);
nor U3719 (N_3719,In_754,In_168);
and U3720 (N_3720,In_1452,In_41);
and U3721 (N_3721,In_1131,In_669);
nand U3722 (N_3722,In_62,In_628);
nor U3723 (N_3723,In_327,In_229);
or U3724 (N_3724,In_659,In_78);
or U3725 (N_3725,In_110,In_314);
and U3726 (N_3726,In_11,In_1038);
and U3727 (N_3727,In_1392,In_1422);
or U3728 (N_3728,In_488,In_494);
nor U3729 (N_3729,In_1197,In_237);
or U3730 (N_3730,In_294,In_754);
nor U3731 (N_3731,In_776,In_73);
and U3732 (N_3732,In_1144,In_1062);
and U3733 (N_3733,In_124,In_1228);
and U3734 (N_3734,In_47,In_95);
nand U3735 (N_3735,In_1388,In_211);
nand U3736 (N_3736,In_95,In_1020);
or U3737 (N_3737,In_536,In_684);
nand U3738 (N_3738,In_213,In_1317);
nor U3739 (N_3739,In_694,In_1444);
nor U3740 (N_3740,In_351,In_827);
and U3741 (N_3741,In_1228,In_400);
nor U3742 (N_3742,In_909,In_580);
and U3743 (N_3743,In_582,In_1266);
and U3744 (N_3744,In_479,In_513);
nor U3745 (N_3745,In_615,In_1279);
and U3746 (N_3746,In_1347,In_753);
or U3747 (N_3747,In_458,In_1103);
or U3748 (N_3748,In_1124,In_1199);
nor U3749 (N_3749,In_1025,In_767);
and U3750 (N_3750,In_150,In_351);
and U3751 (N_3751,In_99,In_122);
or U3752 (N_3752,In_1373,In_732);
nor U3753 (N_3753,In_990,In_661);
nand U3754 (N_3754,In_123,In_226);
nor U3755 (N_3755,In_184,In_653);
and U3756 (N_3756,In_713,In_643);
or U3757 (N_3757,In_832,In_842);
nor U3758 (N_3758,In_239,In_1431);
nand U3759 (N_3759,In_1233,In_278);
nand U3760 (N_3760,In_1027,In_833);
or U3761 (N_3761,In_831,In_753);
or U3762 (N_3762,In_1364,In_739);
and U3763 (N_3763,In_1127,In_785);
or U3764 (N_3764,In_471,In_534);
and U3765 (N_3765,In_1037,In_81);
nand U3766 (N_3766,In_7,In_1472);
or U3767 (N_3767,In_1401,In_456);
nand U3768 (N_3768,In_1357,In_1071);
nor U3769 (N_3769,In_1363,In_1390);
or U3770 (N_3770,In_1010,In_1077);
and U3771 (N_3771,In_726,In_1315);
nor U3772 (N_3772,In_1199,In_1446);
nor U3773 (N_3773,In_429,In_1383);
and U3774 (N_3774,In_1269,In_679);
nor U3775 (N_3775,In_587,In_873);
nor U3776 (N_3776,In_1053,In_254);
or U3777 (N_3777,In_1085,In_336);
nor U3778 (N_3778,In_1035,In_759);
and U3779 (N_3779,In_855,In_555);
nand U3780 (N_3780,In_1266,In_887);
and U3781 (N_3781,In_1353,In_213);
or U3782 (N_3782,In_818,In_1281);
nand U3783 (N_3783,In_1426,In_262);
nor U3784 (N_3784,In_54,In_1417);
nand U3785 (N_3785,In_483,In_389);
nor U3786 (N_3786,In_1029,In_414);
or U3787 (N_3787,In_537,In_740);
nand U3788 (N_3788,In_1150,In_205);
nand U3789 (N_3789,In_811,In_270);
nand U3790 (N_3790,In_537,In_320);
or U3791 (N_3791,In_1490,In_482);
and U3792 (N_3792,In_1312,In_139);
or U3793 (N_3793,In_1221,In_578);
and U3794 (N_3794,In_34,In_299);
or U3795 (N_3795,In_1149,In_639);
nand U3796 (N_3796,In_1136,In_353);
or U3797 (N_3797,In_572,In_1498);
nand U3798 (N_3798,In_318,In_566);
xor U3799 (N_3799,In_1493,In_897);
nand U3800 (N_3800,In_883,In_727);
nand U3801 (N_3801,In_1006,In_944);
or U3802 (N_3802,In_499,In_982);
nor U3803 (N_3803,In_723,In_278);
xor U3804 (N_3804,In_1057,In_203);
and U3805 (N_3805,In_173,In_537);
nor U3806 (N_3806,In_1272,In_448);
nor U3807 (N_3807,In_665,In_1253);
and U3808 (N_3808,In_651,In_26);
and U3809 (N_3809,In_108,In_1332);
nand U3810 (N_3810,In_459,In_51);
nor U3811 (N_3811,In_273,In_1122);
nor U3812 (N_3812,In_1453,In_1316);
and U3813 (N_3813,In_247,In_1183);
and U3814 (N_3814,In_311,In_989);
nand U3815 (N_3815,In_1327,In_702);
or U3816 (N_3816,In_895,In_366);
nand U3817 (N_3817,In_185,In_1097);
nor U3818 (N_3818,In_511,In_576);
nand U3819 (N_3819,In_1067,In_840);
or U3820 (N_3820,In_181,In_511);
nand U3821 (N_3821,In_798,In_481);
nand U3822 (N_3822,In_254,In_1291);
or U3823 (N_3823,In_475,In_128);
and U3824 (N_3824,In_1383,In_148);
xnor U3825 (N_3825,In_847,In_749);
or U3826 (N_3826,In_427,In_699);
or U3827 (N_3827,In_1263,In_1264);
nor U3828 (N_3828,In_1075,In_838);
and U3829 (N_3829,In_553,In_324);
nand U3830 (N_3830,In_824,In_981);
nand U3831 (N_3831,In_935,In_159);
nand U3832 (N_3832,In_1303,In_1342);
nand U3833 (N_3833,In_1309,In_950);
nor U3834 (N_3834,In_186,In_906);
nand U3835 (N_3835,In_591,In_974);
nor U3836 (N_3836,In_635,In_712);
or U3837 (N_3837,In_901,In_592);
nand U3838 (N_3838,In_770,In_400);
or U3839 (N_3839,In_806,In_757);
nand U3840 (N_3840,In_512,In_1372);
nor U3841 (N_3841,In_934,In_1302);
nand U3842 (N_3842,In_1030,In_1423);
or U3843 (N_3843,In_460,In_66);
or U3844 (N_3844,In_82,In_961);
or U3845 (N_3845,In_1119,In_1052);
and U3846 (N_3846,In_544,In_635);
nand U3847 (N_3847,In_560,In_968);
or U3848 (N_3848,In_451,In_297);
nor U3849 (N_3849,In_177,In_842);
or U3850 (N_3850,In_1239,In_1395);
nand U3851 (N_3851,In_840,In_1101);
or U3852 (N_3852,In_1004,In_1059);
or U3853 (N_3853,In_1333,In_270);
or U3854 (N_3854,In_56,In_763);
nand U3855 (N_3855,In_757,In_656);
or U3856 (N_3856,In_109,In_776);
and U3857 (N_3857,In_951,In_1228);
nor U3858 (N_3858,In_1483,In_88);
nand U3859 (N_3859,In_581,In_786);
nor U3860 (N_3860,In_1418,In_1191);
nand U3861 (N_3861,In_11,In_1022);
or U3862 (N_3862,In_199,In_902);
or U3863 (N_3863,In_1283,In_1125);
nor U3864 (N_3864,In_1213,In_42);
and U3865 (N_3865,In_867,In_803);
xor U3866 (N_3866,In_871,In_1314);
nor U3867 (N_3867,In_489,In_1451);
and U3868 (N_3868,In_1142,In_1411);
and U3869 (N_3869,In_1002,In_1137);
nand U3870 (N_3870,In_1448,In_1226);
xnor U3871 (N_3871,In_1047,In_37);
nor U3872 (N_3872,In_1461,In_1393);
and U3873 (N_3873,In_120,In_272);
nand U3874 (N_3874,In_1368,In_252);
and U3875 (N_3875,In_670,In_1383);
nor U3876 (N_3876,In_656,In_915);
or U3877 (N_3877,In_268,In_1085);
nand U3878 (N_3878,In_620,In_625);
nand U3879 (N_3879,In_1478,In_411);
nand U3880 (N_3880,In_448,In_117);
nor U3881 (N_3881,In_309,In_865);
and U3882 (N_3882,In_1089,In_1487);
nand U3883 (N_3883,In_1136,In_929);
and U3884 (N_3884,In_509,In_1432);
or U3885 (N_3885,In_1299,In_371);
nand U3886 (N_3886,In_152,In_1475);
or U3887 (N_3887,In_1342,In_1324);
and U3888 (N_3888,In_1484,In_24);
nand U3889 (N_3889,In_1089,In_1274);
and U3890 (N_3890,In_202,In_572);
and U3891 (N_3891,In_599,In_787);
and U3892 (N_3892,In_888,In_1307);
and U3893 (N_3893,In_1468,In_463);
and U3894 (N_3894,In_51,In_89);
or U3895 (N_3895,In_1129,In_1123);
and U3896 (N_3896,In_806,In_443);
nor U3897 (N_3897,In_1103,In_608);
or U3898 (N_3898,In_1473,In_1468);
nor U3899 (N_3899,In_32,In_976);
and U3900 (N_3900,In_203,In_395);
nor U3901 (N_3901,In_552,In_1358);
nor U3902 (N_3902,In_708,In_665);
and U3903 (N_3903,In_1055,In_1329);
nor U3904 (N_3904,In_853,In_322);
and U3905 (N_3905,In_1433,In_295);
nor U3906 (N_3906,In_1490,In_1001);
nor U3907 (N_3907,In_871,In_1027);
nor U3908 (N_3908,In_802,In_56);
nor U3909 (N_3909,In_789,In_897);
or U3910 (N_3910,In_1394,In_20);
or U3911 (N_3911,In_1076,In_507);
nor U3912 (N_3912,In_1158,In_895);
nand U3913 (N_3913,In_1234,In_509);
and U3914 (N_3914,In_1206,In_437);
or U3915 (N_3915,In_1343,In_182);
and U3916 (N_3916,In_992,In_1433);
and U3917 (N_3917,In_551,In_749);
and U3918 (N_3918,In_1418,In_116);
and U3919 (N_3919,In_1170,In_1299);
and U3920 (N_3920,In_823,In_625);
xnor U3921 (N_3921,In_1012,In_756);
nor U3922 (N_3922,In_1263,In_1149);
or U3923 (N_3923,In_70,In_1212);
or U3924 (N_3924,In_94,In_131);
or U3925 (N_3925,In_1063,In_794);
nand U3926 (N_3926,In_1407,In_342);
nand U3927 (N_3927,In_551,In_1286);
nand U3928 (N_3928,In_1034,In_328);
nand U3929 (N_3929,In_1159,In_576);
nand U3930 (N_3930,In_700,In_1017);
and U3931 (N_3931,In_966,In_1186);
and U3932 (N_3932,In_252,In_278);
nor U3933 (N_3933,In_582,In_1175);
nand U3934 (N_3934,In_841,In_773);
or U3935 (N_3935,In_870,In_1029);
or U3936 (N_3936,In_248,In_1099);
or U3937 (N_3937,In_1229,In_1395);
nor U3938 (N_3938,In_977,In_559);
nor U3939 (N_3939,In_1229,In_714);
or U3940 (N_3940,In_1459,In_868);
or U3941 (N_3941,In_1363,In_1154);
nor U3942 (N_3942,In_294,In_689);
and U3943 (N_3943,In_479,In_304);
nand U3944 (N_3944,In_344,In_1345);
or U3945 (N_3945,In_949,In_958);
nand U3946 (N_3946,In_1494,In_1106);
nand U3947 (N_3947,In_1380,In_939);
or U3948 (N_3948,In_810,In_1272);
nor U3949 (N_3949,In_1309,In_1030);
nor U3950 (N_3950,In_203,In_82);
nor U3951 (N_3951,In_879,In_561);
or U3952 (N_3952,In_1426,In_211);
and U3953 (N_3953,In_822,In_103);
and U3954 (N_3954,In_129,In_632);
nand U3955 (N_3955,In_723,In_189);
and U3956 (N_3956,In_869,In_1190);
and U3957 (N_3957,In_825,In_148);
nand U3958 (N_3958,In_1009,In_179);
nand U3959 (N_3959,In_687,In_1065);
nand U3960 (N_3960,In_1323,In_1265);
or U3961 (N_3961,In_510,In_869);
or U3962 (N_3962,In_1001,In_890);
and U3963 (N_3963,In_1237,In_46);
and U3964 (N_3964,In_998,In_1467);
nor U3965 (N_3965,In_806,In_404);
and U3966 (N_3966,In_832,In_662);
or U3967 (N_3967,In_938,In_31);
and U3968 (N_3968,In_1189,In_1077);
nor U3969 (N_3969,In_1271,In_265);
and U3970 (N_3970,In_1179,In_598);
nand U3971 (N_3971,In_542,In_1411);
or U3972 (N_3972,In_1443,In_368);
or U3973 (N_3973,In_416,In_1473);
nand U3974 (N_3974,In_54,In_211);
and U3975 (N_3975,In_556,In_962);
or U3976 (N_3976,In_1409,In_414);
nand U3977 (N_3977,In_338,In_179);
nand U3978 (N_3978,In_951,In_1312);
xnor U3979 (N_3979,In_302,In_1213);
and U3980 (N_3980,In_148,In_1334);
and U3981 (N_3981,In_116,In_247);
nor U3982 (N_3982,In_0,In_430);
or U3983 (N_3983,In_138,In_845);
or U3984 (N_3984,In_1053,In_354);
or U3985 (N_3985,In_309,In_721);
xnor U3986 (N_3986,In_1363,In_1432);
and U3987 (N_3987,In_1321,In_746);
and U3988 (N_3988,In_230,In_153);
or U3989 (N_3989,In_934,In_183);
nand U3990 (N_3990,In_1242,In_1042);
nor U3991 (N_3991,In_1070,In_1301);
nor U3992 (N_3992,In_209,In_250);
and U3993 (N_3993,In_1083,In_34);
and U3994 (N_3994,In_635,In_947);
nand U3995 (N_3995,In_789,In_1229);
and U3996 (N_3996,In_797,In_29);
xnor U3997 (N_3997,In_915,In_55);
or U3998 (N_3998,In_521,In_1087);
or U3999 (N_3999,In_500,In_1101);
and U4000 (N_4000,In_799,In_891);
nand U4001 (N_4001,In_1006,In_878);
nand U4002 (N_4002,In_1303,In_677);
or U4003 (N_4003,In_764,In_1490);
nand U4004 (N_4004,In_13,In_1302);
nor U4005 (N_4005,In_479,In_1303);
xor U4006 (N_4006,In_1456,In_1257);
and U4007 (N_4007,In_83,In_270);
nand U4008 (N_4008,In_163,In_170);
and U4009 (N_4009,In_185,In_1359);
or U4010 (N_4010,In_918,In_65);
and U4011 (N_4011,In_1232,In_915);
and U4012 (N_4012,In_1451,In_550);
and U4013 (N_4013,In_492,In_671);
nand U4014 (N_4014,In_1499,In_145);
nor U4015 (N_4015,In_193,In_251);
or U4016 (N_4016,In_996,In_1072);
nand U4017 (N_4017,In_226,In_1037);
nor U4018 (N_4018,In_706,In_1319);
nor U4019 (N_4019,In_371,In_1391);
nand U4020 (N_4020,In_691,In_667);
nand U4021 (N_4021,In_67,In_1359);
nor U4022 (N_4022,In_1047,In_71);
nor U4023 (N_4023,In_648,In_304);
and U4024 (N_4024,In_967,In_481);
nor U4025 (N_4025,In_69,In_1219);
and U4026 (N_4026,In_313,In_615);
nor U4027 (N_4027,In_820,In_637);
nand U4028 (N_4028,In_188,In_519);
and U4029 (N_4029,In_651,In_828);
nor U4030 (N_4030,In_888,In_119);
and U4031 (N_4031,In_819,In_92);
or U4032 (N_4032,In_1146,In_1061);
and U4033 (N_4033,In_685,In_546);
nand U4034 (N_4034,In_904,In_1067);
or U4035 (N_4035,In_1484,In_1390);
or U4036 (N_4036,In_1474,In_102);
nand U4037 (N_4037,In_200,In_971);
or U4038 (N_4038,In_1221,In_29);
nor U4039 (N_4039,In_427,In_1193);
nand U4040 (N_4040,In_362,In_363);
nor U4041 (N_4041,In_1174,In_299);
nor U4042 (N_4042,In_933,In_661);
or U4043 (N_4043,In_1021,In_1169);
xor U4044 (N_4044,In_1317,In_1413);
nand U4045 (N_4045,In_211,In_1076);
and U4046 (N_4046,In_1096,In_629);
and U4047 (N_4047,In_245,In_1467);
and U4048 (N_4048,In_895,In_731);
nand U4049 (N_4049,In_330,In_1104);
nor U4050 (N_4050,In_228,In_1180);
nand U4051 (N_4051,In_608,In_988);
and U4052 (N_4052,In_30,In_174);
nor U4053 (N_4053,In_226,In_674);
nor U4054 (N_4054,In_877,In_383);
and U4055 (N_4055,In_1422,In_756);
or U4056 (N_4056,In_864,In_672);
and U4057 (N_4057,In_451,In_1467);
and U4058 (N_4058,In_247,In_663);
xor U4059 (N_4059,In_819,In_221);
nand U4060 (N_4060,In_391,In_343);
and U4061 (N_4061,In_170,In_1350);
nor U4062 (N_4062,In_1472,In_1159);
nand U4063 (N_4063,In_1397,In_837);
nor U4064 (N_4064,In_185,In_1327);
or U4065 (N_4065,In_650,In_748);
and U4066 (N_4066,In_1332,In_1154);
and U4067 (N_4067,In_630,In_68);
nand U4068 (N_4068,In_1413,In_1436);
nand U4069 (N_4069,In_705,In_756);
nor U4070 (N_4070,In_1161,In_461);
nor U4071 (N_4071,In_871,In_518);
nand U4072 (N_4072,In_1320,In_860);
or U4073 (N_4073,In_887,In_1494);
and U4074 (N_4074,In_1340,In_1438);
and U4075 (N_4075,In_769,In_246);
and U4076 (N_4076,In_205,In_73);
nor U4077 (N_4077,In_655,In_1361);
and U4078 (N_4078,In_252,In_1058);
and U4079 (N_4079,In_704,In_11);
or U4080 (N_4080,In_87,In_593);
nand U4081 (N_4081,In_1172,In_931);
nand U4082 (N_4082,In_1172,In_564);
and U4083 (N_4083,In_1356,In_307);
nand U4084 (N_4084,In_1000,In_316);
and U4085 (N_4085,In_274,In_357);
and U4086 (N_4086,In_449,In_149);
nand U4087 (N_4087,In_19,In_617);
nor U4088 (N_4088,In_881,In_1222);
nand U4089 (N_4089,In_1082,In_491);
and U4090 (N_4090,In_114,In_1094);
and U4091 (N_4091,In_175,In_1078);
nand U4092 (N_4092,In_885,In_1282);
nor U4093 (N_4093,In_1328,In_574);
nor U4094 (N_4094,In_1090,In_120);
nor U4095 (N_4095,In_706,In_1101);
and U4096 (N_4096,In_228,In_237);
nor U4097 (N_4097,In_1328,In_535);
or U4098 (N_4098,In_1357,In_31);
and U4099 (N_4099,In_475,In_1148);
and U4100 (N_4100,In_855,In_231);
nor U4101 (N_4101,In_0,In_220);
or U4102 (N_4102,In_1169,In_378);
or U4103 (N_4103,In_1420,In_597);
or U4104 (N_4104,In_1208,In_36);
xnor U4105 (N_4105,In_1231,In_1003);
nand U4106 (N_4106,In_1162,In_1334);
nand U4107 (N_4107,In_270,In_588);
and U4108 (N_4108,In_1201,In_68);
or U4109 (N_4109,In_355,In_1363);
or U4110 (N_4110,In_73,In_701);
nand U4111 (N_4111,In_442,In_876);
nand U4112 (N_4112,In_1099,In_622);
nand U4113 (N_4113,In_970,In_500);
and U4114 (N_4114,In_404,In_392);
nor U4115 (N_4115,In_882,In_337);
or U4116 (N_4116,In_34,In_11);
nor U4117 (N_4117,In_88,In_82);
or U4118 (N_4118,In_960,In_114);
nor U4119 (N_4119,In_940,In_808);
or U4120 (N_4120,In_1206,In_631);
nand U4121 (N_4121,In_357,In_1189);
nor U4122 (N_4122,In_394,In_1479);
or U4123 (N_4123,In_988,In_722);
or U4124 (N_4124,In_35,In_291);
xor U4125 (N_4125,In_374,In_1255);
nor U4126 (N_4126,In_229,In_803);
nand U4127 (N_4127,In_390,In_1306);
and U4128 (N_4128,In_146,In_440);
and U4129 (N_4129,In_97,In_916);
nor U4130 (N_4130,In_1234,In_629);
nor U4131 (N_4131,In_476,In_1116);
or U4132 (N_4132,In_691,In_1032);
and U4133 (N_4133,In_347,In_179);
nor U4134 (N_4134,In_1255,In_1329);
or U4135 (N_4135,In_52,In_947);
or U4136 (N_4136,In_273,In_733);
xor U4137 (N_4137,In_103,In_1254);
or U4138 (N_4138,In_209,In_141);
or U4139 (N_4139,In_1385,In_964);
nor U4140 (N_4140,In_1084,In_1404);
and U4141 (N_4141,In_702,In_629);
and U4142 (N_4142,In_635,In_905);
nand U4143 (N_4143,In_1394,In_746);
or U4144 (N_4144,In_439,In_8);
nor U4145 (N_4145,In_47,In_998);
or U4146 (N_4146,In_1490,In_969);
and U4147 (N_4147,In_4,In_42);
or U4148 (N_4148,In_1239,In_933);
nand U4149 (N_4149,In_769,In_956);
or U4150 (N_4150,In_444,In_24);
or U4151 (N_4151,In_1368,In_753);
nor U4152 (N_4152,In_1445,In_654);
nand U4153 (N_4153,In_1447,In_1448);
and U4154 (N_4154,In_1014,In_810);
nand U4155 (N_4155,In_195,In_770);
or U4156 (N_4156,In_257,In_951);
or U4157 (N_4157,In_137,In_589);
nand U4158 (N_4158,In_425,In_604);
or U4159 (N_4159,In_827,In_455);
nand U4160 (N_4160,In_1150,In_616);
and U4161 (N_4161,In_953,In_1493);
nor U4162 (N_4162,In_430,In_1467);
nor U4163 (N_4163,In_734,In_86);
nor U4164 (N_4164,In_1037,In_230);
nor U4165 (N_4165,In_1159,In_50);
nor U4166 (N_4166,In_1243,In_645);
or U4167 (N_4167,In_918,In_1399);
and U4168 (N_4168,In_942,In_532);
or U4169 (N_4169,In_120,In_81);
xor U4170 (N_4170,In_1021,In_1337);
nand U4171 (N_4171,In_91,In_328);
or U4172 (N_4172,In_418,In_1433);
nand U4173 (N_4173,In_1324,In_493);
nor U4174 (N_4174,In_1047,In_1313);
nor U4175 (N_4175,In_1483,In_929);
or U4176 (N_4176,In_1437,In_662);
nand U4177 (N_4177,In_401,In_1313);
and U4178 (N_4178,In_386,In_702);
or U4179 (N_4179,In_377,In_424);
nor U4180 (N_4180,In_1009,In_335);
nand U4181 (N_4181,In_855,In_1189);
or U4182 (N_4182,In_195,In_76);
or U4183 (N_4183,In_495,In_357);
or U4184 (N_4184,In_772,In_357);
nor U4185 (N_4185,In_1138,In_1283);
or U4186 (N_4186,In_888,In_1396);
and U4187 (N_4187,In_860,In_1328);
nor U4188 (N_4188,In_315,In_460);
nand U4189 (N_4189,In_1169,In_1436);
nor U4190 (N_4190,In_769,In_1132);
nand U4191 (N_4191,In_244,In_509);
or U4192 (N_4192,In_780,In_158);
nand U4193 (N_4193,In_1414,In_766);
and U4194 (N_4194,In_1211,In_791);
and U4195 (N_4195,In_1498,In_1006);
and U4196 (N_4196,In_30,In_1311);
nor U4197 (N_4197,In_924,In_478);
nand U4198 (N_4198,In_813,In_846);
nand U4199 (N_4199,In_1428,In_888);
nand U4200 (N_4200,In_21,In_1141);
and U4201 (N_4201,In_1295,In_1167);
or U4202 (N_4202,In_1237,In_273);
nand U4203 (N_4203,In_445,In_1221);
nand U4204 (N_4204,In_1196,In_535);
nor U4205 (N_4205,In_157,In_373);
nand U4206 (N_4206,In_1087,In_995);
or U4207 (N_4207,In_1381,In_1223);
or U4208 (N_4208,In_825,In_1132);
or U4209 (N_4209,In_360,In_614);
and U4210 (N_4210,In_667,In_1326);
nand U4211 (N_4211,In_1458,In_164);
nand U4212 (N_4212,In_562,In_1355);
nand U4213 (N_4213,In_25,In_727);
nand U4214 (N_4214,In_1371,In_226);
nor U4215 (N_4215,In_406,In_289);
nor U4216 (N_4216,In_470,In_1331);
nor U4217 (N_4217,In_555,In_876);
nand U4218 (N_4218,In_64,In_1216);
or U4219 (N_4219,In_1270,In_218);
or U4220 (N_4220,In_781,In_876);
and U4221 (N_4221,In_436,In_453);
or U4222 (N_4222,In_58,In_842);
or U4223 (N_4223,In_25,In_470);
nand U4224 (N_4224,In_1455,In_578);
nor U4225 (N_4225,In_1424,In_57);
or U4226 (N_4226,In_1054,In_1344);
nor U4227 (N_4227,In_1448,In_722);
nor U4228 (N_4228,In_517,In_274);
and U4229 (N_4229,In_1120,In_1253);
and U4230 (N_4230,In_242,In_248);
nand U4231 (N_4231,In_112,In_659);
or U4232 (N_4232,In_438,In_72);
nand U4233 (N_4233,In_573,In_1194);
nand U4234 (N_4234,In_457,In_66);
and U4235 (N_4235,In_838,In_968);
or U4236 (N_4236,In_1274,In_897);
nor U4237 (N_4237,In_643,In_1367);
nor U4238 (N_4238,In_1001,In_1327);
nand U4239 (N_4239,In_487,In_277);
nor U4240 (N_4240,In_944,In_1103);
nor U4241 (N_4241,In_326,In_965);
nor U4242 (N_4242,In_915,In_156);
or U4243 (N_4243,In_508,In_1149);
nor U4244 (N_4244,In_481,In_726);
nor U4245 (N_4245,In_719,In_1450);
and U4246 (N_4246,In_140,In_1321);
and U4247 (N_4247,In_927,In_1188);
nand U4248 (N_4248,In_611,In_653);
nand U4249 (N_4249,In_1284,In_1061);
or U4250 (N_4250,In_249,In_466);
nand U4251 (N_4251,In_106,In_898);
xor U4252 (N_4252,In_241,In_1165);
or U4253 (N_4253,In_1498,In_755);
and U4254 (N_4254,In_890,In_633);
or U4255 (N_4255,In_1443,In_396);
nor U4256 (N_4256,In_1434,In_595);
nand U4257 (N_4257,In_566,In_287);
nand U4258 (N_4258,In_1258,In_1396);
nand U4259 (N_4259,In_1238,In_1190);
nor U4260 (N_4260,In_783,In_619);
nor U4261 (N_4261,In_472,In_608);
nor U4262 (N_4262,In_1049,In_202);
and U4263 (N_4263,In_693,In_435);
nor U4264 (N_4264,In_96,In_1479);
or U4265 (N_4265,In_1273,In_21);
or U4266 (N_4266,In_78,In_586);
or U4267 (N_4267,In_1216,In_1150);
nand U4268 (N_4268,In_1128,In_1102);
nand U4269 (N_4269,In_1469,In_429);
or U4270 (N_4270,In_937,In_312);
or U4271 (N_4271,In_550,In_1212);
nor U4272 (N_4272,In_1347,In_413);
nor U4273 (N_4273,In_1289,In_210);
nand U4274 (N_4274,In_286,In_523);
or U4275 (N_4275,In_1077,In_835);
or U4276 (N_4276,In_367,In_1459);
and U4277 (N_4277,In_1491,In_977);
nor U4278 (N_4278,In_882,In_8);
nand U4279 (N_4279,In_1268,In_348);
nor U4280 (N_4280,In_760,In_631);
nand U4281 (N_4281,In_919,In_136);
or U4282 (N_4282,In_354,In_1397);
nand U4283 (N_4283,In_1194,In_332);
nor U4284 (N_4284,In_867,In_83);
nor U4285 (N_4285,In_6,In_0);
xor U4286 (N_4286,In_1151,In_958);
or U4287 (N_4287,In_1146,In_747);
nor U4288 (N_4288,In_427,In_214);
and U4289 (N_4289,In_310,In_437);
xnor U4290 (N_4290,In_1385,In_969);
and U4291 (N_4291,In_1119,In_944);
or U4292 (N_4292,In_677,In_905);
nor U4293 (N_4293,In_70,In_909);
and U4294 (N_4294,In_1344,In_507);
nor U4295 (N_4295,In_900,In_57);
and U4296 (N_4296,In_32,In_344);
nor U4297 (N_4297,In_491,In_1379);
nor U4298 (N_4298,In_1125,In_494);
nand U4299 (N_4299,In_519,In_1353);
and U4300 (N_4300,In_1499,In_322);
nand U4301 (N_4301,In_672,In_1411);
and U4302 (N_4302,In_1425,In_794);
or U4303 (N_4303,In_1264,In_41);
nand U4304 (N_4304,In_276,In_193);
nand U4305 (N_4305,In_776,In_1039);
nor U4306 (N_4306,In_348,In_842);
nand U4307 (N_4307,In_857,In_1385);
or U4308 (N_4308,In_1351,In_987);
nand U4309 (N_4309,In_1307,In_1215);
nand U4310 (N_4310,In_993,In_1075);
or U4311 (N_4311,In_1262,In_1014);
nor U4312 (N_4312,In_92,In_449);
or U4313 (N_4313,In_293,In_412);
and U4314 (N_4314,In_903,In_1108);
and U4315 (N_4315,In_1133,In_545);
or U4316 (N_4316,In_348,In_1227);
nand U4317 (N_4317,In_1439,In_237);
or U4318 (N_4318,In_236,In_723);
nor U4319 (N_4319,In_159,In_985);
nor U4320 (N_4320,In_829,In_1033);
xnor U4321 (N_4321,In_938,In_802);
nand U4322 (N_4322,In_511,In_388);
and U4323 (N_4323,In_1250,In_1194);
nand U4324 (N_4324,In_579,In_95);
nand U4325 (N_4325,In_814,In_600);
and U4326 (N_4326,In_739,In_994);
and U4327 (N_4327,In_401,In_209);
nor U4328 (N_4328,In_1395,In_388);
nor U4329 (N_4329,In_408,In_1041);
or U4330 (N_4330,In_49,In_376);
nand U4331 (N_4331,In_934,In_1054);
or U4332 (N_4332,In_375,In_1270);
nor U4333 (N_4333,In_235,In_52);
and U4334 (N_4334,In_1468,In_1459);
and U4335 (N_4335,In_977,In_592);
or U4336 (N_4336,In_155,In_993);
nor U4337 (N_4337,In_1243,In_120);
and U4338 (N_4338,In_605,In_1234);
nand U4339 (N_4339,In_1209,In_304);
nand U4340 (N_4340,In_932,In_792);
nor U4341 (N_4341,In_1214,In_832);
or U4342 (N_4342,In_273,In_1214);
nand U4343 (N_4343,In_945,In_384);
or U4344 (N_4344,In_499,In_1451);
nand U4345 (N_4345,In_1171,In_1181);
nor U4346 (N_4346,In_51,In_1240);
nor U4347 (N_4347,In_241,In_785);
nor U4348 (N_4348,In_507,In_770);
nand U4349 (N_4349,In_748,In_319);
nand U4350 (N_4350,In_905,In_957);
or U4351 (N_4351,In_282,In_1169);
nand U4352 (N_4352,In_975,In_1230);
or U4353 (N_4353,In_582,In_396);
or U4354 (N_4354,In_389,In_471);
and U4355 (N_4355,In_6,In_469);
or U4356 (N_4356,In_1040,In_863);
nand U4357 (N_4357,In_203,In_1405);
or U4358 (N_4358,In_307,In_1250);
nor U4359 (N_4359,In_1419,In_304);
nor U4360 (N_4360,In_851,In_1144);
nand U4361 (N_4361,In_1448,In_1430);
and U4362 (N_4362,In_47,In_94);
nor U4363 (N_4363,In_208,In_799);
and U4364 (N_4364,In_475,In_712);
nor U4365 (N_4365,In_1468,In_168);
or U4366 (N_4366,In_1238,In_937);
or U4367 (N_4367,In_1319,In_218);
nor U4368 (N_4368,In_90,In_760);
and U4369 (N_4369,In_1019,In_1498);
and U4370 (N_4370,In_775,In_883);
nand U4371 (N_4371,In_93,In_53);
and U4372 (N_4372,In_1098,In_4);
and U4373 (N_4373,In_838,In_1063);
nand U4374 (N_4374,In_1270,In_1337);
nand U4375 (N_4375,In_737,In_555);
and U4376 (N_4376,In_1114,In_599);
nor U4377 (N_4377,In_578,In_57);
and U4378 (N_4378,In_964,In_1188);
nand U4379 (N_4379,In_272,In_267);
nand U4380 (N_4380,In_1261,In_18);
nor U4381 (N_4381,In_517,In_398);
and U4382 (N_4382,In_306,In_183);
nor U4383 (N_4383,In_885,In_1428);
nor U4384 (N_4384,In_1384,In_626);
xor U4385 (N_4385,In_985,In_974);
and U4386 (N_4386,In_1214,In_568);
nand U4387 (N_4387,In_1050,In_937);
or U4388 (N_4388,In_1425,In_1399);
or U4389 (N_4389,In_366,In_1234);
nor U4390 (N_4390,In_1070,In_1351);
and U4391 (N_4391,In_1070,In_929);
nor U4392 (N_4392,In_141,In_423);
and U4393 (N_4393,In_1013,In_622);
nand U4394 (N_4394,In_531,In_1178);
and U4395 (N_4395,In_217,In_973);
or U4396 (N_4396,In_627,In_41);
nand U4397 (N_4397,In_1471,In_405);
nand U4398 (N_4398,In_681,In_755);
and U4399 (N_4399,In_292,In_1354);
or U4400 (N_4400,In_417,In_103);
and U4401 (N_4401,In_1274,In_1140);
or U4402 (N_4402,In_1046,In_1059);
and U4403 (N_4403,In_1396,In_904);
and U4404 (N_4404,In_472,In_1071);
or U4405 (N_4405,In_1460,In_445);
or U4406 (N_4406,In_903,In_749);
and U4407 (N_4407,In_439,In_290);
and U4408 (N_4408,In_857,In_912);
nor U4409 (N_4409,In_939,In_278);
or U4410 (N_4410,In_1346,In_1171);
nor U4411 (N_4411,In_736,In_98);
nand U4412 (N_4412,In_1385,In_57);
and U4413 (N_4413,In_990,In_378);
and U4414 (N_4414,In_1221,In_1285);
and U4415 (N_4415,In_1079,In_795);
nor U4416 (N_4416,In_1477,In_211);
or U4417 (N_4417,In_170,In_506);
nor U4418 (N_4418,In_1446,In_1075);
nor U4419 (N_4419,In_309,In_1088);
and U4420 (N_4420,In_101,In_1109);
or U4421 (N_4421,In_218,In_650);
nand U4422 (N_4422,In_1173,In_1110);
or U4423 (N_4423,In_380,In_1152);
xnor U4424 (N_4424,In_1165,In_1029);
nor U4425 (N_4425,In_668,In_329);
and U4426 (N_4426,In_1074,In_321);
nand U4427 (N_4427,In_1163,In_954);
nor U4428 (N_4428,In_537,In_1274);
nand U4429 (N_4429,In_30,In_830);
nand U4430 (N_4430,In_1115,In_923);
nor U4431 (N_4431,In_143,In_404);
and U4432 (N_4432,In_516,In_937);
nor U4433 (N_4433,In_26,In_1426);
nand U4434 (N_4434,In_411,In_454);
nand U4435 (N_4435,In_1421,In_641);
nor U4436 (N_4436,In_482,In_488);
and U4437 (N_4437,In_1450,In_1323);
nor U4438 (N_4438,In_266,In_824);
and U4439 (N_4439,In_1078,In_1496);
or U4440 (N_4440,In_47,In_948);
nand U4441 (N_4441,In_21,In_122);
nor U4442 (N_4442,In_382,In_1440);
nand U4443 (N_4443,In_288,In_1067);
or U4444 (N_4444,In_1167,In_197);
and U4445 (N_4445,In_941,In_1281);
nor U4446 (N_4446,In_1375,In_284);
or U4447 (N_4447,In_5,In_1247);
nand U4448 (N_4448,In_1306,In_467);
nor U4449 (N_4449,In_486,In_259);
or U4450 (N_4450,In_466,In_110);
and U4451 (N_4451,In_440,In_49);
and U4452 (N_4452,In_969,In_1249);
or U4453 (N_4453,In_32,In_740);
nor U4454 (N_4454,In_558,In_1440);
nand U4455 (N_4455,In_1045,In_557);
or U4456 (N_4456,In_548,In_1114);
and U4457 (N_4457,In_62,In_308);
nand U4458 (N_4458,In_306,In_534);
and U4459 (N_4459,In_1041,In_222);
and U4460 (N_4460,In_113,In_821);
nor U4461 (N_4461,In_976,In_1185);
nand U4462 (N_4462,In_615,In_64);
or U4463 (N_4463,In_951,In_1447);
and U4464 (N_4464,In_298,In_646);
or U4465 (N_4465,In_625,In_1221);
or U4466 (N_4466,In_761,In_369);
nor U4467 (N_4467,In_571,In_910);
and U4468 (N_4468,In_973,In_388);
and U4469 (N_4469,In_58,In_281);
nor U4470 (N_4470,In_359,In_1128);
or U4471 (N_4471,In_49,In_1078);
nor U4472 (N_4472,In_238,In_943);
nand U4473 (N_4473,In_524,In_274);
or U4474 (N_4474,In_853,In_1186);
and U4475 (N_4475,In_1025,In_1335);
or U4476 (N_4476,In_616,In_202);
and U4477 (N_4477,In_254,In_944);
or U4478 (N_4478,In_668,In_1236);
nand U4479 (N_4479,In_1376,In_822);
and U4480 (N_4480,In_1085,In_113);
and U4481 (N_4481,In_8,In_38);
nor U4482 (N_4482,In_1433,In_1069);
nand U4483 (N_4483,In_200,In_920);
nor U4484 (N_4484,In_904,In_198);
or U4485 (N_4485,In_866,In_508);
nor U4486 (N_4486,In_441,In_1051);
and U4487 (N_4487,In_672,In_515);
nand U4488 (N_4488,In_196,In_24);
or U4489 (N_4489,In_413,In_1373);
and U4490 (N_4490,In_1165,In_637);
nor U4491 (N_4491,In_1448,In_696);
nand U4492 (N_4492,In_1381,In_768);
nor U4493 (N_4493,In_302,In_61);
nor U4494 (N_4494,In_895,In_164);
nor U4495 (N_4495,In_1488,In_1372);
and U4496 (N_4496,In_1251,In_289);
or U4497 (N_4497,In_165,In_923);
nor U4498 (N_4498,In_909,In_296);
nor U4499 (N_4499,In_77,In_728);
and U4500 (N_4500,In_336,In_1095);
and U4501 (N_4501,In_261,In_1414);
or U4502 (N_4502,In_456,In_867);
nor U4503 (N_4503,In_1355,In_937);
nand U4504 (N_4504,In_1214,In_599);
or U4505 (N_4505,In_1040,In_372);
and U4506 (N_4506,In_1361,In_1411);
nand U4507 (N_4507,In_283,In_610);
and U4508 (N_4508,In_1333,In_454);
or U4509 (N_4509,In_1055,In_1419);
or U4510 (N_4510,In_19,In_456);
nand U4511 (N_4511,In_790,In_414);
and U4512 (N_4512,In_1483,In_853);
nand U4513 (N_4513,In_557,In_1014);
nand U4514 (N_4514,In_1246,In_637);
and U4515 (N_4515,In_1447,In_1340);
and U4516 (N_4516,In_226,In_1222);
nor U4517 (N_4517,In_600,In_672);
and U4518 (N_4518,In_574,In_831);
and U4519 (N_4519,In_537,In_1442);
or U4520 (N_4520,In_998,In_1249);
or U4521 (N_4521,In_72,In_723);
nand U4522 (N_4522,In_1323,In_991);
nand U4523 (N_4523,In_435,In_1014);
and U4524 (N_4524,In_1458,In_1288);
nor U4525 (N_4525,In_764,In_210);
nor U4526 (N_4526,In_142,In_494);
or U4527 (N_4527,In_964,In_712);
nand U4528 (N_4528,In_1448,In_1446);
nand U4529 (N_4529,In_807,In_1125);
and U4530 (N_4530,In_85,In_94);
nor U4531 (N_4531,In_668,In_642);
nand U4532 (N_4532,In_182,In_1155);
nor U4533 (N_4533,In_1122,In_729);
nor U4534 (N_4534,In_853,In_685);
and U4535 (N_4535,In_1005,In_804);
or U4536 (N_4536,In_633,In_621);
nand U4537 (N_4537,In_679,In_238);
nor U4538 (N_4538,In_274,In_507);
and U4539 (N_4539,In_99,In_743);
and U4540 (N_4540,In_846,In_1001);
or U4541 (N_4541,In_1021,In_1361);
or U4542 (N_4542,In_848,In_1396);
nand U4543 (N_4543,In_744,In_1037);
nand U4544 (N_4544,In_1044,In_115);
or U4545 (N_4545,In_1037,In_315);
or U4546 (N_4546,In_1050,In_243);
or U4547 (N_4547,In_220,In_831);
xnor U4548 (N_4548,In_177,In_573);
nand U4549 (N_4549,In_403,In_677);
and U4550 (N_4550,In_1310,In_1298);
nand U4551 (N_4551,In_1182,In_1072);
and U4552 (N_4552,In_972,In_314);
nor U4553 (N_4553,In_1200,In_1013);
and U4554 (N_4554,In_736,In_1364);
or U4555 (N_4555,In_1473,In_610);
and U4556 (N_4556,In_864,In_77);
and U4557 (N_4557,In_919,In_958);
and U4558 (N_4558,In_488,In_1405);
nand U4559 (N_4559,In_1487,In_792);
or U4560 (N_4560,In_45,In_1146);
nor U4561 (N_4561,In_264,In_480);
nor U4562 (N_4562,In_583,In_676);
and U4563 (N_4563,In_880,In_339);
nand U4564 (N_4564,In_1131,In_1317);
nand U4565 (N_4565,In_1175,In_288);
and U4566 (N_4566,In_193,In_283);
or U4567 (N_4567,In_1112,In_110);
nor U4568 (N_4568,In_661,In_921);
or U4569 (N_4569,In_475,In_314);
nand U4570 (N_4570,In_561,In_699);
xor U4571 (N_4571,In_1113,In_1112);
nand U4572 (N_4572,In_1030,In_748);
xnor U4573 (N_4573,In_236,In_381);
or U4574 (N_4574,In_463,In_1310);
nand U4575 (N_4575,In_12,In_792);
and U4576 (N_4576,In_1232,In_1017);
and U4577 (N_4577,In_565,In_1433);
and U4578 (N_4578,In_790,In_787);
or U4579 (N_4579,In_45,In_1384);
nor U4580 (N_4580,In_17,In_943);
and U4581 (N_4581,In_882,In_785);
or U4582 (N_4582,In_839,In_68);
nor U4583 (N_4583,In_754,In_596);
nor U4584 (N_4584,In_1446,In_1326);
nor U4585 (N_4585,In_1289,In_1198);
nand U4586 (N_4586,In_339,In_1377);
nand U4587 (N_4587,In_1032,In_814);
nand U4588 (N_4588,In_1057,In_1033);
nand U4589 (N_4589,In_1378,In_368);
nor U4590 (N_4590,In_1117,In_315);
nand U4591 (N_4591,In_1351,In_310);
nor U4592 (N_4592,In_511,In_63);
and U4593 (N_4593,In_1319,In_1162);
nor U4594 (N_4594,In_725,In_39);
nand U4595 (N_4595,In_753,In_1181);
nand U4596 (N_4596,In_943,In_1403);
nor U4597 (N_4597,In_717,In_1272);
nor U4598 (N_4598,In_649,In_1377);
nor U4599 (N_4599,In_1087,In_504);
nor U4600 (N_4600,In_418,In_1105);
nand U4601 (N_4601,In_1382,In_773);
nand U4602 (N_4602,In_913,In_33);
nand U4603 (N_4603,In_464,In_744);
nor U4604 (N_4604,In_244,In_1157);
and U4605 (N_4605,In_287,In_782);
or U4606 (N_4606,In_923,In_427);
nand U4607 (N_4607,In_804,In_966);
nor U4608 (N_4608,In_1438,In_1);
nor U4609 (N_4609,In_408,In_691);
and U4610 (N_4610,In_1471,In_79);
and U4611 (N_4611,In_469,In_1412);
or U4612 (N_4612,In_739,In_1342);
nor U4613 (N_4613,In_352,In_616);
or U4614 (N_4614,In_156,In_229);
or U4615 (N_4615,In_282,In_1174);
nand U4616 (N_4616,In_520,In_27);
and U4617 (N_4617,In_265,In_429);
and U4618 (N_4618,In_1461,In_305);
nand U4619 (N_4619,In_972,In_510);
or U4620 (N_4620,In_425,In_941);
nand U4621 (N_4621,In_1319,In_1260);
and U4622 (N_4622,In_1234,In_660);
xnor U4623 (N_4623,In_1334,In_1380);
nand U4624 (N_4624,In_177,In_354);
nor U4625 (N_4625,In_803,In_590);
and U4626 (N_4626,In_1466,In_357);
nor U4627 (N_4627,In_1215,In_1039);
nor U4628 (N_4628,In_631,In_1054);
and U4629 (N_4629,In_1026,In_850);
xor U4630 (N_4630,In_1135,In_1096);
and U4631 (N_4631,In_550,In_388);
nand U4632 (N_4632,In_1201,In_283);
and U4633 (N_4633,In_1488,In_1416);
and U4634 (N_4634,In_646,In_129);
or U4635 (N_4635,In_550,In_577);
nand U4636 (N_4636,In_543,In_1462);
nor U4637 (N_4637,In_1183,In_186);
nor U4638 (N_4638,In_221,In_886);
nand U4639 (N_4639,In_393,In_905);
nor U4640 (N_4640,In_167,In_772);
or U4641 (N_4641,In_698,In_193);
and U4642 (N_4642,In_312,In_683);
nor U4643 (N_4643,In_1491,In_1272);
and U4644 (N_4644,In_1272,In_1299);
nor U4645 (N_4645,In_871,In_1049);
and U4646 (N_4646,In_237,In_1224);
nor U4647 (N_4647,In_512,In_1336);
nor U4648 (N_4648,In_175,In_1024);
and U4649 (N_4649,In_1141,In_927);
or U4650 (N_4650,In_338,In_450);
nand U4651 (N_4651,In_233,In_819);
nand U4652 (N_4652,In_239,In_36);
and U4653 (N_4653,In_301,In_1227);
or U4654 (N_4654,In_1357,In_1437);
or U4655 (N_4655,In_338,In_45);
and U4656 (N_4656,In_177,In_1181);
or U4657 (N_4657,In_970,In_1229);
and U4658 (N_4658,In_216,In_1321);
and U4659 (N_4659,In_35,In_62);
nand U4660 (N_4660,In_1132,In_1057);
and U4661 (N_4661,In_759,In_965);
nand U4662 (N_4662,In_1384,In_686);
or U4663 (N_4663,In_233,In_210);
or U4664 (N_4664,In_960,In_1185);
and U4665 (N_4665,In_1440,In_1426);
nand U4666 (N_4666,In_535,In_1437);
nor U4667 (N_4667,In_785,In_1174);
nand U4668 (N_4668,In_849,In_789);
nand U4669 (N_4669,In_1115,In_147);
nand U4670 (N_4670,In_539,In_410);
nand U4671 (N_4671,In_710,In_330);
nor U4672 (N_4672,In_335,In_79);
or U4673 (N_4673,In_1286,In_999);
and U4674 (N_4674,In_939,In_337);
xnor U4675 (N_4675,In_737,In_304);
nand U4676 (N_4676,In_694,In_793);
or U4677 (N_4677,In_1343,In_739);
and U4678 (N_4678,In_560,In_686);
nor U4679 (N_4679,In_1341,In_44);
nand U4680 (N_4680,In_253,In_792);
or U4681 (N_4681,In_1289,In_1334);
or U4682 (N_4682,In_1263,In_1376);
and U4683 (N_4683,In_1222,In_1104);
and U4684 (N_4684,In_889,In_318);
and U4685 (N_4685,In_663,In_1388);
or U4686 (N_4686,In_389,In_213);
nor U4687 (N_4687,In_600,In_271);
nor U4688 (N_4688,In_742,In_798);
nand U4689 (N_4689,In_1281,In_1392);
nor U4690 (N_4690,In_529,In_993);
nand U4691 (N_4691,In_430,In_387);
and U4692 (N_4692,In_259,In_915);
nand U4693 (N_4693,In_696,In_297);
or U4694 (N_4694,In_1043,In_21);
nand U4695 (N_4695,In_542,In_5);
or U4696 (N_4696,In_1482,In_667);
nor U4697 (N_4697,In_1088,In_611);
nand U4698 (N_4698,In_971,In_763);
nand U4699 (N_4699,In_320,In_491);
nor U4700 (N_4700,In_130,In_985);
or U4701 (N_4701,In_1020,In_1145);
nand U4702 (N_4702,In_704,In_740);
nor U4703 (N_4703,In_1213,In_1076);
nand U4704 (N_4704,In_498,In_1442);
and U4705 (N_4705,In_1012,In_357);
or U4706 (N_4706,In_249,In_1149);
and U4707 (N_4707,In_1207,In_485);
nor U4708 (N_4708,In_596,In_1425);
and U4709 (N_4709,In_838,In_1428);
and U4710 (N_4710,In_1445,In_524);
and U4711 (N_4711,In_84,In_1448);
nor U4712 (N_4712,In_1444,In_498);
or U4713 (N_4713,In_1308,In_890);
nand U4714 (N_4714,In_1433,In_44);
and U4715 (N_4715,In_1212,In_626);
or U4716 (N_4716,In_928,In_27);
or U4717 (N_4717,In_1419,In_1142);
xor U4718 (N_4718,In_1358,In_289);
nor U4719 (N_4719,In_227,In_1312);
nor U4720 (N_4720,In_269,In_1329);
and U4721 (N_4721,In_490,In_408);
nand U4722 (N_4722,In_1089,In_492);
and U4723 (N_4723,In_1133,In_1278);
and U4724 (N_4724,In_1237,In_992);
nor U4725 (N_4725,In_284,In_200);
nand U4726 (N_4726,In_281,In_766);
nor U4727 (N_4727,In_30,In_510);
or U4728 (N_4728,In_82,In_488);
and U4729 (N_4729,In_372,In_825);
and U4730 (N_4730,In_26,In_296);
or U4731 (N_4731,In_326,In_730);
nand U4732 (N_4732,In_1130,In_1478);
and U4733 (N_4733,In_1284,In_269);
and U4734 (N_4734,In_1012,In_780);
nand U4735 (N_4735,In_1424,In_831);
nand U4736 (N_4736,In_1050,In_979);
nor U4737 (N_4737,In_689,In_237);
nand U4738 (N_4738,In_1188,In_348);
or U4739 (N_4739,In_1330,In_1371);
nor U4740 (N_4740,In_1043,In_115);
or U4741 (N_4741,In_1268,In_88);
nand U4742 (N_4742,In_817,In_1339);
or U4743 (N_4743,In_1273,In_81);
nor U4744 (N_4744,In_901,In_903);
or U4745 (N_4745,In_1416,In_53);
and U4746 (N_4746,In_86,In_1264);
nor U4747 (N_4747,In_378,In_291);
and U4748 (N_4748,In_1422,In_382);
nand U4749 (N_4749,In_228,In_473);
or U4750 (N_4750,In_1318,In_1228);
nor U4751 (N_4751,In_493,In_1460);
and U4752 (N_4752,In_1342,In_401);
and U4753 (N_4753,In_839,In_854);
nand U4754 (N_4754,In_1145,In_341);
and U4755 (N_4755,In_671,In_835);
nor U4756 (N_4756,In_148,In_385);
nand U4757 (N_4757,In_303,In_468);
nand U4758 (N_4758,In_53,In_1111);
nand U4759 (N_4759,In_789,In_1011);
and U4760 (N_4760,In_1403,In_1151);
and U4761 (N_4761,In_880,In_199);
or U4762 (N_4762,In_462,In_1407);
and U4763 (N_4763,In_1440,In_396);
nand U4764 (N_4764,In_1361,In_719);
nand U4765 (N_4765,In_829,In_1468);
and U4766 (N_4766,In_1044,In_772);
nor U4767 (N_4767,In_668,In_1395);
or U4768 (N_4768,In_1475,In_239);
and U4769 (N_4769,In_1276,In_1264);
or U4770 (N_4770,In_238,In_712);
nand U4771 (N_4771,In_900,In_1411);
or U4772 (N_4772,In_1302,In_566);
nor U4773 (N_4773,In_612,In_724);
nor U4774 (N_4774,In_833,In_773);
nor U4775 (N_4775,In_1003,In_518);
xor U4776 (N_4776,In_559,In_1362);
nand U4777 (N_4777,In_1321,In_586);
nor U4778 (N_4778,In_432,In_1103);
nand U4779 (N_4779,In_402,In_730);
and U4780 (N_4780,In_711,In_979);
nor U4781 (N_4781,In_1377,In_1458);
nor U4782 (N_4782,In_99,In_483);
or U4783 (N_4783,In_1281,In_861);
or U4784 (N_4784,In_1177,In_620);
and U4785 (N_4785,In_131,In_839);
or U4786 (N_4786,In_190,In_127);
and U4787 (N_4787,In_1410,In_761);
nand U4788 (N_4788,In_223,In_1493);
and U4789 (N_4789,In_995,In_677);
and U4790 (N_4790,In_1356,In_592);
nor U4791 (N_4791,In_102,In_998);
nand U4792 (N_4792,In_1015,In_585);
nor U4793 (N_4793,In_1289,In_1312);
and U4794 (N_4794,In_975,In_1433);
nand U4795 (N_4795,In_1377,In_683);
nor U4796 (N_4796,In_666,In_673);
and U4797 (N_4797,In_1040,In_595);
nor U4798 (N_4798,In_1058,In_342);
nand U4799 (N_4799,In_1025,In_1394);
or U4800 (N_4800,In_234,In_1201);
or U4801 (N_4801,In_939,In_808);
nand U4802 (N_4802,In_402,In_667);
or U4803 (N_4803,In_1373,In_1166);
or U4804 (N_4804,In_446,In_1362);
nor U4805 (N_4805,In_514,In_1151);
or U4806 (N_4806,In_1071,In_1163);
nand U4807 (N_4807,In_324,In_1231);
nand U4808 (N_4808,In_812,In_391);
and U4809 (N_4809,In_1172,In_594);
or U4810 (N_4810,In_285,In_1241);
nor U4811 (N_4811,In_902,In_617);
xor U4812 (N_4812,In_740,In_1097);
or U4813 (N_4813,In_973,In_949);
nand U4814 (N_4814,In_740,In_138);
nand U4815 (N_4815,In_972,In_1038);
or U4816 (N_4816,In_1026,In_704);
and U4817 (N_4817,In_735,In_288);
nand U4818 (N_4818,In_636,In_222);
and U4819 (N_4819,In_339,In_443);
or U4820 (N_4820,In_219,In_43);
and U4821 (N_4821,In_811,In_1001);
and U4822 (N_4822,In_1405,In_1301);
nor U4823 (N_4823,In_1090,In_317);
nor U4824 (N_4824,In_1160,In_515);
nor U4825 (N_4825,In_1182,In_21);
nor U4826 (N_4826,In_1498,In_1422);
nor U4827 (N_4827,In_831,In_1385);
and U4828 (N_4828,In_28,In_1193);
nor U4829 (N_4829,In_296,In_1160);
or U4830 (N_4830,In_707,In_1477);
nand U4831 (N_4831,In_603,In_1474);
nor U4832 (N_4832,In_1166,In_19);
or U4833 (N_4833,In_44,In_94);
nor U4834 (N_4834,In_227,In_460);
or U4835 (N_4835,In_634,In_13);
nor U4836 (N_4836,In_477,In_304);
nand U4837 (N_4837,In_221,In_97);
or U4838 (N_4838,In_860,In_854);
nand U4839 (N_4839,In_919,In_1463);
nor U4840 (N_4840,In_95,In_919);
nand U4841 (N_4841,In_1150,In_1172);
and U4842 (N_4842,In_436,In_1103);
nor U4843 (N_4843,In_1479,In_648);
nand U4844 (N_4844,In_764,In_1213);
and U4845 (N_4845,In_938,In_312);
nand U4846 (N_4846,In_935,In_455);
nor U4847 (N_4847,In_929,In_971);
or U4848 (N_4848,In_753,In_354);
nand U4849 (N_4849,In_553,In_700);
nand U4850 (N_4850,In_554,In_210);
or U4851 (N_4851,In_1331,In_610);
and U4852 (N_4852,In_481,In_1348);
nand U4853 (N_4853,In_1158,In_813);
and U4854 (N_4854,In_1112,In_307);
and U4855 (N_4855,In_908,In_252);
or U4856 (N_4856,In_1370,In_292);
or U4857 (N_4857,In_76,In_1043);
nor U4858 (N_4858,In_581,In_778);
or U4859 (N_4859,In_1278,In_121);
or U4860 (N_4860,In_618,In_163);
or U4861 (N_4861,In_1480,In_126);
nand U4862 (N_4862,In_399,In_131);
nor U4863 (N_4863,In_439,In_606);
and U4864 (N_4864,In_1014,In_1267);
or U4865 (N_4865,In_1479,In_1123);
nor U4866 (N_4866,In_731,In_1346);
and U4867 (N_4867,In_1232,In_1433);
and U4868 (N_4868,In_213,In_1440);
or U4869 (N_4869,In_1466,In_112);
or U4870 (N_4870,In_1320,In_570);
and U4871 (N_4871,In_505,In_97);
or U4872 (N_4872,In_683,In_591);
nand U4873 (N_4873,In_114,In_675);
or U4874 (N_4874,In_774,In_1460);
nor U4875 (N_4875,In_1219,In_1391);
or U4876 (N_4876,In_676,In_433);
nor U4877 (N_4877,In_1398,In_40);
or U4878 (N_4878,In_1148,In_282);
and U4879 (N_4879,In_453,In_650);
or U4880 (N_4880,In_957,In_1390);
and U4881 (N_4881,In_1386,In_575);
nor U4882 (N_4882,In_1264,In_1094);
and U4883 (N_4883,In_1060,In_1151);
and U4884 (N_4884,In_1313,In_1326);
nand U4885 (N_4885,In_693,In_184);
or U4886 (N_4886,In_1249,In_1402);
and U4887 (N_4887,In_1386,In_683);
or U4888 (N_4888,In_1431,In_709);
nand U4889 (N_4889,In_77,In_1463);
nor U4890 (N_4890,In_699,In_1393);
nor U4891 (N_4891,In_1225,In_771);
or U4892 (N_4892,In_1477,In_1112);
nand U4893 (N_4893,In_891,In_1464);
nand U4894 (N_4894,In_643,In_484);
nor U4895 (N_4895,In_1248,In_462);
nand U4896 (N_4896,In_213,In_624);
or U4897 (N_4897,In_740,In_1124);
and U4898 (N_4898,In_472,In_720);
or U4899 (N_4899,In_553,In_223);
and U4900 (N_4900,In_60,In_1282);
nand U4901 (N_4901,In_1308,In_595);
nand U4902 (N_4902,In_335,In_191);
nand U4903 (N_4903,In_22,In_747);
nor U4904 (N_4904,In_625,In_813);
nand U4905 (N_4905,In_1241,In_1400);
nand U4906 (N_4906,In_1391,In_510);
and U4907 (N_4907,In_690,In_173);
or U4908 (N_4908,In_518,In_1351);
nand U4909 (N_4909,In_866,In_1086);
nor U4910 (N_4910,In_1236,In_930);
and U4911 (N_4911,In_584,In_1474);
nor U4912 (N_4912,In_473,In_938);
nand U4913 (N_4913,In_217,In_1294);
nand U4914 (N_4914,In_1414,In_423);
nor U4915 (N_4915,In_68,In_896);
nand U4916 (N_4916,In_1066,In_905);
nor U4917 (N_4917,In_613,In_1079);
nand U4918 (N_4918,In_40,In_816);
or U4919 (N_4919,In_736,In_1078);
nand U4920 (N_4920,In_1232,In_255);
nor U4921 (N_4921,In_914,In_560);
and U4922 (N_4922,In_417,In_297);
or U4923 (N_4923,In_736,In_748);
or U4924 (N_4924,In_1419,In_1189);
and U4925 (N_4925,In_842,In_1407);
nand U4926 (N_4926,In_195,In_241);
and U4927 (N_4927,In_197,In_167);
or U4928 (N_4928,In_783,In_1014);
nand U4929 (N_4929,In_541,In_1321);
nand U4930 (N_4930,In_743,In_445);
or U4931 (N_4931,In_5,In_725);
xnor U4932 (N_4932,In_744,In_403);
nor U4933 (N_4933,In_1358,In_229);
nand U4934 (N_4934,In_1267,In_1466);
xnor U4935 (N_4935,In_491,In_151);
and U4936 (N_4936,In_1340,In_1077);
or U4937 (N_4937,In_219,In_1465);
nand U4938 (N_4938,In_831,In_375);
nand U4939 (N_4939,In_1005,In_971);
nand U4940 (N_4940,In_1454,In_1182);
and U4941 (N_4941,In_1143,In_1264);
nand U4942 (N_4942,In_1238,In_1125);
nor U4943 (N_4943,In_108,In_1054);
nand U4944 (N_4944,In_677,In_140);
or U4945 (N_4945,In_620,In_896);
or U4946 (N_4946,In_209,In_1214);
and U4947 (N_4947,In_143,In_187);
and U4948 (N_4948,In_1008,In_901);
and U4949 (N_4949,In_427,In_406);
nor U4950 (N_4950,In_1213,In_1439);
and U4951 (N_4951,In_788,In_1047);
xor U4952 (N_4952,In_639,In_1110);
or U4953 (N_4953,In_477,In_529);
or U4954 (N_4954,In_76,In_86);
nand U4955 (N_4955,In_1064,In_260);
nor U4956 (N_4956,In_1001,In_987);
and U4957 (N_4957,In_1055,In_1132);
and U4958 (N_4958,In_646,In_334);
nor U4959 (N_4959,In_125,In_661);
nand U4960 (N_4960,In_259,In_1000);
nor U4961 (N_4961,In_1024,In_1365);
nand U4962 (N_4962,In_682,In_1201);
or U4963 (N_4963,In_761,In_544);
nand U4964 (N_4964,In_1187,In_1376);
or U4965 (N_4965,In_1346,In_715);
or U4966 (N_4966,In_538,In_1128);
and U4967 (N_4967,In_1414,In_1241);
nor U4968 (N_4968,In_573,In_1443);
nand U4969 (N_4969,In_1499,In_1403);
and U4970 (N_4970,In_388,In_111);
nand U4971 (N_4971,In_211,In_1103);
and U4972 (N_4972,In_417,In_162);
nor U4973 (N_4973,In_1075,In_1188);
nor U4974 (N_4974,In_1035,In_53);
nor U4975 (N_4975,In_530,In_632);
or U4976 (N_4976,In_808,In_628);
and U4977 (N_4977,In_391,In_1280);
or U4978 (N_4978,In_1373,In_834);
and U4979 (N_4979,In_1397,In_253);
or U4980 (N_4980,In_668,In_891);
or U4981 (N_4981,In_1169,In_901);
nand U4982 (N_4982,In_1087,In_1450);
nor U4983 (N_4983,In_1289,In_843);
nor U4984 (N_4984,In_1301,In_950);
or U4985 (N_4985,In_1231,In_172);
or U4986 (N_4986,In_723,In_34);
nor U4987 (N_4987,In_232,In_694);
or U4988 (N_4988,In_1186,In_1237);
and U4989 (N_4989,In_1270,In_1321);
and U4990 (N_4990,In_263,In_1037);
and U4991 (N_4991,In_1445,In_12);
or U4992 (N_4992,In_1483,In_482);
nor U4993 (N_4993,In_937,In_761);
or U4994 (N_4994,In_723,In_1440);
and U4995 (N_4995,In_630,In_1199);
and U4996 (N_4996,In_1281,In_59);
nor U4997 (N_4997,In_691,In_1171);
nor U4998 (N_4998,In_377,In_691);
nor U4999 (N_4999,In_1265,In_714);
or U5000 (N_5000,N_2247,N_1314);
nand U5001 (N_5001,N_4819,N_3065);
nor U5002 (N_5002,N_3322,N_2179);
or U5003 (N_5003,N_3189,N_875);
or U5004 (N_5004,N_889,N_4828);
or U5005 (N_5005,N_3527,N_4098);
nand U5006 (N_5006,N_4724,N_3645);
or U5007 (N_5007,N_3644,N_4435);
and U5008 (N_5008,N_1562,N_2602);
and U5009 (N_5009,N_1865,N_39);
nor U5010 (N_5010,N_1615,N_1952);
xor U5011 (N_5011,N_2155,N_2612);
nor U5012 (N_5012,N_807,N_2005);
nand U5013 (N_5013,N_1520,N_3425);
nand U5014 (N_5014,N_3746,N_3966);
or U5015 (N_5015,N_420,N_4348);
nand U5016 (N_5016,N_3837,N_1488);
nand U5017 (N_5017,N_3371,N_4984);
nand U5018 (N_5018,N_2882,N_2771);
nor U5019 (N_5019,N_2153,N_4167);
or U5020 (N_5020,N_203,N_2885);
and U5021 (N_5021,N_2654,N_3346);
nor U5022 (N_5022,N_1713,N_2187);
nor U5023 (N_5023,N_3175,N_4970);
nor U5024 (N_5024,N_3859,N_3506);
nand U5025 (N_5025,N_4558,N_4257);
and U5026 (N_5026,N_4561,N_1547);
or U5027 (N_5027,N_3730,N_2734);
nor U5028 (N_5028,N_852,N_295);
and U5029 (N_5029,N_1738,N_558);
nand U5030 (N_5030,N_2923,N_3305);
nor U5031 (N_5031,N_4459,N_1822);
and U5032 (N_5032,N_2942,N_3142);
nor U5033 (N_5033,N_3570,N_1475);
nor U5034 (N_5034,N_4507,N_1681);
or U5035 (N_5035,N_4996,N_2931);
nor U5036 (N_5036,N_3917,N_7);
and U5037 (N_5037,N_1332,N_3135);
or U5038 (N_5038,N_2954,N_1744);
nor U5039 (N_5039,N_4600,N_3113);
or U5040 (N_5040,N_1984,N_1135);
nor U5041 (N_5041,N_416,N_4947);
nand U5042 (N_5042,N_974,N_2304);
nand U5043 (N_5043,N_929,N_4519);
nand U5044 (N_5044,N_4451,N_4656);
nor U5045 (N_5045,N_1431,N_2755);
nand U5046 (N_5046,N_4915,N_42);
or U5047 (N_5047,N_3407,N_3347);
nor U5048 (N_5048,N_2126,N_3035);
nor U5049 (N_5049,N_2108,N_1981);
nand U5050 (N_5050,N_3126,N_2461);
or U5051 (N_5051,N_4699,N_1381);
or U5052 (N_5052,N_3516,N_2386);
and U5053 (N_5053,N_615,N_4412);
nor U5054 (N_5054,N_4126,N_1651);
nor U5055 (N_5055,N_973,N_3653);
or U5056 (N_5056,N_4368,N_4843);
nand U5057 (N_5057,N_759,N_1491);
and U5058 (N_5058,N_4616,N_3446);
nand U5059 (N_5059,N_1495,N_3424);
nand U5060 (N_5060,N_391,N_3463);
or U5061 (N_5061,N_898,N_2902);
and U5062 (N_5062,N_347,N_583);
nor U5063 (N_5063,N_4580,N_4246);
nand U5064 (N_5064,N_4465,N_2392);
or U5065 (N_5065,N_3615,N_1468);
nor U5066 (N_5066,N_2395,N_658);
or U5067 (N_5067,N_471,N_4695);
or U5068 (N_5068,N_1511,N_1494);
or U5069 (N_5069,N_1800,N_3833);
or U5070 (N_5070,N_1899,N_2312);
nand U5071 (N_5071,N_1466,N_3408);
and U5072 (N_5072,N_2117,N_341);
and U5073 (N_5073,N_156,N_2029);
nand U5074 (N_5074,N_2008,N_4491);
or U5075 (N_5075,N_1712,N_4788);
nand U5076 (N_5076,N_1594,N_3103);
nand U5077 (N_5077,N_1557,N_4867);
xnor U5078 (N_5078,N_1105,N_3010);
or U5079 (N_5079,N_329,N_4881);
nor U5080 (N_5080,N_590,N_4954);
and U5081 (N_5081,N_2663,N_1196);
nand U5082 (N_5082,N_2977,N_2678);
nor U5083 (N_5083,N_3637,N_1008);
and U5084 (N_5084,N_3068,N_1656);
nor U5085 (N_5085,N_163,N_1815);
nand U5086 (N_5086,N_4234,N_4887);
or U5087 (N_5087,N_530,N_3318);
nor U5088 (N_5088,N_3665,N_4419);
or U5089 (N_5089,N_1393,N_953);
or U5090 (N_5090,N_4055,N_736);
and U5091 (N_5091,N_57,N_433);
nor U5092 (N_5092,N_3695,N_1913);
nand U5093 (N_5093,N_2082,N_1757);
nor U5094 (N_5094,N_3490,N_527);
nor U5095 (N_5095,N_4601,N_1686);
nor U5096 (N_5096,N_2614,N_4801);
nand U5097 (N_5097,N_4012,N_3051);
and U5098 (N_5098,N_1746,N_2397);
nand U5099 (N_5099,N_2537,N_3817);
nor U5100 (N_5100,N_4693,N_4502);
or U5101 (N_5101,N_2487,N_3526);
nand U5102 (N_5102,N_1229,N_4050);
nand U5103 (N_5103,N_3763,N_2100);
and U5104 (N_5104,N_3043,N_3206);
and U5105 (N_5105,N_3134,N_1405);
and U5106 (N_5106,N_1385,N_89);
nand U5107 (N_5107,N_1352,N_3816);
nand U5108 (N_5108,N_2957,N_2698);
nor U5109 (N_5109,N_2054,N_2809);
and U5110 (N_5110,N_4595,N_3618);
xor U5111 (N_5111,N_3078,N_1602);
nand U5112 (N_5112,N_1638,N_1931);
and U5113 (N_5113,N_2789,N_2267);
nor U5114 (N_5114,N_1817,N_303);
nand U5115 (N_5115,N_1426,N_1764);
and U5116 (N_5116,N_4906,N_2798);
and U5117 (N_5117,N_2225,N_4065);
nand U5118 (N_5118,N_33,N_2509);
or U5119 (N_5119,N_3053,N_79);
or U5120 (N_5120,N_2582,N_1218);
or U5121 (N_5121,N_2571,N_2518);
nor U5122 (N_5122,N_2050,N_3168);
and U5123 (N_5123,N_171,N_3931);
and U5124 (N_5124,N_950,N_2817);
and U5125 (N_5125,N_1222,N_3964);
nand U5126 (N_5126,N_584,N_4909);
or U5127 (N_5127,N_3772,N_3231);
or U5128 (N_5128,N_1804,N_2619);
nor U5129 (N_5129,N_2114,N_2468);
nand U5130 (N_5130,N_49,N_3520);
or U5131 (N_5131,N_3034,N_3604);
nor U5132 (N_5132,N_964,N_4272);
or U5133 (N_5133,N_4883,N_575);
or U5134 (N_5134,N_4112,N_1964);
or U5135 (N_5135,N_1716,N_2198);
or U5136 (N_5136,N_4453,N_4344);
and U5137 (N_5137,N_2209,N_1958);
nor U5138 (N_5138,N_826,N_747);
nor U5139 (N_5139,N_3421,N_3088);
and U5140 (N_5140,N_1851,N_1917);
or U5141 (N_5141,N_1502,N_3442);
nor U5142 (N_5142,N_2097,N_513);
nand U5143 (N_5143,N_458,N_1489);
nor U5144 (N_5144,N_991,N_348);
or U5145 (N_5145,N_1787,N_236);
nor U5146 (N_5146,N_2900,N_144);
nor U5147 (N_5147,N_3555,N_582);
nor U5148 (N_5148,N_1420,N_1048);
and U5149 (N_5149,N_1776,N_4751);
or U5150 (N_5150,N_3148,N_4575);
nand U5151 (N_5151,N_2642,N_1191);
and U5152 (N_5152,N_790,N_2206);
or U5153 (N_5153,N_4783,N_1953);
nand U5154 (N_5154,N_967,N_3070);
nand U5155 (N_5155,N_2166,N_1663);
nor U5156 (N_5156,N_714,N_4109);
and U5157 (N_5157,N_1038,N_4389);
and U5158 (N_5158,N_2903,N_309);
or U5159 (N_5159,N_971,N_834);
and U5160 (N_5160,N_4455,N_3758);
or U5161 (N_5161,N_2963,N_2924);
and U5162 (N_5162,N_4392,N_3419);
nand U5163 (N_5163,N_2528,N_1625);
and U5164 (N_5164,N_4129,N_2914);
or U5165 (N_5165,N_2713,N_4586);
xnor U5166 (N_5166,N_3416,N_3119);
nand U5167 (N_5167,N_4152,N_997);
and U5168 (N_5168,N_3578,N_1544);
or U5169 (N_5169,N_3389,N_3289);
nor U5170 (N_5170,N_3215,N_105);
nand U5171 (N_5171,N_4622,N_4629);
nor U5172 (N_5172,N_3806,N_4681);
nand U5173 (N_5173,N_4054,N_3650);
nand U5174 (N_5174,N_2779,N_2139);
nand U5175 (N_5175,N_4767,N_4840);
and U5176 (N_5176,N_4937,N_4916);
or U5177 (N_5177,N_2142,N_2735);
or U5178 (N_5178,N_3176,N_4140);
and U5179 (N_5179,N_2877,N_1448);
nor U5180 (N_5180,N_1153,N_4671);
or U5181 (N_5181,N_4748,N_4525);
and U5182 (N_5182,N_778,N_2157);
nor U5183 (N_5183,N_77,N_4426);
nor U5184 (N_5184,N_267,N_1487);
and U5185 (N_5185,N_436,N_2913);
nor U5186 (N_5186,N_1202,N_849);
nor U5187 (N_5187,N_32,N_3487);
or U5188 (N_5188,N_2937,N_4070);
and U5189 (N_5189,N_2884,N_4479);
nor U5190 (N_5190,N_861,N_3828);
nand U5191 (N_5191,N_2405,N_4544);
nor U5192 (N_5192,N_2423,N_1704);
nor U5193 (N_5193,N_4277,N_36);
or U5194 (N_5194,N_3836,N_1792);
or U5195 (N_5195,N_73,N_1181);
nor U5196 (N_5196,N_1666,N_37);
nand U5197 (N_5197,N_4939,N_2736);
nor U5198 (N_5198,N_1,N_4838);
nor U5199 (N_5199,N_4706,N_1234);
and U5200 (N_5200,N_4709,N_2580);
nand U5201 (N_5201,N_2857,N_760);
nor U5202 (N_5202,N_2645,N_804);
nor U5203 (N_5203,N_389,N_3197);
or U5204 (N_5204,N_625,N_4149);
or U5205 (N_5205,N_4897,N_2228);
and U5206 (N_5206,N_913,N_3157);
and U5207 (N_5207,N_1252,N_3703);
nand U5208 (N_5208,N_638,N_187);
and U5209 (N_5209,N_1015,N_3685);
or U5210 (N_5210,N_1465,N_3085);
nand U5211 (N_5211,N_2714,N_498);
or U5212 (N_5212,N_4036,N_3447);
and U5213 (N_5213,N_453,N_3395);
nor U5214 (N_5214,N_2001,N_2411);
nand U5215 (N_5215,N_4279,N_2687);
nand U5216 (N_5216,N_1144,N_226);
xnor U5217 (N_5217,N_4638,N_4998);
or U5218 (N_5218,N_2432,N_2434);
or U5219 (N_5219,N_1344,N_2607);
or U5220 (N_5220,N_881,N_3659);
or U5221 (N_5221,N_659,N_933);
and U5222 (N_5222,N_4085,N_4782);
nand U5223 (N_5223,N_3845,N_3500);
xnor U5224 (N_5224,N_2065,N_4002);
and U5225 (N_5225,N_3723,N_2326);
or U5226 (N_5226,N_4742,N_4566);
or U5227 (N_5227,N_4687,N_1988);
nand U5228 (N_5228,N_4677,N_721);
or U5229 (N_5229,N_3954,N_312);
and U5230 (N_5230,N_4193,N_845);
nor U5231 (N_5231,N_1578,N_99);
or U5232 (N_5232,N_3603,N_3803);
nor U5233 (N_5233,N_4361,N_3584);
nor U5234 (N_5234,N_3023,N_4933);
nand U5235 (N_5235,N_4532,N_160);
nor U5236 (N_5236,N_3542,N_3856);
or U5237 (N_5237,N_992,N_1652);
nand U5238 (N_5238,N_2699,N_763);
and U5239 (N_5239,N_2656,N_1831);
nor U5240 (N_5240,N_2465,N_2115);
nor U5241 (N_5241,N_3907,N_4164);
and U5242 (N_5242,N_2149,N_2623);
and U5243 (N_5243,N_2071,N_3654);
nor U5244 (N_5244,N_2904,N_4541);
xnor U5245 (N_5245,N_543,N_4370);
or U5246 (N_5246,N_1622,N_3064);
nand U5247 (N_5247,N_3409,N_1205);
nand U5248 (N_5248,N_3171,N_961);
nand U5249 (N_5249,N_637,N_4688);
or U5250 (N_5250,N_3108,N_4609);
nand U5251 (N_5251,N_3201,N_1143);
nor U5252 (N_5252,N_428,N_2995);
nor U5253 (N_5253,N_4860,N_1493);
and U5254 (N_5254,N_266,N_2055);
nand U5255 (N_5255,N_2803,N_633);
and U5256 (N_5256,N_3292,N_1537);
nor U5257 (N_5257,N_1437,N_2310);
nor U5258 (N_5258,N_699,N_3750);
nand U5259 (N_5259,N_446,N_2451);
or U5260 (N_5260,N_4318,N_579);
nor U5261 (N_5261,N_2868,N_1347);
xnor U5262 (N_5262,N_3272,N_3412);
or U5263 (N_5263,N_2987,N_4833);
nand U5264 (N_5264,N_4343,N_1149);
and U5265 (N_5265,N_905,N_4325);
and U5266 (N_5266,N_3307,N_4878);
nand U5267 (N_5267,N_3749,N_4614);
or U5268 (N_5268,N_231,N_1640);
nor U5269 (N_5269,N_2673,N_406);
or U5270 (N_5270,N_3473,N_544);
nand U5271 (N_5271,N_4991,N_4127);
nor U5272 (N_5272,N_1406,N_2940);
nor U5273 (N_5273,N_4401,N_1159);
nand U5274 (N_5274,N_3699,N_2210);
or U5275 (N_5275,N_4730,N_3461);
nor U5276 (N_5276,N_4295,N_2674);
and U5277 (N_5277,N_4873,N_529);
or U5278 (N_5278,N_2638,N_1337);
nand U5279 (N_5279,N_2060,N_3698);
and U5280 (N_5280,N_3511,N_4224);
nand U5281 (N_5281,N_2738,N_4356);
nand U5282 (N_5282,N_1902,N_2222);
or U5283 (N_5283,N_4846,N_4205);
nand U5284 (N_5284,N_1858,N_1490);
nor U5285 (N_5285,N_2531,N_3296);
nor U5286 (N_5286,N_2791,N_3259);
and U5287 (N_5287,N_176,N_1932);
nor U5288 (N_5288,N_3054,N_2551);
or U5289 (N_5289,N_3980,N_2066);
nor U5290 (N_5290,N_2109,N_2358);
nor U5291 (N_5291,N_151,N_1797);
or U5292 (N_5292,N_4766,N_3988);
nor U5293 (N_5293,N_577,N_2070);
or U5294 (N_5294,N_2390,N_4326);
and U5295 (N_5295,N_724,N_92);
and U5296 (N_5296,N_1777,N_3913);
nand U5297 (N_5297,N_573,N_3592);
and U5298 (N_5298,N_1221,N_940);
or U5299 (N_5299,N_2579,N_3013);
or U5300 (N_5300,N_3912,N_4265);
nand U5301 (N_5301,N_1390,N_4090);
nand U5302 (N_5302,N_1302,N_1325);
or U5303 (N_5303,N_1660,N_4570);
or U5304 (N_5304,N_1855,N_3634);
or U5305 (N_5305,N_2154,N_2372);
and U5306 (N_5306,N_1694,N_3969);
and U5307 (N_5307,N_1854,N_536);
or U5308 (N_5308,N_2846,N_521);
and U5309 (N_5309,N_1910,N_4147);
nand U5310 (N_5310,N_2536,N_635);
nor U5311 (N_5311,N_2554,N_4869);
and U5312 (N_5312,N_3846,N_2403);
nor U5313 (N_5313,N_1965,N_2521);
nor U5314 (N_5314,N_1410,N_2766);
nor U5315 (N_5315,N_3312,N_4627);
or U5316 (N_5316,N_677,N_4437);
nand U5317 (N_5317,N_3945,N_2681);
and U5318 (N_5318,N_35,N_2319);
and U5319 (N_5319,N_4832,N_3309);
and U5320 (N_5320,N_3338,N_4274);
and U5321 (N_5321,N_3378,N_382);
nand U5322 (N_5322,N_3809,N_1190);
and U5323 (N_5323,N_434,N_1146);
or U5324 (N_5324,N_2804,N_610);
nor U5325 (N_5325,N_142,N_2653);
nand U5326 (N_5326,N_2493,N_2724);
and U5327 (N_5327,N_4702,N_1481);
and U5328 (N_5328,N_123,N_1185);
nand U5329 (N_5329,N_1457,N_4300);
nand U5330 (N_5330,N_3124,N_4817);
nand U5331 (N_5331,N_3715,N_4088);
and U5332 (N_5332,N_3748,N_4539);
nor U5333 (N_5333,N_3679,N_762);
and U5334 (N_5334,N_3939,N_2233);
or U5335 (N_5335,N_3232,N_3741);
or U5336 (N_5336,N_2510,N_2786);
and U5337 (N_5337,N_1513,N_4245);
nand U5338 (N_5338,N_1977,N_4722);
nand U5339 (N_5339,N_2159,N_3742);
nand U5340 (N_5340,N_4836,N_3218);
or U5341 (N_5341,N_3514,N_1691);
and U5342 (N_5342,N_3936,N_702);
nand U5343 (N_5343,N_3165,N_4146);
or U5344 (N_5344,N_505,N_1606);
nand U5345 (N_5345,N_4000,N_2839);
nor U5346 (N_5346,N_2701,N_1152);
and U5347 (N_5347,N_3989,N_4094);
or U5348 (N_5348,N_3569,N_1950);
and U5349 (N_5349,N_361,N_3680);
nor U5350 (N_5350,N_4841,N_2106);
or U5351 (N_5351,N_1951,N_1091);
or U5352 (N_5352,N_3766,N_645);
nand U5353 (N_5353,N_4095,N_1345);
and U5354 (N_5354,N_3100,N_4449);
nand U5355 (N_5355,N_3564,N_3160);
and U5356 (N_5356,N_3496,N_4689);
and U5357 (N_5357,N_1673,N_1267);
nor U5358 (N_5358,N_2934,N_2123);
nand U5359 (N_5359,N_631,N_4241);
or U5360 (N_5360,N_469,N_3812);
nand U5361 (N_5361,N_2966,N_3897);
nor U5362 (N_5362,N_1469,N_96);
or U5363 (N_5363,N_1005,N_3243);
nand U5364 (N_5364,N_4639,N_1370);
nor U5365 (N_5365,N_1549,N_4930);
or U5366 (N_5366,N_2852,N_3454);
nand U5367 (N_5367,N_2428,N_2000);
xor U5368 (N_5368,N_3965,N_580);
nand U5369 (N_5369,N_2746,N_2460);
nand U5370 (N_5370,N_3001,N_1862);
nand U5371 (N_5371,N_4045,N_1912);
nor U5372 (N_5372,N_88,N_2811);
nand U5373 (N_5373,N_1654,N_657);
and U5374 (N_5374,N_3994,N_4131);
xnor U5375 (N_5375,N_1526,N_235);
or U5376 (N_5376,N_4630,N_2258);
or U5377 (N_5377,N_1085,N_2031);
nand U5378 (N_5378,N_765,N_4642);
and U5379 (N_5379,N_983,N_545);
or U5380 (N_5380,N_2671,N_2637);
or U5381 (N_5381,N_738,N_4776);
and U5382 (N_5382,N_4189,N_825);
and U5383 (N_5383,N_4905,N_3890);
or U5384 (N_5384,N_3428,N_3952);
nand U5385 (N_5385,N_2611,N_2784);
nor U5386 (N_5386,N_3238,N_1885);
xnor U5387 (N_5387,N_1446,N_506);
and U5388 (N_5388,N_1035,N_3074);
or U5389 (N_5389,N_3513,N_1591);
nand U5390 (N_5390,N_4168,N_4078);
and U5391 (N_5391,N_2519,N_4211);
nand U5392 (N_5392,N_4966,N_651);
and U5393 (N_5393,N_1053,N_4461);
or U5394 (N_5394,N_2053,N_553);
and U5395 (N_5395,N_2245,N_2767);
nor U5396 (N_5396,N_3785,N_1546);
or U5397 (N_5397,N_429,N_565);
or U5398 (N_5398,N_3501,N_218);
or U5399 (N_5399,N_387,N_1067);
nand U5400 (N_5400,N_334,N_4963);
and U5401 (N_5401,N_2776,N_4120);
nand U5402 (N_5402,N_1366,N_3867);
nand U5403 (N_5403,N_4548,N_3609);
or U5404 (N_5404,N_3303,N_4750);
or U5405 (N_5405,N_4014,N_4402);
nand U5406 (N_5406,N_1721,N_415);
or U5407 (N_5407,N_192,N_2613);
nor U5408 (N_5408,N_2028,N_398);
and U5409 (N_5409,N_2476,N_1768);
nand U5410 (N_5410,N_261,N_1667);
nor U5411 (N_5411,N_2315,N_4135);
and U5412 (N_5412,N_116,N_3476);
nand U5413 (N_5413,N_4394,N_492);
nor U5414 (N_5414,N_2124,N_481);
nand U5415 (N_5415,N_2418,N_239);
nor U5416 (N_5416,N_4114,N_1975);
nand U5417 (N_5417,N_3063,N_379);
nand U5418 (N_5418,N_1263,N_1970);
nand U5419 (N_5419,N_4068,N_2928);
nand U5420 (N_5420,N_3862,N_1641);
and U5421 (N_5421,N_706,N_3884);
or U5422 (N_5422,N_1772,N_2533);
nand U5423 (N_5423,N_1158,N_1324);
nand U5424 (N_5424,N_1432,N_2978);
and U5425 (N_5425,N_3217,N_1948);
nand U5426 (N_5426,N_856,N_4810);
nor U5427 (N_5427,N_3342,N_3082);
nor U5428 (N_5428,N_2834,N_1046);
nand U5429 (N_5429,N_4229,N_1006);
and U5430 (N_5430,N_3102,N_161);
nand U5431 (N_5431,N_1901,N_846);
and U5432 (N_5432,N_2158,N_4864);
and U5433 (N_5433,N_1188,N_3136);
nor U5434 (N_5434,N_2458,N_3277);
nor U5435 (N_5435,N_468,N_4529);
and U5436 (N_5436,N_1639,N_2262);
or U5437 (N_5437,N_3616,N_4569);
nand U5438 (N_5438,N_1259,N_2442);
nor U5439 (N_5439,N_4369,N_2912);
and U5440 (N_5440,N_2601,N_4852);
and U5441 (N_5441,N_806,N_177);
nand U5442 (N_5442,N_3387,N_4926);
nor U5443 (N_5443,N_4849,N_1371);
nand U5444 (N_5444,N_3237,N_735);
and U5445 (N_5445,N_3125,N_3686);
and U5446 (N_5446,N_15,N_2865);
and U5447 (N_5447,N_4631,N_1269);
nand U5448 (N_5448,N_4943,N_1171);
nor U5449 (N_5449,N_1456,N_3694);
and U5450 (N_5450,N_2345,N_2086);
and U5451 (N_5451,N_1102,N_655);
and U5452 (N_5452,N_2726,N_894);
nand U5453 (N_5453,N_4433,N_2200);
xor U5454 (N_5454,N_3904,N_3398);
nand U5455 (N_5455,N_1076,N_4587);
nor U5456 (N_5456,N_4212,N_4781);
nand U5457 (N_5457,N_4200,N_299);
and U5458 (N_5458,N_3707,N_3090);
or U5459 (N_5459,N_2965,N_883);
or U5460 (N_5460,N_1966,N_4216);
nor U5461 (N_5461,N_2858,N_535);
or U5462 (N_5462,N_3976,N_3820);
and U5463 (N_5463,N_130,N_2953);
or U5464 (N_5464,N_2705,N_3316);
nor U5465 (N_5465,N_906,N_3340);
nor U5466 (N_5466,N_126,N_1524);
and U5467 (N_5467,N_4907,N_485);
or U5468 (N_5468,N_3799,N_3839);
nand U5469 (N_5469,N_3778,N_1329);
and U5470 (N_5470,N_740,N_548);
nand U5471 (N_5471,N_1206,N_31);
nand U5472 (N_5472,N_3236,N_586);
or U5473 (N_5473,N_1870,N_4307);
or U5474 (N_5474,N_355,N_817);
and U5475 (N_5475,N_3401,N_4624);
or U5476 (N_5476,N_3978,N_4927);
or U5477 (N_5477,N_2552,N_1200);
and U5478 (N_5478,N_118,N_1924);
or U5479 (N_5479,N_1725,N_1552);
nor U5480 (N_5480,N_4740,N_1223);
and U5481 (N_5481,N_431,N_1353);
nand U5482 (N_5482,N_3345,N_1014);
and U5483 (N_5483,N_514,N_3492);
nor U5484 (N_5484,N_2983,N_3561);
or U5485 (N_5485,N_3355,N_4238);
nor U5486 (N_5486,N_164,N_3574);
nand U5487 (N_5487,N_2318,N_85);
and U5488 (N_5488,N_133,N_4005);
or U5489 (N_5489,N_3098,N_4559);
nor U5490 (N_5490,N_2414,N_4715);
nor U5491 (N_5491,N_3747,N_1799);
and U5492 (N_5492,N_3629,N_776);
and U5493 (N_5493,N_1589,N_3911);
or U5494 (N_5494,N_915,N_540);
nand U5495 (N_5495,N_2491,N_3497);
nand U5496 (N_5496,N_1750,N_4469);
nand U5497 (N_5497,N_3842,N_4266);
and U5498 (N_5498,N_4008,N_4117);
or U5499 (N_5499,N_4514,N_3678);
or U5500 (N_5500,N_3619,N_1438);
or U5501 (N_5501,N_914,N_851);
nand U5502 (N_5502,N_1396,N_380);
or U5503 (N_5503,N_2078,N_1170);
nand U5504 (N_5504,N_2747,N_2780);
or U5505 (N_5505,N_2249,N_3111);
nor U5506 (N_5506,N_4009,N_3223);
nand U5507 (N_5507,N_1927,N_1464);
nor U5508 (N_5508,N_1189,N_557);
nand U5509 (N_5509,N_1786,N_1790);
and U5510 (N_5510,N_4591,N_4184);
nor U5511 (N_5511,N_1919,N_4145);
nor U5512 (N_5512,N_3866,N_2168);
or U5513 (N_5513,N_4406,N_4560);
or U5514 (N_5514,N_1213,N_2860);
and U5515 (N_5515,N_3529,N_1291);
or U5516 (N_5516,N_4230,N_3953);
nand U5517 (N_5517,N_26,N_2204);
nand U5518 (N_5518,N_1089,N_14);
nor U5519 (N_5519,N_62,N_2842);
or U5520 (N_5520,N_788,N_2478);
or U5521 (N_5521,N_435,N_4317);
nor U5522 (N_5522,N_3733,N_827);
nor U5523 (N_5523,N_1753,N_711);
nand U5524 (N_5524,N_1732,N_848);
and U5525 (N_5525,N_2644,N_1873);
nor U5526 (N_5526,N_2297,N_1895);
and U5527 (N_5527,N_1203,N_960);
nor U5528 (N_5528,N_1982,N_3823);
or U5529 (N_5529,N_4248,N_4105);
nor U5530 (N_5530,N_3595,N_2152);
or U5531 (N_5531,N_621,N_2085);
nand U5532 (N_5532,N_4132,N_799);
and U5533 (N_5533,N_4093,N_3179);
or U5534 (N_5534,N_4208,N_3754);
and U5535 (N_5535,N_712,N_1482);
and U5536 (N_5536,N_197,N_4253);
nand U5537 (N_5537,N_927,N_761);
nand U5538 (N_5538,N_2349,N_1634);
and U5539 (N_5539,N_56,N_2263);
or U5540 (N_5540,N_2757,N_1943);
or U5541 (N_5541,N_4312,N_3692);
and U5542 (N_5542,N_2183,N_1619);
nand U5543 (N_5543,N_4651,N_746);
or U5544 (N_5544,N_3267,N_3721);
or U5545 (N_5545,N_3478,N_3959);
nor U5546 (N_5546,N_2584,N_3523);
nor U5547 (N_5547,N_3056,N_4510);
nor U5548 (N_5548,N_641,N_1018);
and U5549 (N_5549,N_4983,N_4288);
nand U5550 (N_5550,N_1316,N_3080);
and U5551 (N_5551,N_2300,N_794);
nand U5552 (N_5552,N_432,N_4304);
and U5553 (N_5553,N_2294,N_4110);
or U5554 (N_5554,N_51,N_1239);
nor U5555 (N_5555,N_858,N_2039);
and U5556 (N_5556,N_4269,N_2541);
nor U5557 (N_5557,N_4201,N_4495);
or U5558 (N_5558,N_3893,N_1199);
nand U5559 (N_5559,N_3724,N_1391);
and U5560 (N_5560,N_2052,N_2131);
and U5561 (N_5561,N_1754,N_1268);
nand U5562 (N_5562,N_3613,N_2221);
and U5563 (N_5563,N_59,N_4958);
nand U5564 (N_5564,N_4682,N_570);
or U5565 (N_5565,N_1416,N_21);
nor U5566 (N_5566,N_148,N_1364);
nor U5567 (N_5567,N_3872,N_2121);
nor U5568 (N_5568,N_3112,N_707);
nand U5569 (N_5569,N_1477,N_4708);
nand U5570 (N_5570,N_4125,N_3568);
and U5571 (N_5571,N_1421,N_516);
nand U5572 (N_5572,N_4025,N_597);
nand U5573 (N_5573,N_1845,N_2847);
and U5574 (N_5574,N_302,N_1703);
nand U5575 (N_5575,N_2772,N_671);
nand U5576 (N_5576,N_3605,N_3026);
and U5577 (N_5577,N_3174,N_3755);
nor U5578 (N_5578,N_3577,N_4340);
nand U5579 (N_5579,N_4118,N_4381);
nand U5580 (N_5580,N_3301,N_319);
nand U5581 (N_5581,N_270,N_417);
nand U5582 (N_5582,N_482,N_1253);
or U5583 (N_5583,N_644,N_4703);
or U5584 (N_5584,N_4710,N_2009);
nor U5585 (N_5585,N_1842,N_1058);
nand U5586 (N_5586,N_2988,N_225);
or U5587 (N_5587,N_3282,N_3532);
and U5588 (N_5588,N_3288,N_539);
nor U5589 (N_5589,N_1318,N_2925);
and U5590 (N_5590,N_2360,N_1823);
and U5591 (N_5591,N_2084,N_2344);
and U5592 (N_5592,N_1847,N_4143);
nor U5593 (N_5593,N_74,N_3400);
nor U5594 (N_5594,N_3187,N_2651);
or U5595 (N_5595,N_1467,N_4771);
or U5596 (N_5596,N_1621,N_2303);
or U5597 (N_5597,N_4604,N_2658);
nor U5598 (N_5598,N_4470,N_385);
and U5599 (N_5599,N_2668,N_2566);
nand U5600 (N_5600,N_3229,N_41);
and U5601 (N_5601,N_1834,N_2195);
and U5602 (N_5602,N_3633,N_3127);
nor U5603 (N_5603,N_3055,N_4711);
and U5604 (N_5604,N_4263,N_2019);
nor U5605 (N_5605,N_3363,N_4407);
nor U5606 (N_5606,N_3586,N_2760);
and U5607 (N_5607,N_588,N_3071);
or U5608 (N_5608,N_487,N_206);
nand U5609 (N_5609,N_2347,N_280);
nor U5610 (N_5610,N_3434,N_2007);
nand U5611 (N_5611,N_2901,N_2592);
nor U5612 (N_5612,N_3729,N_3752);
nor U5613 (N_5613,N_4815,N_4945);
or U5614 (N_5614,N_2393,N_2301);
or U5615 (N_5615,N_4768,N_4610);
nor U5616 (N_5616,N_4366,N_1543);
or U5617 (N_5617,N_3199,N_1078);
nor U5618 (N_5618,N_3360,N_3367);
and U5619 (N_5619,N_1947,N_4557);
or U5620 (N_5620,N_1990,N_3017);
nand U5621 (N_5621,N_652,N_2631);
nor U5622 (N_5622,N_3058,N_4418);
nor U5623 (N_5623,N_962,N_4082);
or U5624 (N_5624,N_3562,N_1596);
nor U5625 (N_5625,N_1803,N_27);
and U5626 (N_5626,N_4504,N_4476);
nand U5627 (N_5627,N_4424,N_3287);
and U5628 (N_5628,N_1297,N_322);
nor U5629 (N_5629,N_662,N_1963);
or U5630 (N_5630,N_1244,N_2507);
nor U5631 (N_5631,N_1664,N_2715);
and U5632 (N_5632,N_2696,N_1459);
nand U5633 (N_5633,N_1131,N_227);
nand U5634 (N_5634,N_4798,N_2445);
and U5635 (N_5635,N_3517,N_976);
nor U5636 (N_5636,N_3131,N_770);
and U5637 (N_5637,N_2560,N_2211);
and U5638 (N_5638,N_667,N_1232);
nor U5639 (N_5639,N_3800,N_1439);
nand U5640 (N_5640,N_4886,N_3008);
nand U5641 (N_5641,N_963,N_2266);
nor U5642 (N_5642,N_2639,N_410);
and U5643 (N_5643,N_1305,N_2635);
and U5644 (N_5644,N_3682,N_129);
nand U5645 (N_5645,N_4292,N_442);
nor U5646 (N_5646,N_4123,N_3805);
or U5647 (N_5647,N_1307,N_4444);
or U5648 (N_5648,N_673,N_1812);
nor U5649 (N_5649,N_2649,N_1499);
nand U5650 (N_5650,N_4925,N_2753);
and U5651 (N_5651,N_2720,N_4006);
nand U5652 (N_5652,N_3970,N_1486);
nand U5653 (N_5653,N_3726,N_853);
nor U5654 (N_5654,N_409,N_2993);
nand U5655 (N_5655,N_3515,N_217);
nor U5656 (N_5656,N_768,N_4171);
or U5657 (N_5657,N_70,N_4298);
or U5658 (N_5658,N_3007,N_4562);
and U5659 (N_5659,N_2337,N_1108);
and U5660 (N_5660,N_4967,N_4337);
and U5661 (N_5661,N_1281,N_4196);
and U5662 (N_5662,N_675,N_4481);
and U5663 (N_5663,N_3745,N_3159);
and U5664 (N_5664,N_232,N_3025);
and U5665 (N_5665,N_1474,N_4209);
and U5666 (N_5666,N_978,N_360);
or U5667 (N_5667,N_3278,N_3565);
nor U5668 (N_5668,N_98,N_2104);
or U5669 (N_5669,N_3898,N_4030);
and U5670 (N_5670,N_2464,N_1079);
or U5671 (N_5671,N_2597,N_243);
nand U5672 (N_5672,N_413,N_1534);
nand U5673 (N_5673,N_4430,N_3302);
nand U5674 (N_5674,N_1451,N_1559);
nand U5675 (N_5675,N_3681,N_2048);
nor U5676 (N_5676,N_4204,N_4342);
nor U5677 (N_5677,N_2741,N_305);
or U5678 (N_5678,N_4816,N_3652);
nor U5679 (N_5679,N_3255,N_975);
or U5680 (N_5680,N_4870,N_1055);
or U5681 (N_5681,N_4305,N_3982);
nor U5682 (N_5682,N_672,N_174);
nand U5683 (N_5683,N_4267,N_3036);
nand U5684 (N_5684,N_4291,N_2967);
or U5685 (N_5685,N_1125,N_2994);
and U5686 (N_5686,N_134,N_2284);
or U5687 (N_5687,N_1273,N_3308);
nor U5688 (N_5688,N_1516,N_3372);
and U5689 (N_5689,N_1247,N_3731);
nand U5690 (N_5690,N_283,N_3956);
nor U5691 (N_5691,N_3329,N_1249);
nor U5692 (N_5692,N_4973,N_4830);
or U5693 (N_5693,N_1082,N_3589);
or U5694 (N_5694,N_4075,N_626);
nor U5695 (N_5695,N_193,N_1896);
nor U5696 (N_5696,N_281,N_3596);
and U5697 (N_5697,N_2174,N_2133);
nor U5698 (N_5698,N_3559,N_2702);
or U5699 (N_5699,N_2783,N_4791);
or U5700 (N_5700,N_3865,N_2343);
nor U5701 (N_5701,N_1617,N_2915);
or U5702 (N_5702,N_4446,N_968);
nor U5703 (N_5703,N_3986,N_2083);
or U5704 (N_5704,N_224,N_1723);
xnor U5705 (N_5705,N_3351,N_3622);
or U5706 (N_5706,N_1517,N_4468);
nand U5707 (N_5707,N_4237,N_1309);
xnor U5708 (N_5708,N_143,N_72);
and U5709 (N_5709,N_2293,N_1711);
nor U5710 (N_5710,N_2542,N_1114);
nand U5711 (N_5711,N_4845,N_2437);
and U5712 (N_5712,N_926,N_127);
or U5713 (N_5713,N_2207,N_3519);
nor U5714 (N_5714,N_4753,N_4654);
and U5715 (N_5715,N_1308,N_2352);
and U5716 (N_5716,N_4231,N_3798);
nand U5717 (N_5717,N_563,N_567);
and U5718 (N_5718,N_4992,N_1360);
nor U5719 (N_5719,N_3333,N_466);
nand U5720 (N_5720,N_2196,N_1914);
and U5721 (N_5721,N_3958,N_263);
or U5722 (N_5722,N_58,N_3581);
nand U5723 (N_5723,N_4415,N_378);
and U5724 (N_5724,N_4334,N_2033);
and U5725 (N_5725,N_3431,N_121);
and U5726 (N_5726,N_456,N_298);
or U5727 (N_5727,N_2540,N_1928);
nor U5728 (N_5728,N_2997,N_2457);
nand U5729 (N_5729,N_1905,N_3221);
or U5730 (N_5730,N_2336,N_2659);
nor U5731 (N_5731,N_3689,N_4372);
and U5732 (N_5732,N_3245,N_1068);
or U5733 (N_5733,N_293,N_4013);
nand U5734 (N_5734,N_1120,N_1174);
nor U5735 (N_5735,N_4543,N_2129);
nand U5736 (N_5736,N_3202,N_4919);
nor U5737 (N_5737,N_2689,N_866);
xnor U5738 (N_5738,N_1689,N_3498);
nand U5739 (N_5739,N_2939,N_4185);
or U5740 (N_5740,N_3759,N_3639);
nand U5741 (N_5741,N_3402,N_4524);
nor U5742 (N_5742,N_4148,N_649);
or U5743 (N_5743,N_3949,N_4061);
or U5744 (N_5744,N_1881,N_884);
or U5745 (N_5745,N_3894,N_2383);
nor U5746 (N_5746,N_276,N_1785);
nor U5747 (N_5747,N_3000,N_147);
and U5748 (N_5748,N_2632,N_1303);
and U5749 (N_5749,N_1906,N_1506);
and U5750 (N_5750,N_3041,N_3256);
nand U5751 (N_5751,N_4928,N_3829);
nor U5752 (N_5752,N_3957,N_3524);
nor U5753 (N_5753,N_2941,N_4290);
and U5754 (N_5754,N_91,N_323);
nor U5755 (N_5755,N_288,N_1702);
or U5756 (N_5756,N_2729,N_4540);
nand U5757 (N_5757,N_1128,N_2870);
and U5758 (N_5758,N_3920,N_880);
and U5759 (N_5759,N_1550,N_2814);
nor U5760 (N_5760,N_3099,N_4803);
nor U5761 (N_5761,N_3002,N_3048);
nand U5762 (N_5762,N_3611,N_512);
nand U5763 (N_5763,N_2508,N_4278);
nand U5764 (N_5764,N_4329,N_2710);
or U5765 (N_5765,N_3553,N_1134);
nor U5766 (N_5766,N_691,N_2013);
or U5767 (N_5767,N_3433,N_2694);
nor U5768 (N_5768,N_3757,N_1911);
nor U5769 (N_5769,N_2339,N_4101);
nand U5770 (N_5770,N_2832,N_813);
nand U5771 (N_5771,N_850,N_4717);
nor U5772 (N_5772,N_3188,N_4232);
and U5773 (N_5773,N_3863,N_3332);
nand U5774 (N_5774,N_4416,N_3996);
nor U5775 (N_5775,N_45,N_4605);
or U5776 (N_5776,N_4787,N_4198);
nor U5777 (N_5777,N_1237,N_1856);
or U5778 (N_5778,N_3323,N_4400);
and U5779 (N_5779,N_4015,N_4080);
and U5780 (N_5780,N_2459,N_3888);
nand U5781 (N_5781,N_2038,N_2292);
or U5782 (N_5782,N_251,N_4303);
nor U5783 (N_5783,N_3607,N_1001);
or U5784 (N_5784,N_3795,N_3504);
and U5785 (N_5785,N_1755,N_3250);
nand U5786 (N_5786,N_3882,N_4626);
nor U5787 (N_5787,N_1765,N_3535);
and U5788 (N_5788,N_3183,N_170);
or U5789 (N_5789,N_1978,N_4420);
and U5790 (N_5790,N_3011,N_1653);
or U5791 (N_5791,N_948,N_3673);
and U5792 (N_5792,N_3508,N_3926);
nor U5793 (N_5793,N_1626,N_1528);
and U5794 (N_5794,N_4770,N_2666);
nor U5795 (N_5795,N_782,N_3163);
nand U5796 (N_5796,N_3709,N_508);
nand U5797 (N_5797,N_979,N_860);
or U5798 (N_5798,N_3548,N_4155);
and U5799 (N_5799,N_71,N_890);
or U5800 (N_5800,N_3330,N_700);
nand U5801 (N_5801,N_569,N_3300);
nand U5802 (N_5802,N_4417,N_4197);
and U5803 (N_5803,N_1270,N_4741);
nor U5804 (N_5804,N_3868,N_3797);
or U5805 (N_5805,N_326,N_4790);
or U5806 (N_5806,N_3552,N_3076);
or U5807 (N_5807,N_1404,N_2074);
or U5808 (N_5808,N_816,N_3801);
nor U5809 (N_5809,N_708,N_4287);
and U5810 (N_5810,N_4138,N_1649);
and U5811 (N_5811,N_3625,N_394);
nand U5812 (N_5812,N_2692,N_2778);
or U5813 (N_5813,N_4327,N_4262);
nand U5814 (N_5814,N_1743,N_4373);
nand U5815 (N_5815,N_1699,N_1398);
and U5816 (N_5816,N_369,N_247);
nor U5817 (N_5817,N_798,N_196);
and U5818 (N_5818,N_3549,N_2227);
or U5819 (N_5819,N_3486,N_3732);
nor U5820 (N_5820,N_525,N_2557);
nor U5821 (N_5821,N_4102,N_2888);
and U5822 (N_5822,N_4663,N_430);
nand U5823 (N_5823,N_4520,N_2388);
nand U5824 (N_5824,N_2891,N_2469);
nand U5825 (N_5825,N_104,N_1340);
nand U5826 (N_5826,N_3331,N_4621);
or U5827 (N_5827,N_1047,N_4632);
nor U5828 (N_5828,N_3990,N_180);
nand U5829 (N_5829,N_4376,N_4341);
nor U5830 (N_5830,N_1400,N_871);
or U5831 (N_5831,N_4723,N_1354);
nor U5832 (N_5832,N_3901,N_3184);
and U5833 (N_5833,N_4665,N_1235);
and U5834 (N_5834,N_2709,N_3495);
nor U5835 (N_5835,N_209,N_3854);
nand U5836 (N_5836,N_2833,N_2960);
nand U5837 (N_5837,N_705,N_54);
nand U5838 (N_5838,N_1193,N_1087);
nor U5839 (N_5839,N_2272,N_4979);
nand U5840 (N_5840,N_1751,N_2516);
nand U5841 (N_5841,N_1301,N_4745);
and U5842 (N_5842,N_2328,N_183);
nor U5843 (N_5843,N_4989,N_2449);
or U5844 (N_5844,N_1814,N_2273);
and U5845 (N_5845,N_3479,N_820);
nand U5846 (N_5846,N_748,N_423);
or U5847 (N_5847,N_2217,N_4076);
nor U5848 (N_5848,N_578,N_3246);
nor U5849 (N_5849,N_1063,N_3162);
xor U5850 (N_5850,N_2918,N_3147);
and U5851 (N_5851,N_337,N_3802);
nand U5852 (N_5852,N_653,N_3925);
nor U5853 (N_5853,N_3435,N_2598);
nor U5854 (N_5854,N_3831,N_4482);
nor U5855 (N_5855,N_2110,N_450);
nor U5856 (N_5856,N_1844,N_4021);
nand U5857 (N_5857,N_199,N_4280);
nor U5858 (N_5858,N_2711,N_29);
or U5859 (N_5859,N_2374,N_3031);
nor U5860 (N_5860,N_1077,N_1358);
nand U5861 (N_5861,N_2250,N_253);
or U5862 (N_5862,N_1735,N_4182);
or U5863 (N_5863,N_4390,N_2951);
nor U5864 (N_5864,N_2981,N_1624);
nand U5865 (N_5865,N_2010,N_4403);
or U5866 (N_5866,N_2421,N_3878);
and U5867 (N_5867,N_4062,N_1414);
nand U5868 (N_5868,N_3998,N_4106);
nor U5869 (N_5869,N_4289,N_1402);
nand U5870 (N_5870,N_4685,N_3046);
nor U5871 (N_5871,N_3276,N_4720);
nand U5872 (N_5872,N_2622,N_1819);
and U5873 (N_5873,N_1088,N_287);
nor U5874 (N_5874,N_4345,N_166);
or U5875 (N_5875,N_184,N_2474);
or U5876 (N_5876,N_4084,N_1551);
and U5877 (N_5877,N_4914,N_307);
and U5878 (N_5878,N_185,N_639);
or U5879 (N_5879,N_3620,N_3094);
and U5880 (N_5880,N_363,N_3137);
or U5881 (N_5881,N_784,N_3362);
and U5882 (N_5882,N_3710,N_240);
nor U5883 (N_5883,N_2391,N_4904);
nand U5884 (N_5884,N_1867,N_4215);
and U5885 (N_5885,N_1539,N_4911);
and U5886 (N_5886,N_1295,N_3962);
or U5887 (N_5887,N_384,N_4579);
or U5888 (N_5888,N_970,N_494);
or U5889 (N_5889,N_3104,N_82);
nor U5890 (N_5890,N_2762,N_1644);
or U5891 (N_5891,N_2633,N_4250);
or U5892 (N_5892,N_2563,N_1592);
nor U5893 (N_5893,N_208,N_78);
or U5894 (N_5894,N_1080,N_1957);
and U5895 (N_5895,N_3546,N_4923);
or U5896 (N_5896,N_4764,N_4731);
nand U5897 (N_5897,N_2577,N_4936);
nor U5898 (N_5898,N_480,N_2203);
nand U5899 (N_5899,N_4214,N_1040);
nand U5900 (N_5900,N_3427,N_2976);
and U5901 (N_5901,N_2586,N_331);
or U5902 (N_5902,N_1778,N_1849);
or U5903 (N_5903,N_2933,N_2880);
and U5904 (N_5904,N_10,N_4328);
nor U5905 (N_5905,N_1938,N_28);
and U5906 (N_5906,N_1384,N_4737);
or U5907 (N_5907,N_1260,N_3192);
and U5908 (N_5908,N_4634,N_1110);
nor U5909 (N_5909,N_685,N_2742);
nor U5910 (N_5910,N_1908,N_709);
and U5911 (N_5911,N_1554,N_407);
nor U5912 (N_5912,N_532,N_3792);
nand U5913 (N_5913,N_321,N_114);
nor U5914 (N_5914,N_4678,N_4503);
nor U5915 (N_5915,N_4884,N_661);
nor U5916 (N_5916,N_2205,N_4357);
nor U5917 (N_5917,N_3943,N_2216);
and U5918 (N_5918,N_3921,N_4463);
nor U5919 (N_5919,N_3660,N_888);
nand U5920 (N_5920,N_839,N_4611);
nand U5921 (N_5921,N_3825,N_4448);
nor U5922 (N_5922,N_3210,N_2409);
nand U5923 (N_5923,N_1821,N_4777);
and U5924 (N_5924,N_3406,N_533);
nor U5925 (N_5925,N_1279,N_2756);
nor U5926 (N_5926,N_2073,N_1215);
and U5927 (N_5927,N_1887,N_1194);
nor U5928 (N_5928,N_2489,N_887);
or U5929 (N_5929,N_623,N_3582);
nand U5930 (N_5930,N_4526,N_3062);
nor U5931 (N_5931,N_4553,N_4484);
or U5932 (N_5932,N_3204,N_2351);
and U5933 (N_5933,N_4023,N_3350);
and U5934 (N_5934,N_1827,N_4802);
or U5935 (N_5935,N_4445,N_212);
and U5936 (N_5936,N_1372,N_4893);
and U5937 (N_5937,N_16,N_3177);
nand U5938 (N_5938,N_3024,N_2150);
nor U5939 (N_5939,N_4736,N_4169);
or U5940 (N_5940,N_3185,N_4754);
and U5941 (N_5941,N_4077,N_4918);
nand U5942 (N_5942,N_1240,N_989);
nand U5943 (N_5943,N_2984,N_766);
and U5944 (N_5944,N_808,N_1604);
or U5945 (N_5945,N_2974,N_4641);
or U5946 (N_5946,N_405,N_2704);
nand U5947 (N_5947,N_60,N_496);
nor U5948 (N_5948,N_3004,N_1326);
or U5949 (N_5949,N_2394,N_2943);
or U5950 (N_5950,N_2911,N_3314);
and U5951 (N_5951,N_628,N_2185);
and U5952 (N_5952,N_1092,N_1556);
and U5953 (N_5953,N_3258,N_1479);
and U5954 (N_5954,N_1132,N_1706);
nand U5955 (N_5955,N_4260,N_2122);
and U5956 (N_5956,N_426,N_4859);
and U5957 (N_5957,N_687,N_600);
and U5958 (N_5958,N_3610,N_395);
nand U5959 (N_5959,N_4206,N_1460);
nor U5960 (N_5960,N_4976,N_4038);
nor U5961 (N_5961,N_2268,N_257);
xnor U5962 (N_5962,N_1415,N_4725);
nor U5963 (N_5963,N_2120,N_3410);
nor U5964 (N_5964,N_938,N_3086);
and U5965 (N_5965,N_2188,N_4957);
and U5966 (N_5966,N_2908,N_2189);
nand U5967 (N_5967,N_3460,N_2886);
and U5968 (N_5968,N_1010,N_1424);
or U5969 (N_5969,N_4242,N_1566);
nor U5970 (N_5970,N_4901,N_3780);
or U5971 (N_5971,N_2555,N_3656);
nand U5972 (N_5972,N_1629,N_2190);
or U5973 (N_5973,N_2096,N_4285);
nor U5974 (N_5974,N_935,N_2801);
nor U5975 (N_5975,N_3667,N_4697);
nor U5976 (N_5976,N_3015,N_1628);
or U5977 (N_5977,N_2456,N_2325);
nand U5978 (N_5978,N_697,N_2385);
nand U5979 (N_5979,N_2677,N_4396);
and U5980 (N_5980,N_2667,N_2413);
nand U5981 (N_5981,N_2496,N_4414);
nor U5982 (N_5982,N_1137,N_2119);
nor U5983 (N_5983,N_399,N_3826);
or U5984 (N_5984,N_317,N_1401);
and U5985 (N_5985,N_942,N_1019);
and U5986 (N_5986,N_1262,N_3438);
nor U5987 (N_5987,N_1671,N_1878);
or U5988 (N_5988,N_642,N_1348);
or U5989 (N_5989,N_1290,N_2454);
and U5990 (N_5990,N_3935,N_878);
nor U5991 (N_5991,N_2433,N_210);
or U5992 (N_5992,N_717,N_4554);
and U5993 (N_5993,N_2593,N_3522);
nand U5994 (N_5994,N_3631,N_4877);
nand U5995 (N_5995,N_3040,N_3325);
nand U5996 (N_5996,N_3815,N_4733);
nand U5997 (N_5997,N_857,N_904);
nor U5998 (N_5998,N_2815,N_1581);
nor U5999 (N_5999,N_4522,N_4411);
nor U6000 (N_6000,N_1586,N_393);
or U6001 (N_6001,N_358,N_4067);
nor U6002 (N_6002,N_603,N_2426);
nor U6003 (N_6003,N_1127,N_3606);
nand U6004 (N_6004,N_754,N_2558);
nand U6005 (N_6005,N_4640,N_4565);
and U6006 (N_6006,N_1944,N_234);
and U6007 (N_6007,N_4496,N_3543);
or U6008 (N_6008,N_2947,N_1271);
nor U6009 (N_6009,N_3450,N_1342);
or U6010 (N_6010,N_3997,N_3874);
nor U6011 (N_6011,N_4619,N_2118);
nand U6012 (N_6012,N_1802,N_2648);
and U6013 (N_6013,N_943,N_2307);
or U6014 (N_6014,N_4259,N_68);
and U6015 (N_6015,N_4698,N_734);
or U6016 (N_6016,N_1781,N_2851);
and U6017 (N_6017,N_2348,N_3640);
nand U6018 (N_6018,N_2199,N_213);
nand U6019 (N_6019,N_2830,N_2522);
and U6020 (N_6020,N_1882,N_3381);
or U6021 (N_6021,N_419,N_2897);
and U6022 (N_6022,N_1242,N_837);
nand U6023 (N_6023,N_4228,N_1256);
or U6024 (N_6024,N_3544,N_4673);
and U6025 (N_6025,N_472,N_1553);
nor U6026 (N_6026,N_215,N_3630);
nor U6027 (N_6027,N_396,N_980);
nor U6028 (N_6028,N_1636,N_11);
or U6029 (N_6029,N_985,N_2675);
and U6030 (N_6030,N_2399,N_2751);
nor U6031 (N_6031,N_2305,N_3955);
nand U6032 (N_6032,N_2165,N_3813);
nor U6033 (N_6033,N_3771,N_230);
nor U6034 (N_6034,N_2125,N_1563);
nand U6035 (N_6035,N_4664,N_4019);
nand U6036 (N_6036,N_618,N_2218);
and U6037 (N_6037,N_2810,N_1016);
nor U6038 (N_6038,N_2062,N_4137);
nand U6039 (N_6039,N_805,N_2092);
nand U6040 (N_6040,N_3875,N_3209);
or U6041 (N_6041,N_2718,N_3161);
or U6042 (N_6042,N_1052,N_351);
or U6043 (N_6043,N_2549,N_3489);
nand U6044 (N_6044,N_1584,N_1141);
or U6045 (N_6045,N_1678,N_1061);
or U6046 (N_6046,N_1284,N_810);
and U6047 (N_6047,N_2561,N_1427);
or U6048 (N_6048,N_1522,N_1722);
and U6049 (N_6049,N_2972,N_2945);
and U6050 (N_6050,N_847,N_191);
nand U6051 (N_6051,N_2450,N_2708);
nor U6052 (N_6052,N_1949,N_2302);
nor U6053 (N_6053,N_1130,N_2545);
and U6054 (N_6054,N_1869,N_289);
nand U6055 (N_6055,N_3528,N_3791);
or U6056 (N_6056,N_1763,N_542);
nand U6057 (N_6057,N_695,N_50);
nor U6058 (N_6058,N_1374,N_1368);
or U6059 (N_6059,N_1029,N_3674);
and U6060 (N_6060,N_325,N_743);
nor U6061 (N_6061,N_519,N_1265);
nand U6062 (N_6062,N_589,N_2916);
nand U6063 (N_6063,N_1136,N_284);
nor U6064 (N_6064,N_371,N_3472);
or U6065 (N_6065,N_891,N_159);
or U6066 (N_6066,N_1888,N_4551);
and U6067 (N_6067,N_4941,N_120);
or U6068 (N_6068,N_2502,N_3014);
nand U6069 (N_6069,N_3294,N_4177);
nand U6070 (N_6070,N_952,N_3983);
nor U6071 (N_6071,N_4377,N_993);
or U6072 (N_6072,N_3765,N_4960);
nor U6073 (N_6073,N_2684,N_2596);
or U6074 (N_6074,N_4121,N_2670);
nor U6075 (N_6075,N_486,N_297);
and U6076 (N_6076,N_2242,N_524);
or U6077 (N_6077,N_4784,N_1536);
and U6078 (N_6078,N_4183,N_3158);
nand U6079 (N_6079,N_4920,N_3178);
or U6080 (N_6080,N_1692,N_2788);
nand U6081 (N_6081,N_4261,N_3775);
and U6082 (N_6082,N_3819,N_425);
nor U6083 (N_6083,N_1991,N_4103);
nand U6084 (N_6084,N_1717,N_3452);
nor U6085 (N_6085,N_2812,N_4538);
and U6086 (N_6086,N_1186,N_1109);
or U6087 (N_6087,N_1929,N_2045);
or U6088 (N_6088,N_1916,N_3711);
nor U6089 (N_6089,N_4903,N_1996);
and U6090 (N_6090,N_4743,N_3077);
nor U6091 (N_6091,N_3827,N_3538);
and U6092 (N_6092,N_4391,N_660);
nand U6093 (N_6093,N_350,N_2163);
or U6094 (N_6094,N_3359,N_214);
nand U6095 (N_6095,N_3601,N_1567);
nor U6096 (N_6096,N_24,N_3474);
nor U6097 (N_6097,N_1876,N_3264);
nor U6098 (N_6098,N_2761,N_2167);
and U6099 (N_6099,N_4789,N_2864);
and U6100 (N_6100,N_422,N_2412);
nand U6101 (N_6101,N_2697,N_155);
and U6102 (N_6102,N_2027,N_2161);
nand U6103 (N_6103,N_370,N_1734);
nand U6104 (N_6104,N_4807,N_2481);
or U6105 (N_6105,N_1369,N_2378);
or U6106 (N_6106,N_1012,N_3704);
nand U6107 (N_6107,N_2999,N_3353);
and U6108 (N_6108,N_1113,N_877);
nand U6109 (N_6109,N_4756,N_1417);
and U6110 (N_6110,N_1684,N_1618);
and U6111 (N_6111,N_3290,N_2194);
or U6112 (N_6112,N_4744,N_4405);
nor U6113 (N_6113,N_676,N_682);
nor U6114 (N_6114,N_3475,N_981);
nand U6115 (N_6115,N_4046,N_1832);
nand U6116 (N_6116,N_2482,N_1762);
nor U6117 (N_6117,N_3905,N_476);
nand U6118 (N_6118,N_1933,N_4175);
nand U6119 (N_6119,N_2883,N_2289);
nor U6120 (N_6120,N_2717,N_3445);
nor U6121 (N_6121,N_2026,N_354);
and U6122 (N_6122,N_1355,N_1719);
nand U6123 (N_6123,N_4436,N_2905);
nor U6124 (N_6124,N_666,N_1962);
and U6125 (N_6125,N_1985,N_2369);
and U6126 (N_6126,N_2261,N_4505);
nand U6127 (N_6127,N_2455,N_2808);
or U6128 (N_6128,N_1361,N_3233);
or U6129 (N_6129,N_269,N_2240);
and U6130 (N_6130,N_3037,N_2323);
nor U6131 (N_6131,N_4378,N_4746);
or U6132 (N_6132,N_4191,N_2826);
nand U6133 (N_6133,N_925,N_4100);
nor U6134 (N_6134,N_4309,N_3254);
nor U6135 (N_6135,N_1771,N_19);
nor U6136 (N_6136,N_1225,N_1992);
and U6137 (N_6137,N_491,N_4686);
nor U6138 (N_6138,N_3571,N_3087);
and U6139 (N_6139,N_2364,N_4949);
nand U6140 (N_6140,N_1571,N_3636);
nand U6141 (N_6141,N_83,N_4385);
nor U6142 (N_6142,N_4475,N_3337);
nand U6143 (N_6143,N_670,N_4506);
or U6144 (N_6144,N_3770,N_727);
nand U6145 (N_6145,N_2254,N_824);
and U6146 (N_6146,N_1409,N_2148);
and U6147 (N_6147,N_4494,N_3284);
nor U6148 (N_6148,N_1643,N_2881);
or U6149 (N_6149,N_4339,N_1389);
nor U6150 (N_6150,N_882,N_3999);
nand U6151 (N_6151,N_1336,N_3934);
or U6152 (N_6152,N_3702,N_2017);
and U6153 (N_6153,N_4568,N_2462);
or U6154 (N_6154,N_2683,N_1363);
nor U6155 (N_6155,N_1533,N_561);
or U6156 (N_6156,N_1810,N_1004);
or U6157 (N_6157,N_404,N_3655);
nor U6158 (N_6158,N_4968,N_2173);
nand U6159 (N_6159,N_3016,N_3767);
and U6160 (N_6160,N_4590,N_1696);
and U6161 (N_6161,N_4765,N_1840);
and U6162 (N_6162,N_1954,N_2990);
or U6163 (N_6163,N_1587,N_4443);
or U6164 (N_6164,N_4868,N_1642);
or U6165 (N_6165,N_3279,N_4064);
nor U6166 (N_6166,N_732,N_4834);
and U6167 (N_6167,N_1250,N_617);
nand U6168 (N_6168,N_4456,N_1335);
or U6169 (N_6169,N_773,N_789);
nand U6170 (N_6170,N_893,N_3786);
nor U6171 (N_6171,N_493,N_4513);
or U6172 (N_6172,N_2485,N_3456);
nand U6173 (N_6173,N_2362,N_2271);
and U6174 (N_6174,N_1507,N_4612);
nand U6175 (N_6175,N_4946,N_25);
nand U6176 (N_6176,N_1007,N_2843);
nor U6177 (N_6177,N_2059,N_1960);
nor U6178 (N_6178,N_1351,N_1731);
or U6179 (N_6179,N_2095,N_2051);
nand U6180 (N_6180,N_3861,N_3635);
and U6181 (N_6181,N_1809,N_2920);
xnor U6182 (N_6182,N_2134,N_2137);
nor U6183 (N_6183,N_3317,N_1519);
nand U6184 (N_6184,N_4594,N_859);
or U6185 (N_6185,N_4179,N_2620);
and U6186 (N_6186,N_4297,N_2749);
and U6187 (N_6187,N_594,N_4249);
and U6188 (N_6188,N_2213,N_3768);
nand U6189 (N_6189,N_4029,N_1292);
or U6190 (N_6190,N_3150,N_3155);
nor U6191 (N_6191,N_1429,N_4170);
nor U6192 (N_6192,N_3992,N_2515);
or U6193 (N_6193,N_4805,N_1498);
nand U6194 (N_6194,N_1164,N_3539);
and U6195 (N_6195,N_2890,N_2665);
and U6196 (N_6196,N_4033,N_4371);
and U6197 (N_6197,N_246,N_1156);
and U6198 (N_6198,N_3599,N_1044);
or U6199 (N_6199,N_4666,N_1119);
nor U6200 (N_6200,N_2396,N_2224);
nand U6201 (N_6201,N_3892,N_131);
or U6202 (N_6202,N_4959,N_1165);
or U6203 (N_6203,N_753,N_2964);
or U6204 (N_6204,N_4150,N_4240);
nand U6205 (N_6205,N_386,N_3885);
nand U6206 (N_6206,N_932,N_1846);
or U6207 (N_6207,N_1635,N_844);
and U6208 (N_6208,N_4533,N_4818);
and U6209 (N_6209,N_271,N_4861);
nor U6210 (N_6210,N_4119,N_3789);
and U6211 (N_6211,N_1485,N_3248);
and U6212 (N_6212,N_3393,N_4199);
or U6213 (N_6213,N_4202,N_1705);
or U6214 (N_6214,N_3649,N_1848);
and U6215 (N_6215,N_1245,N_1321);
nand U6216 (N_6216,N_275,N_4322);
or U6217 (N_6217,N_219,N_3143);
nor U6218 (N_6218,N_1241,N_1805);
nand U6219 (N_6219,N_373,N_802);
and U6220 (N_6220,N_1022,N_874);
nand U6221 (N_6221,N_2111,N_2532);
and U6222 (N_6222,N_412,N_4951);
or U6223 (N_6223,N_4273,N_1893);
nor U6224 (N_6224,N_119,N_2695);
or U6225 (N_6225,N_1728,N_769);
and U6226 (N_6226,N_1121,N_2156);
and U6227 (N_6227,N_668,N_2624);
or U6228 (N_6228,N_2075,N_2243);
and U6229 (N_6229,N_2599,N_2501);
or U6230 (N_6230,N_4809,N_1852);
or U6231 (N_6231,N_2719,N_3477);
and U6232 (N_6232,N_392,N_377);
nor U6233 (N_6233,N_2661,N_223);
xor U6234 (N_6234,N_1670,N_4934);
nor U6235 (N_6235,N_2700,N_3275);
nor U6236 (N_6236,N_1538,N_534);
and U6237 (N_6237,N_1056,N_4346);
and U6238 (N_6238,N_2604,N_4268);
nand U6239 (N_6239,N_2313,N_455);
or U6240 (N_6240,N_4111,N_650);
nand U6241 (N_6241,N_619,N_4690);
nor U6242 (N_6242,N_2311,N_1747);
or U6243 (N_6243,N_4487,N_3914);
or U6244 (N_6244,N_1357,N_3203);
and U6245 (N_6245,N_4556,N_3214);
or U6246 (N_6246,N_501,N_1616);
or U6247 (N_6247,N_2444,N_2170);
or U6248 (N_6248,N_683,N_1730);
nor U6249 (N_6249,N_2408,N_3382);
nor U6250 (N_6250,N_2949,N_1081);
nor U6251 (N_6251,N_2280,N_1580);
nor U6252 (N_6252,N_461,N_1813);
nor U6253 (N_6253,N_2298,N_4058);
and U6254 (N_6254,N_1220,N_3432);
nand U6255 (N_6255,N_4721,N_2424);
nor U6256 (N_6256,N_1122,N_4608);
or U6257 (N_6257,N_3521,N_939);
and U6258 (N_6258,N_4172,N_656);
and U6259 (N_6259,N_2787,N_752);
nor U6260 (N_6260,N_3583,N_2962);
nor U6261 (N_6261,N_2556,N_122);
nor U6262 (N_6262,N_4555,N_3944);
and U6263 (N_6263,N_2825,N_900);
and U6264 (N_6264,N_3366,N_1687);
or U6265 (N_6265,N_2127,N_1039);
and U6266 (N_6266,N_286,N_2707);
nor U6267 (N_6267,N_1890,N_4073);
or U6268 (N_6268,N_2014,N_822);
nand U6269 (N_6269,N_1286,N_3822);
and U6270 (N_6270,N_1535,N_3590);
and U6271 (N_6271,N_2495,N_374);
and U6272 (N_6272,N_2252,N_2514);
nand U6273 (N_6273,N_2296,N_1935);
nand U6274 (N_6274,N_3343,N_2077);
nand U6275 (N_6275,N_2237,N_2980);
nand U6276 (N_6276,N_2565,N_1320);
nand U6277 (N_6277,N_1676,N_2570);
or U6278 (N_6278,N_4236,N_1936);
nand U6279 (N_6279,N_1413,N_353);
nand U6280 (N_6280,N_4203,N_4509);
nand U6281 (N_6281,N_3483,N_1024);
and U6282 (N_6282,N_2287,N_2553);
nand U6283 (N_6283,N_2796,N_4001);
nand U6284 (N_6284,N_3271,N_4398);
or U6285 (N_6285,N_4166,N_1521);
or U6286 (N_6286,N_1677,N_2248);
or U6287 (N_6287,N_3458,N_1383);
nand U6288 (N_6288,N_2685,N_2342);
or U6289 (N_6289,N_3871,N_4016);
nand U6290 (N_6290,N_2479,N_728);
or U6291 (N_6291,N_1623,N_2146);
and U6292 (N_6292,N_254,N_1531);
or U6293 (N_6293,N_3853,N_4655);
and U6294 (N_6294,N_1737,N_3810);
or U6295 (N_6295,N_3744,N_3180);
and U6296 (N_6296,N_3449,N_783);
nor U6297 (N_6297,N_1573,N_2878);
and U6298 (N_6298,N_2079,N_1710);
nand U6299 (N_6299,N_3414,N_2806);
nand U6300 (N_6300,N_2022,N_2061);
nand U6301 (N_6301,N_2863,N_3422);
nor U6302 (N_6302,N_172,N_3283);
or U6303 (N_6303,N_2740,N_3219);
nor U6304 (N_6304,N_2087,N_1115);
or U6305 (N_6305,N_189,N_2959);
and U6306 (N_6306,N_2641,N_872);
nor U6307 (N_6307,N_1904,N_1331);
nand U6308 (N_6308,N_2484,N_4956);
and U6309 (N_6309,N_4395,N_3608);
nand U6310 (N_6310,N_3641,N_2679);
xnor U6311 (N_6311,N_2299,N_4026);
and U6312 (N_6312,N_2576,N_1162);
or U6313 (N_6313,N_1248,N_2441);
and U6314 (N_6314,N_1313,N_3784);
and U6315 (N_6315,N_1230,N_739);
nor U6316 (N_6316,N_2682,N_1112);
nand U6317 (N_6317,N_4778,N_1599);
nor U6318 (N_6318,N_3208,N_3200);
nor U6319 (N_6319,N_2279,N_3688);
and U6320 (N_6320,N_1184,N_314);
nand U6321 (N_6321,N_3743,N_4567);
nand U6322 (N_6322,N_640,N_457);
and U6323 (N_6323,N_97,N_4217);
nor U6324 (N_6324,N_4728,N_1449);
and U6325 (N_6325,N_1837,N_522);
nand U6326 (N_6326,N_346,N_4964);
or U6327 (N_6327,N_1959,N_1903);
or U6328 (N_6328,N_101,N_3937);
nand U6329 (N_6329,N_4800,N_2909);
or U6330 (N_6330,N_2377,N_4646);
or U6331 (N_6331,N_4159,N_572);
and U6332 (N_6332,N_2470,N_1341);
nand U6333 (N_6333,N_2259,N_381);
nor U6334 (N_6334,N_1782,N_3573);
nor U6335 (N_6335,N_2546,N_1447);
and U6336 (N_6336,N_40,N_4473);
nand U6337 (N_6337,N_2650,N_4596);
nand U6338 (N_6338,N_1073,N_1423);
nand U6339 (N_6339,N_4040,N_4219);
nor U6340 (N_6340,N_503,N_797);
or U6341 (N_6341,N_3657,N_928);
nor U6342 (N_6342,N_2436,N_1296);
and U6343 (N_6343,N_1979,N_499);
and U6344 (N_6344,N_2178,N_304);
or U6345 (N_6345,N_1898,N_917);
or U6346 (N_6346,N_2056,N_2662);
nand U6347 (N_6347,N_4549,N_502);
nand U6348 (N_6348,N_198,N_1527);
and U6349 (N_6349,N_1154,N_1972);
or U6350 (N_6350,N_4041,N_3975);
nor U6351 (N_6351,N_356,N_1555);
or U6352 (N_6352,N_3216,N_613);
or U6353 (N_6353,N_4151,N_612);
or U6354 (N_6354,N_3671,N_344);
nand U6355 (N_6355,N_3628,N_1168);
or U6356 (N_6356,N_1026,N_4825);
nor U6357 (N_6357,N_2407,N_4413);
nand U6358 (N_6358,N_2099,N_2567);
nand U6359 (N_6359,N_4319,N_902);
or U6360 (N_6360,N_4128,N_3235);
and U6361 (N_6361,N_2985,N_1645);
and U6362 (N_6362,N_2246,N_2265);
or U6363 (N_6363,N_3646,N_1661);
nand U6364 (N_6364,N_4162,N_3140);
nand U6365 (N_6365,N_1422,N_2805);
nor U6366 (N_6366,N_1894,N_2777);
nor U6367 (N_6367,N_4680,N_1440);
nand U6368 (N_6368,N_1169,N_3915);
nor U6369 (N_6369,N_818,N_1841);
or U6370 (N_6370,N_2848,N_1668);
and U6371 (N_6371,N_3190,N_449);
nor U6372 (N_6372,N_3556,N_562);
nand U6373 (N_6373,N_911,N_1796);
nand U6374 (N_6374,N_4332,N_4347);
nand U6375 (N_6375,N_2745,N_3971);
nand U6376 (N_6376,N_2691,N_315);
or U6377 (N_6377,N_4122,N_1542);
and U6378 (N_6378,N_4063,N_4349);
or U6379 (N_6379,N_3567,N_3439);
and U6380 (N_6380,N_2853,N_2023);
nor U6381 (N_6381,N_3751,N_4726);
and U6382 (N_6382,N_4732,N_2887);
and U6383 (N_6383,N_4835,N_1798);
nand U6384 (N_6384,N_1967,N_764);
or U6385 (N_6385,N_2035,N_1124);
or U6386 (N_6386,N_464,N_2844);
and U6387 (N_6387,N_3891,N_3651);
and U6388 (N_6388,N_3364,N_1872);
and U6389 (N_6389,N_2850,N_4382);
or U6390 (N_6390,N_1084,N_4338);
nor U6391 (N_6391,N_1501,N_2363);
or U6392 (N_6392,N_3170,N_12);
and U6393 (N_6393,N_4364,N_1251);
nor U6394 (N_6394,N_3840,N_840);
nor U6395 (N_6395,N_1690,N_2430);
nor U6396 (N_6396,N_2402,N_630);
and U6397 (N_6397,N_3084,N_301);
nor U6398 (N_6398,N_2002,N_2524);
nor U6399 (N_6399,N_4144,N_4879);
nand U6400 (N_6400,N_3850,N_689);
nor U6401 (N_6401,N_2770,N_2136);
nor U6402 (N_6402,N_772,N_4813);
or U6403 (N_6403,N_4498,N_115);
nand U6404 (N_6404,N_2431,N_3769);
or U6405 (N_6405,N_2603,N_1294);
nor U6406 (N_6406,N_2214,N_445);
nor U6407 (N_6407,N_1216,N_3121);
nor U6408 (N_6408,N_165,N_4489);
and U6409 (N_6409,N_2236,N_4653);
or U6410 (N_6410,N_4027,N_3830);
nand U6411 (N_6411,N_4439,N_1207);
and U6412 (N_6412,N_1577,N_4423);
or U6413 (N_6413,N_173,N_1074);
xor U6414 (N_6414,N_194,N_4981);
nor U6415 (N_6415,N_4944,N_4856);
or U6416 (N_6416,N_4615,N_2235);
and U6417 (N_6417,N_2899,N_2876);
nand U6418 (N_6418,N_2316,N_3038);
or U6419 (N_6419,N_2818,N_2859);
nor U6420 (N_6420,N_1151,N_2535);
or U6421 (N_6421,N_609,N_1987);
nand U6422 (N_6422,N_4994,N_4447);
nand U6423 (N_6423,N_4480,N_554);
and U6424 (N_6424,N_3518,N_972);
or U6425 (N_6425,N_3405,N_66);
or U6426 (N_6426,N_4427,N_2583);
nand U6427 (N_6427,N_774,N_3675);
and U6428 (N_6428,N_1930,N_886);
or U6429 (N_6429,N_3927,N_3096);
or U6430 (N_6430,N_1444,N_3948);
nand U6431 (N_6431,N_1811,N_955);
nor U6432 (N_6432,N_3152,N_910);
and U6433 (N_6433,N_1172,N_1036);
nor U6434 (N_6434,N_75,N_167);
nor U6435 (N_6435,N_1900,N_3503);
nor U6436 (N_6436,N_1277,N_4659);
nand U6437 (N_6437,N_328,N_1701);
nand U6438 (N_6438,N_2012,N_4133);
nand U6439 (N_6439,N_1679,N_4301);
or U6440 (N_6440,N_1394,N_2406);
nor U6441 (N_6441,N_1441,N_216);
nand U6442 (N_6442,N_3386,N_2429);
nor U6443 (N_6443,N_1148,N_3021);
or U6444 (N_6444,N_3005,N_3251);
nor U6445 (N_6445,N_4315,N_3712);
or U6446 (N_6446,N_1157,N_2286);
and U6447 (N_6447,N_3341,N_3697);
or U6448 (N_6448,N_3313,N_103);
nand U6449 (N_6449,N_3441,N_4097);
nor U6450 (N_6450,N_1816,N_4847);
nor U6451 (N_6451,N_4452,N_4222);
or U6452 (N_6452,N_3818,N_526);
nand U6453 (N_6453,N_4714,N_3032);
and U6454 (N_6454,N_3368,N_2467);
nor U6455 (N_6455,N_1140,N_2676);
and U6456 (N_6456,N_2011,N_4518);
nand U6457 (N_6457,N_2693,N_2628);
or U6458 (N_6458,N_80,N_4896);
nor U6459 (N_6459,N_4306,N_4912);
or U6460 (N_6460,N_4264,N_1041);
nor U6461 (N_6461,N_140,N_4576);
and U6462 (N_6462,N_4669,N_3484);
and U6463 (N_6463,N_20,N_4142);
nor U6464 (N_6464,N_710,N_2955);
nor U6465 (N_6465,N_3172,N_3257);
and U6466 (N_6466,N_1945,N_2256);
or U6467 (N_6467,N_2232,N_4793);
or U6468 (N_6468,N_3857,N_1450);
or U6469 (N_6469,N_46,N_4464);
and U6470 (N_6470,N_2617,N_3109);
nand U6471 (N_6471,N_336,N_1999);
and U6472 (N_6472,N_1276,N_1574);
or U6473 (N_6473,N_3739,N_365);
and U6474 (N_6474,N_2497,N_636);
and U6475 (N_6475,N_3860,N_3902);
nand U6476 (N_6476,N_2748,N_448);
or U6477 (N_6477,N_188,N_3459);
xor U6478 (N_6478,N_3194,N_2513);
nand U6479 (N_6479,N_4844,N_3130);
or U6480 (N_6480,N_1343,N_2003);
nand U6481 (N_6481,N_949,N_2792);
and U6482 (N_6482,N_2452,N_473);
nand U6483 (N_6483,N_22,N_831);
nand U6484 (N_6484,N_2439,N_1362);
and U6485 (N_6485,N_842,N_4950);
and U6486 (N_6486,N_2171,N_4429);
and U6487 (N_6487,N_2539,N_441);
xnor U6488 (N_6488,N_2795,N_3621);
or U6489 (N_6489,N_367,N_4521);
and U6490 (N_6490,N_3525,N_4235);
nor U6491 (N_6491,N_3115,N_2952);
nor U6492 (N_6492,N_507,N_1883);
nor U6493 (N_6493,N_2589,N_795);
or U6494 (N_6494,N_2361,N_1375);
nand U6495 (N_6495,N_4477,N_3560);
and U6496 (N_6496,N_3876,N_2276);
nor U6497 (N_6497,N_2979,N_150);
nor U6498 (N_6498,N_478,N_2440);
and U6499 (N_6499,N_1770,N_2660);
and U6500 (N_6500,N_237,N_1178);
or U6501 (N_6501,N_244,N_2094);
and U6502 (N_6502,N_3169,N_1934);
nor U6503 (N_6503,N_3404,N_4083);
and U6504 (N_6504,N_111,N_462);
nand U6505 (N_6505,N_1266,N_4613);
nand U6506 (N_6506,N_2147,N_1289);
or U6507 (N_6507,N_2800,N_3985);
nor U6508 (N_6508,N_2164,N_1072);
or U6509 (N_6509,N_2606,N_999);
and U6510 (N_6510,N_4458,N_1212);
or U6511 (N_6511,N_4700,N_546);
or U6512 (N_6512,N_1889,N_402);
nor U6513 (N_6513,N_3033,N_2629);
nand U6514 (N_6514,N_4431,N_4694);
nand U6515 (N_6515,N_1198,N_1570);
nand U6516 (N_6516,N_3642,N_2032);
nand U6517 (N_6517,N_1274,N_1339);
nand U6518 (N_6518,N_3879,N_3761);
xor U6519 (N_6519,N_2837,N_1163);
nor U6520 (N_6520,N_4779,N_3028);
nand U6521 (N_6521,N_1525,N_2588);
nand U6522 (N_6522,N_3356,N_1891);
or U6523 (N_6523,N_4225,N_181);
or U6524 (N_6524,N_2855,N_3485);
or U6525 (N_6525,N_599,N_1350);
or U6526 (N_6526,N_3182,N_1231);
nand U6527 (N_6527,N_397,N_3491);
and U6528 (N_6528,N_3263,N_4749);
and U6529 (N_6529,N_4704,N_4987);
nand U6530 (N_6530,N_1090,N_1756);
or U6531 (N_6531,N_1373,N_4386);
or U6532 (N_6532,N_1545,N_342);
or U6533 (N_6533,N_4885,N_495);
or U6534 (N_6534,N_2618,N_2759);
nor U6535 (N_6535,N_2141,N_1745);
nand U6536 (N_6536,N_1333,N_146);
or U6537 (N_6537,N_4174,N_1002);
or U6538 (N_6538,N_3575,N_3851);
and U6539 (N_6539,N_1210,N_3211);
or U6540 (N_6540,N_3247,N_4308);
nand U6541 (N_6541,N_4032,N_2422);
xnor U6542 (N_6542,N_947,N_1254);
xnor U6543 (N_6543,N_1328,N_895);
and U6544 (N_6544,N_821,N_726);
nor U6545 (N_6545,N_3128,N_2854);
or U6546 (N_6546,N_4952,N_969);
nor U6547 (N_6547,N_1071,N_2572);
and U6548 (N_6548,N_4908,N_3662);
and U6549 (N_6549,N_1646,N_951);
or U6550 (N_6550,N_424,N_4938);
nand U6551 (N_6551,N_2971,N_3968);
nor U6552 (N_6552,N_52,N_1150);
and U6553 (N_6553,N_1287,N_4178);
and U6554 (N_6554,N_3299,N_4034);
nand U6555 (N_6555,N_1515,N_696);
nand U6556 (N_6556,N_757,N_3782);
or U6557 (N_6557,N_3494,N_2655);
nand U6558 (N_6558,N_855,N_694);
or U6559 (N_6559,N_3092,N_4310);
nand U6560 (N_6560,N_440,N_3814);
nand U6561 (N_6561,N_2180,N_4729);
and U6562 (N_6562,N_3858,N_3864);
nor U6563 (N_6563,N_2335,N_3734);
nand U6564 (N_6564,N_713,N_3647);
nand U6565 (N_6565,N_4316,N_4379);
nor U6566 (N_6566,N_1462,N_2333);
and U6567 (N_6567,N_2530,N_2922);
or U6568 (N_6568,N_1956,N_1590);
nor U6569 (N_6569,N_2288,N_4163);
and U6570 (N_6570,N_835,N_3572);
and U6571 (N_6571,N_1727,N_2956);
nand U6572 (N_6572,N_1892,N_4255);
and U6573 (N_6573,N_2105,N_220);
nand U6574 (N_6574,N_1866,N_2138);
and U6575 (N_6575,N_3095,N_3612);
or U6576 (N_6576,N_3776,N_4534);
and U6577 (N_6577,N_2220,N_4719);
or U6578 (N_6578,N_3677,N_1334);
nor U6579 (N_6579,N_2042,N_2512);
and U6580 (N_6580,N_414,N_537);
nor U6581 (N_6581,N_4472,N_2004);
nor U6582 (N_6582,N_1541,N_1909);
nand U6583 (N_6583,N_4829,N_439);
and U6584 (N_6584,N_3738,N_4516);
nand U6585 (N_6585,N_3069,N_4022);
nor U6586 (N_6586,N_1529,N_4769);
or U6587 (N_6587,N_4354,N_867);
nor U6588 (N_6588,N_259,N_945);
nor U6589 (N_6589,N_3661,N_4592);
nor U6590 (N_6590,N_912,N_1123);
and U6591 (N_6591,N_13,N_4831);
and U6592 (N_6592,N_3714,N_211);
nand U6593 (N_6593,N_2907,N_556);
or U6594 (N_6594,N_2573,N_504);
nor U6595 (N_6595,N_338,N_4658);
nor U6596 (N_6596,N_1435,N_755);
or U6597 (N_6597,N_3052,N_1857);
and U6598 (N_6598,N_2874,N_2821);
or U6599 (N_6599,N_1595,N_785);
and U6600 (N_6600,N_2324,N_3720);
nor U6601 (N_6601,N_4582,N_607);
or U6602 (N_6602,N_3220,N_4866);
and U6603 (N_6603,N_1877,N_4902);
nor U6604 (N_6604,N_2926,N_228);
nor U6605 (N_6605,N_383,N_3995);
or U6606 (N_6606,N_2253,N_107);
nor U6607 (N_6607,N_4792,N_2526);
nor U6608 (N_6608,N_2591,N_128);
or U6609 (N_6609,N_1214,N_1133);
nor U6610 (N_6610,N_2006,N_1155);
or U6611 (N_6611,N_1879,N_3696);
and U6612 (N_6612,N_2946,N_2782);
nor U6613 (N_6613,N_4161,N_1659);
nand U6614 (N_6614,N_3270,N_1983);
and U6615 (N_6615,N_1319,N_2816);
nand U6616 (N_6616,N_3448,N_779);
and U6617 (N_6617,N_2208,N_1037);
and U6618 (N_6618,N_531,N_2350);
or U6619 (N_6619,N_3593,N_4578);
and U6620 (N_6620,N_3886,N_4628);
nor U6621 (N_6621,N_324,N_977);
and U6622 (N_6622,N_3030,N_1611);
and U6623 (N_6623,N_132,N_3832);
nand U6624 (N_6624,N_4115,N_771);
or U6625 (N_6625,N_3787,N_3198);
or U6626 (N_6626,N_4679,N_4074);
or U6627 (N_6627,N_1680,N_4660);
nor U6628 (N_6628,N_3377,N_145);
nand U6629 (N_6629,N_157,N_48);
nor U6630 (N_6630,N_2030,N_2564);
nor U6631 (N_6631,N_4637,N_1961);
nor U6632 (N_6632,N_3437,N_4471);
nand U6633 (N_6633,N_966,N_2415);
nor U6634 (N_6634,N_190,N_1568);
nor U6635 (N_6635,N_34,N_1478);
and U6636 (N_6636,N_2621,N_1688);
or U6637 (N_6637,N_352,N_2827);
nand U6638 (N_6638,N_3951,N_1278);
or U6639 (N_6639,N_4882,N_934);
nand U6640 (N_6640,N_809,N_2290);
and U6641 (N_6641,N_3870,N_576);
and U6642 (N_6642,N_4797,N_1630);
or U6643 (N_6643,N_1033,N_1720);
nand U6644 (N_6644,N_679,N_3967);
nand U6645 (N_6645,N_2401,N_3262);
nor U6646 (N_6646,N_1104,N_444);
or U6647 (N_6647,N_4577,N_2067);
and U6648 (N_6648,N_1195,N_1418);
and U6649 (N_6649,N_3196,N_692);
nand U6650 (N_6650,N_1759,N_3922);
nand U6651 (N_6651,N_4017,N_459);
nor U6652 (N_6652,N_3295,N_2961);
and U6653 (N_6653,N_1801,N_2416);
nor U6654 (N_6654,N_4186,N_720);
and U6655 (N_6655,N_3727,N_601);
nand U6656 (N_6656,N_2640,N_1783);
nor U6657 (N_6657,N_2427,N_3591);
and U6658 (N_6658,N_1780,N_484);
nor U6659 (N_6659,N_634,N_3547);
nor U6660 (N_6660,N_3281,N_2893);
nor U6661 (N_6661,N_2627,N_4990);
nor U6662 (N_6662,N_1925,N_4644);
and U6663 (N_6663,N_3241,N_1020);
or U6664 (N_6664,N_1032,N_1500);
and U6665 (N_6665,N_2802,N_4602);
nor U6666 (N_6666,N_1503,N_1013);
or U6667 (N_6667,N_282,N_1243);
nand U6668 (N_6668,N_2410,N_330);
nor U6669 (N_6669,N_2036,N_320);
or U6670 (N_6670,N_585,N_786);
and U6671 (N_6671,N_2058,N_4924);
nand U6672 (N_6672,N_3145,N_4421);
nor U6673 (N_6673,N_2991,N_245);
and U6674 (N_6674,N_3252,N_1051);
nand U6675 (N_6675,N_4359,N_1859);
or U6676 (N_6676,N_4512,N_87);
and U6677 (N_6677,N_2636,N_4442);
and U6678 (N_6678,N_3889,N_749);
nor U6679 (N_6679,N_1648,N_1065);
and U6680 (N_6680,N_892,N_2568);
and U6681 (N_6681,N_1637,N_3669);
or U6682 (N_6682,N_3981,N_2807);
and U6683 (N_6683,N_836,N_3153);
and U6684 (N_6684,N_4668,N_2982);
nand U6685 (N_6685,N_3348,N_3910);
nand U6686 (N_6686,N_3376,N_1672);
or U6687 (N_6687,N_4874,N_195);
or U6688 (N_6688,N_411,N_622);
nor U6689 (N_6689,N_2229,N_873);
or U6690 (N_6690,N_4814,N_2219);
and U6691 (N_6691,N_3808,N_3728);
nand U6692 (N_6692,N_1791,N_568);
and U6693 (N_6693,N_2630,N_3916);
or U6694 (N_6694,N_2889,N_919);
nand U6695 (N_6695,N_4011,N_4645);
and U6696 (N_6696,N_2728,N_4850);
nor U6697 (N_6697,N_4889,N_4141);
nand U6698 (N_6698,N_3838,N_4488);
nand U6699 (N_6699,N_23,N_781);
nor U6700 (N_6700,N_1922,N_1973);
and U6701 (N_6701,N_796,N_2201);
nand U6702 (N_6702,N_2365,N_488);
nand U6703 (N_6703,N_2370,N_718);
nand U6704 (N_6704,N_2472,N_3166);
nor U6705 (N_6705,N_897,N_3324);
and U6706 (N_6706,N_2544,N_1588);
nor U6707 (N_6707,N_3693,N_1023);
and U6708 (N_6708,N_2643,N_4986);
or U6709 (N_6709,N_3139,N_4942);
xor U6710 (N_6710,N_1736,N_2898);
or U6711 (N_6711,N_2822,N_1989);
nor U6712 (N_6712,N_64,N_3903);
nor U6713 (N_6713,N_1208,N_4239);
nor U6714 (N_6714,N_4210,N_4997);
nor U6715 (N_6715,N_44,N_792);
nand U6716 (N_6716,N_3554,N_4647);
nor U6717 (N_6717,N_862,N_988);
or U6718 (N_6718,N_2373,N_47);
and U6719 (N_6719,N_3321,N_2354);
nor U6720 (N_6720,N_3848,N_3587);
and U6721 (N_6721,N_510,N_907);
and U6722 (N_6722,N_4048,N_3594);
and U6723 (N_6723,N_4384,N_3361);
nand U6724 (N_6724,N_4948,N_3807);
and U6725 (N_6725,N_4527,N_918);
or U6726 (N_6726,N_1923,N_4839);
nand U6727 (N_6727,N_1530,N_1941);
nor U6728 (N_6728,N_3873,N_3545);
and U6729 (N_6729,N_3339,N_3794);
nor U6730 (N_6730,N_596,N_4462);
xnor U6731 (N_6731,N_2477,N_2037);
nor U6732 (N_6732,N_179,N_3617);
nand U6733 (N_6733,N_339,N_3269);
nand U6734 (N_6734,N_4059,N_4858);
and U6735 (N_6735,N_1718,N_139);
and U6736 (N_6736,N_4755,N_135);
and U6737 (N_6737,N_1758,N_3895);
nor U6738 (N_6738,N_2016,N_1455);
nor U6739 (N_6739,N_4060,N_3380);
nor U6740 (N_6740,N_4441,N_4393);
or U6741 (N_6741,N_2547,N_3440);
nor U6742 (N_6742,N_1483,N_2282);
or U6743 (N_6743,N_2,N_479);
nand U6744 (N_6744,N_1760,N_202);
or U6745 (N_6745,N_4104,N_1356);
and U6746 (N_6746,N_43,N_2872);
nand U6747 (N_6747,N_4086,N_1204);
nand U6748 (N_6748,N_117,N_1282);
nand U6749 (N_6749,N_2819,N_2823);
and U6750 (N_6750,N_2829,N_4738);
nand U6751 (N_6751,N_1003,N_2320);
and U6752 (N_6752,N_3110,N_4713);
nand U6753 (N_6753,N_3455,N_3906);
or U6754 (N_6754,N_4955,N_3852);
and U6755 (N_6755,N_3762,N_924);
nand U6756 (N_6756,N_965,N_3114);
or U6757 (N_6757,N_318,N_2473);
nor U6758 (N_6758,N_2548,N_1980);
and U6759 (N_6759,N_359,N_4187);
and U6760 (N_6760,N_1197,N_2690);
nor U6761 (N_6761,N_1097,N_1669);
or U6762 (N_6762,N_1257,N_3690);
or U6763 (N_6763,N_3044,N_3499);
or U6764 (N_6764,N_2996,N_279);
and U6765 (N_6765,N_2932,N_1853);
and U6766 (N_6766,N_2750,N_3261);
nand U6767 (N_6767,N_3370,N_76);
xnor U6768 (N_6768,N_2443,N_2504);
nand U6769 (N_6769,N_2929,N_3390);
nand U6770 (N_6770,N_3764,N_3541);
nor U6771 (N_6771,N_830,N_956);
nand U6772 (N_6772,N_688,N_1582);
nor U6773 (N_6773,N_3116,N_868);
nand U6774 (N_6774,N_3396,N_3533);
and U6775 (N_6775,N_451,N_954);
or U6776 (N_6776,N_2910,N_1920);
and U6777 (N_6777,N_3117,N_84);
xor U6778 (N_6778,N_2257,N_0);
or U6779 (N_6779,N_3336,N_2081);
or U6780 (N_6780,N_3793,N_3777);
nor U6781 (N_6781,N_1425,N_1907);
nand U6782 (N_6782,N_2647,N_4270);
nand U6783 (N_6783,N_1103,N_500);
nand U6784 (N_6784,N_1275,N_3009);
or U6785 (N_6785,N_3234,N_3672);
and U6786 (N_6786,N_4293,N_1609);
and U6787 (N_6787,N_1226,N_4092);
nor U6788 (N_6788,N_1794,N_2400);
and U6789 (N_6789,N_2090,N_4872);
nor U6790 (N_6790,N_1860,N_2969);
nor U6791 (N_6791,N_3466,N_958);
nand U6792 (N_6792,N_2765,N_1766);
or U6793 (N_6793,N_3146,N_1773);
nand U6794 (N_6794,N_1612,N_3273);
nand U6795 (N_6795,N_3227,N_4661);
or U6796 (N_6796,N_1064,N_3429);
nand U6797 (N_6797,N_4233,N_4974);
nand U6798 (N_6798,N_95,N_152);
nor U6799 (N_6799,N_1839,N_3045);
and U6800 (N_6800,N_1246,N_2277);
nand U6801 (N_6801,N_2725,N_182);
or U6802 (N_6802,N_559,N_2744);
nand U6803 (N_6803,N_2151,N_2944);
and U6804 (N_6804,N_864,N_3722);
or U6805 (N_6805,N_1099,N_4773);
nand U6806 (N_6806,N_3253,N_2935);
nor U6807 (N_6807,N_1397,N_102);
and U6808 (N_6808,N_1613,N_2376);
nand U6809 (N_6809,N_3941,N_3824);
or U6810 (N_6810,N_67,N_4643);
nand U6811 (N_6811,N_2813,N_1492);
nand U6812 (N_6812,N_2764,N_65);
or U6813 (N_6813,N_3896,N_3083);
nand U6814 (N_6814,N_141,N_3436);
or U6815 (N_6815,N_3918,N_3664);
nand U6816 (N_6816,N_3451,N_4511);
nor U6817 (N_6817,N_2625,N_4018);
nand U6818 (N_6818,N_4450,N_4508);
or U6819 (N_6819,N_1561,N_4786);
nand U6820 (N_6820,N_3003,N_313);
and U6821 (N_6821,N_4485,N_4454);
nor U6822 (N_6822,N_4761,N_1884);
or U6823 (N_6823,N_3222,N_2181);
nand U6824 (N_6824,N_4618,N_663);
or U6825 (N_6825,N_1272,N_1011);
nand U6826 (N_6826,N_2063,N_3899);
nor U6827 (N_6827,N_437,N_552);
nand U6828 (N_6828,N_3057,N_2917);
or U6829 (N_6829,N_343,N_4799);
nand U6830 (N_6830,N_624,N_3144);
or U6831 (N_6831,N_4281,N_3708);
nand U6832 (N_6832,N_3950,N_1049);
and U6833 (N_6833,N_3919,N_3019);
and U6834 (N_6834,N_4727,N_2936);
nand U6835 (N_6835,N_3507,N_3471);
or U6836 (N_6836,N_1695,N_3018);
and U6837 (N_6837,N_1138,N_1540);
or U6838 (N_6838,N_3240,N_168);
and U6839 (N_6839,N_1106,N_490);
or U6840 (N_6840,N_4598,N_3413);
or U6841 (N_6841,N_4718,N_4087);
and U6842 (N_6842,N_4352,N_1632);
or U6843 (N_6843,N_3365,N_2664);
nand U6844 (N_6844,N_3097,N_408);
and U6845 (N_6845,N_4195,N_2241);
nand U6846 (N_6846,N_4024,N_1161);
nor U6847 (N_6847,N_2239,N_1700);
nor U6848 (N_6848,N_4043,N_3122);
xor U6849 (N_6849,N_1835,N_162);
and U6850 (N_6850,N_4220,N_3334);
nor U6851 (N_6851,N_3081,N_1160);
or U6852 (N_6852,N_4535,N_3394);
and U6853 (N_6853,N_4313,N_922);
and U6854 (N_6854,N_2132,N_1850);
nand U6855 (N_6855,N_1505,N_149);
nor U6856 (N_6856,N_1789,N_3462);
or U6857 (N_6857,N_2523,N_9);
nor U6858 (N_6858,N_1075,N_2794);
or U6859 (N_6859,N_3107,N_941);
nor U6860 (N_6860,N_3154,N_4213);
nor U6861 (N_6861,N_124,N_2680);
nor U6862 (N_6862,N_4650,N_2646);
and U6863 (N_6863,N_869,N_1042);
nand U6864 (N_6864,N_2230,N_4331);
nor U6865 (N_6865,N_1830,N_4895);
or U6866 (N_6866,N_3563,N_2140);
nand U6867 (N_6867,N_1009,N_4283);
or U6868 (N_6868,N_1597,N_4978);
nand U6869 (N_6869,N_876,N_2387);
nor U6870 (N_6870,N_4980,N_2534);
or U6871 (N_6871,N_4497,N_819);
nand U6872 (N_6872,N_222,N_4808);
or U6873 (N_6873,N_2486,N_2103);
nor U6874 (N_6874,N_61,N_2453);
or U6875 (N_6875,N_4004,N_841);
or U6876 (N_6876,N_4047,N_3042);
and U6877 (N_6877,N_4683,N_2989);
nor U6878 (N_6878,N_833,N_260);
and U6879 (N_6879,N_4853,N_465);
and U6880 (N_6880,N_3453,N_729);
nand U6881 (N_6881,N_1633,N_3352);
nor U6882 (N_6882,N_2308,N_4675);
nor U6883 (N_6883,N_4333,N_1224);
or U6884 (N_6884,N_2797,N_984);
or U6885 (N_6885,N_815,N_2511);
and U6886 (N_6886,N_332,N_996);
or U6887 (N_6887,N_4330,N_3293);
and U6888 (N_6888,N_1380,N_3298);
or U6889 (N_6889,N_4857,N_595);
and U6890 (N_6890,N_1509,N_931);
nor U6891 (N_6891,N_957,N_2538);
or U6892 (N_6892,N_401,N_4258);
and U6893 (N_6893,N_3469,N_4932);
or U6894 (N_6894,N_2896,N_4042);
and U6895 (N_6895,N_4890,N_3430);
nand U6896 (N_6896,N_1937,N_4324);
and U6897 (N_6897,N_4483,N_364);
and U6898 (N_6898,N_2743,N_3306);
and U6899 (N_6899,N_1217,N_3658);
nor U6900 (N_6900,N_3676,N_53);
nand U6901 (N_6901,N_4935,N_4985);
nand U6902 (N_6902,N_2093,N_923);
nor U6903 (N_6903,N_1512,N_4190);
nor U6904 (N_6904,N_106,N_1579);
nor U6905 (N_6905,N_4536,N_4921);
nand U6906 (N_6906,N_3550,N_1293);
xnor U6907 (N_6907,N_175,N_550);
nand U6908 (N_6908,N_4181,N_1300);
and U6909 (N_6909,N_3869,N_903);
nor U6910 (N_6910,N_1861,N_3614);
nand U6911 (N_6911,N_4530,N_110);
nand U6912 (N_6912,N_1236,N_3067);
and U6913 (N_6913,N_207,N_3072);
and U6914 (N_6914,N_4888,N_1657);
nand U6915 (N_6915,N_1338,N_3963);
nand U6916 (N_6916,N_1173,N_1129);
nand U6917 (N_6917,N_982,N_4052);
or U6918 (N_6918,N_920,N_811);
nand U6919 (N_6919,N_3470,N_4739);
nor U6920 (N_6920,N_3457,N_4636);
nor U6921 (N_6921,N_4071,N_136);
and U6922 (N_6922,N_1280,N_1050);
and U6923 (N_6923,N_777,N_3713);
or U6924 (N_6924,N_3773,N_308);
nor U6925 (N_6925,N_4672,N_3493);
nand U6926 (N_6926,N_3973,N_1986);
nand U6927 (N_6927,N_4276,N_2404);
nand U6928 (N_6928,N_2306,N_1829);
and U6929 (N_6929,N_4099,N_3213);
nor U6930 (N_6930,N_4564,N_3089);
or U6931 (N_6931,N_1836,N_3066);
nor U6932 (N_6932,N_4572,N_2948);
or U6933 (N_6933,N_4876,N_4107);
nand U6934 (N_6934,N_3933,N_1461);
and U6935 (N_6935,N_801,N_1585);
nand U6936 (N_6936,N_1030,N_3285);
nor U6937 (N_6937,N_1921,N_4517);
and U6938 (N_6938,N_290,N_4633);
and U6939 (N_6939,N_255,N_4617);
nor U6940 (N_6940,N_4490,N_4363);
or U6941 (N_6941,N_3091,N_2238);
nand U6942 (N_6942,N_2828,N_1322);
nor U6943 (N_6943,N_256,N_812);
nor U6944 (N_6944,N_438,N_3417);
or U6945 (N_6945,N_3663,N_2578);
nand U6946 (N_6946,N_3260,N_3597);
nand U6947 (N_6947,N_4194,N_832);
nand U6948 (N_6948,N_1315,N_2894);
nand U6949 (N_6949,N_1428,N_2269);
or U6950 (N_6950,N_2172,N_300);
and U6951 (N_6951,N_2186,N_4355);
nor U6952 (N_6952,N_4499,N_3908);
nand U6953 (N_6953,N_1000,N_3796);
nor U6954 (N_6954,N_2799,N_3512);
nor U6955 (N_6955,N_1614,N_4158);
and U6956 (N_6956,N_2590,N_264);
nand U6957 (N_6957,N_758,N_571);
nand U6958 (N_6958,N_1864,N_3666);
or U6959 (N_6959,N_3701,N_4705);
nand U6960 (N_6960,N_2463,N_1993);
nor U6961 (N_6961,N_2490,N_4271);
and U6962 (N_6962,N_2973,N_1484);
nand U6963 (N_6963,N_2024,N_3626);
and U6964 (N_6964,N_3881,N_1306);
and U6965 (N_6965,N_2652,N_4157);
nand U6966 (N_6966,N_489,N_2733);
nor U6967 (N_6967,N_684,N_3049);
or U6968 (N_6968,N_452,N_2046);
and U6969 (N_6969,N_1433,N_2244);
nand U6970 (N_6970,N_3790,N_1376);
and U6971 (N_6971,N_3804,N_4716);
or U6972 (N_6972,N_2285,N_4207);
or U6973 (N_6973,N_1139,N_3510);
and U6974 (N_6974,N_4922,N_4969);
nand U6975 (N_6975,N_4256,N_3191);
nor U6976 (N_6976,N_803,N_2569);
and U6977 (N_6977,N_1824,N_3118);
nor U6978 (N_6978,N_3123,N_483);
and U6979 (N_6979,N_598,N_5);
or U6980 (N_6980,N_2184,N_2047);
and U6981 (N_6981,N_4620,N_3960);
nor U6982 (N_6982,N_541,N_1386);
or U6983 (N_6983,N_4434,N_2291);
and U6984 (N_6984,N_250,N_3226);
nand U6985 (N_6985,N_1382,N_3725);
and U6986 (N_6986,N_3392,N_4811);
or U6987 (N_6987,N_2281,N_3540);
nor U6988 (N_6988,N_467,N_4467);
nand U6989 (N_6989,N_4898,N_4982);
or U6990 (N_6990,N_1808,N_2389);
nand U6991 (N_6991,N_4953,N_946);
and U6992 (N_6992,N_1060,N_4871);
or U6993 (N_6993,N_4752,N_2574);
or U6994 (N_6994,N_4428,N_899);
nand U6995 (N_6995,N_2359,N_1408);
nor U6996 (N_6996,N_4500,N_3632);
nand U6997 (N_6997,N_2610,N_3195);
nand U6998 (N_6998,N_201,N_3984);
and U6999 (N_6999,N_3205,N_2072);
or U7000 (N_7000,N_1430,N_885);
or U7001 (N_7001,N_4039,N_1685);
and U7002 (N_7002,N_4821,N_1454);
nor U7003 (N_7003,N_528,N_4552);
or U7004 (N_7004,N_3509,N_3397);
or U7005 (N_7005,N_4550,N_3779);
nand U7006 (N_7006,N_3181,N_2775);
nand U7007 (N_7007,N_1774,N_1683);
xnor U7008 (N_7008,N_730,N_1083);
nor U7009 (N_7009,N_285,N_4531);
nor U7010 (N_7010,N_2634,N_221);
nand U7011 (N_7011,N_1349,N_3600);
nand U7012 (N_7012,N_3737,N_1167);
and U7013 (N_7013,N_390,N_4362);
nand U7014 (N_7014,N_2192,N_4282);
or U7015 (N_7015,N_1442,N_94);
nand U7016 (N_7016,N_1177,N_2543);
or U7017 (N_7017,N_698,N_930);
nand U7018 (N_7018,N_474,N_4350);
and U7019 (N_7019,N_463,N_901);
nor U7020 (N_7020,N_1377,N_4804);
or U7021 (N_7021,N_4003,N_4425);
and U7022 (N_7022,N_4460,N_3249);
or U7023 (N_7023,N_497,N_4284);
nor U7024 (N_7024,N_400,N_1807);
or U7025 (N_7025,N_2906,N_3482);
or U7026 (N_7026,N_3821,N_4432);
or U7027 (N_7027,N_1650,N_4625);
or U7028 (N_7028,N_2107,N_750);
or U7029 (N_7029,N_178,N_2605);
nand U7030 (N_7030,N_2840,N_262);
and U7031 (N_7031,N_3029,N_2384);
nor U7032 (N_7032,N_2752,N_2475);
nor U7033 (N_7033,N_1387,N_3887);
and U7034 (N_7034,N_690,N_1227);
nand U7035 (N_7035,N_1658,N_3265);
and U7036 (N_7036,N_4335,N_3418);
nor U7037 (N_7037,N_4855,N_2754);
nor U7038 (N_7038,N_1769,N_100);
or U7039 (N_7039,N_4286,N_2041);
nand U7040 (N_7040,N_4563,N_3388);
and U7041 (N_7041,N_643,N_200);
nor U7042 (N_7042,N_1698,N_879);
and U7043 (N_7043,N_205,N_1101);
nand U7044 (N_7044,N_1238,N_1693);
and U7045 (N_7045,N_3244,N_3993);
or U7046 (N_7046,N_2020,N_2867);
or U7047 (N_7047,N_515,N_745);
or U7048 (N_7048,N_3588,N_1182);
or U7049 (N_7049,N_1826,N_4676);
and U7050 (N_7050,N_3928,N_4079);
nand U7051 (N_7051,N_632,N_4775);
nor U7052 (N_7052,N_4780,N_1886);
nand U7053 (N_7053,N_1436,N_4583);
nor U7054 (N_7054,N_937,N_3923);
or U7055 (N_7055,N_2862,N_843);
nor U7056 (N_7056,N_1403,N_614);
nor U7057 (N_7057,N_3328,N_703);
nand U7058 (N_7058,N_4635,N_4360);
and U7059 (N_7059,N_4794,N_2143);
or U7060 (N_7060,N_4031,N_375);
and U7061 (N_7061,N_4176,N_4474);
nor U7062 (N_7062,N_1818,N_4367);
and U7063 (N_7063,N_2346,N_2367);
or U7064 (N_7064,N_2018,N_3354);
or U7065 (N_7065,N_3946,N_1662);
or U7066 (N_7066,N_138,N_3706);
nand U7067 (N_7067,N_3138,N_4975);
nand U7068 (N_7068,N_2562,N_4940);
and U7069 (N_7069,N_4035,N_1748);
or U7070 (N_7070,N_1183,N_1093);
or U7071 (N_7071,N_944,N_1434);
or U7072 (N_7072,N_1395,N_1031);
or U7073 (N_7073,N_3883,N_4823);
nor U7074 (N_7074,N_1117,N_4299);
nand U7075 (N_7075,N_4573,N_2076);
or U7076 (N_7076,N_2112,N_3536);
nand U7077 (N_7077,N_3373,N_2879);
nand U7078 (N_7078,N_4321,N_2835);
nor U7079 (N_7079,N_1471,N_3900);
nor U7080 (N_7080,N_4848,N_3311);
nor U7081 (N_7081,N_4387,N_2356);
and U7082 (N_7082,N_511,N_55);
xnor U7083 (N_7083,N_1463,N_3444);
nand U7084 (N_7084,N_3977,N_647);
nor U7085 (N_7085,N_112,N_3502);
or U7086 (N_7086,N_3481,N_4774);
nand U7087 (N_7087,N_2169,N_767);
nand U7088 (N_7088,N_3383,N_2382);
nand U7089 (N_7089,N_2992,N_704);
nand U7090 (N_7090,N_2435,N_4053);
nand U7091 (N_7091,N_2505,N_701);
and U7092 (N_7092,N_693,N_896);
or U7093 (N_7093,N_2135,N_1825);
nand U7094 (N_7094,N_2234,N_3580);
or U7095 (N_7095,N_780,N_3310);
nor U7096 (N_7096,N_3239,N_1795);
nor U7097 (N_7097,N_4820,N_3855);
or U7098 (N_7098,N_4696,N_555);
or U7099 (N_7099,N_4862,N_335);
or U7100 (N_7100,N_3326,N_908);
nand U7101 (N_7101,N_2255,N_1497);
nor U7102 (N_7102,N_4037,N_4758);
and U7103 (N_7103,N_1569,N_1452);
nand U7104 (N_7104,N_3924,N_4854);
or U7105 (N_7105,N_564,N_987);
nand U7106 (N_7106,N_268,N_2015);
and U7107 (N_7107,N_4827,N_1564);
nor U7108 (N_7108,N_242,N_4173);
nand U7109 (N_7109,N_427,N_2820);
or U7110 (N_7110,N_4785,N_814);
or U7111 (N_7111,N_1025,N_3844);
nand U7112 (N_7112,N_3558,N_1066);
nand U7113 (N_7113,N_2831,N_2113);
or U7114 (N_7114,N_2068,N_1875);
and U7115 (N_7115,N_2774,N_2498);
nor U7116 (N_7116,N_4735,N_722);
and U7117 (N_7117,N_3947,N_3717);
or U7118 (N_7118,N_109,N_4842);
or U7119 (N_7119,N_154,N_2575);
or U7120 (N_7120,N_2723,N_3531);
nor U7121 (N_7121,N_2278,N_1176);
xnor U7122 (N_7122,N_2609,N_680);
nor U7123 (N_7123,N_1558,N_1175);
or U7124 (N_7124,N_4409,N_1458);
and U7125 (N_7125,N_2866,N_3101);
nand U7126 (N_7126,N_4028,N_3468);
nand U7127 (N_7127,N_1998,N_2357);
or U7128 (N_7128,N_4648,N_3670);
nor U7129 (N_7129,N_2091,N_4056);
nor U7130 (N_7130,N_4096,N_1166);
or U7131 (N_7131,N_2130,N_4165);
and U7132 (N_7132,N_1942,N_2338);
and U7133 (N_7133,N_3834,N_376);
and U7134 (N_7134,N_4374,N_3320);
and U7135 (N_7135,N_1576,N_4336);
and U7136 (N_7136,N_2116,N_2873);
nand U7137 (N_7137,N_1784,N_3648);
nand U7138 (N_7138,N_686,N_3585);
and U7139 (N_7139,N_3530,N_2417);
nor U7140 (N_7140,N_3909,N_1631);
nor U7141 (N_7141,N_2089,N_2368);
and U7142 (N_7142,N_1560,N_2102);
and U7143 (N_7143,N_593,N_1327);
and U7144 (N_7144,N_1045,N_1868);
nand U7145 (N_7145,N_2587,N_4707);
nand U7146 (N_7146,N_2585,N_4478);
nor U7147 (N_7147,N_1057,N_4607);
nor U7148 (N_7148,N_4251,N_1070);
nor U7149 (N_7149,N_3027,N_2251);
or U7150 (N_7150,N_1976,N_3465);
or U7151 (N_7151,N_4965,N_2970);
and U7152 (N_7152,N_3225,N_3132);
nor U7153 (N_7153,N_443,N_1627);
nor U7154 (N_7154,N_3423,N_1940);
or U7155 (N_7155,N_2930,N_2160);
nand U7156 (N_7156,N_3480,N_368);
nor U7157 (N_7157,N_2480,N_4227);
and U7158 (N_7158,N_2875,N_4192);
or U7159 (N_7159,N_4603,N_2446);
nand U7160 (N_7160,N_716,N_4574);
and U7161 (N_7161,N_2340,N_2494);
or U7162 (N_7162,N_229,N_731);
and U7163 (N_7163,N_1514,N_1365);
nand U7164 (N_7164,N_3880,N_2758);
or U7165 (N_7165,N_3106,N_3420);
or U7166 (N_7166,N_2737,N_1926);
and U7167 (N_7167,N_723,N_2730);
nor U7168 (N_7168,N_2657,N_4492);
or U7169 (N_7169,N_3020,N_1312);
and U7170 (N_7170,N_63,N_854);
and U7171 (N_7171,N_3932,N_233);
and U7172 (N_7172,N_4875,N_3602);
nor U7173 (N_7173,N_681,N_2044);
or U7174 (N_7174,N_4323,N_3716);
nand U7175 (N_7175,N_296,N_1793);
nand U7176 (N_7176,N_4044,N_3684);
or U7177 (N_7177,N_4072,N_125);
or U7178 (N_7178,N_4320,N_3987);
or U7179 (N_7179,N_2559,N_2892);
nand U7180 (N_7180,N_3719,N_3940);
nand U7181 (N_7181,N_4571,N_1523);
nand U7182 (N_7182,N_3379,N_4806);
or U7183 (N_7183,N_2332,N_986);
and U7184 (N_7184,N_3705,N_3991);
and U7185 (N_7185,N_4314,N_3384);
and U7186 (N_7186,N_3403,N_1359);
and U7187 (N_7187,N_3760,N_3415);
and U7188 (N_7188,N_1310,N_4358);
nand U7189 (N_7189,N_4188,N_2769);
nor U7190 (N_7190,N_4351,N_4545);
nand U7191 (N_7191,N_1740,N_169);
and U7192 (N_7192,N_551,N_2721);
or U7193 (N_7193,N_2763,N_733);
nand U7194 (N_7194,N_2049,N_1472);
nand U7195 (N_7195,N_1367,N_4057);
nand U7196 (N_7196,N_3335,N_744);
nor U7197 (N_7197,N_4020,N_719);
and U7198 (N_7198,N_1379,N_4081);
nor U7199 (N_7199,N_4007,N_509);
or U7200 (N_7200,N_316,N_310);
nor U7201 (N_7201,N_2375,N_648);
or U7202 (N_7202,N_2021,N_828);
nor U7203 (N_7203,N_1939,N_241);
nand U7204 (N_7204,N_1788,N_3375);
or U7205 (N_7205,N_591,N_204);
or U7206 (N_7206,N_265,N_3443);
nor U7207 (N_7207,N_475,N_292);
nand U7208 (N_7208,N_3551,N_1399);
and U7209 (N_7209,N_664,N_791);
and U7210 (N_7210,N_4993,N_3700);
or U7211 (N_7211,N_566,N_4136);
or U7212 (N_7212,N_3061,N_3624);
or U7213 (N_7213,N_238,N_2716);
nand U7214 (N_7214,N_4091,N_2790);
or U7215 (N_7215,N_606,N_2921);
nor U7216 (N_7216,N_1647,N_1142);
or U7217 (N_7217,N_4010,N_2838);
and U7218 (N_7218,N_1510,N_3242);
or U7219 (N_7219,N_403,N_2871);
nand U7220 (N_7220,N_1775,N_3979);
nor U7221 (N_7221,N_646,N_4296);
or U7222 (N_7222,N_1749,N_1504);
nor U7223 (N_7223,N_4375,N_838);
and U7224 (N_7224,N_327,N_1288);
nor U7225 (N_7225,N_4623,N_2600);
or U7226 (N_7226,N_1697,N_3668);
nor U7227 (N_7227,N_2550,N_2527);
and U7228 (N_7228,N_1742,N_3974);
nand U7229 (N_7229,N_620,N_349);
or U7230 (N_7230,N_4995,N_4747);
nor U7231 (N_7231,N_4762,N_4977);
and U7232 (N_7232,N_1708,N_278);
nor U7233 (N_7233,N_608,N_1111);
or U7234 (N_7234,N_1062,N_581);
nor U7235 (N_7235,N_592,N_3186);
or U7236 (N_7236,N_4069,N_3623);
nor U7237 (N_7237,N_4593,N_2998);
and U7238 (N_7238,N_1378,N_3735);
or U7239 (N_7239,N_2447,N_1179);
nor U7240 (N_7240,N_2731,N_4584);
and U7241 (N_7241,N_3638,N_1330);
nand U7242 (N_7242,N_2483,N_2419);
or U7243 (N_7243,N_3120,N_1043);
nand U7244 (N_7244,N_1974,N_3358);
or U7245 (N_7245,N_4542,N_1346);
and U7246 (N_7246,N_1095,N_2330);
or U7247 (N_7247,N_2353,N_1871);
nand U7248 (N_7248,N_4988,N_4865);
and U7249 (N_7249,N_2520,N_3039);
or U7250 (N_7250,N_1017,N_3534);
or U7251 (N_7251,N_2626,N_1021);
or U7252 (N_7252,N_252,N_4134);
and U7253 (N_7253,N_517,N_1034);
xnor U7254 (N_7254,N_3141,N_549);
and U7255 (N_7255,N_306,N_6);
and U7256 (N_7256,N_725,N_4108);
nor U7257 (N_7257,N_3557,N_1126);
nand U7258 (N_7258,N_560,N_3006);
nand U7259 (N_7259,N_909,N_1820);
or U7260 (N_7260,N_1607,N_916);
and U7261 (N_7261,N_1968,N_3781);
nor U7262 (N_7262,N_2506,N_518);
nor U7263 (N_7263,N_3788,N_1714);
and U7264 (N_7264,N_3467,N_2849);
and U7265 (N_7265,N_2322,N_3327);
nor U7266 (N_7266,N_1575,N_4684);
nand U7267 (N_7267,N_3783,N_2616);
nand U7268 (N_7268,N_1470,N_654);
or U7269 (N_7269,N_936,N_1600);
nand U7270 (N_7270,N_2785,N_345);
nor U7271 (N_7271,N_158,N_1741);
nor U7272 (N_7272,N_1729,N_3149);
or U7273 (N_7273,N_30,N_2317);
nor U7274 (N_7274,N_108,N_4712);
and U7275 (N_7275,N_81,N_2773);
or U7276 (N_7276,N_3938,N_2581);
nand U7277 (N_7277,N_1995,N_4156);
and U7278 (N_7278,N_3505,N_1147);
and U7279 (N_7279,N_2264,N_1572);
or U7280 (N_7280,N_3073,N_4763);
and U7281 (N_7281,N_793,N_4547);
or U7282 (N_7282,N_4691,N_2722);
or U7283 (N_7283,N_2295,N_870);
and U7284 (N_7284,N_4247,N_1258);
nor U7285 (N_7285,N_4051,N_3627);
or U7286 (N_7286,N_18,N_4701);
and U7287 (N_7287,N_2088,N_2841);
nor U7288 (N_7288,N_4139,N_4880);
or U7289 (N_7289,N_4999,N_2366);
and U7290 (N_7290,N_4667,N_2309);
and U7291 (N_7291,N_4049,N_678);
xnor U7292 (N_7292,N_3683,N_4113);
nand U7293 (N_7293,N_4962,N_1897);
or U7294 (N_7294,N_470,N_1201);
or U7295 (N_7295,N_998,N_2080);
and U7296 (N_7296,N_741,N_4670);
nand U7297 (N_7297,N_674,N_3079);
and U7298 (N_7298,N_2425,N_3488);
or U7299 (N_7299,N_1779,N_2275);
nor U7300 (N_7300,N_372,N_2503);
or U7301 (N_7301,N_1603,N_4440);
nand U7302 (N_7302,N_1094,N_2380);
and U7303 (N_7303,N_2615,N_2594);
or U7304 (N_7304,N_2064,N_3929);
nor U7305 (N_7305,N_153,N_3093);
nand U7306 (N_7306,N_4153,N_4254);
xor U7307 (N_7307,N_4759,N_775);
nor U7308 (N_7308,N_3930,N_3060);
or U7309 (N_7309,N_1610,N_4244);
nor U7310 (N_7310,N_2144,N_1605);
nor U7311 (N_7311,N_1709,N_2958);
or U7312 (N_7312,N_4353,N_2845);
nand U7313 (N_7313,N_421,N_3537);
nand U7314 (N_7314,N_1388,N_1593);
or U7315 (N_7315,N_865,N_1880);
or U7316 (N_7316,N_4218,N_742);
nand U7317 (N_7317,N_2869,N_1707);
nor U7318 (N_7318,N_737,N_3228);
nand U7319 (N_7319,N_4588,N_627);
or U7320 (N_7320,N_520,N_3212);
or U7321 (N_7321,N_113,N_1445);
and U7322 (N_7322,N_3942,N_829);
nand U7323 (N_7323,N_1971,N_4546);
or U7324 (N_7324,N_1192,N_2379);
nand U7325 (N_7325,N_3075,N_1583);
or U7326 (N_7326,N_3811,N_2420);
nor U7327 (N_7327,N_3050,N_1767);
nand U7328 (N_7328,N_2202,N_3129);
nand U7329 (N_7329,N_4311,N_1608);
nor U7330 (N_7330,N_2128,N_4397);
nand U7331 (N_7331,N_2034,N_1180);
nor U7332 (N_7332,N_2327,N_2499);
and U7333 (N_7333,N_1027,N_366);
nor U7334 (N_7334,N_994,N_4599);
and U7335 (N_7335,N_3576,N_4124);
and U7336 (N_7336,N_3841,N_3193);
nor U7337 (N_7337,N_2836,N_4466);
and U7338 (N_7338,N_2768,N_1419);
nand U7339 (N_7339,N_258,N_4223);
nand U7340 (N_7340,N_340,N_273);
nor U7341 (N_7341,N_1761,N_38);
and U7342 (N_7342,N_2025,N_3391);
and U7343 (N_7343,N_2098,N_3156);
or U7344 (N_7344,N_4824,N_2260);
or U7345 (N_7345,N_611,N_3718);
nor U7346 (N_7346,N_2175,N_1508);
nor U7347 (N_7347,N_1145,N_1955);
or U7348 (N_7348,N_1098,N_3224);
or U7349 (N_7349,N_4537,N_4404);
nor U7350 (N_7350,N_602,N_1317);
or U7351 (N_7351,N_2895,N_3304);
and U7352 (N_7352,N_1298,N_3280);
nand U7353 (N_7353,N_3059,N_3207);
nor U7354 (N_7354,N_1059,N_3268);
nand U7355 (N_7355,N_418,N_4899);
nand U7356 (N_7356,N_4892,N_3151);
or U7357 (N_7357,N_2355,N_1674);
nand U7358 (N_7358,N_2145,N_3164);
nor U7359 (N_7359,N_574,N_4252);
or U7360 (N_7360,N_2950,N_800);
nand U7361 (N_7361,N_605,N_4493);
nor U7362 (N_7362,N_2043,N_1264);
nand U7363 (N_7363,N_2732,N_2314);
or U7364 (N_7364,N_2861,N_4894);
nand U7365 (N_7365,N_3374,N_2176);
nand U7366 (N_7366,N_4380,N_751);
nor U7367 (N_7367,N_294,N_1518);
and U7368 (N_7368,N_959,N_2975);
and U7369 (N_7369,N_2595,N_4180);
nor U7370 (N_7370,N_547,N_477);
and U7371 (N_7371,N_1473,N_1675);
or U7372 (N_7372,N_587,N_2466);
nand U7373 (N_7373,N_2381,N_3691);
nand U7374 (N_7374,N_4457,N_629);
nor U7375 (N_7375,N_1997,N_249);
nor U7376 (N_7376,N_4528,N_362);
nor U7377 (N_7377,N_4365,N_311);
nand U7378 (N_7378,N_1411,N_4826);
and U7379 (N_7379,N_4226,N_3736);
and U7380 (N_7380,N_186,N_86);
or U7381 (N_7381,N_4961,N_90);
nor U7382 (N_7382,N_4408,N_3369);
and U7383 (N_7383,N_3598,N_2781);
or U7384 (N_7384,N_2283,N_2688);
nor U7385 (N_7385,N_3411,N_2193);
nor U7386 (N_7386,N_4657,N_2968);
or U7387 (N_7387,N_333,N_1299);
and U7388 (N_7388,N_3266,N_1453);
and U7389 (N_7389,N_4422,N_4772);
nand U7390 (N_7390,N_4294,N_1028);
nand U7391 (N_7391,N_1118,N_4917);
and U7392 (N_7392,N_1620,N_1806);
nor U7393 (N_7393,N_2162,N_3012);
or U7394 (N_7394,N_2215,N_1412);
nor U7395 (N_7395,N_2197,N_2182);
nand U7396 (N_7396,N_3756,N_2057);
nand U7397 (N_7397,N_2329,N_1304);
or U7398 (N_7398,N_4760,N_272);
and U7399 (N_7399,N_4243,N_4581);
nand U7400 (N_7400,N_4891,N_3687);
and U7401 (N_7401,N_4089,N_4606);
and U7402 (N_7402,N_4692,N_2321);
nand U7403 (N_7403,N_2398,N_4501);
nand U7404 (N_7404,N_1682,N_4486);
nor U7405 (N_7405,N_3344,N_863);
nand U7406 (N_7406,N_2069,N_4972);
or U7407 (N_7407,N_2488,N_93);
or U7408 (N_7408,N_1261,N_2824);
nor U7409 (N_7409,N_715,N_1187);
nor U7410 (N_7410,N_388,N_1532);
or U7411 (N_7411,N_3291,N_665);
nand U7412 (N_7412,N_3315,N_4837);
nor U7413 (N_7413,N_2529,N_4438);
nand U7414 (N_7414,N_1233,N_2177);
nand U7415 (N_7415,N_4649,N_1994);
and U7416 (N_7416,N_604,N_1724);
or U7417 (N_7417,N_4388,N_4589);
nor U7418 (N_7418,N_1918,N_3847);
and U7419 (N_7419,N_1107,N_4221);
nand U7420 (N_7420,N_3579,N_2448);
and U7421 (N_7421,N_538,N_921);
nand U7422 (N_7422,N_3357,N_787);
or U7423 (N_7423,N_1283,N_1219);
or U7424 (N_7424,N_3643,N_1733);
nand U7425 (N_7425,N_1565,N_3426);
nand U7426 (N_7426,N_2331,N_137);
or U7427 (N_7427,N_69,N_1665);
and U7428 (N_7428,N_4913,N_4734);
and U7429 (N_7429,N_1739,N_2500);
or U7430 (N_7430,N_1476,N_2793);
nor U7431 (N_7431,N_4523,N_4662);
and U7432 (N_7432,N_1863,N_3319);
nand U7433 (N_7433,N_3961,N_3464);
nor U7434 (N_7434,N_1715,N_2669);
nand U7435 (N_7435,N_669,N_3399);
nor U7436 (N_7436,N_3022,N_1086);
or U7437 (N_7437,N_2672,N_2471);
nor U7438 (N_7438,N_990,N_1443);
nand U7439 (N_7439,N_4066,N_2191);
or U7440 (N_7440,N_447,N_4585);
nand U7441 (N_7441,N_3774,N_3877);
nor U7442 (N_7442,N_2223,N_3753);
and U7443 (N_7443,N_4795,N_1096);
or U7444 (N_7444,N_4383,N_616);
and U7445 (N_7445,N_3385,N_4910);
and U7446 (N_7446,N_3349,N_4302);
nand U7447 (N_7447,N_3843,N_1874);
or U7448 (N_7448,N_2525,N_4929);
nor U7449 (N_7449,N_1228,N_4822);
and U7450 (N_7450,N_1392,N_2706);
xnor U7451 (N_7451,N_4863,N_4971);
or U7452 (N_7452,N_1480,N_4160);
nor U7453 (N_7453,N_4652,N_823);
or U7454 (N_7454,N_8,N_4130);
nand U7455 (N_7455,N_1209,N_1655);
or U7456 (N_7456,N_1548,N_2341);
or U7457 (N_7457,N_3566,N_2492);
or U7458 (N_7458,N_3972,N_2101);
nor U7459 (N_7459,N_1915,N_4674);
nand U7460 (N_7460,N_1601,N_2270);
nand U7461 (N_7461,N_4757,N_2703);
nand U7462 (N_7462,N_1323,N_1407);
nor U7463 (N_7463,N_2938,N_2334);
and U7464 (N_7464,N_4275,N_2856);
nand U7465 (N_7465,N_2231,N_1054);
or U7466 (N_7466,N_3274,N_277);
nor U7467 (N_7467,N_2212,N_2371);
nand U7468 (N_7468,N_4931,N_1726);
nand U7469 (N_7469,N_1255,N_460);
and U7470 (N_7470,N_2517,N_1069);
and U7471 (N_7471,N_3,N_3173);
or U7472 (N_7472,N_1833,N_1969);
nand U7473 (N_7473,N_1285,N_4515);
and U7474 (N_7474,N_2919,N_2274);
nor U7475 (N_7475,N_3230,N_2438);
nor U7476 (N_7476,N_3286,N_4154);
or U7477 (N_7477,N_1598,N_3849);
or U7478 (N_7478,N_2927,N_17);
or U7479 (N_7479,N_1843,N_3133);
xnor U7480 (N_7480,N_4597,N_2040);
nand U7481 (N_7481,N_2986,N_1211);
nor U7482 (N_7482,N_1311,N_1116);
or U7483 (N_7483,N_1100,N_4851);
or U7484 (N_7484,N_2686,N_2727);
nor U7485 (N_7485,N_357,N_2712);
nor U7486 (N_7486,N_1838,N_4);
nand U7487 (N_7487,N_1946,N_1752);
nand U7488 (N_7488,N_523,N_4116);
or U7489 (N_7489,N_1496,N_248);
or U7490 (N_7490,N_3297,N_3835);
or U7491 (N_7491,N_291,N_1828);
and U7492 (N_7492,N_995,N_3740);
xor U7493 (N_7493,N_4410,N_4399);
or U7494 (N_7494,N_4812,N_454);
nand U7495 (N_7495,N_2739,N_756);
nand U7496 (N_7496,N_2226,N_3167);
and U7497 (N_7497,N_2608,N_3047);
nand U7498 (N_7498,N_3105,N_274);
and U7499 (N_7499,N_4900,N_4796);
nand U7500 (N_7500,N_395,N_959);
nand U7501 (N_7501,N_3825,N_2243);
or U7502 (N_7502,N_44,N_4095);
nor U7503 (N_7503,N_3081,N_1907);
or U7504 (N_7504,N_4889,N_3984);
nor U7505 (N_7505,N_1471,N_654);
or U7506 (N_7506,N_2331,N_4943);
nand U7507 (N_7507,N_2178,N_2697);
and U7508 (N_7508,N_3671,N_304);
and U7509 (N_7509,N_842,N_2729);
and U7510 (N_7510,N_840,N_1801);
nand U7511 (N_7511,N_254,N_3911);
and U7512 (N_7512,N_3187,N_1278);
or U7513 (N_7513,N_2260,N_1895);
or U7514 (N_7514,N_2547,N_3586);
nand U7515 (N_7515,N_3221,N_1201);
nor U7516 (N_7516,N_4855,N_3903);
nand U7517 (N_7517,N_582,N_4378);
nand U7518 (N_7518,N_3064,N_77);
and U7519 (N_7519,N_3707,N_3629);
nand U7520 (N_7520,N_634,N_3266);
nor U7521 (N_7521,N_3630,N_4158);
or U7522 (N_7522,N_102,N_2138);
nor U7523 (N_7523,N_3709,N_4399);
or U7524 (N_7524,N_2983,N_3110);
or U7525 (N_7525,N_2047,N_1351);
nor U7526 (N_7526,N_1039,N_155);
nand U7527 (N_7527,N_4086,N_3075);
nor U7528 (N_7528,N_4472,N_3721);
and U7529 (N_7529,N_4838,N_2418);
nand U7530 (N_7530,N_4512,N_186);
nor U7531 (N_7531,N_3092,N_1578);
and U7532 (N_7532,N_4087,N_97);
and U7533 (N_7533,N_853,N_1377);
or U7534 (N_7534,N_4882,N_2892);
or U7535 (N_7535,N_3449,N_3600);
nand U7536 (N_7536,N_4930,N_907);
nor U7537 (N_7537,N_2277,N_1738);
nand U7538 (N_7538,N_4888,N_1055);
nor U7539 (N_7539,N_4415,N_4825);
nand U7540 (N_7540,N_1701,N_564);
nand U7541 (N_7541,N_1315,N_2304);
and U7542 (N_7542,N_4877,N_1826);
or U7543 (N_7543,N_2046,N_3158);
nand U7544 (N_7544,N_3270,N_4678);
or U7545 (N_7545,N_4428,N_1033);
or U7546 (N_7546,N_515,N_729);
nand U7547 (N_7547,N_541,N_1188);
and U7548 (N_7548,N_3654,N_507);
nor U7549 (N_7549,N_3709,N_440);
and U7550 (N_7550,N_917,N_2530);
and U7551 (N_7551,N_512,N_1848);
xnor U7552 (N_7552,N_1391,N_3631);
nand U7553 (N_7553,N_2337,N_1239);
and U7554 (N_7554,N_1112,N_4904);
or U7555 (N_7555,N_154,N_2439);
and U7556 (N_7556,N_4769,N_57);
or U7557 (N_7557,N_4038,N_3258);
nand U7558 (N_7558,N_1388,N_2341);
nor U7559 (N_7559,N_2028,N_4426);
nand U7560 (N_7560,N_590,N_3692);
and U7561 (N_7561,N_1921,N_1808);
xnor U7562 (N_7562,N_4504,N_227);
and U7563 (N_7563,N_1638,N_705);
or U7564 (N_7564,N_977,N_2406);
nor U7565 (N_7565,N_4138,N_4518);
and U7566 (N_7566,N_4095,N_1294);
nand U7567 (N_7567,N_4547,N_1428);
nand U7568 (N_7568,N_3696,N_4065);
nand U7569 (N_7569,N_1173,N_1233);
and U7570 (N_7570,N_2374,N_454);
and U7571 (N_7571,N_658,N_4873);
nor U7572 (N_7572,N_4422,N_4387);
or U7573 (N_7573,N_909,N_835);
or U7574 (N_7574,N_1750,N_188);
and U7575 (N_7575,N_1332,N_3165);
nand U7576 (N_7576,N_1139,N_4724);
or U7577 (N_7577,N_2902,N_2719);
nand U7578 (N_7578,N_3391,N_77);
nand U7579 (N_7579,N_3410,N_3161);
nand U7580 (N_7580,N_2269,N_3635);
or U7581 (N_7581,N_3119,N_735);
or U7582 (N_7582,N_3107,N_134);
xnor U7583 (N_7583,N_2262,N_4980);
nand U7584 (N_7584,N_4021,N_1274);
or U7585 (N_7585,N_1008,N_2409);
nor U7586 (N_7586,N_1470,N_2132);
nor U7587 (N_7587,N_3248,N_4831);
and U7588 (N_7588,N_4986,N_561);
and U7589 (N_7589,N_3949,N_3208);
nor U7590 (N_7590,N_547,N_4888);
or U7591 (N_7591,N_2642,N_509);
and U7592 (N_7592,N_1137,N_469);
nor U7593 (N_7593,N_2323,N_4710);
and U7594 (N_7594,N_2503,N_3955);
or U7595 (N_7595,N_3593,N_1832);
nor U7596 (N_7596,N_3471,N_437);
nand U7597 (N_7597,N_366,N_1188);
nor U7598 (N_7598,N_280,N_1204);
nand U7599 (N_7599,N_1287,N_928);
xnor U7600 (N_7600,N_4938,N_303);
or U7601 (N_7601,N_1673,N_2919);
and U7602 (N_7602,N_1814,N_2285);
nor U7603 (N_7603,N_1658,N_2293);
nand U7604 (N_7604,N_2001,N_4311);
or U7605 (N_7605,N_296,N_1365);
nand U7606 (N_7606,N_3513,N_4622);
nor U7607 (N_7607,N_1938,N_4485);
and U7608 (N_7608,N_2579,N_1399);
nand U7609 (N_7609,N_4107,N_4381);
nand U7610 (N_7610,N_2980,N_1014);
nor U7611 (N_7611,N_3683,N_1010);
and U7612 (N_7612,N_875,N_2880);
nand U7613 (N_7613,N_295,N_3007);
nand U7614 (N_7614,N_1885,N_1783);
and U7615 (N_7615,N_1040,N_767);
nor U7616 (N_7616,N_3178,N_4719);
nand U7617 (N_7617,N_1226,N_1522);
nand U7618 (N_7618,N_1662,N_1900);
or U7619 (N_7619,N_4452,N_717);
nor U7620 (N_7620,N_3821,N_4132);
and U7621 (N_7621,N_3077,N_2206);
or U7622 (N_7622,N_1762,N_1026);
nor U7623 (N_7623,N_3263,N_2479);
or U7624 (N_7624,N_397,N_4082);
or U7625 (N_7625,N_1918,N_1082);
nor U7626 (N_7626,N_588,N_3564);
and U7627 (N_7627,N_3012,N_2497);
or U7628 (N_7628,N_1277,N_2231);
xor U7629 (N_7629,N_2758,N_1651);
or U7630 (N_7630,N_2654,N_3359);
nand U7631 (N_7631,N_4418,N_1181);
and U7632 (N_7632,N_951,N_931);
and U7633 (N_7633,N_2414,N_3859);
or U7634 (N_7634,N_3605,N_3741);
and U7635 (N_7635,N_4583,N_3936);
and U7636 (N_7636,N_2729,N_2234);
nor U7637 (N_7637,N_3597,N_3943);
nor U7638 (N_7638,N_2133,N_3292);
and U7639 (N_7639,N_4932,N_4293);
nand U7640 (N_7640,N_1111,N_368);
nor U7641 (N_7641,N_1469,N_374);
and U7642 (N_7642,N_3391,N_3454);
nand U7643 (N_7643,N_3484,N_1031);
nor U7644 (N_7644,N_3803,N_303);
or U7645 (N_7645,N_4979,N_12);
and U7646 (N_7646,N_4289,N_1294);
or U7647 (N_7647,N_4563,N_4386);
nand U7648 (N_7648,N_3144,N_4631);
nor U7649 (N_7649,N_3372,N_1888);
or U7650 (N_7650,N_3414,N_627);
nand U7651 (N_7651,N_4689,N_2794);
nor U7652 (N_7652,N_2435,N_2252);
nand U7653 (N_7653,N_2740,N_1792);
nand U7654 (N_7654,N_4494,N_606);
xor U7655 (N_7655,N_2300,N_3409);
and U7656 (N_7656,N_4710,N_846);
nand U7657 (N_7657,N_1296,N_3359);
nor U7658 (N_7658,N_486,N_4818);
and U7659 (N_7659,N_813,N_2631);
nand U7660 (N_7660,N_274,N_1479);
nand U7661 (N_7661,N_3532,N_3081);
nand U7662 (N_7662,N_2431,N_1715);
and U7663 (N_7663,N_3774,N_4904);
nand U7664 (N_7664,N_3511,N_1178);
nand U7665 (N_7665,N_2483,N_2896);
nand U7666 (N_7666,N_4227,N_4756);
nand U7667 (N_7667,N_724,N_728);
nand U7668 (N_7668,N_4435,N_3772);
nor U7669 (N_7669,N_1955,N_3471);
and U7670 (N_7670,N_2364,N_4832);
or U7671 (N_7671,N_1140,N_3771);
or U7672 (N_7672,N_4526,N_2898);
and U7673 (N_7673,N_4445,N_1140);
or U7674 (N_7674,N_2318,N_3198);
and U7675 (N_7675,N_1960,N_3155);
nor U7676 (N_7676,N_685,N_2729);
or U7677 (N_7677,N_1514,N_3123);
nor U7678 (N_7678,N_4310,N_3810);
or U7679 (N_7679,N_3087,N_1079);
or U7680 (N_7680,N_3366,N_1506);
or U7681 (N_7681,N_4478,N_1521);
and U7682 (N_7682,N_665,N_298);
and U7683 (N_7683,N_1085,N_4625);
and U7684 (N_7684,N_1332,N_4270);
xor U7685 (N_7685,N_1930,N_148);
nand U7686 (N_7686,N_1024,N_4220);
and U7687 (N_7687,N_2812,N_4822);
nor U7688 (N_7688,N_3253,N_4670);
nand U7689 (N_7689,N_30,N_2182);
nand U7690 (N_7690,N_1539,N_95);
nor U7691 (N_7691,N_2696,N_989);
nor U7692 (N_7692,N_3929,N_1949);
and U7693 (N_7693,N_2023,N_1322);
or U7694 (N_7694,N_2936,N_1969);
and U7695 (N_7695,N_1260,N_4030);
or U7696 (N_7696,N_4885,N_3016);
and U7697 (N_7697,N_2031,N_4157);
nor U7698 (N_7698,N_1667,N_2484);
nor U7699 (N_7699,N_997,N_905);
nor U7700 (N_7700,N_4181,N_6);
or U7701 (N_7701,N_3965,N_2372);
nand U7702 (N_7702,N_1304,N_4167);
nand U7703 (N_7703,N_3518,N_4274);
or U7704 (N_7704,N_70,N_778);
and U7705 (N_7705,N_3924,N_236);
and U7706 (N_7706,N_614,N_1782);
nand U7707 (N_7707,N_2490,N_2198);
and U7708 (N_7708,N_1346,N_3703);
nand U7709 (N_7709,N_4550,N_346);
or U7710 (N_7710,N_2701,N_4201);
or U7711 (N_7711,N_4430,N_4062);
and U7712 (N_7712,N_4331,N_3109);
or U7713 (N_7713,N_458,N_1804);
nand U7714 (N_7714,N_1792,N_4626);
nor U7715 (N_7715,N_3746,N_2598);
or U7716 (N_7716,N_1684,N_1208);
nand U7717 (N_7717,N_2835,N_3656);
nor U7718 (N_7718,N_1096,N_13);
nor U7719 (N_7719,N_409,N_1254);
xnor U7720 (N_7720,N_927,N_353);
nand U7721 (N_7721,N_745,N_2747);
or U7722 (N_7722,N_1783,N_3487);
nand U7723 (N_7723,N_4711,N_2207);
nand U7724 (N_7724,N_3668,N_4377);
and U7725 (N_7725,N_2286,N_4372);
or U7726 (N_7726,N_308,N_4584);
nor U7727 (N_7727,N_229,N_1623);
nand U7728 (N_7728,N_3655,N_3708);
or U7729 (N_7729,N_2788,N_3512);
and U7730 (N_7730,N_3559,N_3358);
nand U7731 (N_7731,N_3595,N_1506);
nand U7732 (N_7732,N_276,N_4394);
nand U7733 (N_7733,N_3711,N_957);
nand U7734 (N_7734,N_3272,N_3071);
nand U7735 (N_7735,N_3514,N_3891);
or U7736 (N_7736,N_2870,N_3515);
nand U7737 (N_7737,N_1336,N_2016);
or U7738 (N_7738,N_2287,N_2317);
or U7739 (N_7739,N_44,N_3609);
nor U7740 (N_7740,N_4639,N_4138);
nand U7741 (N_7741,N_2375,N_4529);
or U7742 (N_7742,N_3866,N_1298);
and U7743 (N_7743,N_3130,N_4613);
xor U7744 (N_7744,N_4765,N_1689);
nand U7745 (N_7745,N_1507,N_2879);
nand U7746 (N_7746,N_1869,N_994);
or U7747 (N_7747,N_637,N_1901);
nor U7748 (N_7748,N_343,N_1044);
nand U7749 (N_7749,N_173,N_1845);
or U7750 (N_7750,N_1884,N_3527);
and U7751 (N_7751,N_1202,N_4730);
nand U7752 (N_7752,N_1715,N_4145);
nor U7753 (N_7753,N_1235,N_4420);
nand U7754 (N_7754,N_3597,N_3323);
or U7755 (N_7755,N_4682,N_3824);
and U7756 (N_7756,N_563,N_3195);
or U7757 (N_7757,N_4012,N_1719);
nor U7758 (N_7758,N_2136,N_2379);
nand U7759 (N_7759,N_314,N_1647);
and U7760 (N_7760,N_4638,N_2746);
nand U7761 (N_7761,N_971,N_3325);
or U7762 (N_7762,N_1007,N_2157);
and U7763 (N_7763,N_4594,N_457);
and U7764 (N_7764,N_4321,N_3888);
or U7765 (N_7765,N_66,N_3615);
or U7766 (N_7766,N_2385,N_4368);
and U7767 (N_7767,N_2820,N_4446);
nor U7768 (N_7768,N_2147,N_4227);
nor U7769 (N_7769,N_1033,N_1127);
nor U7770 (N_7770,N_4817,N_2995);
and U7771 (N_7771,N_93,N_3490);
and U7772 (N_7772,N_2006,N_4736);
and U7773 (N_7773,N_315,N_4275);
nor U7774 (N_7774,N_1294,N_881);
and U7775 (N_7775,N_3157,N_2512);
or U7776 (N_7776,N_1091,N_2449);
nor U7777 (N_7777,N_3895,N_2989);
nor U7778 (N_7778,N_3438,N_3169);
nor U7779 (N_7779,N_737,N_575);
and U7780 (N_7780,N_3137,N_2858);
nand U7781 (N_7781,N_2671,N_850);
and U7782 (N_7782,N_4635,N_920);
nor U7783 (N_7783,N_4632,N_1562);
or U7784 (N_7784,N_3692,N_4803);
nand U7785 (N_7785,N_785,N_1154);
nand U7786 (N_7786,N_4233,N_684);
and U7787 (N_7787,N_3464,N_4874);
nor U7788 (N_7788,N_4863,N_3717);
nand U7789 (N_7789,N_1851,N_4026);
or U7790 (N_7790,N_1540,N_573);
and U7791 (N_7791,N_4374,N_3995);
or U7792 (N_7792,N_660,N_339);
nor U7793 (N_7793,N_859,N_3222);
and U7794 (N_7794,N_876,N_2608);
nand U7795 (N_7795,N_1932,N_2025);
and U7796 (N_7796,N_1782,N_4630);
or U7797 (N_7797,N_4436,N_2199);
or U7798 (N_7798,N_255,N_3653);
nor U7799 (N_7799,N_4342,N_758);
or U7800 (N_7800,N_686,N_587);
nor U7801 (N_7801,N_2364,N_3891);
nor U7802 (N_7802,N_1132,N_2976);
or U7803 (N_7803,N_1366,N_1362);
nor U7804 (N_7804,N_1279,N_1819);
nor U7805 (N_7805,N_639,N_626);
nand U7806 (N_7806,N_4047,N_2164);
nand U7807 (N_7807,N_1715,N_2769);
nand U7808 (N_7808,N_3752,N_3562);
and U7809 (N_7809,N_2290,N_674);
nand U7810 (N_7810,N_3638,N_683);
nor U7811 (N_7811,N_445,N_440);
and U7812 (N_7812,N_4936,N_2830);
nand U7813 (N_7813,N_4454,N_1760);
or U7814 (N_7814,N_101,N_987);
or U7815 (N_7815,N_4329,N_1196);
nor U7816 (N_7816,N_1000,N_3520);
or U7817 (N_7817,N_4457,N_1963);
nand U7818 (N_7818,N_4175,N_4017);
nand U7819 (N_7819,N_3319,N_26);
or U7820 (N_7820,N_2627,N_1671);
nand U7821 (N_7821,N_4226,N_3221);
nand U7822 (N_7822,N_3744,N_354);
nor U7823 (N_7823,N_2034,N_742);
and U7824 (N_7824,N_3609,N_1010);
nor U7825 (N_7825,N_3837,N_1674);
nand U7826 (N_7826,N_661,N_3863);
and U7827 (N_7827,N_4748,N_1205);
nor U7828 (N_7828,N_1142,N_825);
and U7829 (N_7829,N_366,N_1925);
or U7830 (N_7830,N_2859,N_1573);
and U7831 (N_7831,N_2856,N_3085);
nand U7832 (N_7832,N_3765,N_2169);
or U7833 (N_7833,N_4062,N_1788);
nor U7834 (N_7834,N_3649,N_743);
nor U7835 (N_7835,N_1344,N_4690);
xor U7836 (N_7836,N_4953,N_4436);
and U7837 (N_7837,N_977,N_3256);
and U7838 (N_7838,N_2322,N_2698);
nor U7839 (N_7839,N_3355,N_620);
nand U7840 (N_7840,N_131,N_1525);
nor U7841 (N_7841,N_3237,N_4005);
and U7842 (N_7842,N_4253,N_451);
nand U7843 (N_7843,N_4627,N_1587);
nor U7844 (N_7844,N_3051,N_3022);
or U7845 (N_7845,N_1796,N_17);
nand U7846 (N_7846,N_1780,N_2675);
nand U7847 (N_7847,N_3869,N_2033);
nor U7848 (N_7848,N_110,N_459);
or U7849 (N_7849,N_4676,N_2265);
and U7850 (N_7850,N_2262,N_3210);
nor U7851 (N_7851,N_1764,N_461);
or U7852 (N_7852,N_1161,N_3279);
and U7853 (N_7853,N_236,N_3282);
nor U7854 (N_7854,N_2760,N_3219);
or U7855 (N_7855,N_613,N_4377);
or U7856 (N_7856,N_570,N_3108);
and U7857 (N_7857,N_2907,N_1755);
and U7858 (N_7858,N_1843,N_3615);
nand U7859 (N_7859,N_4351,N_3010);
or U7860 (N_7860,N_3369,N_305);
and U7861 (N_7861,N_583,N_3452);
and U7862 (N_7862,N_2446,N_1505);
nand U7863 (N_7863,N_4688,N_3503);
nor U7864 (N_7864,N_4383,N_525);
or U7865 (N_7865,N_2386,N_4737);
or U7866 (N_7866,N_4085,N_3110);
and U7867 (N_7867,N_467,N_2940);
and U7868 (N_7868,N_4132,N_1682);
or U7869 (N_7869,N_261,N_4319);
nand U7870 (N_7870,N_19,N_2819);
nor U7871 (N_7871,N_289,N_4565);
nand U7872 (N_7872,N_3690,N_1272);
nand U7873 (N_7873,N_3017,N_1201);
and U7874 (N_7874,N_1518,N_1138);
or U7875 (N_7875,N_2764,N_3708);
nand U7876 (N_7876,N_3137,N_2285);
and U7877 (N_7877,N_3607,N_1545);
or U7878 (N_7878,N_2255,N_3468);
nand U7879 (N_7879,N_1345,N_3513);
or U7880 (N_7880,N_1153,N_2041);
nand U7881 (N_7881,N_685,N_655);
or U7882 (N_7882,N_2696,N_4930);
and U7883 (N_7883,N_3158,N_4733);
nor U7884 (N_7884,N_4458,N_3010);
nand U7885 (N_7885,N_4478,N_385);
nand U7886 (N_7886,N_4631,N_2874);
nor U7887 (N_7887,N_3225,N_904);
nand U7888 (N_7888,N_4120,N_3285);
and U7889 (N_7889,N_888,N_4363);
nor U7890 (N_7890,N_418,N_1740);
nor U7891 (N_7891,N_4338,N_3120);
or U7892 (N_7892,N_4624,N_4837);
or U7893 (N_7893,N_3802,N_2551);
or U7894 (N_7894,N_829,N_194);
nand U7895 (N_7895,N_492,N_2566);
nor U7896 (N_7896,N_1677,N_4405);
and U7897 (N_7897,N_3430,N_815);
or U7898 (N_7898,N_3140,N_889);
or U7899 (N_7899,N_1612,N_3887);
nand U7900 (N_7900,N_4196,N_829);
nor U7901 (N_7901,N_4145,N_4706);
and U7902 (N_7902,N_3452,N_1101);
nor U7903 (N_7903,N_2262,N_1291);
nor U7904 (N_7904,N_3351,N_3796);
nor U7905 (N_7905,N_153,N_242);
nand U7906 (N_7906,N_4107,N_1542);
nor U7907 (N_7907,N_1913,N_520);
and U7908 (N_7908,N_3891,N_1703);
nor U7909 (N_7909,N_1570,N_3161);
and U7910 (N_7910,N_4831,N_2994);
nand U7911 (N_7911,N_1528,N_3832);
nand U7912 (N_7912,N_2869,N_4855);
or U7913 (N_7913,N_3214,N_3377);
nor U7914 (N_7914,N_1354,N_1191);
nor U7915 (N_7915,N_4362,N_3166);
or U7916 (N_7916,N_3468,N_218);
or U7917 (N_7917,N_2435,N_3230);
and U7918 (N_7918,N_998,N_1228);
or U7919 (N_7919,N_1161,N_3002);
nor U7920 (N_7920,N_27,N_294);
nand U7921 (N_7921,N_2162,N_519);
nand U7922 (N_7922,N_2793,N_4413);
nor U7923 (N_7923,N_1693,N_1003);
nor U7924 (N_7924,N_1497,N_2807);
nor U7925 (N_7925,N_4545,N_2470);
or U7926 (N_7926,N_22,N_621);
nand U7927 (N_7927,N_3193,N_1377);
and U7928 (N_7928,N_1258,N_4227);
or U7929 (N_7929,N_206,N_3052);
or U7930 (N_7930,N_2466,N_2379);
and U7931 (N_7931,N_867,N_662);
nand U7932 (N_7932,N_4156,N_3653);
xnor U7933 (N_7933,N_1038,N_3183);
and U7934 (N_7934,N_2406,N_192);
nor U7935 (N_7935,N_4897,N_1687);
nor U7936 (N_7936,N_1471,N_776);
nand U7937 (N_7937,N_793,N_3506);
nor U7938 (N_7938,N_734,N_1017);
nor U7939 (N_7939,N_1188,N_2688);
and U7940 (N_7940,N_4551,N_1558);
or U7941 (N_7941,N_4438,N_4354);
and U7942 (N_7942,N_2615,N_4119);
nor U7943 (N_7943,N_725,N_993);
nand U7944 (N_7944,N_959,N_2775);
and U7945 (N_7945,N_4278,N_1661);
nor U7946 (N_7946,N_3111,N_4809);
and U7947 (N_7947,N_4742,N_480);
and U7948 (N_7948,N_2302,N_3137);
nor U7949 (N_7949,N_2699,N_1079);
nand U7950 (N_7950,N_722,N_4995);
nor U7951 (N_7951,N_46,N_4915);
nor U7952 (N_7952,N_1727,N_3294);
nor U7953 (N_7953,N_196,N_3336);
or U7954 (N_7954,N_4692,N_341);
or U7955 (N_7955,N_3229,N_4549);
or U7956 (N_7956,N_698,N_3772);
and U7957 (N_7957,N_3051,N_4398);
nor U7958 (N_7958,N_3197,N_2399);
and U7959 (N_7959,N_1078,N_3707);
or U7960 (N_7960,N_4353,N_4165);
or U7961 (N_7961,N_4781,N_2604);
and U7962 (N_7962,N_4797,N_2262);
nand U7963 (N_7963,N_1577,N_29);
or U7964 (N_7964,N_2174,N_1779);
and U7965 (N_7965,N_4885,N_2727);
and U7966 (N_7966,N_1505,N_219);
nor U7967 (N_7967,N_94,N_4169);
and U7968 (N_7968,N_1264,N_3100);
or U7969 (N_7969,N_4438,N_4950);
and U7970 (N_7970,N_2608,N_3191);
nand U7971 (N_7971,N_1865,N_4380);
nor U7972 (N_7972,N_911,N_88);
and U7973 (N_7973,N_3336,N_2041);
nor U7974 (N_7974,N_3719,N_2051);
nor U7975 (N_7975,N_1024,N_3759);
nand U7976 (N_7976,N_2791,N_301);
nand U7977 (N_7977,N_446,N_1306);
or U7978 (N_7978,N_364,N_2293);
and U7979 (N_7979,N_2807,N_4711);
or U7980 (N_7980,N_4528,N_2128);
or U7981 (N_7981,N_4723,N_4733);
or U7982 (N_7982,N_1039,N_3577);
and U7983 (N_7983,N_687,N_4304);
and U7984 (N_7984,N_311,N_2823);
and U7985 (N_7985,N_2857,N_1192);
or U7986 (N_7986,N_2480,N_3419);
nor U7987 (N_7987,N_1447,N_1729);
nor U7988 (N_7988,N_3645,N_1632);
nor U7989 (N_7989,N_4791,N_4046);
or U7990 (N_7990,N_3492,N_3265);
and U7991 (N_7991,N_1584,N_2509);
and U7992 (N_7992,N_4133,N_3197);
nand U7993 (N_7993,N_3518,N_363);
or U7994 (N_7994,N_185,N_1580);
or U7995 (N_7995,N_999,N_3683);
nand U7996 (N_7996,N_2872,N_615);
or U7997 (N_7997,N_3768,N_3802);
nand U7998 (N_7998,N_3330,N_507);
nor U7999 (N_7999,N_4554,N_3223);
or U8000 (N_8000,N_4590,N_3752);
nor U8001 (N_8001,N_2595,N_3301);
nor U8002 (N_8002,N_442,N_233);
nand U8003 (N_8003,N_3990,N_2214);
and U8004 (N_8004,N_4129,N_2847);
nand U8005 (N_8005,N_3635,N_2272);
nor U8006 (N_8006,N_3264,N_4381);
or U8007 (N_8007,N_4431,N_3797);
or U8008 (N_8008,N_2186,N_2506);
nand U8009 (N_8009,N_3722,N_1907);
or U8010 (N_8010,N_1915,N_2169);
nor U8011 (N_8011,N_1211,N_3164);
nand U8012 (N_8012,N_2063,N_4023);
or U8013 (N_8013,N_1336,N_2099);
xor U8014 (N_8014,N_3422,N_3345);
nor U8015 (N_8015,N_1215,N_2462);
or U8016 (N_8016,N_2796,N_4476);
or U8017 (N_8017,N_3459,N_2489);
or U8018 (N_8018,N_202,N_3230);
nor U8019 (N_8019,N_2130,N_1647);
nand U8020 (N_8020,N_2589,N_4722);
nor U8021 (N_8021,N_184,N_3737);
or U8022 (N_8022,N_2613,N_1778);
or U8023 (N_8023,N_2941,N_1807);
nand U8024 (N_8024,N_1728,N_4505);
nor U8025 (N_8025,N_441,N_1582);
or U8026 (N_8026,N_3802,N_4303);
xnor U8027 (N_8027,N_1786,N_1482);
xor U8028 (N_8028,N_1753,N_1828);
nand U8029 (N_8029,N_3745,N_1749);
nor U8030 (N_8030,N_2463,N_2764);
nand U8031 (N_8031,N_4853,N_620);
or U8032 (N_8032,N_4873,N_141);
nand U8033 (N_8033,N_1650,N_4439);
and U8034 (N_8034,N_1055,N_2065);
nor U8035 (N_8035,N_3492,N_1837);
and U8036 (N_8036,N_2499,N_880);
nor U8037 (N_8037,N_345,N_4057);
and U8038 (N_8038,N_2570,N_2142);
nor U8039 (N_8039,N_297,N_2976);
nand U8040 (N_8040,N_147,N_2181);
and U8041 (N_8041,N_2529,N_2870);
or U8042 (N_8042,N_1436,N_4681);
nand U8043 (N_8043,N_3906,N_1281);
nand U8044 (N_8044,N_2907,N_4996);
nand U8045 (N_8045,N_4066,N_4887);
nor U8046 (N_8046,N_785,N_2801);
and U8047 (N_8047,N_1079,N_2416);
nor U8048 (N_8048,N_4510,N_3869);
and U8049 (N_8049,N_4595,N_200);
nand U8050 (N_8050,N_4838,N_4433);
nor U8051 (N_8051,N_3900,N_4073);
nor U8052 (N_8052,N_2669,N_4095);
nor U8053 (N_8053,N_3147,N_4285);
nand U8054 (N_8054,N_3655,N_751);
nand U8055 (N_8055,N_2781,N_2818);
or U8056 (N_8056,N_1031,N_3717);
nand U8057 (N_8057,N_1164,N_3481);
and U8058 (N_8058,N_3552,N_298);
and U8059 (N_8059,N_500,N_520);
or U8060 (N_8060,N_482,N_267);
and U8061 (N_8061,N_2588,N_4620);
and U8062 (N_8062,N_235,N_1380);
and U8063 (N_8063,N_4472,N_3091);
or U8064 (N_8064,N_422,N_1798);
and U8065 (N_8065,N_674,N_265);
and U8066 (N_8066,N_2787,N_4034);
and U8067 (N_8067,N_3046,N_3578);
and U8068 (N_8068,N_4399,N_1307);
nand U8069 (N_8069,N_2036,N_1631);
or U8070 (N_8070,N_3320,N_1680);
xnor U8071 (N_8071,N_3899,N_1922);
nand U8072 (N_8072,N_4264,N_1184);
nor U8073 (N_8073,N_434,N_2711);
and U8074 (N_8074,N_1794,N_2949);
and U8075 (N_8075,N_2338,N_4709);
nor U8076 (N_8076,N_1406,N_1914);
or U8077 (N_8077,N_4484,N_4917);
nor U8078 (N_8078,N_3410,N_304);
nand U8079 (N_8079,N_2475,N_3708);
and U8080 (N_8080,N_58,N_1410);
and U8081 (N_8081,N_4039,N_2989);
and U8082 (N_8082,N_4988,N_828);
and U8083 (N_8083,N_4341,N_4818);
and U8084 (N_8084,N_328,N_4909);
and U8085 (N_8085,N_2367,N_4851);
and U8086 (N_8086,N_3719,N_3343);
or U8087 (N_8087,N_2304,N_3060);
and U8088 (N_8088,N_3395,N_1194);
nand U8089 (N_8089,N_1842,N_1493);
nor U8090 (N_8090,N_1505,N_2524);
or U8091 (N_8091,N_204,N_184);
nor U8092 (N_8092,N_2021,N_1524);
nor U8093 (N_8093,N_2389,N_3154);
and U8094 (N_8094,N_4447,N_4107);
nor U8095 (N_8095,N_1737,N_1803);
and U8096 (N_8096,N_744,N_2709);
or U8097 (N_8097,N_2081,N_2408);
or U8098 (N_8098,N_4227,N_1562);
nand U8099 (N_8099,N_168,N_1737);
or U8100 (N_8100,N_1310,N_1939);
and U8101 (N_8101,N_1038,N_3035);
or U8102 (N_8102,N_1637,N_1840);
and U8103 (N_8103,N_2117,N_2490);
or U8104 (N_8104,N_2975,N_3816);
nor U8105 (N_8105,N_38,N_3971);
nand U8106 (N_8106,N_3583,N_1097);
nor U8107 (N_8107,N_710,N_1140);
nor U8108 (N_8108,N_3132,N_2038);
nand U8109 (N_8109,N_4467,N_4346);
and U8110 (N_8110,N_4605,N_2422);
nand U8111 (N_8111,N_494,N_599);
nor U8112 (N_8112,N_1585,N_3903);
nand U8113 (N_8113,N_2305,N_3007);
or U8114 (N_8114,N_4761,N_3896);
nand U8115 (N_8115,N_4806,N_4318);
nand U8116 (N_8116,N_2586,N_837);
nor U8117 (N_8117,N_37,N_4113);
or U8118 (N_8118,N_4333,N_1016);
nor U8119 (N_8119,N_2548,N_2965);
and U8120 (N_8120,N_834,N_16);
and U8121 (N_8121,N_2660,N_1014);
and U8122 (N_8122,N_4792,N_2186);
nor U8123 (N_8123,N_4924,N_4310);
and U8124 (N_8124,N_3705,N_258);
or U8125 (N_8125,N_3390,N_210);
nand U8126 (N_8126,N_1074,N_1623);
nand U8127 (N_8127,N_1658,N_801);
nor U8128 (N_8128,N_2859,N_122);
nand U8129 (N_8129,N_4306,N_4441);
nand U8130 (N_8130,N_1800,N_2808);
nor U8131 (N_8131,N_1497,N_2766);
nor U8132 (N_8132,N_3385,N_1162);
nor U8133 (N_8133,N_4903,N_1410);
nor U8134 (N_8134,N_4294,N_3804);
or U8135 (N_8135,N_3832,N_323);
nor U8136 (N_8136,N_3547,N_903);
and U8137 (N_8137,N_2650,N_2302);
or U8138 (N_8138,N_213,N_1958);
nor U8139 (N_8139,N_1644,N_2300);
and U8140 (N_8140,N_284,N_617);
and U8141 (N_8141,N_3184,N_1472);
or U8142 (N_8142,N_4030,N_2798);
nand U8143 (N_8143,N_2999,N_644);
and U8144 (N_8144,N_622,N_1281);
nand U8145 (N_8145,N_3532,N_313);
nand U8146 (N_8146,N_3189,N_3990);
or U8147 (N_8147,N_1581,N_2789);
nor U8148 (N_8148,N_3651,N_3422);
nor U8149 (N_8149,N_2364,N_2136);
nor U8150 (N_8150,N_1444,N_2521);
nor U8151 (N_8151,N_4714,N_516);
nand U8152 (N_8152,N_3468,N_2451);
and U8153 (N_8153,N_4920,N_2690);
or U8154 (N_8154,N_3780,N_1730);
nor U8155 (N_8155,N_2473,N_2465);
and U8156 (N_8156,N_4029,N_3192);
nand U8157 (N_8157,N_578,N_1728);
nand U8158 (N_8158,N_4315,N_699);
nand U8159 (N_8159,N_3692,N_511);
and U8160 (N_8160,N_4936,N_3318);
and U8161 (N_8161,N_1886,N_3078);
nand U8162 (N_8162,N_2611,N_4963);
nor U8163 (N_8163,N_1861,N_3489);
and U8164 (N_8164,N_2893,N_1950);
nor U8165 (N_8165,N_222,N_3266);
nand U8166 (N_8166,N_4301,N_2859);
nand U8167 (N_8167,N_4357,N_4957);
and U8168 (N_8168,N_40,N_2388);
nor U8169 (N_8169,N_4703,N_1208);
or U8170 (N_8170,N_3810,N_2223);
or U8171 (N_8171,N_4310,N_4783);
nand U8172 (N_8172,N_4164,N_2517);
nand U8173 (N_8173,N_13,N_4646);
and U8174 (N_8174,N_4682,N_4956);
or U8175 (N_8175,N_654,N_4225);
and U8176 (N_8176,N_1646,N_3544);
nor U8177 (N_8177,N_2673,N_302);
nand U8178 (N_8178,N_266,N_2179);
nand U8179 (N_8179,N_1649,N_4979);
or U8180 (N_8180,N_231,N_4644);
nand U8181 (N_8181,N_331,N_245);
nor U8182 (N_8182,N_1622,N_2237);
nor U8183 (N_8183,N_4984,N_4239);
or U8184 (N_8184,N_2327,N_3597);
nor U8185 (N_8185,N_628,N_59);
nor U8186 (N_8186,N_767,N_2456);
or U8187 (N_8187,N_3298,N_4764);
nand U8188 (N_8188,N_3427,N_3511);
or U8189 (N_8189,N_2540,N_662);
nor U8190 (N_8190,N_3573,N_126);
nand U8191 (N_8191,N_444,N_906);
nand U8192 (N_8192,N_4801,N_621);
and U8193 (N_8193,N_2355,N_2695);
or U8194 (N_8194,N_4670,N_4083);
xnor U8195 (N_8195,N_772,N_429);
or U8196 (N_8196,N_3069,N_727);
and U8197 (N_8197,N_3955,N_173);
nand U8198 (N_8198,N_3105,N_4154);
nor U8199 (N_8199,N_4554,N_2232);
and U8200 (N_8200,N_768,N_2111);
and U8201 (N_8201,N_558,N_184);
or U8202 (N_8202,N_1657,N_665);
nor U8203 (N_8203,N_4301,N_1873);
nor U8204 (N_8204,N_4542,N_504);
nand U8205 (N_8205,N_3382,N_1088);
or U8206 (N_8206,N_4159,N_1781);
and U8207 (N_8207,N_4350,N_666);
nand U8208 (N_8208,N_1017,N_3168);
and U8209 (N_8209,N_334,N_1365);
and U8210 (N_8210,N_2934,N_1946);
and U8211 (N_8211,N_4844,N_909);
nor U8212 (N_8212,N_2107,N_2506);
nor U8213 (N_8213,N_4546,N_49);
and U8214 (N_8214,N_1330,N_3858);
nand U8215 (N_8215,N_756,N_3855);
nand U8216 (N_8216,N_2864,N_3996);
nor U8217 (N_8217,N_3141,N_1624);
nand U8218 (N_8218,N_1977,N_3986);
nand U8219 (N_8219,N_2048,N_1223);
or U8220 (N_8220,N_631,N_1761);
or U8221 (N_8221,N_364,N_2384);
nand U8222 (N_8222,N_4668,N_1991);
or U8223 (N_8223,N_724,N_3620);
or U8224 (N_8224,N_3029,N_1656);
nand U8225 (N_8225,N_4280,N_3231);
and U8226 (N_8226,N_2760,N_2254);
or U8227 (N_8227,N_997,N_3177);
nor U8228 (N_8228,N_4945,N_3901);
nand U8229 (N_8229,N_1106,N_1472);
nor U8230 (N_8230,N_4113,N_905);
and U8231 (N_8231,N_2016,N_278);
and U8232 (N_8232,N_184,N_2590);
and U8233 (N_8233,N_350,N_2280);
or U8234 (N_8234,N_1530,N_226);
or U8235 (N_8235,N_4188,N_2956);
and U8236 (N_8236,N_972,N_4440);
nand U8237 (N_8237,N_4799,N_3592);
nor U8238 (N_8238,N_1476,N_3100);
nand U8239 (N_8239,N_1600,N_1399);
nor U8240 (N_8240,N_4233,N_1961);
and U8241 (N_8241,N_3411,N_2265);
nor U8242 (N_8242,N_2892,N_170);
or U8243 (N_8243,N_274,N_4413);
or U8244 (N_8244,N_3130,N_2163);
or U8245 (N_8245,N_1154,N_3672);
and U8246 (N_8246,N_1645,N_1148);
nor U8247 (N_8247,N_1127,N_4686);
and U8248 (N_8248,N_3786,N_4405);
nor U8249 (N_8249,N_2333,N_1543);
or U8250 (N_8250,N_4642,N_4293);
nor U8251 (N_8251,N_4998,N_519);
or U8252 (N_8252,N_4477,N_548);
nor U8253 (N_8253,N_4244,N_833);
or U8254 (N_8254,N_1137,N_1965);
nand U8255 (N_8255,N_2391,N_23);
nand U8256 (N_8256,N_3763,N_3215);
or U8257 (N_8257,N_1986,N_1391);
nor U8258 (N_8258,N_745,N_3147);
or U8259 (N_8259,N_1751,N_761);
nor U8260 (N_8260,N_3701,N_1225);
or U8261 (N_8261,N_2242,N_2223);
nor U8262 (N_8262,N_3745,N_3950);
nand U8263 (N_8263,N_3169,N_2956);
or U8264 (N_8264,N_955,N_126);
nand U8265 (N_8265,N_2699,N_1679);
nor U8266 (N_8266,N_4551,N_4659);
nand U8267 (N_8267,N_190,N_3386);
nand U8268 (N_8268,N_2202,N_3889);
or U8269 (N_8269,N_83,N_142);
nand U8270 (N_8270,N_2689,N_3006);
nor U8271 (N_8271,N_3472,N_2320);
or U8272 (N_8272,N_3275,N_3947);
nor U8273 (N_8273,N_994,N_2152);
or U8274 (N_8274,N_4786,N_3304);
or U8275 (N_8275,N_477,N_2900);
or U8276 (N_8276,N_4580,N_1607);
nor U8277 (N_8277,N_1157,N_4963);
or U8278 (N_8278,N_4835,N_2681);
nor U8279 (N_8279,N_503,N_2057);
nor U8280 (N_8280,N_230,N_4149);
nand U8281 (N_8281,N_3892,N_4523);
nand U8282 (N_8282,N_1532,N_1751);
and U8283 (N_8283,N_3519,N_4918);
and U8284 (N_8284,N_3542,N_1063);
and U8285 (N_8285,N_2097,N_2);
and U8286 (N_8286,N_511,N_840);
nor U8287 (N_8287,N_4206,N_2460);
nand U8288 (N_8288,N_3658,N_2494);
and U8289 (N_8289,N_1730,N_1969);
or U8290 (N_8290,N_2813,N_3823);
nand U8291 (N_8291,N_2634,N_1782);
nor U8292 (N_8292,N_4528,N_1276);
and U8293 (N_8293,N_1243,N_4582);
and U8294 (N_8294,N_571,N_4675);
nor U8295 (N_8295,N_4547,N_1395);
or U8296 (N_8296,N_224,N_3439);
and U8297 (N_8297,N_2619,N_2320);
nor U8298 (N_8298,N_1639,N_2028);
nor U8299 (N_8299,N_1624,N_3455);
or U8300 (N_8300,N_4838,N_3808);
or U8301 (N_8301,N_2942,N_2860);
or U8302 (N_8302,N_4145,N_1853);
or U8303 (N_8303,N_494,N_3134);
nor U8304 (N_8304,N_960,N_4169);
or U8305 (N_8305,N_62,N_3026);
nand U8306 (N_8306,N_3657,N_3857);
and U8307 (N_8307,N_672,N_645);
nand U8308 (N_8308,N_3471,N_972);
and U8309 (N_8309,N_4669,N_4822);
nor U8310 (N_8310,N_4387,N_731);
nand U8311 (N_8311,N_2965,N_4005);
nor U8312 (N_8312,N_3674,N_924);
and U8313 (N_8313,N_3381,N_4382);
nand U8314 (N_8314,N_2975,N_63);
or U8315 (N_8315,N_465,N_3074);
nand U8316 (N_8316,N_2728,N_3839);
and U8317 (N_8317,N_2539,N_3217);
nor U8318 (N_8318,N_1986,N_3137);
or U8319 (N_8319,N_3568,N_3028);
and U8320 (N_8320,N_4842,N_3493);
nor U8321 (N_8321,N_4606,N_4529);
nand U8322 (N_8322,N_4554,N_3410);
or U8323 (N_8323,N_1199,N_2389);
nand U8324 (N_8324,N_1452,N_1046);
nand U8325 (N_8325,N_4161,N_1115);
or U8326 (N_8326,N_3591,N_1981);
and U8327 (N_8327,N_693,N_1760);
nand U8328 (N_8328,N_2943,N_366);
or U8329 (N_8329,N_4838,N_4980);
and U8330 (N_8330,N_2012,N_1562);
nor U8331 (N_8331,N_2037,N_630);
and U8332 (N_8332,N_3640,N_2933);
or U8333 (N_8333,N_1917,N_4920);
nor U8334 (N_8334,N_1560,N_2938);
and U8335 (N_8335,N_3516,N_4450);
or U8336 (N_8336,N_4785,N_2512);
nand U8337 (N_8337,N_3209,N_192);
xor U8338 (N_8338,N_4043,N_3590);
nand U8339 (N_8339,N_885,N_4818);
nand U8340 (N_8340,N_1076,N_3636);
xor U8341 (N_8341,N_522,N_2424);
and U8342 (N_8342,N_1845,N_4700);
or U8343 (N_8343,N_3148,N_2287);
and U8344 (N_8344,N_390,N_1661);
and U8345 (N_8345,N_1230,N_2413);
nor U8346 (N_8346,N_2651,N_2539);
or U8347 (N_8347,N_398,N_2131);
and U8348 (N_8348,N_4914,N_3375);
nand U8349 (N_8349,N_1379,N_649);
and U8350 (N_8350,N_2285,N_3232);
nor U8351 (N_8351,N_2973,N_1847);
and U8352 (N_8352,N_688,N_4621);
nand U8353 (N_8353,N_2177,N_3691);
or U8354 (N_8354,N_611,N_1106);
or U8355 (N_8355,N_3246,N_648);
and U8356 (N_8356,N_141,N_461);
nand U8357 (N_8357,N_3342,N_3662);
and U8358 (N_8358,N_837,N_1387);
nor U8359 (N_8359,N_2319,N_1080);
and U8360 (N_8360,N_4692,N_1581);
nor U8361 (N_8361,N_3760,N_2992);
or U8362 (N_8362,N_4518,N_3879);
and U8363 (N_8363,N_748,N_2568);
nand U8364 (N_8364,N_2505,N_977);
or U8365 (N_8365,N_1263,N_4341);
nor U8366 (N_8366,N_1713,N_797);
and U8367 (N_8367,N_4095,N_1053);
and U8368 (N_8368,N_2258,N_3880);
and U8369 (N_8369,N_2139,N_4756);
nand U8370 (N_8370,N_4867,N_4615);
nor U8371 (N_8371,N_4744,N_3006);
nor U8372 (N_8372,N_2751,N_4787);
or U8373 (N_8373,N_642,N_859);
nor U8374 (N_8374,N_1179,N_755);
or U8375 (N_8375,N_4036,N_4733);
and U8376 (N_8376,N_4075,N_4607);
nor U8377 (N_8377,N_3407,N_3713);
or U8378 (N_8378,N_2183,N_819);
or U8379 (N_8379,N_3013,N_4340);
and U8380 (N_8380,N_4257,N_4191);
nor U8381 (N_8381,N_4004,N_3372);
nor U8382 (N_8382,N_1142,N_204);
or U8383 (N_8383,N_1197,N_2375);
or U8384 (N_8384,N_3708,N_1124);
nor U8385 (N_8385,N_223,N_1339);
nand U8386 (N_8386,N_676,N_2183);
or U8387 (N_8387,N_3994,N_197);
nor U8388 (N_8388,N_1585,N_3585);
nand U8389 (N_8389,N_4781,N_616);
nand U8390 (N_8390,N_164,N_3822);
nand U8391 (N_8391,N_2547,N_582);
nor U8392 (N_8392,N_852,N_4905);
and U8393 (N_8393,N_1907,N_334);
and U8394 (N_8394,N_728,N_4867);
and U8395 (N_8395,N_3740,N_2436);
and U8396 (N_8396,N_2765,N_2436);
nand U8397 (N_8397,N_1838,N_4869);
nor U8398 (N_8398,N_2025,N_1684);
and U8399 (N_8399,N_492,N_1100);
nor U8400 (N_8400,N_2131,N_4544);
and U8401 (N_8401,N_3117,N_2774);
nor U8402 (N_8402,N_2605,N_3937);
or U8403 (N_8403,N_4723,N_2134);
nor U8404 (N_8404,N_3951,N_4039);
or U8405 (N_8405,N_3257,N_1844);
and U8406 (N_8406,N_1728,N_3350);
and U8407 (N_8407,N_2946,N_1427);
nand U8408 (N_8408,N_1427,N_1446);
and U8409 (N_8409,N_2636,N_921);
or U8410 (N_8410,N_2533,N_4134);
and U8411 (N_8411,N_4142,N_3916);
nand U8412 (N_8412,N_4741,N_4898);
nor U8413 (N_8413,N_2530,N_3965);
nor U8414 (N_8414,N_4640,N_4615);
or U8415 (N_8415,N_4726,N_1807);
nand U8416 (N_8416,N_3131,N_2925);
or U8417 (N_8417,N_3069,N_1497);
nor U8418 (N_8418,N_427,N_3641);
or U8419 (N_8419,N_4010,N_683);
and U8420 (N_8420,N_3216,N_535);
and U8421 (N_8421,N_1431,N_4712);
or U8422 (N_8422,N_753,N_2960);
nor U8423 (N_8423,N_657,N_3242);
nand U8424 (N_8424,N_4842,N_3375);
nand U8425 (N_8425,N_4360,N_1401);
or U8426 (N_8426,N_3034,N_316);
nor U8427 (N_8427,N_1777,N_4705);
nand U8428 (N_8428,N_776,N_4501);
or U8429 (N_8429,N_28,N_553);
and U8430 (N_8430,N_3075,N_3502);
or U8431 (N_8431,N_3788,N_219);
or U8432 (N_8432,N_1004,N_2349);
and U8433 (N_8433,N_4168,N_1978);
or U8434 (N_8434,N_3950,N_3287);
or U8435 (N_8435,N_1940,N_2245);
and U8436 (N_8436,N_1071,N_3097);
nor U8437 (N_8437,N_2858,N_1446);
nor U8438 (N_8438,N_1087,N_1361);
or U8439 (N_8439,N_3355,N_4230);
or U8440 (N_8440,N_2162,N_816);
and U8441 (N_8441,N_3351,N_1644);
nand U8442 (N_8442,N_3016,N_1829);
and U8443 (N_8443,N_214,N_1933);
nor U8444 (N_8444,N_1999,N_2575);
nand U8445 (N_8445,N_3702,N_405);
or U8446 (N_8446,N_2290,N_3259);
or U8447 (N_8447,N_4069,N_3862);
or U8448 (N_8448,N_3110,N_1658);
or U8449 (N_8449,N_2020,N_961);
nor U8450 (N_8450,N_3216,N_1099);
or U8451 (N_8451,N_4748,N_1335);
nand U8452 (N_8452,N_1426,N_4851);
nor U8453 (N_8453,N_1069,N_537);
or U8454 (N_8454,N_921,N_832);
and U8455 (N_8455,N_1313,N_4741);
nand U8456 (N_8456,N_1098,N_1517);
or U8457 (N_8457,N_4071,N_3892);
and U8458 (N_8458,N_4809,N_1330);
nand U8459 (N_8459,N_4618,N_2448);
nand U8460 (N_8460,N_1245,N_1962);
or U8461 (N_8461,N_1764,N_4410);
or U8462 (N_8462,N_3914,N_1643);
nor U8463 (N_8463,N_4025,N_1501);
nand U8464 (N_8464,N_4374,N_166);
nor U8465 (N_8465,N_672,N_3317);
and U8466 (N_8466,N_3139,N_2156);
nand U8467 (N_8467,N_3482,N_3399);
nand U8468 (N_8468,N_1752,N_4204);
or U8469 (N_8469,N_3428,N_770);
nand U8470 (N_8470,N_248,N_4983);
nor U8471 (N_8471,N_4895,N_1391);
and U8472 (N_8472,N_4519,N_296);
and U8473 (N_8473,N_1458,N_346);
and U8474 (N_8474,N_905,N_3314);
and U8475 (N_8475,N_551,N_946);
or U8476 (N_8476,N_3119,N_205);
xnor U8477 (N_8477,N_338,N_3368);
or U8478 (N_8478,N_4172,N_693);
nor U8479 (N_8479,N_103,N_3463);
nand U8480 (N_8480,N_3568,N_3869);
nand U8481 (N_8481,N_3487,N_124);
and U8482 (N_8482,N_2650,N_3140);
nor U8483 (N_8483,N_1465,N_174);
nand U8484 (N_8484,N_3415,N_4380);
nand U8485 (N_8485,N_2416,N_4149);
nand U8486 (N_8486,N_4863,N_3723);
nor U8487 (N_8487,N_4138,N_1276);
and U8488 (N_8488,N_2004,N_2715);
and U8489 (N_8489,N_2664,N_4898);
nor U8490 (N_8490,N_1883,N_4987);
nand U8491 (N_8491,N_4861,N_2848);
or U8492 (N_8492,N_203,N_1763);
nand U8493 (N_8493,N_4262,N_2147);
nand U8494 (N_8494,N_3302,N_3078);
nand U8495 (N_8495,N_1820,N_3915);
nor U8496 (N_8496,N_998,N_1085);
nor U8497 (N_8497,N_4126,N_4797);
or U8498 (N_8498,N_1243,N_956);
nand U8499 (N_8499,N_3704,N_1894);
nand U8500 (N_8500,N_1302,N_4755);
nor U8501 (N_8501,N_4543,N_33);
nand U8502 (N_8502,N_988,N_3808);
and U8503 (N_8503,N_2336,N_646);
nand U8504 (N_8504,N_224,N_2641);
or U8505 (N_8505,N_1034,N_3213);
or U8506 (N_8506,N_801,N_3471);
and U8507 (N_8507,N_2026,N_250);
and U8508 (N_8508,N_2010,N_1476);
nor U8509 (N_8509,N_2288,N_4639);
and U8510 (N_8510,N_2445,N_2307);
and U8511 (N_8511,N_4534,N_629);
and U8512 (N_8512,N_1949,N_1353);
or U8513 (N_8513,N_374,N_3932);
nor U8514 (N_8514,N_1580,N_4753);
or U8515 (N_8515,N_4,N_2139);
or U8516 (N_8516,N_4112,N_2799);
or U8517 (N_8517,N_1574,N_233);
nor U8518 (N_8518,N_3519,N_2706);
or U8519 (N_8519,N_816,N_3637);
or U8520 (N_8520,N_2857,N_2702);
nor U8521 (N_8521,N_4465,N_2076);
nor U8522 (N_8522,N_1850,N_3485);
nor U8523 (N_8523,N_137,N_3090);
or U8524 (N_8524,N_3452,N_3071);
or U8525 (N_8525,N_4103,N_1272);
nor U8526 (N_8526,N_4348,N_3338);
and U8527 (N_8527,N_4007,N_4955);
nor U8528 (N_8528,N_261,N_2346);
nand U8529 (N_8529,N_1005,N_1498);
nor U8530 (N_8530,N_575,N_2574);
nor U8531 (N_8531,N_2317,N_1319);
and U8532 (N_8532,N_1510,N_1439);
nand U8533 (N_8533,N_412,N_3916);
nand U8534 (N_8534,N_1641,N_192);
nor U8535 (N_8535,N_3480,N_1228);
nor U8536 (N_8536,N_3472,N_78);
or U8537 (N_8537,N_1506,N_3152);
nor U8538 (N_8538,N_2828,N_2848);
and U8539 (N_8539,N_3549,N_3238);
or U8540 (N_8540,N_3590,N_3076);
nor U8541 (N_8541,N_2074,N_4123);
or U8542 (N_8542,N_3045,N_3865);
or U8543 (N_8543,N_1268,N_3877);
and U8544 (N_8544,N_2500,N_4922);
nand U8545 (N_8545,N_2243,N_1115);
nand U8546 (N_8546,N_4498,N_2109);
nor U8547 (N_8547,N_1760,N_4755);
nor U8548 (N_8548,N_3256,N_296);
nor U8549 (N_8549,N_4747,N_4540);
and U8550 (N_8550,N_2883,N_162);
and U8551 (N_8551,N_2884,N_988);
nor U8552 (N_8552,N_1861,N_4817);
or U8553 (N_8553,N_1683,N_2049);
and U8554 (N_8554,N_314,N_4158);
or U8555 (N_8555,N_4008,N_106);
nand U8556 (N_8556,N_703,N_4469);
nand U8557 (N_8557,N_45,N_699);
and U8558 (N_8558,N_2573,N_293);
nor U8559 (N_8559,N_3693,N_4688);
nor U8560 (N_8560,N_1364,N_2532);
and U8561 (N_8561,N_4088,N_170);
and U8562 (N_8562,N_4880,N_3987);
nor U8563 (N_8563,N_4310,N_887);
nor U8564 (N_8564,N_1293,N_1961);
nand U8565 (N_8565,N_165,N_1151);
nor U8566 (N_8566,N_3193,N_3350);
or U8567 (N_8567,N_2847,N_1786);
nand U8568 (N_8568,N_3959,N_2708);
nor U8569 (N_8569,N_355,N_3039);
nor U8570 (N_8570,N_3748,N_94);
and U8571 (N_8571,N_1310,N_2500);
nor U8572 (N_8572,N_4267,N_2030);
or U8573 (N_8573,N_1305,N_4744);
nand U8574 (N_8574,N_2579,N_1243);
nor U8575 (N_8575,N_3289,N_2569);
or U8576 (N_8576,N_1150,N_2252);
nand U8577 (N_8577,N_544,N_1048);
and U8578 (N_8578,N_3879,N_413);
nand U8579 (N_8579,N_1950,N_376);
and U8580 (N_8580,N_3454,N_3688);
nand U8581 (N_8581,N_4258,N_3648);
and U8582 (N_8582,N_3537,N_3354);
or U8583 (N_8583,N_3200,N_3965);
nand U8584 (N_8584,N_723,N_3334);
nand U8585 (N_8585,N_562,N_1590);
and U8586 (N_8586,N_1115,N_1143);
and U8587 (N_8587,N_326,N_565);
nor U8588 (N_8588,N_2597,N_4015);
nand U8589 (N_8589,N_1584,N_1317);
nand U8590 (N_8590,N_2653,N_262);
nor U8591 (N_8591,N_1069,N_955);
nor U8592 (N_8592,N_1544,N_4938);
or U8593 (N_8593,N_2523,N_3236);
nand U8594 (N_8594,N_3703,N_2442);
nand U8595 (N_8595,N_3418,N_3032);
and U8596 (N_8596,N_4191,N_3135);
or U8597 (N_8597,N_412,N_1125);
nor U8598 (N_8598,N_4676,N_4705);
and U8599 (N_8599,N_3986,N_290);
nand U8600 (N_8600,N_1210,N_2068);
or U8601 (N_8601,N_718,N_3702);
nand U8602 (N_8602,N_385,N_222);
or U8603 (N_8603,N_3409,N_392);
nand U8604 (N_8604,N_2876,N_31);
and U8605 (N_8605,N_2880,N_162);
and U8606 (N_8606,N_1175,N_1280);
nor U8607 (N_8607,N_2665,N_4528);
or U8608 (N_8608,N_4280,N_1870);
or U8609 (N_8609,N_1327,N_3010);
and U8610 (N_8610,N_4390,N_2924);
nor U8611 (N_8611,N_638,N_2527);
or U8612 (N_8612,N_466,N_1086);
nor U8613 (N_8613,N_1635,N_1782);
nand U8614 (N_8614,N_1969,N_2380);
nand U8615 (N_8615,N_1008,N_408);
nor U8616 (N_8616,N_3679,N_1080);
nor U8617 (N_8617,N_532,N_1115);
nand U8618 (N_8618,N_1176,N_4817);
or U8619 (N_8619,N_4631,N_3820);
or U8620 (N_8620,N_1385,N_1244);
nand U8621 (N_8621,N_2955,N_3930);
nand U8622 (N_8622,N_2196,N_2580);
nand U8623 (N_8623,N_662,N_796);
nand U8624 (N_8624,N_1324,N_1110);
and U8625 (N_8625,N_105,N_925);
nor U8626 (N_8626,N_3681,N_4446);
nor U8627 (N_8627,N_100,N_2896);
nand U8628 (N_8628,N_4529,N_3184);
nand U8629 (N_8629,N_4347,N_490);
nor U8630 (N_8630,N_4045,N_4718);
nand U8631 (N_8631,N_531,N_2384);
or U8632 (N_8632,N_1722,N_3112);
nand U8633 (N_8633,N_1767,N_535);
nor U8634 (N_8634,N_3019,N_1507);
nand U8635 (N_8635,N_1379,N_1112);
or U8636 (N_8636,N_2419,N_4337);
nand U8637 (N_8637,N_4902,N_3894);
or U8638 (N_8638,N_2912,N_3632);
nand U8639 (N_8639,N_959,N_4091);
and U8640 (N_8640,N_3376,N_2164);
nor U8641 (N_8641,N_2138,N_607);
nor U8642 (N_8642,N_4742,N_1852);
or U8643 (N_8643,N_2533,N_3602);
or U8644 (N_8644,N_3821,N_58);
and U8645 (N_8645,N_4402,N_51);
nor U8646 (N_8646,N_267,N_1084);
and U8647 (N_8647,N_3226,N_370);
nand U8648 (N_8648,N_863,N_3191);
nand U8649 (N_8649,N_4863,N_4276);
nor U8650 (N_8650,N_4370,N_3651);
and U8651 (N_8651,N_3659,N_4344);
and U8652 (N_8652,N_1339,N_2089);
and U8653 (N_8653,N_3220,N_53);
or U8654 (N_8654,N_768,N_2073);
and U8655 (N_8655,N_1413,N_3279);
nor U8656 (N_8656,N_3904,N_138);
and U8657 (N_8657,N_2304,N_3075);
or U8658 (N_8658,N_568,N_2798);
xor U8659 (N_8659,N_89,N_3410);
or U8660 (N_8660,N_797,N_4764);
nand U8661 (N_8661,N_1207,N_3854);
nand U8662 (N_8662,N_3833,N_782);
or U8663 (N_8663,N_492,N_4881);
and U8664 (N_8664,N_343,N_1730);
nor U8665 (N_8665,N_122,N_4925);
and U8666 (N_8666,N_406,N_2888);
nand U8667 (N_8667,N_4930,N_1723);
nor U8668 (N_8668,N_4102,N_2679);
nor U8669 (N_8669,N_425,N_3703);
or U8670 (N_8670,N_1264,N_4809);
and U8671 (N_8671,N_2550,N_2395);
nand U8672 (N_8672,N_3768,N_3897);
nor U8673 (N_8673,N_1304,N_1457);
and U8674 (N_8674,N_3654,N_4255);
nor U8675 (N_8675,N_4965,N_3307);
or U8676 (N_8676,N_2135,N_567);
or U8677 (N_8677,N_959,N_3670);
nor U8678 (N_8678,N_4987,N_4308);
or U8679 (N_8679,N_771,N_4095);
and U8680 (N_8680,N_1418,N_1078);
nand U8681 (N_8681,N_3321,N_3743);
or U8682 (N_8682,N_2058,N_746);
or U8683 (N_8683,N_148,N_559);
nand U8684 (N_8684,N_4543,N_2157);
or U8685 (N_8685,N_1814,N_3981);
and U8686 (N_8686,N_95,N_144);
or U8687 (N_8687,N_3227,N_2599);
nand U8688 (N_8688,N_807,N_4375);
nor U8689 (N_8689,N_4682,N_4583);
and U8690 (N_8690,N_1103,N_2427);
and U8691 (N_8691,N_4663,N_167);
nand U8692 (N_8692,N_475,N_699);
nor U8693 (N_8693,N_2882,N_4187);
nand U8694 (N_8694,N_4305,N_1079);
and U8695 (N_8695,N_4593,N_3007);
nand U8696 (N_8696,N_997,N_1099);
nor U8697 (N_8697,N_1426,N_2637);
nor U8698 (N_8698,N_141,N_4629);
nor U8699 (N_8699,N_4597,N_2941);
or U8700 (N_8700,N_4015,N_4919);
nand U8701 (N_8701,N_872,N_3785);
or U8702 (N_8702,N_1987,N_2654);
nand U8703 (N_8703,N_3177,N_4167);
nor U8704 (N_8704,N_4837,N_4829);
or U8705 (N_8705,N_2596,N_1405);
nand U8706 (N_8706,N_1061,N_2495);
or U8707 (N_8707,N_1722,N_752);
and U8708 (N_8708,N_1231,N_1784);
and U8709 (N_8709,N_2702,N_2665);
and U8710 (N_8710,N_4594,N_812);
nor U8711 (N_8711,N_2348,N_2377);
and U8712 (N_8712,N_2808,N_699);
nor U8713 (N_8713,N_2175,N_1195);
nor U8714 (N_8714,N_3280,N_321);
and U8715 (N_8715,N_1509,N_4568);
nor U8716 (N_8716,N_3361,N_1208);
and U8717 (N_8717,N_3868,N_3991);
or U8718 (N_8718,N_2860,N_3774);
xor U8719 (N_8719,N_388,N_1606);
or U8720 (N_8720,N_1511,N_2381);
nand U8721 (N_8721,N_913,N_1866);
or U8722 (N_8722,N_1755,N_2073);
or U8723 (N_8723,N_4223,N_3364);
nor U8724 (N_8724,N_1093,N_3594);
or U8725 (N_8725,N_320,N_3111);
nand U8726 (N_8726,N_3148,N_2435);
and U8727 (N_8727,N_3302,N_2295);
or U8728 (N_8728,N_2572,N_1192);
and U8729 (N_8729,N_4242,N_4405);
nor U8730 (N_8730,N_2472,N_244);
or U8731 (N_8731,N_3244,N_4713);
or U8732 (N_8732,N_683,N_4661);
xor U8733 (N_8733,N_1128,N_4356);
nor U8734 (N_8734,N_716,N_4933);
or U8735 (N_8735,N_3703,N_950);
nor U8736 (N_8736,N_4849,N_1408);
and U8737 (N_8737,N_3708,N_618);
and U8738 (N_8738,N_715,N_3302);
or U8739 (N_8739,N_214,N_146);
or U8740 (N_8740,N_4272,N_1028);
or U8741 (N_8741,N_3157,N_1360);
or U8742 (N_8742,N_2687,N_770);
or U8743 (N_8743,N_2486,N_3348);
nor U8744 (N_8744,N_4044,N_1195);
and U8745 (N_8745,N_557,N_805);
and U8746 (N_8746,N_1896,N_3231);
nand U8747 (N_8747,N_3477,N_2338);
or U8748 (N_8748,N_4323,N_3444);
and U8749 (N_8749,N_563,N_2744);
or U8750 (N_8750,N_3545,N_2649);
nand U8751 (N_8751,N_64,N_4397);
or U8752 (N_8752,N_323,N_2846);
nor U8753 (N_8753,N_2390,N_522);
or U8754 (N_8754,N_1888,N_1086);
and U8755 (N_8755,N_3009,N_1333);
nor U8756 (N_8756,N_1929,N_902);
nor U8757 (N_8757,N_3684,N_80);
nor U8758 (N_8758,N_4449,N_4177);
nand U8759 (N_8759,N_1295,N_2425);
or U8760 (N_8760,N_376,N_4258);
nand U8761 (N_8761,N_4545,N_3160);
nand U8762 (N_8762,N_3702,N_342);
and U8763 (N_8763,N_4286,N_861);
or U8764 (N_8764,N_853,N_782);
or U8765 (N_8765,N_1742,N_2737);
nand U8766 (N_8766,N_3797,N_4962);
and U8767 (N_8767,N_3584,N_456);
and U8768 (N_8768,N_4282,N_58);
or U8769 (N_8769,N_4175,N_404);
nand U8770 (N_8770,N_3941,N_563);
and U8771 (N_8771,N_2821,N_40);
or U8772 (N_8772,N_7,N_1671);
and U8773 (N_8773,N_3021,N_642);
or U8774 (N_8774,N_4007,N_4239);
nor U8775 (N_8775,N_2456,N_4695);
and U8776 (N_8776,N_3759,N_3182);
and U8777 (N_8777,N_4192,N_1277);
and U8778 (N_8778,N_788,N_3447);
and U8779 (N_8779,N_4747,N_3507);
nor U8780 (N_8780,N_4099,N_2680);
nand U8781 (N_8781,N_4214,N_3603);
or U8782 (N_8782,N_3235,N_4300);
nor U8783 (N_8783,N_3948,N_3681);
and U8784 (N_8784,N_166,N_2174);
or U8785 (N_8785,N_1152,N_4916);
nand U8786 (N_8786,N_1695,N_701);
and U8787 (N_8787,N_1843,N_3310);
or U8788 (N_8788,N_52,N_4996);
or U8789 (N_8789,N_606,N_1660);
and U8790 (N_8790,N_3485,N_1817);
xor U8791 (N_8791,N_2176,N_101);
or U8792 (N_8792,N_4775,N_4860);
and U8793 (N_8793,N_3367,N_1569);
nor U8794 (N_8794,N_2733,N_2351);
nand U8795 (N_8795,N_3911,N_1817);
and U8796 (N_8796,N_4554,N_2133);
or U8797 (N_8797,N_1347,N_4641);
nand U8798 (N_8798,N_3105,N_4797);
and U8799 (N_8799,N_3312,N_4260);
or U8800 (N_8800,N_4479,N_4886);
and U8801 (N_8801,N_4439,N_297);
or U8802 (N_8802,N_2887,N_3475);
and U8803 (N_8803,N_2127,N_3672);
nand U8804 (N_8804,N_4354,N_1254);
or U8805 (N_8805,N_3519,N_3163);
nand U8806 (N_8806,N_2836,N_125);
nand U8807 (N_8807,N_2386,N_4796);
or U8808 (N_8808,N_1706,N_259);
or U8809 (N_8809,N_827,N_4545);
nor U8810 (N_8810,N_4662,N_4062);
and U8811 (N_8811,N_3183,N_3776);
nor U8812 (N_8812,N_681,N_907);
nor U8813 (N_8813,N_149,N_67);
or U8814 (N_8814,N_1274,N_2285);
or U8815 (N_8815,N_1799,N_3225);
nand U8816 (N_8816,N_2869,N_3966);
or U8817 (N_8817,N_2055,N_2109);
and U8818 (N_8818,N_4250,N_4786);
or U8819 (N_8819,N_404,N_1481);
and U8820 (N_8820,N_2046,N_2248);
nor U8821 (N_8821,N_1426,N_2783);
nor U8822 (N_8822,N_1050,N_2686);
nor U8823 (N_8823,N_1598,N_4849);
nand U8824 (N_8824,N_3107,N_2980);
nand U8825 (N_8825,N_1200,N_3859);
nand U8826 (N_8826,N_4775,N_2575);
nor U8827 (N_8827,N_3524,N_2791);
and U8828 (N_8828,N_1509,N_4053);
and U8829 (N_8829,N_503,N_1307);
nor U8830 (N_8830,N_1018,N_2862);
nand U8831 (N_8831,N_4285,N_2917);
nor U8832 (N_8832,N_4343,N_175);
nor U8833 (N_8833,N_4476,N_1213);
nand U8834 (N_8834,N_274,N_1041);
nand U8835 (N_8835,N_1258,N_2339);
nand U8836 (N_8836,N_4896,N_279);
or U8837 (N_8837,N_2502,N_1427);
and U8838 (N_8838,N_2337,N_3487);
and U8839 (N_8839,N_360,N_414);
and U8840 (N_8840,N_739,N_801);
or U8841 (N_8841,N_494,N_1763);
or U8842 (N_8842,N_1975,N_2655);
nor U8843 (N_8843,N_3675,N_2465);
nand U8844 (N_8844,N_4038,N_4624);
nand U8845 (N_8845,N_2757,N_1813);
nor U8846 (N_8846,N_3536,N_4975);
or U8847 (N_8847,N_1789,N_2461);
nand U8848 (N_8848,N_4187,N_3546);
or U8849 (N_8849,N_407,N_2264);
nand U8850 (N_8850,N_975,N_772);
nand U8851 (N_8851,N_2677,N_488);
and U8852 (N_8852,N_3422,N_3848);
and U8853 (N_8853,N_794,N_3013);
nor U8854 (N_8854,N_187,N_1183);
nor U8855 (N_8855,N_3075,N_1890);
and U8856 (N_8856,N_2170,N_3572);
and U8857 (N_8857,N_4452,N_48);
and U8858 (N_8858,N_3576,N_4696);
nand U8859 (N_8859,N_388,N_1341);
or U8860 (N_8860,N_1026,N_620);
nand U8861 (N_8861,N_1687,N_3128);
and U8862 (N_8862,N_3781,N_1119);
or U8863 (N_8863,N_127,N_2477);
or U8864 (N_8864,N_3706,N_4512);
nor U8865 (N_8865,N_1056,N_1406);
and U8866 (N_8866,N_566,N_3081);
and U8867 (N_8867,N_2235,N_2943);
nor U8868 (N_8868,N_2716,N_2105);
and U8869 (N_8869,N_4045,N_3055);
and U8870 (N_8870,N_4150,N_1230);
or U8871 (N_8871,N_1048,N_1695);
or U8872 (N_8872,N_1840,N_4648);
and U8873 (N_8873,N_4890,N_4073);
and U8874 (N_8874,N_3288,N_1818);
nor U8875 (N_8875,N_585,N_38);
nand U8876 (N_8876,N_4881,N_3683);
nor U8877 (N_8877,N_1640,N_3939);
or U8878 (N_8878,N_4656,N_3496);
and U8879 (N_8879,N_3909,N_740);
nor U8880 (N_8880,N_2298,N_2104);
nand U8881 (N_8881,N_942,N_470);
or U8882 (N_8882,N_2007,N_4366);
and U8883 (N_8883,N_1785,N_1775);
and U8884 (N_8884,N_877,N_4585);
nor U8885 (N_8885,N_1538,N_1621);
or U8886 (N_8886,N_3484,N_499);
nor U8887 (N_8887,N_4030,N_3664);
nand U8888 (N_8888,N_444,N_3570);
nand U8889 (N_8889,N_119,N_4521);
nor U8890 (N_8890,N_3655,N_1157);
or U8891 (N_8891,N_2332,N_4495);
nor U8892 (N_8892,N_747,N_577);
and U8893 (N_8893,N_4763,N_1837);
or U8894 (N_8894,N_3918,N_4491);
nor U8895 (N_8895,N_1985,N_2306);
or U8896 (N_8896,N_357,N_1733);
nor U8897 (N_8897,N_398,N_1570);
or U8898 (N_8898,N_4002,N_1202);
nand U8899 (N_8899,N_2640,N_1603);
nor U8900 (N_8900,N_15,N_4356);
or U8901 (N_8901,N_1057,N_3042);
nand U8902 (N_8902,N_3808,N_3746);
nor U8903 (N_8903,N_1165,N_1731);
nor U8904 (N_8904,N_4926,N_4032);
or U8905 (N_8905,N_4967,N_3284);
or U8906 (N_8906,N_4638,N_2559);
and U8907 (N_8907,N_2931,N_1629);
or U8908 (N_8908,N_3041,N_870);
and U8909 (N_8909,N_4153,N_3386);
nor U8910 (N_8910,N_3640,N_2924);
or U8911 (N_8911,N_4120,N_1795);
or U8912 (N_8912,N_1675,N_2752);
nand U8913 (N_8913,N_380,N_4907);
nand U8914 (N_8914,N_2591,N_2555);
nand U8915 (N_8915,N_2983,N_2887);
nand U8916 (N_8916,N_3471,N_4562);
and U8917 (N_8917,N_3253,N_1609);
and U8918 (N_8918,N_1528,N_3367);
and U8919 (N_8919,N_490,N_335);
or U8920 (N_8920,N_283,N_3813);
and U8921 (N_8921,N_2806,N_396);
and U8922 (N_8922,N_340,N_192);
and U8923 (N_8923,N_4366,N_1900);
xor U8924 (N_8924,N_2048,N_460);
nand U8925 (N_8925,N_2292,N_86);
and U8926 (N_8926,N_2968,N_1499);
nand U8927 (N_8927,N_4837,N_2951);
nand U8928 (N_8928,N_4661,N_2286);
or U8929 (N_8929,N_857,N_673);
nor U8930 (N_8930,N_2860,N_1766);
and U8931 (N_8931,N_3524,N_806);
nand U8932 (N_8932,N_3973,N_2623);
nand U8933 (N_8933,N_2789,N_385);
nor U8934 (N_8934,N_1598,N_3314);
or U8935 (N_8935,N_2137,N_4052);
nand U8936 (N_8936,N_568,N_777);
and U8937 (N_8937,N_4846,N_2870);
nor U8938 (N_8938,N_1950,N_1994);
and U8939 (N_8939,N_610,N_4785);
and U8940 (N_8940,N_2691,N_1438);
and U8941 (N_8941,N_3034,N_3762);
or U8942 (N_8942,N_2654,N_1967);
and U8943 (N_8943,N_1429,N_1610);
or U8944 (N_8944,N_4025,N_358);
nand U8945 (N_8945,N_3241,N_432);
or U8946 (N_8946,N_651,N_4689);
nor U8947 (N_8947,N_1661,N_1463);
and U8948 (N_8948,N_4868,N_1122);
and U8949 (N_8949,N_1307,N_2949);
and U8950 (N_8950,N_4077,N_4709);
or U8951 (N_8951,N_1406,N_3115);
or U8952 (N_8952,N_710,N_2736);
or U8953 (N_8953,N_143,N_2888);
or U8954 (N_8954,N_1176,N_1808);
and U8955 (N_8955,N_1008,N_4475);
and U8956 (N_8956,N_4224,N_2133);
nor U8957 (N_8957,N_2445,N_3454);
xnor U8958 (N_8958,N_504,N_1702);
nor U8959 (N_8959,N_750,N_2339);
or U8960 (N_8960,N_372,N_4408);
and U8961 (N_8961,N_2565,N_3509);
nand U8962 (N_8962,N_1304,N_2726);
nor U8963 (N_8963,N_3933,N_2158);
and U8964 (N_8964,N_3267,N_214);
nor U8965 (N_8965,N_1212,N_1414);
and U8966 (N_8966,N_1928,N_2875);
and U8967 (N_8967,N_816,N_4434);
nor U8968 (N_8968,N_4945,N_495);
nor U8969 (N_8969,N_516,N_2697);
or U8970 (N_8970,N_4832,N_1103);
nor U8971 (N_8971,N_3019,N_1847);
and U8972 (N_8972,N_4982,N_1928);
or U8973 (N_8973,N_1424,N_3027);
and U8974 (N_8974,N_4719,N_428);
or U8975 (N_8975,N_2600,N_1664);
nand U8976 (N_8976,N_1861,N_1292);
nor U8977 (N_8977,N_2979,N_4410);
nor U8978 (N_8978,N_2980,N_4394);
nor U8979 (N_8979,N_1516,N_3573);
nand U8980 (N_8980,N_3103,N_1712);
nand U8981 (N_8981,N_1779,N_657);
and U8982 (N_8982,N_1308,N_2321);
or U8983 (N_8983,N_1263,N_760);
and U8984 (N_8984,N_3310,N_4090);
nor U8985 (N_8985,N_4019,N_2466);
or U8986 (N_8986,N_4906,N_1974);
nor U8987 (N_8987,N_4429,N_4906);
or U8988 (N_8988,N_4269,N_3903);
nand U8989 (N_8989,N_2571,N_1210);
or U8990 (N_8990,N_2399,N_1136);
or U8991 (N_8991,N_4661,N_3606);
or U8992 (N_8992,N_3871,N_3195);
nor U8993 (N_8993,N_3609,N_214);
nor U8994 (N_8994,N_581,N_3865);
nor U8995 (N_8995,N_890,N_2971);
and U8996 (N_8996,N_1671,N_2829);
or U8997 (N_8997,N_1791,N_973);
and U8998 (N_8998,N_3205,N_265);
or U8999 (N_8999,N_3927,N_2085);
and U9000 (N_9000,N_2579,N_500);
and U9001 (N_9001,N_1120,N_2153);
nand U9002 (N_9002,N_1738,N_3470);
or U9003 (N_9003,N_3111,N_2299);
or U9004 (N_9004,N_3133,N_2188);
and U9005 (N_9005,N_4364,N_91);
nor U9006 (N_9006,N_2177,N_4885);
nor U9007 (N_9007,N_181,N_2394);
nor U9008 (N_9008,N_342,N_825);
and U9009 (N_9009,N_4968,N_3993);
and U9010 (N_9010,N_1468,N_1482);
or U9011 (N_9011,N_709,N_3116);
nand U9012 (N_9012,N_3773,N_4144);
nor U9013 (N_9013,N_3311,N_3726);
and U9014 (N_9014,N_1138,N_140);
and U9015 (N_9015,N_3326,N_793);
and U9016 (N_9016,N_1465,N_2201);
nor U9017 (N_9017,N_864,N_3153);
nor U9018 (N_9018,N_2580,N_1619);
nor U9019 (N_9019,N_1518,N_1277);
nand U9020 (N_9020,N_1279,N_3433);
and U9021 (N_9021,N_2570,N_3239);
and U9022 (N_9022,N_245,N_2989);
and U9023 (N_9023,N_762,N_2548);
and U9024 (N_9024,N_1743,N_3530);
nand U9025 (N_9025,N_4937,N_3466);
nand U9026 (N_9026,N_4346,N_3230);
and U9027 (N_9027,N_815,N_2292);
and U9028 (N_9028,N_4620,N_375);
and U9029 (N_9029,N_2058,N_4583);
nand U9030 (N_9030,N_3535,N_2006);
and U9031 (N_9031,N_1535,N_55);
nor U9032 (N_9032,N_2309,N_586);
nand U9033 (N_9033,N_70,N_4055);
and U9034 (N_9034,N_3209,N_1111);
and U9035 (N_9035,N_3645,N_2221);
or U9036 (N_9036,N_190,N_4596);
nand U9037 (N_9037,N_953,N_1422);
nor U9038 (N_9038,N_4960,N_2525);
nand U9039 (N_9039,N_485,N_2567);
nand U9040 (N_9040,N_3663,N_2196);
nand U9041 (N_9041,N_2165,N_3785);
nand U9042 (N_9042,N_3556,N_3681);
nor U9043 (N_9043,N_2145,N_919);
nor U9044 (N_9044,N_1895,N_4080);
and U9045 (N_9045,N_4233,N_1736);
or U9046 (N_9046,N_3080,N_4861);
nand U9047 (N_9047,N_3401,N_647);
nand U9048 (N_9048,N_4010,N_4368);
or U9049 (N_9049,N_236,N_3938);
nor U9050 (N_9050,N_682,N_3821);
and U9051 (N_9051,N_2989,N_1511);
xnor U9052 (N_9052,N_2514,N_4069);
or U9053 (N_9053,N_1877,N_2161);
and U9054 (N_9054,N_4131,N_3760);
nand U9055 (N_9055,N_3531,N_4111);
and U9056 (N_9056,N_3436,N_4789);
xor U9057 (N_9057,N_3461,N_724);
or U9058 (N_9058,N_1485,N_3368);
nand U9059 (N_9059,N_1967,N_2928);
and U9060 (N_9060,N_3261,N_3002);
nor U9061 (N_9061,N_4133,N_2128);
nand U9062 (N_9062,N_1685,N_110);
nand U9063 (N_9063,N_1057,N_3503);
nor U9064 (N_9064,N_557,N_354);
nor U9065 (N_9065,N_877,N_2451);
nand U9066 (N_9066,N_4632,N_4073);
or U9067 (N_9067,N_2942,N_4109);
nor U9068 (N_9068,N_2586,N_594);
and U9069 (N_9069,N_3292,N_1418);
nor U9070 (N_9070,N_480,N_224);
and U9071 (N_9071,N_3247,N_4070);
nor U9072 (N_9072,N_2925,N_168);
nor U9073 (N_9073,N_4816,N_1833);
and U9074 (N_9074,N_1342,N_1403);
nand U9075 (N_9075,N_4455,N_3876);
or U9076 (N_9076,N_3708,N_1235);
and U9077 (N_9077,N_600,N_4258);
nand U9078 (N_9078,N_1517,N_2034);
and U9079 (N_9079,N_1591,N_1537);
nand U9080 (N_9080,N_2112,N_846);
nand U9081 (N_9081,N_4361,N_17);
nand U9082 (N_9082,N_2449,N_3700);
and U9083 (N_9083,N_2720,N_2339);
or U9084 (N_9084,N_3694,N_2209);
or U9085 (N_9085,N_4525,N_3075);
nand U9086 (N_9086,N_1090,N_4327);
or U9087 (N_9087,N_3134,N_2177);
nor U9088 (N_9088,N_3633,N_366);
nor U9089 (N_9089,N_4847,N_2497);
or U9090 (N_9090,N_4253,N_3781);
or U9091 (N_9091,N_4879,N_2863);
nor U9092 (N_9092,N_3988,N_4236);
or U9093 (N_9093,N_161,N_1849);
nor U9094 (N_9094,N_3945,N_3053);
nand U9095 (N_9095,N_1231,N_3908);
or U9096 (N_9096,N_1115,N_1153);
or U9097 (N_9097,N_4161,N_2837);
and U9098 (N_9098,N_4846,N_4739);
nand U9099 (N_9099,N_3678,N_201);
or U9100 (N_9100,N_4337,N_916);
or U9101 (N_9101,N_3998,N_2315);
and U9102 (N_9102,N_2705,N_3593);
nand U9103 (N_9103,N_1880,N_3010);
and U9104 (N_9104,N_2852,N_756);
nand U9105 (N_9105,N_4710,N_3115);
nand U9106 (N_9106,N_855,N_2097);
or U9107 (N_9107,N_4985,N_723);
or U9108 (N_9108,N_1888,N_217);
nor U9109 (N_9109,N_511,N_4177);
or U9110 (N_9110,N_59,N_1439);
and U9111 (N_9111,N_190,N_4582);
nor U9112 (N_9112,N_964,N_2125);
nor U9113 (N_9113,N_1359,N_2041);
or U9114 (N_9114,N_1417,N_1043);
and U9115 (N_9115,N_244,N_1449);
or U9116 (N_9116,N_1038,N_4433);
nand U9117 (N_9117,N_470,N_618);
or U9118 (N_9118,N_3949,N_1224);
nor U9119 (N_9119,N_694,N_723);
nor U9120 (N_9120,N_4835,N_2592);
and U9121 (N_9121,N_2607,N_1541);
nand U9122 (N_9122,N_1963,N_3436);
or U9123 (N_9123,N_2393,N_3442);
and U9124 (N_9124,N_3375,N_4439);
or U9125 (N_9125,N_4292,N_4131);
nor U9126 (N_9126,N_1972,N_2208);
and U9127 (N_9127,N_2873,N_547);
or U9128 (N_9128,N_2444,N_3659);
or U9129 (N_9129,N_1180,N_3433);
nand U9130 (N_9130,N_2092,N_3776);
nor U9131 (N_9131,N_4358,N_1939);
or U9132 (N_9132,N_2821,N_1215);
or U9133 (N_9133,N_2217,N_3751);
or U9134 (N_9134,N_813,N_3865);
nand U9135 (N_9135,N_3501,N_2959);
and U9136 (N_9136,N_1637,N_2176);
and U9137 (N_9137,N_1916,N_3790);
and U9138 (N_9138,N_4138,N_1545);
and U9139 (N_9139,N_2260,N_4597);
nand U9140 (N_9140,N_3429,N_1597);
nor U9141 (N_9141,N_4857,N_4011);
or U9142 (N_9142,N_2211,N_4765);
nor U9143 (N_9143,N_1945,N_1154);
nand U9144 (N_9144,N_3032,N_3897);
nand U9145 (N_9145,N_592,N_2369);
nand U9146 (N_9146,N_4470,N_1240);
and U9147 (N_9147,N_4839,N_3302);
nand U9148 (N_9148,N_2636,N_2533);
or U9149 (N_9149,N_311,N_4693);
and U9150 (N_9150,N_283,N_1062);
nor U9151 (N_9151,N_2121,N_4483);
or U9152 (N_9152,N_4818,N_4183);
nand U9153 (N_9153,N_3342,N_2890);
and U9154 (N_9154,N_2165,N_4251);
nand U9155 (N_9155,N_2774,N_1756);
and U9156 (N_9156,N_3694,N_3422);
nor U9157 (N_9157,N_2259,N_1948);
or U9158 (N_9158,N_4661,N_3851);
and U9159 (N_9159,N_4515,N_2820);
nand U9160 (N_9160,N_2103,N_626);
and U9161 (N_9161,N_1955,N_535);
nor U9162 (N_9162,N_894,N_2919);
or U9163 (N_9163,N_3899,N_1016);
nor U9164 (N_9164,N_3592,N_770);
nand U9165 (N_9165,N_2664,N_3574);
nor U9166 (N_9166,N_4601,N_484);
or U9167 (N_9167,N_2493,N_3229);
xnor U9168 (N_9168,N_1707,N_4329);
nor U9169 (N_9169,N_4731,N_3940);
nand U9170 (N_9170,N_4713,N_916);
nor U9171 (N_9171,N_4610,N_913);
nand U9172 (N_9172,N_1568,N_30);
or U9173 (N_9173,N_4373,N_1704);
nand U9174 (N_9174,N_1937,N_4071);
nor U9175 (N_9175,N_854,N_1817);
and U9176 (N_9176,N_1875,N_4968);
and U9177 (N_9177,N_4162,N_2922);
and U9178 (N_9178,N_3790,N_4890);
nor U9179 (N_9179,N_144,N_1590);
nand U9180 (N_9180,N_3510,N_746);
nor U9181 (N_9181,N_3016,N_698);
and U9182 (N_9182,N_113,N_3678);
nor U9183 (N_9183,N_4924,N_2860);
nand U9184 (N_9184,N_868,N_2005);
xnor U9185 (N_9185,N_4528,N_1177);
or U9186 (N_9186,N_175,N_1884);
and U9187 (N_9187,N_1279,N_2012);
xor U9188 (N_9188,N_2738,N_3327);
and U9189 (N_9189,N_666,N_2282);
or U9190 (N_9190,N_363,N_1979);
nand U9191 (N_9191,N_1557,N_890);
or U9192 (N_9192,N_602,N_2850);
nand U9193 (N_9193,N_4547,N_4766);
nand U9194 (N_9194,N_3260,N_3865);
nand U9195 (N_9195,N_1359,N_4570);
and U9196 (N_9196,N_2230,N_7);
nand U9197 (N_9197,N_4407,N_1616);
and U9198 (N_9198,N_908,N_784);
nand U9199 (N_9199,N_2487,N_4615);
nand U9200 (N_9200,N_2206,N_4512);
or U9201 (N_9201,N_2879,N_4994);
and U9202 (N_9202,N_4635,N_662);
nand U9203 (N_9203,N_2867,N_4190);
nor U9204 (N_9204,N_2320,N_3813);
or U9205 (N_9205,N_3445,N_2095);
nand U9206 (N_9206,N_4785,N_3212);
or U9207 (N_9207,N_4776,N_2233);
nor U9208 (N_9208,N_4123,N_3373);
nor U9209 (N_9209,N_2131,N_805);
and U9210 (N_9210,N_2298,N_4391);
or U9211 (N_9211,N_4692,N_2963);
nand U9212 (N_9212,N_3974,N_1060);
nand U9213 (N_9213,N_1291,N_1039);
nor U9214 (N_9214,N_680,N_1186);
and U9215 (N_9215,N_2434,N_1443);
or U9216 (N_9216,N_1186,N_2771);
and U9217 (N_9217,N_1405,N_1943);
or U9218 (N_9218,N_426,N_2221);
and U9219 (N_9219,N_940,N_3522);
nor U9220 (N_9220,N_2408,N_4716);
or U9221 (N_9221,N_1400,N_3122);
and U9222 (N_9222,N_2897,N_764);
and U9223 (N_9223,N_735,N_1991);
or U9224 (N_9224,N_2004,N_1046);
and U9225 (N_9225,N_1666,N_4732);
or U9226 (N_9226,N_3229,N_3606);
nand U9227 (N_9227,N_828,N_4576);
or U9228 (N_9228,N_399,N_1260);
or U9229 (N_9229,N_4671,N_1148);
nor U9230 (N_9230,N_3521,N_92);
and U9231 (N_9231,N_1891,N_799);
nor U9232 (N_9232,N_1434,N_527);
and U9233 (N_9233,N_878,N_739);
nor U9234 (N_9234,N_3115,N_2454);
and U9235 (N_9235,N_2273,N_4159);
nor U9236 (N_9236,N_155,N_4950);
nor U9237 (N_9237,N_1429,N_4862);
or U9238 (N_9238,N_415,N_4182);
nor U9239 (N_9239,N_3596,N_758);
or U9240 (N_9240,N_2590,N_2458);
nand U9241 (N_9241,N_2433,N_1831);
or U9242 (N_9242,N_703,N_3440);
or U9243 (N_9243,N_39,N_3311);
nand U9244 (N_9244,N_74,N_3421);
or U9245 (N_9245,N_2351,N_3129);
nand U9246 (N_9246,N_2564,N_796);
and U9247 (N_9247,N_4809,N_3205);
nand U9248 (N_9248,N_3739,N_1294);
nand U9249 (N_9249,N_982,N_3370);
nor U9250 (N_9250,N_679,N_837);
nor U9251 (N_9251,N_3066,N_503);
nor U9252 (N_9252,N_978,N_2812);
xor U9253 (N_9253,N_4362,N_2699);
and U9254 (N_9254,N_4085,N_3403);
nand U9255 (N_9255,N_380,N_3493);
nand U9256 (N_9256,N_4686,N_1730);
and U9257 (N_9257,N_1404,N_883);
nor U9258 (N_9258,N_1439,N_4496);
and U9259 (N_9259,N_3184,N_3107);
nand U9260 (N_9260,N_1304,N_2759);
nor U9261 (N_9261,N_4877,N_984);
and U9262 (N_9262,N_3377,N_957);
and U9263 (N_9263,N_1685,N_2135);
nand U9264 (N_9264,N_990,N_2213);
nand U9265 (N_9265,N_785,N_3574);
nor U9266 (N_9266,N_70,N_806);
or U9267 (N_9267,N_192,N_2484);
nand U9268 (N_9268,N_1818,N_1309);
and U9269 (N_9269,N_4930,N_4673);
xor U9270 (N_9270,N_845,N_2530);
nor U9271 (N_9271,N_3080,N_1517);
and U9272 (N_9272,N_1455,N_2088);
and U9273 (N_9273,N_2703,N_4411);
nor U9274 (N_9274,N_4059,N_3818);
nor U9275 (N_9275,N_4981,N_977);
nand U9276 (N_9276,N_4747,N_4263);
nor U9277 (N_9277,N_4938,N_1026);
and U9278 (N_9278,N_3027,N_4340);
and U9279 (N_9279,N_1115,N_2293);
and U9280 (N_9280,N_2625,N_3915);
nor U9281 (N_9281,N_1333,N_3088);
or U9282 (N_9282,N_2360,N_3325);
or U9283 (N_9283,N_1345,N_4420);
nand U9284 (N_9284,N_2070,N_3091);
nor U9285 (N_9285,N_3943,N_4086);
or U9286 (N_9286,N_1408,N_2541);
and U9287 (N_9287,N_2806,N_1303);
or U9288 (N_9288,N_4177,N_1766);
nor U9289 (N_9289,N_2102,N_592);
nor U9290 (N_9290,N_1773,N_1786);
nand U9291 (N_9291,N_4471,N_4858);
nor U9292 (N_9292,N_4131,N_408);
or U9293 (N_9293,N_1726,N_3525);
or U9294 (N_9294,N_3984,N_610);
or U9295 (N_9295,N_4232,N_320);
and U9296 (N_9296,N_128,N_3021);
nor U9297 (N_9297,N_3765,N_2599);
and U9298 (N_9298,N_3826,N_711);
or U9299 (N_9299,N_4804,N_4556);
or U9300 (N_9300,N_1888,N_734);
nor U9301 (N_9301,N_4477,N_4855);
and U9302 (N_9302,N_2708,N_2619);
nand U9303 (N_9303,N_4808,N_3505);
or U9304 (N_9304,N_581,N_973);
nand U9305 (N_9305,N_3562,N_566);
nand U9306 (N_9306,N_2893,N_3201);
and U9307 (N_9307,N_3589,N_1105);
or U9308 (N_9308,N_3332,N_4865);
nor U9309 (N_9309,N_1093,N_4865);
nand U9310 (N_9310,N_4023,N_3460);
nor U9311 (N_9311,N_1779,N_3420);
nand U9312 (N_9312,N_4538,N_2324);
nand U9313 (N_9313,N_3028,N_1421);
and U9314 (N_9314,N_1857,N_2895);
nor U9315 (N_9315,N_1612,N_4104);
nand U9316 (N_9316,N_4739,N_3098);
and U9317 (N_9317,N_2302,N_4948);
nor U9318 (N_9318,N_4506,N_1668);
or U9319 (N_9319,N_2272,N_4992);
nand U9320 (N_9320,N_1868,N_531);
nand U9321 (N_9321,N_23,N_432);
nor U9322 (N_9322,N_3293,N_4905);
nand U9323 (N_9323,N_4053,N_4673);
and U9324 (N_9324,N_656,N_1550);
or U9325 (N_9325,N_230,N_4085);
nor U9326 (N_9326,N_1424,N_2039);
nand U9327 (N_9327,N_450,N_4855);
or U9328 (N_9328,N_3919,N_3052);
nor U9329 (N_9329,N_4838,N_3518);
nor U9330 (N_9330,N_4386,N_3335);
and U9331 (N_9331,N_1774,N_436);
and U9332 (N_9332,N_1759,N_522);
nand U9333 (N_9333,N_4066,N_2743);
and U9334 (N_9334,N_3397,N_30);
or U9335 (N_9335,N_2415,N_1190);
or U9336 (N_9336,N_2752,N_2571);
and U9337 (N_9337,N_4935,N_1938);
or U9338 (N_9338,N_1685,N_804);
nand U9339 (N_9339,N_4648,N_3261);
or U9340 (N_9340,N_4498,N_1852);
and U9341 (N_9341,N_530,N_120);
nand U9342 (N_9342,N_2108,N_191);
or U9343 (N_9343,N_570,N_2546);
nor U9344 (N_9344,N_344,N_2856);
and U9345 (N_9345,N_1505,N_2977);
nor U9346 (N_9346,N_4466,N_929);
and U9347 (N_9347,N_4923,N_3401);
or U9348 (N_9348,N_1831,N_3360);
or U9349 (N_9349,N_4946,N_3941);
nand U9350 (N_9350,N_2303,N_496);
nand U9351 (N_9351,N_3909,N_3214);
nand U9352 (N_9352,N_2501,N_1327);
or U9353 (N_9353,N_3063,N_4916);
nor U9354 (N_9354,N_1626,N_1531);
nor U9355 (N_9355,N_4757,N_952);
nor U9356 (N_9356,N_1437,N_4814);
nor U9357 (N_9357,N_2246,N_2771);
or U9358 (N_9358,N_1181,N_2301);
nand U9359 (N_9359,N_2513,N_4666);
or U9360 (N_9360,N_2340,N_3797);
and U9361 (N_9361,N_3103,N_3484);
and U9362 (N_9362,N_3497,N_4771);
nor U9363 (N_9363,N_3663,N_2393);
and U9364 (N_9364,N_2826,N_4914);
nor U9365 (N_9365,N_667,N_2825);
and U9366 (N_9366,N_4325,N_2777);
nor U9367 (N_9367,N_4840,N_3031);
or U9368 (N_9368,N_2453,N_31);
or U9369 (N_9369,N_1078,N_3077);
and U9370 (N_9370,N_4665,N_3012);
nor U9371 (N_9371,N_4902,N_2770);
or U9372 (N_9372,N_4112,N_3877);
or U9373 (N_9373,N_3327,N_3897);
or U9374 (N_9374,N_3607,N_2576);
nand U9375 (N_9375,N_4865,N_2511);
or U9376 (N_9376,N_385,N_3275);
and U9377 (N_9377,N_4509,N_2495);
nor U9378 (N_9378,N_2467,N_609);
nor U9379 (N_9379,N_1451,N_1414);
and U9380 (N_9380,N_2894,N_4919);
nor U9381 (N_9381,N_3117,N_1048);
and U9382 (N_9382,N_3573,N_1331);
or U9383 (N_9383,N_36,N_693);
and U9384 (N_9384,N_3238,N_1658);
nand U9385 (N_9385,N_3004,N_3238);
or U9386 (N_9386,N_3802,N_1815);
nand U9387 (N_9387,N_1815,N_3216);
or U9388 (N_9388,N_1421,N_4599);
nand U9389 (N_9389,N_2259,N_1274);
nand U9390 (N_9390,N_1318,N_2199);
or U9391 (N_9391,N_3333,N_4158);
and U9392 (N_9392,N_1023,N_1206);
or U9393 (N_9393,N_700,N_4251);
and U9394 (N_9394,N_2025,N_2328);
or U9395 (N_9395,N_4096,N_2186);
and U9396 (N_9396,N_441,N_3129);
or U9397 (N_9397,N_4631,N_580);
and U9398 (N_9398,N_4390,N_1275);
and U9399 (N_9399,N_3731,N_1942);
nand U9400 (N_9400,N_4664,N_4493);
or U9401 (N_9401,N_3630,N_3446);
and U9402 (N_9402,N_4711,N_4244);
or U9403 (N_9403,N_836,N_3931);
nand U9404 (N_9404,N_1733,N_4773);
and U9405 (N_9405,N_2403,N_4798);
nor U9406 (N_9406,N_3928,N_1265);
or U9407 (N_9407,N_533,N_4909);
or U9408 (N_9408,N_1267,N_848);
nor U9409 (N_9409,N_345,N_2917);
nand U9410 (N_9410,N_2941,N_4428);
nor U9411 (N_9411,N_289,N_3269);
or U9412 (N_9412,N_4040,N_4128);
nand U9413 (N_9413,N_545,N_1467);
xnor U9414 (N_9414,N_4856,N_1616);
nor U9415 (N_9415,N_1374,N_3946);
nor U9416 (N_9416,N_3889,N_2158);
nor U9417 (N_9417,N_4880,N_1407);
or U9418 (N_9418,N_2815,N_490);
and U9419 (N_9419,N_1393,N_2164);
or U9420 (N_9420,N_2970,N_2460);
and U9421 (N_9421,N_3014,N_2457);
nand U9422 (N_9422,N_941,N_2551);
nor U9423 (N_9423,N_2378,N_3601);
nand U9424 (N_9424,N_928,N_2671);
nand U9425 (N_9425,N_3898,N_1147);
nor U9426 (N_9426,N_1033,N_217);
and U9427 (N_9427,N_3555,N_791);
and U9428 (N_9428,N_3584,N_1364);
nand U9429 (N_9429,N_2364,N_2119);
nor U9430 (N_9430,N_1956,N_2461);
nand U9431 (N_9431,N_745,N_1967);
nor U9432 (N_9432,N_4760,N_827);
and U9433 (N_9433,N_360,N_4010);
nand U9434 (N_9434,N_610,N_245);
and U9435 (N_9435,N_4831,N_1953);
xnor U9436 (N_9436,N_3903,N_53);
nand U9437 (N_9437,N_1544,N_999);
or U9438 (N_9438,N_2587,N_169);
or U9439 (N_9439,N_1144,N_4839);
nor U9440 (N_9440,N_2680,N_3593);
or U9441 (N_9441,N_3366,N_4171);
and U9442 (N_9442,N_317,N_50);
nand U9443 (N_9443,N_4634,N_2145);
nor U9444 (N_9444,N_45,N_4275);
or U9445 (N_9445,N_4324,N_1760);
and U9446 (N_9446,N_2924,N_1090);
nor U9447 (N_9447,N_2803,N_1779);
nand U9448 (N_9448,N_934,N_2363);
nor U9449 (N_9449,N_790,N_2903);
and U9450 (N_9450,N_1177,N_680);
nand U9451 (N_9451,N_611,N_3893);
and U9452 (N_9452,N_3137,N_3976);
nor U9453 (N_9453,N_3578,N_2170);
and U9454 (N_9454,N_3751,N_782);
nand U9455 (N_9455,N_997,N_1832);
or U9456 (N_9456,N_2570,N_4970);
or U9457 (N_9457,N_4736,N_4157);
or U9458 (N_9458,N_4571,N_4141);
or U9459 (N_9459,N_3301,N_794);
and U9460 (N_9460,N_716,N_3135);
nor U9461 (N_9461,N_3882,N_3875);
xor U9462 (N_9462,N_2731,N_122);
and U9463 (N_9463,N_4246,N_1099);
nand U9464 (N_9464,N_3740,N_2346);
nand U9465 (N_9465,N_242,N_3866);
and U9466 (N_9466,N_4862,N_1150);
nor U9467 (N_9467,N_4532,N_4924);
nor U9468 (N_9468,N_4992,N_2761);
nand U9469 (N_9469,N_3050,N_2451);
or U9470 (N_9470,N_4905,N_326);
or U9471 (N_9471,N_662,N_1198);
or U9472 (N_9472,N_3554,N_979);
and U9473 (N_9473,N_3462,N_1353);
nor U9474 (N_9474,N_1600,N_2039);
nand U9475 (N_9475,N_3541,N_4127);
and U9476 (N_9476,N_2858,N_1189);
nor U9477 (N_9477,N_1163,N_4015);
or U9478 (N_9478,N_1077,N_214);
or U9479 (N_9479,N_751,N_2374);
nand U9480 (N_9480,N_1294,N_4245);
or U9481 (N_9481,N_4543,N_1811);
nand U9482 (N_9482,N_2094,N_3053);
or U9483 (N_9483,N_10,N_962);
and U9484 (N_9484,N_2430,N_4373);
or U9485 (N_9485,N_2358,N_4043);
nor U9486 (N_9486,N_1116,N_1024);
nor U9487 (N_9487,N_968,N_2287);
nor U9488 (N_9488,N_3657,N_1091);
and U9489 (N_9489,N_4236,N_3798);
nor U9490 (N_9490,N_2420,N_3937);
or U9491 (N_9491,N_4417,N_573);
and U9492 (N_9492,N_4378,N_4655);
and U9493 (N_9493,N_4059,N_1928);
xnor U9494 (N_9494,N_212,N_4701);
nor U9495 (N_9495,N_111,N_2527);
or U9496 (N_9496,N_3867,N_4347);
and U9497 (N_9497,N_178,N_3267);
nor U9498 (N_9498,N_1718,N_1018);
nand U9499 (N_9499,N_1804,N_2895);
nor U9500 (N_9500,N_148,N_3020);
xor U9501 (N_9501,N_1854,N_2314);
and U9502 (N_9502,N_4164,N_2011);
or U9503 (N_9503,N_925,N_4689);
nor U9504 (N_9504,N_4995,N_1801);
and U9505 (N_9505,N_4171,N_4833);
nor U9506 (N_9506,N_1629,N_1804);
and U9507 (N_9507,N_2072,N_4025);
nor U9508 (N_9508,N_1652,N_3232);
nand U9509 (N_9509,N_4538,N_3617);
nand U9510 (N_9510,N_3117,N_1885);
nor U9511 (N_9511,N_4106,N_2991);
or U9512 (N_9512,N_246,N_2087);
nand U9513 (N_9513,N_4684,N_3953);
nand U9514 (N_9514,N_3509,N_1273);
nand U9515 (N_9515,N_2100,N_1738);
nand U9516 (N_9516,N_989,N_4268);
nor U9517 (N_9517,N_4807,N_574);
nand U9518 (N_9518,N_1016,N_2356);
or U9519 (N_9519,N_2368,N_344);
nor U9520 (N_9520,N_3703,N_876);
nand U9521 (N_9521,N_3316,N_2782);
nor U9522 (N_9522,N_4769,N_3692);
xor U9523 (N_9523,N_2651,N_1781);
or U9524 (N_9524,N_3008,N_1439);
and U9525 (N_9525,N_1191,N_4897);
and U9526 (N_9526,N_919,N_4839);
and U9527 (N_9527,N_4559,N_1425);
or U9528 (N_9528,N_4410,N_3507);
nor U9529 (N_9529,N_1081,N_572);
nand U9530 (N_9530,N_4437,N_3863);
or U9531 (N_9531,N_4525,N_1529);
nand U9532 (N_9532,N_4560,N_4883);
or U9533 (N_9533,N_2224,N_1919);
nand U9534 (N_9534,N_4338,N_1253);
and U9535 (N_9535,N_594,N_2632);
and U9536 (N_9536,N_3308,N_1967);
or U9537 (N_9537,N_4124,N_3019);
nor U9538 (N_9538,N_1505,N_4735);
nor U9539 (N_9539,N_1340,N_3732);
nand U9540 (N_9540,N_1158,N_28);
nand U9541 (N_9541,N_1968,N_130);
nor U9542 (N_9542,N_4917,N_4933);
or U9543 (N_9543,N_1921,N_393);
or U9544 (N_9544,N_4417,N_933);
and U9545 (N_9545,N_947,N_3878);
or U9546 (N_9546,N_4724,N_1945);
nand U9547 (N_9547,N_7,N_2779);
or U9548 (N_9548,N_4292,N_4601);
or U9549 (N_9549,N_4302,N_1806);
and U9550 (N_9550,N_2257,N_1767);
nor U9551 (N_9551,N_3767,N_4890);
or U9552 (N_9552,N_4704,N_2383);
nor U9553 (N_9553,N_4562,N_4728);
and U9554 (N_9554,N_4997,N_3568);
nor U9555 (N_9555,N_2476,N_3531);
and U9556 (N_9556,N_4925,N_1249);
nand U9557 (N_9557,N_2075,N_3332);
and U9558 (N_9558,N_4407,N_4415);
nor U9559 (N_9559,N_787,N_1194);
nor U9560 (N_9560,N_1600,N_3282);
and U9561 (N_9561,N_3951,N_3343);
nor U9562 (N_9562,N_1347,N_1360);
nor U9563 (N_9563,N_1033,N_4005);
or U9564 (N_9564,N_4937,N_2186);
and U9565 (N_9565,N_3402,N_4151);
and U9566 (N_9566,N_2958,N_4394);
and U9567 (N_9567,N_750,N_4262);
and U9568 (N_9568,N_882,N_4820);
nand U9569 (N_9569,N_1942,N_517);
nor U9570 (N_9570,N_3213,N_1131);
or U9571 (N_9571,N_413,N_898);
nand U9572 (N_9572,N_4131,N_2312);
nor U9573 (N_9573,N_3864,N_1340);
or U9574 (N_9574,N_4617,N_2964);
or U9575 (N_9575,N_658,N_3912);
or U9576 (N_9576,N_3040,N_2243);
nand U9577 (N_9577,N_1544,N_4866);
nor U9578 (N_9578,N_3028,N_3234);
nand U9579 (N_9579,N_4719,N_2703);
nand U9580 (N_9580,N_458,N_2570);
nand U9581 (N_9581,N_3769,N_724);
and U9582 (N_9582,N_347,N_3862);
xnor U9583 (N_9583,N_2431,N_1827);
and U9584 (N_9584,N_471,N_4224);
nand U9585 (N_9585,N_2623,N_823);
nand U9586 (N_9586,N_585,N_782);
nor U9587 (N_9587,N_2953,N_3788);
nor U9588 (N_9588,N_4973,N_1222);
or U9589 (N_9589,N_1972,N_1839);
nand U9590 (N_9590,N_2250,N_2270);
or U9591 (N_9591,N_2941,N_2133);
nor U9592 (N_9592,N_3935,N_2039);
and U9593 (N_9593,N_317,N_2873);
or U9594 (N_9594,N_806,N_2522);
nor U9595 (N_9595,N_4626,N_2645);
nor U9596 (N_9596,N_245,N_630);
nor U9597 (N_9597,N_2477,N_188);
and U9598 (N_9598,N_1458,N_2190);
nand U9599 (N_9599,N_3483,N_2106);
nor U9600 (N_9600,N_4173,N_4610);
or U9601 (N_9601,N_3435,N_3107);
or U9602 (N_9602,N_2852,N_1547);
nor U9603 (N_9603,N_3731,N_1100);
or U9604 (N_9604,N_2573,N_296);
nand U9605 (N_9605,N_2694,N_2843);
nand U9606 (N_9606,N_3809,N_3232);
nand U9607 (N_9607,N_4206,N_2429);
nor U9608 (N_9608,N_2705,N_668);
or U9609 (N_9609,N_3181,N_4234);
and U9610 (N_9610,N_4505,N_1685);
nor U9611 (N_9611,N_2460,N_4399);
or U9612 (N_9612,N_518,N_1670);
nand U9613 (N_9613,N_2582,N_3138);
nand U9614 (N_9614,N_4832,N_3956);
and U9615 (N_9615,N_3826,N_632);
nor U9616 (N_9616,N_3288,N_2028);
or U9617 (N_9617,N_41,N_2616);
nor U9618 (N_9618,N_2788,N_925);
nor U9619 (N_9619,N_1562,N_4660);
and U9620 (N_9620,N_3557,N_3793);
nand U9621 (N_9621,N_2415,N_1484);
nor U9622 (N_9622,N_699,N_147);
nand U9623 (N_9623,N_2507,N_1718);
nand U9624 (N_9624,N_516,N_3207);
or U9625 (N_9625,N_760,N_3345);
nand U9626 (N_9626,N_3495,N_480);
and U9627 (N_9627,N_4570,N_3437);
or U9628 (N_9628,N_3624,N_907);
nand U9629 (N_9629,N_4793,N_2512);
nor U9630 (N_9630,N_2850,N_1865);
nand U9631 (N_9631,N_4760,N_2667);
nand U9632 (N_9632,N_2068,N_4918);
or U9633 (N_9633,N_1702,N_4692);
or U9634 (N_9634,N_4811,N_2533);
nor U9635 (N_9635,N_2508,N_783);
nor U9636 (N_9636,N_125,N_3424);
nor U9637 (N_9637,N_90,N_80);
and U9638 (N_9638,N_1673,N_2464);
nor U9639 (N_9639,N_4567,N_777);
and U9640 (N_9640,N_1120,N_4110);
or U9641 (N_9641,N_4735,N_2444);
nand U9642 (N_9642,N_1695,N_402);
and U9643 (N_9643,N_2035,N_4009);
or U9644 (N_9644,N_4541,N_913);
nand U9645 (N_9645,N_106,N_2628);
and U9646 (N_9646,N_3284,N_2051);
nand U9647 (N_9647,N_761,N_1930);
or U9648 (N_9648,N_2893,N_1182);
nor U9649 (N_9649,N_4118,N_2991);
nand U9650 (N_9650,N_239,N_3980);
and U9651 (N_9651,N_4553,N_1359);
or U9652 (N_9652,N_4042,N_3197);
or U9653 (N_9653,N_4310,N_737);
and U9654 (N_9654,N_3586,N_936);
nor U9655 (N_9655,N_129,N_1450);
xor U9656 (N_9656,N_3477,N_4264);
nand U9657 (N_9657,N_2246,N_1706);
nand U9658 (N_9658,N_1900,N_773);
nor U9659 (N_9659,N_2104,N_2391);
nor U9660 (N_9660,N_1623,N_2264);
and U9661 (N_9661,N_378,N_4903);
nor U9662 (N_9662,N_3016,N_741);
nand U9663 (N_9663,N_3152,N_1404);
nand U9664 (N_9664,N_1085,N_421);
nor U9665 (N_9665,N_14,N_2621);
nor U9666 (N_9666,N_773,N_869);
nor U9667 (N_9667,N_4529,N_2293);
or U9668 (N_9668,N_1755,N_3529);
and U9669 (N_9669,N_740,N_1325);
nor U9670 (N_9670,N_2749,N_1762);
and U9671 (N_9671,N_3365,N_2907);
nand U9672 (N_9672,N_966,N_2859);
or U9673 (N_9673,N_4836,N_1958);
nor U9674 (N_9674,N_228,N_1862);
nor U9675 (N_9675,N_575,N_4787);
nand U9676 (N_9676,N_4046,N_3401);
or U9677 (N_9677,N_4328,N_2210);
nand U9678 (N_9678,N_4209,N_1202);
nor U9679 (N_9679,N_25,N_4390);
or U9680 (N_9680,N_3841,N_3616);
nor U9681 (N_9681,N_950,N_4554);
and U9682 (N_9682,N_4412,N_3058);
or U9683 (N_9683,N_1037,N_4463);
and U9684 (N_9684,N_2602,N_2270);
and U9685 (N_9685,N_1141,N_4558);
or U9686 (N_9686,N_696,N_3523);
nand U9687 (N_9687,N_4109,N_1354);
nor U9688 (N_9688,N_1424,N_3068);
and U9689 (N_9689,N_1939,N_341);
and U9690 (N_9690,N_877,N_3014);
nor U9691 (N_9691,N_923,N_827);
nor U9692 (N_9692,N_2377,N_2141);
nand U9693 (N_9693,N_4623,N_4252);
nand U9694 (N_9694,N_2525,N_4972);
or U9695 (N_9695,N_1478,N_3399);
nor U9696 (N_9696,N_1747,N_360);
nand U9697 (N_9697,N_4768,N_3678);
and U9698 (N_9698,N_3569,N_3140);
or U9699 (N_9699,N_2017,N_4460);
xor U9700 (N_9700,N_2993,N_2669);
or U9701 (N_9701,N_1275,N_1435);
or U9702 (N_9702,N_3677,N_1431);
or U9703 (N_9703,N_261,N_2177);
and U9704 (N_9704,N_1232,N_3048);
or U9705 (N_9705,N_3737,N_4917);
and U9706 (N_9706,N_2000,N_1967);
nor U9707 (N_9707,N_2426,N_4597);
and U9708 (N_9708,N_2387,N_2910);
nand U9709 (N_9709,N_842,N_70);
and U9710 (N_9710,N_1481,N_4440);
and U9711 (N_9711,N_3326,N_2581);
or U9712 (N_9712,N_589,N_2839);
and U9713 (N_9713,N_4898,N_4077);
nand U9714 (N_9714,N_3835,N_260);
or U9715 (N_9715,N_2592,N_3755);
or U9716 (N_9716,N_2896,N_249);
or U9717 (N_9717,N_1431,N_294);
nand U9718 (N_9718,N_1846,N_4938);
or U9719 (N_9719,N_4313,N_1230);
or U9720 (N_9720,N_853,N_1426);
nor U9721 (N_9721,N_295,N_2420);
and U9722 (N_9722,N_3275,N_32);
or U9723 (N_9723,N_1377,N_2904);
xor U9724 (N_9724,N_4344,N_4719);
nand U9725 (N_9725,N_3273,N_2027);
nor U9726 (N_9726,N_2903,N_1605);
or U9727 (N_9727,N_4676,N_2387);
or U9728 (N_9728,N_3888,N_3470);
nor U9729 (N_9729,N_1194,N_4874);
nor U9730 (N_9730,N_2993,N_4544);
or U9731 (N_9731,N_691,N_1964);
nor U9732 (N_9732,N_2451,N_4640);
nor U9733 (N_9733,N_3665,N_1846);
and U9734 (N_9734,N_3336,N_3839);
and U9735 (N_9735,N_3969,N_3892);
or U9736 (N_9736,N_64,N_4301);
nand U9737 (N_9737,N_4948,N_3984);
nand U9738 (N_9738,N_4415,N_3474);
nor U9739 (N_9739,N_3429,N_4097);
or U9740 (N_9740,N_22,N_4963);
nor U9741 (N_9741,N_4641,N_2345);
or U9742 (N_9742,N_561,N_1616);
nand U9743 (N_9743,N_2893,N_2799);
xnor U9744 (N_9744,N_2588,N_4097);
or U9745 (N_9745,N_2538,N_1627);
nand U9746 (N_9746,N_689,N_1511);
nand U9747 (N_9747,N_1007,N_646);
nand U9748 (N_9748,N_1049,N_2889);
nand U9749 (N_9749,N_3325,N_4087);
nand U9750 (N_9750,N_1840,N_1012);
or U9751 (N_9751,N_4027,N_2931);
or U9752 (N_9752,N_1840,N_197);
nand U9753 (N_9753,N_4394,N_2852);
or U9754 (N_9754,N_2294,N_1265);
and U9755 (N_9755,N_538,N_2153);
nand U9756 (N_9756,N_2388,N_1706);
or U9757 (N_9757,N_3924,N_4216);
or U9758 (N_9758,N_4984,N_3441);
or U9759 (N_9759,N_867,N_4715);
and U9760 (N_9760,N_740,N_3102);
and U9761 (N_9761,N_3616,N_2980);
and U9762 (N_9762,N_1742,N_2081);
or U9763 (N_9763,N_4086,N_3615);
nor U9764 (N_9764,N_4376,N_4483);
or U9765 (N_9765,N_3732,N_1463);
nor U9766 (N_9766,N_3171,N_1378);
or U9767 (N_9767,N_3719,N_616);
nor U9768 (N_9768,N_35,N_2214);
or U9769 (N_9769,N_2267,N_4198);
or U9770 (N_9770,N_700,N_4283);
nand U9771 (N_9771,N_946,N_3615);
nand U9772 (N_9772,N_1110,N_1794);
nor U9773 (N_9773,N_3784,N_2454);
nand U9774 (N_9774,N_1841,N_431);
or U9775 (N_9775,N_2754,N_4588);
nor U9776 (N_9776,N_141,N_1720);
nand U9777 (N_9777,N_1459,N_423);
or U9778 (N_9778,N_381,N_395);
or U9779 (N_9779,N_3398,N_2646);
nand U9780 (N_9780,N_4951,N_15);
and U9781 (N_9781,N_4496,N_4783);
nor U9782 (N_9782,N_1245,N_1560);
and U9783 (N_9783,N_3078,N_1995);
and U9784 (N_9784,N_4199,N_2877);
or U9785 (N_9785,N_452,N_900);
nand U9786 (N_9786,N_1386,N_1775);
or U9787 (N_9787,N_1875,N_4089);
and U9788 (N_9788,N_2557,N_3128);
or U9789 (N_9789,N_3688,N_4274);
or U9790 (N_9790,N_2426,N_2382);
nor U9791 (N_9791,N_2472,N_4635);
nor U9792 (N_9792,N_1451,N_2609);
nand U9793 (N_9793,N_4030,N_1702);
or U9794 (N_9794,N_2794,N_4737);
nand U9795 (N_9795,N_4367,N_4537);
nor U9796 (N_9796,N_3022,N_1182);
nand U9797 (N_9797,N_1274,N_4086);
and U9798 (N_9798,N_2691,N_3233);
nand U9799 (N_9799,N_816,N_1335);
nor U9800 (N_9800,N_3086,N_4953);
nor U9801 (N_9801,N_4617,N_754);
or U9802 (N_9802,N_1817,N_3294);
nand U9803 (N_9803,N_1608,N_4907);
nand U9804 (N_9804,N_1094,N_1305);
nand U9805 (N_9805,N_1799,N_207);
and U9806 (N_9806,N_2048,N_3719);
and U9807 (N_9807,N_4635,N_4946);
nand U9808 (N_9808,N_1255,N_3206);
or U9809 (N_9809,N_352,N_4862);
xor U9810 (N_9810,N_2806,N_4029);
or U9811 (N_9811,N_3282,N_325);
and U9812 (N_9812,N_4665,N_1641);
nand U9813 (N_9813,N_4069,N_165);
and U9814 (N_9814,N_2129,N_3690);
nor U9815 (N_9815,N_3797,N_2248);
nand U9816 (N_9816,N_584,N_4973);
or U9817 (N_9817,N_815,N_4118);
and U9818 (N_9818,N_76,N_673);
xnor U9819 (N_9819,N_2547,N_2911);
and U9820 (N_9820,N_4034,N_3672);
nand U9821 (N_9821,N_4153,N_1092);
nand U9822 (N_9822,N_4790,N_3170);
nand U9823 (N_9823,N_2981,N_924);
nor U9824 (N_9824,N_1692,N_2710);
nand U9825 (N_9825,N_537,N_4524);
nand U9826 (N_9826,N_2226,N_2066);
or U9827 (N_9827,N_624,N_481);
or U9828 (N_9828,N_3305,N_2834);
nor U9829 (N_9829,N_3319,N_1113);
xor U9830 (N_9830,N_3213,N_1672);
or U9831 (N_9831,N_1978,N_1498);
nand U9832 (N_9832,N_2613,N_4868);
and U9833 (N_9833,N_4202,N_1740);
nor U9834 (N_9834,N_989,N_280);
or U9835 (N_9835,N_4678,N_3891);
nand U9836 (N_9836,N_2327,N_709);
nor U9837 (N_9837,N_3605,N_4053);
nor U9838 (N_9838,N_1841,N_4560);
nand U9839 (N_9839,N_659,N_2435);
and U9840 (N_9840,N_1936,N_810);
and U9841 (N_9841,N_2105,N_2704);
and U9842 (N_9842,N_644,N_2802);
or U9843 (N_9843,N_1714,N_4344);
or U9844 (N_9844,N_827,N_4691);
and U9845 (N_9845,N_674,N_621);
and U9846 (N_9846,N_2295,N_4046);
and U9847 (N_9847,N_3553,N_4189);
or U9848 (N_9848,N_409,N_2750);
and U9849 (N_9849,N_2620,N_1141);
and U9850 (N_9850,N_3680,N_1415);
or U9851 (N_9851,N_2695,N_3286);
nand U9852 (N_9852,N_2709,N_3827);
nand U9853 (N_9853,N_1902,N_4968);
nand U9854 (N_9854,N_481,N_3120);
or U9855 (N_9855,N_3431,N_2888);
or U9856 (N_9856,N_3369,N_4937);
and U9857 (N_9857,N_2888,N_1801);
nor U9858 (N_9858,N_4454,N_2306);
nand U9859 (N_9859,N_4227,N_787);
or U9860 (N_9860,N_1619,N_109);
nor U9861 (N_9861,N_1507,N_4591);
or U9862 (N_9862,N_639,N_3022);
nor U9863 (N_9863,N_1553,N_2843);
or U9864 (N_9864,N_686,N_535);
or U9865 (N_9865,N_1010,N_4531);
or U9866 (N_9866,N_1723,N_1041);
nand U9867 (N_9867,N_4498,N_4141);
xnor U9868 (N_9868,N_4503,N_4418);
nor U9869 (N_9869,N_814,N_3422);
nor U9870 (N_9870,N_736,N_2527);
or U9871 (N_9871,N_4588,N_1924);
nor U9872 (N_9872,N_3741,N_4844);
nor U9873 (N_9873,N_2314,N_19);
or U9874 (N_9874,N_4211,N_201);
or U9875 (N_9875,N_519,N_4973);
nor U9876 (N_9876,N_3577,N_2140);
or U9877 (N_9877,N_3222,N_178);
and U9878 (N_9878,N_321,N_2216);
or U9879 (N_9879,N_1653,N_4086);
nor U9880 (N_9880,N_2392,N_3593);
nor U9881 (N_9881,N_2603,N_4731);
or U9882 (N_9882,N_4747,N_1788);
or U9883 (N_9883,N_1854,N_4839);
and U9884 (N_9884,N_4519,N_2860);
nand U9885 (N_9885,N_3163,N_947);
nand U9886 (N_9886,N_4878,N_1858);
and U9887 (N_9887,N_2252,N_3430);
or U9888 (N_9888,N_4552,N_3840);
or U9889 (N_9889,N_4266,N_3882);
nand U9890 (N_9890,N_4038,N_3301);
nor U9891 (N_9891,N_4482,N_4633);
nand U9892 (N_9892,N_215,N_74);
nand U9893 (N_9893,N_3427,N_4728);
nand U9894 (N_9894,N_1343,N_4480);
nor U9895 (N_9895,N_383,N_3603);
nand U9896 (N_9896,N_1152,N_568);
and U9897 (N_9897,N_3221,N_2307);
and U9898 (N_9898,N_1693,N_3492);
or U9899 (N_9899,N_1146,N_1982);
nand U9900 (N_9900,N_1208,N_240);
nor U9901 (N_9901,N_2396,N_1511);
xnor U9902 (N_9902,N_1875,N_664);
nand U9903 (N_9903,N_1935,N_84);
or U9904 (N_9904,N_922,N_2352);
nand U9905 (N_9905,N_356,N_2461);
or U9906 (N_9906,N_833,N_3260);
nor U9907 (N_9907,N_1410,N_4410);
nor U9908 (N_9908,N_3054,N_4565);
nand U9909 (N_9909,N_4314,N_218);
nor U9910 (N_9910,N_1670,N_2695);
nor U9911 (N_9911,N_4085,N_1468);
or U9912 (N_9912,N_1637,N_2856);
nand U9913 (N_9913,N_4300,N_4932);
and U9914 (N_9914,N_3531,N_580);
or U9915 (N_9915,N_3761,N_1544);
nor U9916 (N_9916,N_1207,N_4082);
nor U9917 (N_9917,N_48,N_2819);
nor U9918 (N_9918,N_29,N_1025);
or U9919 (N_9919,N_280,N_1935);
nor U9920 (N_9920,N_1954,N_4585);
or U9921 (N_9921,N_422,N_2100);
nor U9922 (N_9922,N_3132,N_2503);
nand U9923 (N_9923,N_4818,N_4647);
and U9924 (N_9924,N_175,N_2613);
nand U9925 (N_9925,N_1925,N_176);
and U9926 (N_9926,N_2697,N_3738);
or U9927 (N_9927,N_4944,N_3717);
or U9928 (N_9928,N_2200,N_231);
nand U9929 (N_9929,N_3441,N_2144);
nor U9930 (N_9930,N_4987,N_223);
nand U9931 (N_9931,N_4132,N_4964);
and U9932 (N_9932,N_3173,N_4512);
nor U9933 (N_9933,N_4000,N_2195);
and U9934 (N_9934,N_4492,N_69);
nand U9935 (N_9935,N_443,N_1510);
nand U9936 (N_9936,N_1818,N_958);
and U9937 (N_9937,N_3161,N_2412);
nor U9938 (N_9938,N_3594,N_3574);
nand U9939 (N_9939,N_3956,N_3659);
or U9940 (N_9940,N_2958,N_744);
nor U9941 (N_9941,N_3522,N_452);
nor U9942 (N_9942,N_2792,N_348);
or U9943 (N_9943,N_3283,N_2912);
nand U9944 (N_9944,N_3059,N_125);
and U9945 (N_9945,N_4991,N_2270);
nor U9946 (N_9946,N_421,N_965);
or U9947 (N_9947,N_1558,N_2278);
and U9948 (N_9948,N_2022,N_4081);
nand U9949 (N_9949,N_512,N_4361);
nand U9950 (N_9950,N_795,N_3566);
or U9951 (N_9951,N_3528,N_3845);
or U9952 (N_9952,N_2865,N_1560);
nor U9953 (N_9953,N_2964,N_4997);
or U9954 (N_9954,N_506,N_30);
nand U9955 (N_9955,N_3851,N_2908);
nand U9956 (N_9956,N_3244,N_452);
or U9957 (N_9957,N_4937,N_3025);
nor U9958 (N_9958,N_802,N_4358);
and U9959 (N_9959,N_3395,N_4647);
nand U9960 (N_9960,N_974,N_4103);
nor U9961 (N_9961,N_4519,N_316);
or U9962 (N_9962,N_2842,N_3023);
and U9963 (N_9963,N_3472,N_2571);
or U9964 (N_9964,N_4081,N_2271);
and U9965 (N_9965,N_3958,N_3869);
nand U9966 (N_9966,N_4234,N_4952);
nand U9967 (N_9967,N_1223,N_2426);
and U9968 (N_9968,N_4369,N_4231);
nor U9969 (N_9969,N_292,N_3620);
nand U9970 (N_9970,N_4592,N_2110);
and U9971 (N_9971,N_3018,N_4270);
nor U9972 (N_9972,N_3290,N_4302);
or U9973 (N_9973,N_429,N_364);
and U9974 (N_9974,N_2510,N_4834);
nor U9975 (N_9975,N_2460,N_2433);
and U9976 (N_9976,N_2577,N_705);
or U9977 (N_9977,N_208,N_4575);
or U9978 (N_9978,N_3123,N_2778);
and U9979 (N_9979,N_2726,N_4645);
and U9980 (N_9980,N_3186,N_2799);
nand U9981 (N_9981,N_2029,N_770);
nand U9982 (N_9982,N_857,N_184);
or U9983 (N_9983,N_3855,N_2825);
nand U9984 (N_9984,N_287,N_3123);
nor U9985 (N_9985,N_1652,N_1675);
and U9986 (N_9986,N_2412,N_1605);
or U9987 (N_9987,N_2655,N_996);
and U9988 (N_9988,N_3718,N_3725);
or U9989 (N_9989,N_3510,N_2841);
or U9990 (N_9990,N_1722,N_1418);
nand U9991 (N_9991,N_1107,N_4787);
and U9992 (N_9992,N_2777,N_4217);
or U9993 (N_9993,N_1764,N_3571);
and U9994 (N_9994,N_997,N_1427);
or U9995 (N_9995,N_399,N_1673);
nor U9996 (N_9996,N_2738,N_4234);
nand U9997 (N_9997,N_3438,N_2863);
and U9998 (N_9998,N_4837,N_3573);
nor U9999 (N_9999,N_584,N_57);
and U10000 (N_10000,N_9288,N_8970);
nor U10001 (N_10001,N_7421,N_5217);
nand U10002 (N_10002,N_7902,N_7676);
nor U10003 (N_10003,N_9436,N_5313);
and U10004 (N_10004,N_5766,N_8471);
or U10005 (N_10005,N_6558,N_6791);
and U10006 (N_10006,N_8106,N_5604);
nor U10007 (N_10007,N_9695,N_5381);
and U10008 (N_10008,N_7827,N_9928);
and U10009 (N_10009,N_6293,N_7538);
nand U10010 (N_10010,N_7499,N_7179);
nor U10011 (N_10011,N_8846,N_6298);
or U10012 (N_10012,N_6303,N_5938);
nand U10013 (N_10013,N_8632,N_8637);
nor U10014 (N_10014,N_6316,N_7053);
nand U10015 (N_10015,N_9482,N_6081);
and U10016 (N_10016,N_8203,N_8977);
and U10017 (N_10017,N_7699,N_9941);
nand U10018 (N_10018,N_9658,N_7219);
and U10019 (N_10019,N_7960,N_8923);
or U10020 (N_10020,N_8799,N_5507);
nand U10021 (N_10021,N_6227,N_8291);
nor U10022 (N_10022,N_5989,N_5404);
or U10023 (N_10023,N_9652,N_6543);
nand U10024 (N_10024,N_8739,N_6030);
or U10025 (N_10025,N_9660,N_6383);
or U10026 (N_10026,N_8440,N_7974);
nor U10027 (N_10027,N_7181,N_7287);
nor U10028 (N_10028,N_7630,N_7868);
and U10029 (N_10029,N_8925,N_7609);
nor U10030 (N_10030,N_7050,N_9053);
nand U10031 (N_10031,N_5974,N_8720);
or U10032 (N_10032,N_8803,N_7970);
nor U10033 (N_10033,N_6928,N_8378);
nand U10034 (N_10034,N_8123,N_9791);
nand U10035 (N_10035,N_6283,N_5556);
nand U10036 (N_10036,N_7038,N_8549);
and U10037 (N_10037,N_7327,N_9698);
nor U10038 (N_10038,N_5872,N_5657);
and U10039 (N_10039,N_6158,N_8480);
or U10040 (N_10040,N_8772,N_7476);
nand U10041 (N_10041,N_7443,N_5957);
or U10042 (N_10042,N_7469,N_5117);
or U10043 (N_10043,N_7493,N_7062);
nand U10044 (N_10044,N_6003,N_9200);
xnor U10045 (N_10045,N_8577,N_5934);
nand U10046 (N_10046,N_7463,N_6741);
or U10047 (N_10047,N_9082,N_7143);
nand U10048 (N_10048,N_5082,N_9573);
nor U10049 (N_10049,N_7547,N_6175);
and U10050 (N_10050,N_7928,N_9712);
and U10051 (N_10051,N_5294,N_7010);
nor U10052 (N_10052,N_5794,N_8060);
nand U10053 (N_10053,N_7140,N_5401);
and U10054 (N_10054,N_9632,N_8539);
and U10055 (N_10055,N_7404,N_8751);
nor U10056 (N_10056,N_8987,N_8042);
nand U10057 (N_10057,N_9068,N_7718);
nand U10058 (N_10058,N_7317,N_8266);
nor U10059 (N_10059,N_7151,N_7383);
or U10060 (N_10060,N_6872,N_5227);
or U10061 (N_10061,N_8727,N_5838);
nor U10062 (N_10062,N_9372,N_8442);
and U10063 (N_10063,N_9514,N_9891);
nor U10064 (N_10064,N_9285,N_6481);
or U10065 (N_10065,N_9310,N_6955);
and U10066 (N_10066,N_6803,N_5245);
nor U10067 (N_10067,N_8824,N_6944);
and U10068 (N_10068,N_6880,N_8371);
nand U10069 (N_10069,N_5742,N_9459);
nor U10070 (N_10070,N_8244,N_8491);
and U10071 (N_10071,N_7527,N_7119);
or U10072 (N_10072,N_5943,N_5478);
nand U10073 (N_10073,N_5237,N_9052);
or U10074 (N_10074,N_7751,N_7311);
or U10075 (N_10075,N_6152,N_9563);
nor U10076 (N_10076,N_5095,N_8607);
nand U10077 (N_10077,N_5728,N_7516);
and U10078 (N_10078,N_7220,N_6291);
or U10079 (N_10079,N_8761,N_6732);
and U10080 (N_10080,N_8680,N_8779);
and U10081 (N_10081,N_5308,N_6210);
or U10082 (N_10082,N_9401,N_5810);
or U10083 (N_10083,N_8399,N_7435);
nor U10084 (N_10084,N_7703,N_6546);
nor U10085 (N_10085,N_6060,N_8598);
nand U10086 (N_10086,N_5455,N_7820);
nor U10087 (N_10087,N_8307,N_5268);
or U10088 (N_10088,N_7309,N_7821);
nor U10089 (N_10089,N_8974,N_5145);
or U10090 (N_10090,N_5622,N_8520);
or U10091 (N_10091,N_7407,N_7714);
nor U10092 (N_10092,N_9431,N_7056);
or U10093 (N_10093,N_8995,N_5876);
or U10094 (N_10094,N_6666,N_9504);
nand U10095 (N_10095,N_6408,N_7885);
and U10096 (N_10096,N_8855,N_8490);
and U10097 (N_10097,N_9984,N_7625);
and U10098 (N_10098,N_6407,N_8612);
nand U10099 (N_10099,N_7280,N_5012);
or U10100 (N_10100,N_9795,N_6331);
nor U10101 (N_10101,N_5331,N_6179);
nand U10102 (N_10102,N_7526,N_8786);
and U10103 (N_10103,N_8109,N_5707);
and U10104 (N_10104,N_8630,N_6373);
and U10105 (N_10105,N_8650,N_9621);
nor U10106 (N_10106,N_9251,N_9314);
and U10107 (N_10107,N_9510,N_5655);
and U10108 (N_10108,N_9091,N_9432);
and U10109 (N_10109,N_5407,N_5349);
xnor U10110 (N_10110,N_8438,N_7271);
nor U10111 (N_10111,N_6613,N_9766);
nand U10112 (N_10112,N_9533,N_7337);
or U10113 (N_10113,N_6315,N_5521);
or U10114 (N_10114,N_8294,N_7442);
nor U10115 (N_10115,N_8199,N_7835);
or U10116 (N_10116,N_6514,N_6160);
nor U10117 (N_10117,N_6806,N_5686);
nand U10118 (N_10118,N_8578,N_7302);
and U10119 (N_10119,N_5028,N_9722);
nand U10120 (N_10120,N_6345,N_9426);
nor U10121 (N_10121,N_7414,N_5234);
or U10122 (N_10122,N_8516,N_9583);
nor U10123 (N_10123,N_7150,N_9370);
nand U10124 (N_10124,N_6819,N_6773);
or U10125 (N_10125,N_6380,N_5183);
nand U10126 (N_10126,N_9151,N_8777);
nor U10127 (N_10127,N_7784,N_9262);
or U10128 (N_10128,N_5696,N_9168);
and U10129 (N_10129,N_9130,N_5904);
or U10130 (N_10130,N_8953,N_9298);
or U10131 (N_10131,N_8253,N_5474);
nand U10132 (N_10132,N_8104,N_5896);
or U10133 (N_10133,N_7156,N_9815);
and U10134 (N_10134,N_9453,N_7536);
nand U10135 (N_10135,N_7815,N_9341);
and U10136 (N_10136,N_9936,N_5911);
nor U10137 (N_10137,N_5097,N_5466);
or U10138 (N_10138,N_7306,N_6338);
or U10139 (N_10139,N_9065,N_5053);
nand U10140 (N_10140,N_8187,N_9366);
or U10141 (N_10141,N_9116,N_6900);
nor U10142 (N_10142,N_9394,N_9282);
nand U10143 (N_10143,N_6740,N_6846);
and U10144 (N_10144,N_7272,N_5009);
nand U10145 (N_10145,N_6433,N_5491);
nor U10146 (N_10146,N_5787,N_7298);
nand U10147 (N_10147,N_5037,N_5879);
nor U10148 (N_10148,N_7657,N_5855);
and U10149 (N_10149,N_5816,N_9269);
nor U10150 (N_10150,N_5813,N_5506);
and U10151 (N_10151,N_6604,N_7698);
nand U10152 (N_10152,N_6513,N_9931);
nor U10153 (N_10153,N_5475,N_5162);
or U10154 (N_10154,N_7793,N_5251);
nand U10155 (N_10155,N_8069,N_9222);
nand U10156 (N_10156,N_6263,N_5928);
nor U10157 (N_10157,N_6905,N_6082);
nand U10158 (N_10158,N_6930,N_8332);
nand U10159 (N_10159,N_5588,N_7291);
and U10160 (N_10160,N_6190,N_8384);
or U10161 (N_10161,N_6270,N_6463);
nand U10162 (N_10162,N_7859,N_9238);
or U10163 (N_10163,N_5098,N_6568);
and U10164 (N_10164,N_9882,N_8822);
or U10165 (N_10165,N_7637,N_9392);
nor U10166 (N_10166,N_7163,N_6452);
or U10167 (N_10167,N_6685,N_6959);
nand U10168 (N_10168,N_9111,N_5388);
nor U10169 (N_10169,N_6123,N_7899);
nand U10170 (N_10170,N_9989,N_9208);
and U10171 (N_10171,N_9121,N_5607);
nand U10172 (N_10172,N_9085,N_7343);
nor U10173 (N_10173,N_6884,N_7456);
and U10174 (N_10174,N_7632,N_6848);
nand U10175 (N_10175,N_7221,N_7646);
or U10176 (N_10176,N_9646,N_7993);
or U10177 (N_10177,N_5972,N_6101);
and U10178 (N_10178,N_9280,N_5261);
and U10179 (N_10179,N_8073,N_5052);
nor U10180 (N_10180,N_6339,N_9073);
or U10181 (N_10181,N_9544,N_5555);
or U10182 (N_10182,N_8380,N_6785);
nor U10183 (N_10183,N_8210,N_5930);
or U10184 (N_10184,N_5380,N_8991);
or U10185 (N_10185,N_6649,N_5057);
nor U10186 (N_10186,N_8241,N_7350);
nand U10187 (N_10187,N_9843,N_7133);
nand U10188 (N_10188,N_8349,N_5111);
or U10189 (N_10189,N_6562,N_9833);
or U10190 (N_10190,N_9172,N_6322);
or U10191 (N_10191,N_9768,N_6606);
or U10192 (N_10192,N_8949,N_6896);
and U10193 (N_10193,N_8896,N_8536);
and U10194 (N_10194,N_5887,N_6737);
and U10195 (N_10195,N_5460,N_9334);
and U10196 (N_10196,N_8864,N_6120);
nor U10197 (N_10197,N_7356,N_7935);
and U10198 (N_10198,N_6902,N_6775);
and U10199 (N_10199,N_8507,N_8606);
and U10200 (N_10200,N_5371,N_8622);
or U10201 (N_10201,N_8496,N_9872);
and U10202 (N_10202,N_8942,N_5248);
nand U10203 (N_10203,N_5903,N_5005);
nand U10204 (N_10204,N_5590,N_5419);
nand U10205 (N_10205,N_9912,N_7716);
or U10206 (N_10206,N_9373,N_5399);
or U10207 (N_10207,N_5801,N_8082);
nor U10208 (N_10208,N_9273,N_8406);
nor U10209 (N_10209,N_5638,N_5621);
or U10210 (N_10210,N_7576,N_9947);
nand U10211 (N_10211,N_9291,N_9678);
nor U10212 (N_10212,N_6047,N_7213);
and U10213 (N_10213,N_7616,N_9032);
nor U10214 (N_10214,N_6153,N_7748);
nor U10215 (N_10215,N_8363,N_9673);
or U10216 (N_10216,N_7344,N_5266);
and U10217 (N_10217,N_9029,N_8673);
and U10218 (N_10218,N_9910,N_8935);
nand U10219 (N_10219,N_9744,N_5503);
and U10220 (N_10220,N_8039,N_6484);
nor U10221 (N_10221,N_9363,N_7679);
or U10222 (N_10222,N_7838,N_6051);
or U10223 (N_10223,N_8425,N_5583);
and U10224 (N_10224,N_7484,N_5523);
or U10225 (N_10225,N_6108,N_5580);
or U10226 (N_10226,N_5635,N_5471);
and U10227 (N_10227,N_6676,N_9902);
and U10228 (N_10228,N_8508,N_9059);
and U10229 (N_10229,N_7037,N_7077);
and U10230 (N_10230,N_5290,N_8628);
nor U10231 (N_10231,N_8365,N_5884);
and U10232 (N_10232,N_8584,N_7799);
nor U10233 (N_10233,N_7677,N_5436);
and U10234 (N_10234,N_8623,N_6334);
or U10235 (N_10235,N_9279,N_6854);
nand U10236 (N_10236,N_7043,N_6214);
and U10237 (N_10237,N_9518,N_5494);
or U10238 (N_10238,N_7091,N_7408);
nor U10239 (N_10239,N_6639,N_6019);
and U10240 (N_10240,N_5970,N_9747);
nand U10241 (N_10241,N_9127,N_8011);
nand U10242 (N_10242,N_9026,N_6275);
or U10243 (N_10243,N_8838,N_5385);
nand U10244 (N_10244,N_8835,N_8326);
nand U10245 (N_10245,N_6603,N_5403);
nor U10246 (N_10246,N_6539,N_7401);
nor U10247 (N_10247,N_9359,N_9226);
nor U10248 (N_10248,N_8319,N_7845);
or U10249 (N_10249,N_7958,N_7186);
and U10250 (N_10250,N_6583,N_5780);
or U10251 (N_10251,N_6638,N_6501);
or U10252 (N_10252,N_8401,N_5958);
and U10253 (N_10253,N_6779,N_9315);
nor U10254 (N_10254,N_9429,N_6524);
or U10255 (N_10255,N_9227,N_8184);
xnor U10256 (N_10256,N_5739,N_7121);
and U10257 (N_10257,N_9987,N_5786);
nor U10258 (N_10258,N_8752,N_9103);
nand U10259 (N_10259,N_7795,N_6947);
nand U10260 (N_10260,N_8359,N_8770);
nand U10261 (N_10261,N_8028,N_9959);
nand U10262 (N_10262,N_7082,N_8548);
nor U10263 (N_10263,N_8844,N_8046);
nor U10264 (N_10264,N_9350,N_9955);
and U10265 (N_10265,N_7159,N_7438);
nand U10266 (N_10266,N_7125,N_9958);
nand U10267 (N_10267,N_5587,N_5770);
nor U10268 (N_10268,N_5878,N_7021);
and U10269 (N_10269,N_5582,N_7122);
nor U10270 (N_10270,N_5431,N_9433);
and U10271 (N_10271,N_6771,N_5184);
nand U10272 (N_10272,N_7914,N_9344);
and U10273 (N_10273,N_9072,N_9203);
or U10274 (N_10274,N_5917,N_9878);
nand U10275 (N_10275,N_8175,N_6011);
or U10276 (N_10276,N_9758,N_6099);
and U10277 (N_10277,N_8528,N_6278);
and U10278 (N_10278,N_5936,N_8601);
nand U10279 (N_10279,N_9772,N_7172);
or U10280 (N_10280,N_9278,N_9122);
nor U10281 (N_10281,N_6997,N_8968);
or U10282 (N_10282,N_5505,N_7135);
nand U10283 (N_10283,N_7639,N_8735);
nand U10284 (N_10284,N_7319,N_5048);
nand U10285 (N_10285,N_8264,N_9940);
nand U10286 (N_10286,N_6333,N_6274);
or U10287 (N_10287,N_9917,N_9276);
nand U10288 (N_10288,N_7529,N_6103);
or U10289 (N_10289,N_7420,N_5519);
nand U10290 (N_10290,N_6687,N_5714);
nor U10291 (N_10291,N_7146,N_9581);
and U10292 (N_10292,N_8676,N_6037);
nor U10293 (N_10293,N_5716,N_9930);
and U10294 (N_10294,N_6976,N_9977);
nor U10295 (N_10295,N_5026,N_7851);
nand U10296 (N_10296,N_5516,N_7847);
nand U10297 (N_10297,N_8108,N_8408);
or U10298 (N_10298,N_8267,N_6261);
or U10299 (N_10299,N_6913,N_7558);
nand U10300 (N_10300,N_7171,N_7071);
or U10301 (N_10301,N_6001,N_5703);
nand U10302 (N_10302,N_8288,N_5096);
nand U10303 (N_10303,N_6967,N_8213);
nand U10304 (N_10304,N_6960,N_8181);
and U10305 (N_10305,N_7020,N_8724);
and U10306 (N_10306,N_5181,N_8851);
nor U10307 (N_10307,N_8703,N_7480);
or U10308 (N_10308,N_5808,N_7524);
and U10309 (N_10309,N_7923,N_6203);
or U10310 (N_10310,N_8986,N_5230);
and U10311 (N_10311,N_8328,N_7113);
and U10312 (N_10312,N_5546,N_6480);
nor U10313 (N_10313,N_9752,N_5033);
or U10314 (N_10314,N_8809,N_9981);
or U10315 (N_10315,N_8597,N_8122);
nand U10316 (N_10316,N_8570,N_9312);
nand U10317 (N_10317,N_7666,N_6290);
or U10318 (N_10318,N_7013,N_8447);
and U10319 (N_10319,N_7076,N_6474);
and U10320 (N_10320,N_7200,N_9476);
and U10321 (N_10321,N_5612,N_6095);
nor U10322 (N_10322,N_7270,N_7101);
nor U10323 (N_10323,N_7663,N_6061);
and U10324 (N_10324,N_8647,N_9181);
nor U10325 (N_10325,N_5074,N_6735);
and U10326 (N_10326,N_6588,N_6520);
nor U10327 (N_10327,N_6444,N_9503);
and U10328 (N_10328,N_6002,N_9997);
nand U10329 (N_10329,N_8463,N_9040);
nand U10330 (N_10330,N_7505,N_8876);
nand U10331 (N_10331,N_8792,N_7412);
nand U10332 (N_10332,N_5456,N_7279);
nor U10333 (N_10333,N_8712,N_9873);
nor U10334 (N_10334,N_7798,N_8976);
nor U10335 (N_10335,N_5880,N_8097);
nand U10336 (N_10336,N_5791,N_8091);
nand U10337 (N_10337,N_8559,N_7451);
or U10338 (N_10338,N_8860,N_5683);
nand U10339 (N_10339,N_6951,N_8541);
or U10340 (N_10340,N_7587,N_9763);
nor U10341 (N_10341,N_7892,N_7474);
or U10342 (N_10342,N_5561,N_6607);
nand U10343 (N_10343,N_7908,N_9223);
and U10344 (N_10344,N_5156,N_9824);
nor U10345 (N_10345,N_6498,N_5032);
nor U10346 (N_10346,N_8211,N_6795);
and U10347 (N_10347,N_8455,N_6301);
nor U10348 (N_10348,N_7426,N_9598);
and U10349 (N_10349,N_9674,N_6197);
or U10350 (N_10350,N_6516,N_8538);
or U10351 (N_10351,N_9756,N_9641);
and U10352 (N_10352,N_7683,N_9247);
or U10353 (N_10353,N_8793,N_9428);
nor U10354 (N_10354,N_7266,N_8745);
nand U10355 (N_10355,N_8845,N_9662);
nand U10356 (N_10356,N_7046,N_9348);
and U10357 (N_10357,N_5921,N_9450);
nand U10358 (N_10358,N_9663,N_6220);
nor U10359 (N_10359,N_5015,N_8514);
or U10360 (N_10360,N_7345,N_9876);
nand U10361 (N_10361,N_7889,N_5221);
and U10362 (N_10362,N_5821,N_9998);
or U10363 (N_10363,N_9299,N_6821);
and U10364 (N_10364,N_6566,N_5852);
xnor U10365 (N_10365,N_8848,N_9905);
nand U10366 (N_10366,N_7399,N_8512);
and U10367 (N_10367,N_7952,N_7015);
nand U10368 (N_10368,N_6335,N_8988);
nor U10369 (N_10369,N_6849,N_8383);
xor U10370 (N_10370,N_8615,N_8146);
or U10371 (N_10371,N_5106,N_7884);
and U10372 (N_10372,N_9407,N_5065);
nand U10373 (N_10373,N_5215,N_7081);
nand U10374 (N_10374,N_6653,N_6432);
nand U10375 (N_10375,N_6114,N_9743);
and U10376 (N_10376,N_8767,N_8800);
nor U10377 (N_10377,N_6388,N_8978);
and U10378 (N_10378,N_6204,N_6236);
nor U10379 (N_10379,N_6209,N_9018);
and U10380 (N_10380,N_7522,N_5336);
and U10381 (N_10381,N_6704,N_5870);
and U10382 (N_10382,N_6772,N_8144);
nand U10383 (N_10383,N_5263,N_9943);
and U10384 (N_10384,N_7770,N_8639);
nand U10385 (N_10385,N_7987,N_5259);
nor U10386 (N_10386,N_9729,N_8713);
and U10387 (N_10387,N_5204,N_9041);
nor U10388 (N_10388,N_9994,N_6742);
nor U10389 (N_10389,N_9513,N_6843);
and U10390 (N_10390,N_6296,N_9061);
or U10391 (N_10391,N_6752,N_8219);
nand U10392 (N_10392,N_5345,N_9801);
and U10393 (N_10393,N_9534,N_8836);
nand U10394 (N_10394,N_6926,N_8228);
nor U10395 (N_10395,N_9804,N_8556);
nand U10396 (N_10396,N_8907,N_7996);
and U10397 (N_10397,N_7688,N_9252);
or U10398 (N_10398,N_8155,N_5805);
nand U10399 (N_10399,N_6999,N_7961);
nor U10400 (N_10400,N_8128,N_5568);
and U10401 (N_10401,N_5067,N_7903);
nand U10402 (N_10402,N_6479,N_8462);
and U10403 (N_10403,N_9357,N_9665);
nor U10404 (N_10404,N_8814,N_6858);
nor U10405 (N_10405,N_5007,N_8590);
nand U10406 (N_10406,N_5164,N_6958);
nand U10407 (N_10407,N_9439,N_7063);
or U10408 (N_10408,N_7583,N_6054);
and U10409 (N_10409,N_5913,N_7794);
or U10410 (N_10410,N_9317,N_6264);
and U10411 (N_10411,N_6981,N_9080);
nor U10412 (N_10412,N_5443,N_5931);
or U10413 (N_10413,N_7305,N_8224);
nand U10414 (N_10414,N_9270,N_7393);
nor U10415 (N_10415,N_7162,N_6887);
nand U10416 (N_10416,N_6243,N_9754);
nand U10417 (N_10417,N_9733,N_9391);
and U10418 (N_10418,N_8591,N_5611);
nor U10419 (N_10419,N_7814,N_6782);
nand U10420 (N_10420,N_7118,N_9395);
nor U10421 (N_10421,N_7364,N_5323);
and U10422 (N_10422,N_5900,N_5072);
nor U10423 (N_10423,N_8301,N_8944);
nor U10424 (N_10424,N_9165,N_9811);
nand U10425 (N_10425,N_6337,N_8029);
nand U10426 (N_10426,N_5483,N_6512);
nor U10427 (N_10427,N_5562,N_5600);
nor U10428 (N_10428,N_6435,N_6554);
and U10429 (N_10429,N_6937,N_8022);
and U10430 (N_10430,N_5297,N_6332);
nand U10431 (N_10431,N_6211,N_5250);
nor U10432 (N_10432,N_6465,N_9520);
and U10433 (N_10433,N_9051,N_6957);
nand U10434 (N_10434,N_6182,N_7888);
or U10435 (N_10435,N_5526,N_5688);
and U10436 (N_10436,N_7992,N_9530);
nor U10437 (N_10437,N_7965,N_7145);
nand U10438 (N_10438,N_6438,N_7656);
and U10439 (N_10439,N_9779,N_6678);
and U10440 (N_10440,N_7052,N_8295);
and U10441 (N_10441,N_8499,N_8140);
nand U10442 (N_10442,N_5748,N_5848);
and U10443 (N_10443,N_7072,N_6135);
and U10444 (N_10444,N_5724,N_7497);
or U10445 (N_10445,N_6320,N_6411);
nand U10446 (N_10446,N_9832,N_5132);
or U10447 (N_10447,N_8687,N_6269);
nor U10448 (N_10448,N_8856,N_5016);
nor U10449 (N_10449,N_8882,N_9687);
or U10450 (N_10450,N_6744,N_5077);
and U10451 (N_10451,N_8992,N_7453);
and U10452 (N_10452,N_6507,N_8348);
and U10453 (N_10453,N_7202,N_7065);
and U10454 (N_10454,N_8185,N_8188);
or U10455 (N_10455,N_6068,N_6698);
nand U10456 (N_10456,N_8588,N_6126);
and U10457 (N_10457,N_7129,N_5733);
nor U10458 (N_10458,N_5083,N_6075);
nand U10459 (N_10459,N_8327,N_5409);
nor U10460 (N_10460,N_5863,N_9769);
xor U10461 (N_10461,N_9988,N_9720);
or U10462 (N_10462,N_8427,N_9812);
nor U10463 (N_10463,N_7746,N_7907);
and U10464 (N_10464,N_7230,N_5410);
and U10465 (N_10465,N_9126,N_9472);
nand U10466 (N_10466,N_8409,N_6777);
or U10467 (N_10467,N_6788,N_6194);
or U10468 (N_10468,N_9409,N_8675);
nor U10469 (N_10469,N_8441,N_9871);
and U10470 (N_10470,N_8202,N_9979);
and U10471 (N_10471,N_5734,N_7785);
and U10472 (N_10472,N_8034,N_7715);
nand U10473 (N_10473,N_9820,N_8043);
nand U10474 (N_10474,N_6087,N_5087);
nand U10475 (N_10475,N_9538,N_9457);
nor U10476 (N_10476,N_8439,N_8100);
nor U10477 (N_10477,N_6116,N_5743);
and U10478 (N_10478,N_5898,N_6934);
nor U10479 (N_10479,N_5840,N_8503);
and U10480 (N_10480,N_6491,N_8346);
nand U10481 (N_10481,N_6398,N_8481);
nand U10482 (N_10482,N_8892,N_7066);
and U10483 (N_10483,N_5396,N_8467);
nor U10484 (N_10484,N_9494,N_5186);
nor U10485 (N_10485,N_7001,N_8279);
and U10486 (N_10486,N_6144,N_8697);
or U10487 (N_10487,N_8960,N_8054);
or U10488 (N_10488,N_9934,N_9895);
or U10489 (N_10489,N_9656,N_5697);
or U10490 (N_10490,N_8037,N_8718);
nor U10491 (N_10491,N_5301,N_7875);
nand U10492 (N_10492,N_5303,N_8790);
nand U10493 (N_10493,N_6273,N_5937);
and U10494 (N_10494,N_8917,N_6710);
or U10495 (N_10495,N_7944,N_8709);
or U10496 (N_10496,N_5171,N_7957);
and U10497 (N_10497,N_5205,N_8775);
nand U10498 (N_10498,N_5795,N_8200);
and U10499 (N_10499,N_7955,N_5883);
and U10500 (N_10500,N_9264,N_5889);
nand U10501 (N_10501,N_6810,N_9045);
or U10502 (N_10502,N_9693,N_8902);
nand U10503 (N_10503,N_7087,N_8573);
nor U10504 (N_10504,N_9686,N_8260);
nor U10505 (N_10505,N_9739,N_8149);
xor U10506 (N_10506,N_7727,N_9042);
or U10507 (N_10507,N_7501,N_5952);
or U10508 (N_10508,N_8936,N_7029);
nand U10509 (N_10509,N_5271,N_7823);
nand U10510 (N_10510,N_7234,N_8686);
nand U10511 (N_10511,N_8899,N_6036);
or U10512 (N_10512,N_7295,N_7619);
nand U10513 (N_10513,N_9957,N_7132);
nand U10514 (N_10514,N_8643,N_5662);
or U10515 (N_10515,N_7381,N_5322);
nor U10516 (N_10516,N_7500,N_9892);
xor U10517 (N_10517,N_7417,N_9784);
nand U10518 (N_10518,N_5877,N_7890);
nor U10519 (N_10519,N_9189,N_5920);
nand U10520 (N_10520,N_5377,N_5071);
or U10521 (N_10521,N_9420,N_5803);
nand U10522 (N_10522,N_9033,N_5010);
or U10523 (N_10523,N_9177,N_8863);
or U10524 (N_10524,N_8131,N_9322);
or U10525 (N_10525,N_5457,N_5979);
and U10526 (N_10526,N_9109,N_7627);
nand U10527 (N_10527,N_9405,N_5666);
or U10528 (N_10528,N_7602,N_9019);
or U10529 (N_10529,N_9284,N_8915);
or U10530 (N_10530,N_9398,N_8934);
or U10531 (N_10531,N_5778,N_5985);
nor U10532 (N_10532,N_5713,N_9740);
or U10533 (N_10533,N_7913,N_8135);
nand U10534 (N_10534,N_8906,N_8196);
nor U10535 (N_10535,N_5343,N_7492);
or U10536 (N_10536,N_8952,N_9077);
or U10537 (N_10537,N_8257,N_8698);
nor U10538 (N_10538,N_9438,N_5809);
or U10539 (N_10539,N_9113,N_5897);
nor U10540 (N_10540,N_9642,N_5995);
or U10541 (N_10541,N_7946,N_8394);
and U10542 (N_10542,N_8807,N_5375);
nor U10543 (N_10543,N_5275,N_5550);
or U10544 (N_10544,N_9365,N_6375);
and U10545 (N_10545,N_8353,N_6284);
and U10546 (N_10546,N_7288,N_8903);
or U10547 (N_10547,N_5687,N_6007);
nor U10548 (N_10548,N_6894,N_6972);
or U10549 (N_10549,N_7661,N_8087);
nor U10550 (N_10550,N_8449,N_5765);
or U10551 (N_10551,N_7568,N_5790);
nor U10552 (N_10552,N_5826,N_8744);
and U10553 (N_10553,N_9430,N_7207);
nand U10554 (N_10554,N_9465,N_5200);
nor U10555 (N_10555,N_8252,N_9715);
nor U10556 (N_10556,N_6006,N_5045);
and U10557 (N_10557,N_7694,N_8723);
nor U10558 (N_10558,N_6307,N_5839);
nand U10559 (N_10559,N_9787,N_9448);
nand U10560 (N_10560,N_5185,N_8208);
nand U10561 (N_10561,N_8466,N_5459);
and U10562 (N_10562,N_9790,N_7433);
or U10563 (N_10563,N_5745,N_9487);
nand U10564 (N_10564,N_6770,N_9914);
nand U10565 (N_10565,N_7722,N_5213);
or U10566 (N_10566,N_9228,N_7117);
nand U10567 (N_10567,N_9903,N_8024);
nand U10568 (N_10568,N_9942,N_8511);
xor U10569 (N_10569,N_8280,N_7097);
nand U10570 (N_10570,N_9764,N_7355);
nor U10571 (N_10571,N_7904,N_5807);
nand U10572 (N_10572,N_6881,N_7424);
nor U10573 (N_10573,N_7329,N_5685);
and U10574 (N_10574,N_9770,N_5382);
or U10575 (N_10575,N_7411,N_6811);
nand U10576 (N_10576,N_9755,N_9364);
nor U10577 (N_10577,N_5167,N_9788);
nor U10578 (N_10578,N_9417,N_5435);
and U10579 (N_10579,N_9475,N_8052);
and U10580 (N_10580,N_8016,N_8049);
nor U10581 (N_10581,N_8958,N_9574);
nand U10582 (N_10582,N_8811,N_5944);
or U10583 (N_10583,N_5579,N_9010);
and U10584 (N_10584,N_5426,N_9635);
or U10585 (N_10585,N_5835,N_8141);
and U10586 (N_10586,N_9415,N_9064);
or U10587 (N_10587,N_8255,N_6535);
or U10588 (N_10588,N_6840,N_9183);
or U10589 (N_10589,N_8875,N_6385);
and U10590 (N_10590,N_5761,N_9105);
nor U10591 (N_10591,N_5330,N_5669);
and U10592 (N_10592,N_6212,N_7388);
nand U10593 (N_10593,N_5084,N_7014);
nor U10594 (N_10594,N_6029,N_8117);
and U10595 (N_10595,N_8068,N_6798);
and U10596 (N_10596,N_7930,N_6409);
and U10597 (N_10597,N_5493,N_7116);
nand U10598 (N_10598,N_7766,N_7294);
nand U10599 (N_10599,N_6492,N_6244);
nor U10600 (N_10600,N_9753,N_5659);
and U10601 (N_10601,N_6442,N_7927);
nand U10602 (N_10602,N_6419,N_6974);
nor U10603 (N_10603,N_7419,N_8357);
or U10604 (N_10604,N_7614,N_7297);
nand U10605 (N_10605,N_8084,N_6711);
and U10606 (N_10606,N_9995,N_7797);
and U10607 (N_10607,N_6280,N_7155);
and U10608 (N_10608,N_6138,N_8918);
nor U10609 (N_10609,N_6998,N_8857);
nand U10610 (N_10610,N_5317,N_5971);
nand U10611 (N_10611,N_7733,N_7308);
nand U10612 (N_10612,N_5150,N_8003);
or U10613 (N_10613,N_5654,N_8475);
nand U10614 (N_10614,N_7941,N_9501);
and U10615 (N_10615,N_7857,N_7256);
nand U10616 (N_10616,N_9624,N_8370);
or U10617 (N_10617,N_6441,N_5969);
nor U10618 (N_10618,N_7060,N_9379);
and U10619 (N_10619,N_8214,N_8421);
nand U10620 (N_10620,N_5357,N_6000);
xor U10621 (N_10621,N_8956,N_8871);
nand U10622 (N_10622,N_8710,N_6453);
or U10623 (N_10623,N_6648,N_7507);
nand U10624 (N_10624,N_9265,N_6596);
or U10625 (N_10625,N_8079,N_6573);
and U10626 (N_10626,N_7352,N_9837);
nor U10627 (N_10627,N_8000,N_5499);
or U10628 (N_10628,N_5822,N_5412);
nor U10629 (N_10629,N_9071,N_5139);
and U10630 (N_10630,N_8515,N_5667);
or U10631 (N_10631,N_7304,N_5594);
nor U10632 (N_10632,N_6208,N_8030);
xor U10633 (N_10633,N_5030,N_9568);
and U10634 (N_10634,N_7689,N_7301);
nand U10635 (N_10635,N_5831,N_8910);
and U10636 (N_10636,N_7723,N_6199);
and U10637 (N_10637,N_8250,N_7496);
nor U10638 (N_10638,N_9408,N_6620);
nand U10639 (N_10639,N_8336,N_8784);
or U10640 (N_10640,N_9850,N_8768);
nand U10641 (N_10641,N_5581,N_7809);
or U10642 (N_10642,N_5578,N_7246);
nand U10643 (N_10643,N_6133,N_5647);
nor U10644 (N_10644,N_6169,N_9576);
or U10645 (N_10645,N_9342,N_7771);
and U10646 (N_10646,N_7626,N_9838);
and U10647 (N_10647,N_9340,N_8159);
or U10648 (N_10648,N_9968,N_8426);
nor U10649 (N_10649,N_9580,N_6429);
nor U10650 (N_10650,N_6178,N_6556);
and U10651 (N_10651,N_7338,N_9388);
nor U10652 (N_10652,N_7860,N_9147);
nor U10653 (N_10653,N_6495,N_6170);
nor U10654 (N_10654,N_7502,N_6134);
or U10655 (N_10655,N_9561,N_7921);
or U10656 (N_10656,N_7869,N_5773);
nor U10657 (N_10657,N_7739,N_8167);
and U10658 (N_10658,N_8677,N_5557);
and U10659 (N_10659,N_7846,N_5202);
nand U10660 (N_10660,N_6229,N_7669);
nand U10661 (N_10661,N_9206,N_5836);
nor U10662 (N_10662,N_8333,N_9295);
nand U10663 (N_10663,N_5168,N_8435);
nor U10664 (N_10664,N_7849,N_7591);
nor U10665 (N_10665,N_9675,N_9125);
or U10666 (N_10666,N_9009,N_8659);
or U10667 (N_10667,N_7425,N_5094);
nand U10668 (N_10668,N_6893,N_6860);
or U10669 (N_10669,N_9499,N_8021);
or U10670 (N_10670,N_5708,N_7744);
nand U10671 (N_10671,N_9974,N_5360);
and U10672 (N_10672,N_7648,N_9326);
nand U10673 (N_10673,N_8689,N_5434);
or U10674 (N_10674,N_7183,N_5454);
nor U10675 (N_10675,N_8794,N_8932);
or U10676 (N_10676,N_9374,N_9309);
or U10677 (N_10677,N_7585,N_7471);
nand U10678 (N_10678,N_9347,N_5353);
and U10679 (N_10679,N_8656,N_5576);
or U10680 (N_10680,N_5682,N_9700);
nor U10681 (N_10681,N_7111,N_6496);
nand U10682 (N_10682,N_8884,N_8373);
nand U10683 (N_10683,N_9050,N_5486);
and U10684 (N_10684,N_6865,N_8137);
xnor U10685 (N_10685,N_8696,N_6403);
or U10686 (N_10686,N_6372,N_5020);
and U10687 (N_10687,N_8055,N_5368);
nor U10688 (N_10688,N_7969,N_9324);
nor U10689 (N_10689,N_7149,N_5305);
nor U10690 (N_10690,N_8592,N_5141);
or U10691 (N_10691,N_9425,N_5155);
nand U10692 (N_10692,N_6586,N_6629);
and U10693 (N_10693,N_6985,N_8771);
nand U10694 (N_10694,N_9377,N_5130);
nand U10695 (N_10695,N_5929,N_8139);
nand U10696 (N_10696,N_7574,N_5624);
or U10697 (N_10697,N_9798,N_6437);
nand U10698 (N_10698,N_8828,N_9011);
nor U10699 (N_10699,N_9816,N_5287);
or U10700 (N_10700,N_8660,N_8683);
nand U10701 (N_10701,N_6841,N_7829);
and U10702 (N_10702,N_7265,N_5643);
or U10703 (N_10703,N_9375,N_7184);
or U10704 (N_10704,N_8152,N_8605);
or U10705 (N_10705,N_9412,N_6808);
and U10706 (N_10706,N_7670,N_6489);
or U10707 (N_10707,N_6823,N_7105);
or U10708 (N_10708,N_8436,N_5449);
nand U10709 (N_10709,N_8314,N_6056);
or U10710 (N_10710,N_7617,N_5511);
or U10711 (N_10711,N_7989,N_5291);
nand U10712 (N_10712,N_6405,N_5108);
and U10713 (N_10713,N_6309,N_7620);
nor U10714 (N_10714,N_7318,N_6412);
nor U10715 (N_10715,N_8058,N_5529);
nor U10716 (N_10716,N_6633,N_9511);
nor U10717 (N_10717,N_9088,N_5575);
nand U10718 (N_10718,N_6304,N_6106);
and U10719 (N_10719,N_5534,N_8533);
or U10720 (N_10720,N_5195,N_6215);
or U10721 (N_10721,N_7250,N_5107);
nor U10722 (N_10722,N_7441,N_6792);
or U10723 (N_10723,N_8671,N_5061);
and U10724 (N_10724,N_7057,N_7216);
and U10725 (N_10725,N_6221,N_9922);
or U10726 (N_10726,N_9155,N_9240);
nand U10727 (N_10727,N_9777,N_5114);
nand U10728 (N_10728,N_8316,N_7867);
nand U10729 (N_10729,N_8306,N_5109);
and U10730 (N_10730,N_6528,N_8269);
or U10731 (N_10731,N_6448,N_7850);
or U10732 (N_10732,N_5642,N_7662);
nor U10733 (N_10733,N_8599,N_9215);
nor U10734 (N_10734,N_5335,N_9160);
and U10735 (N_10735,N_9158,N_9901);
and U10736 (N_10736,N_7361,N_6689);
nand U10737 (N_10737,N_6063,N_5698);
and U10738 (N_10738,N_9323,N_8389);
nor U10739 (N_10739,N_9650,N_5628);
nor U10740 (N_10740,N_5055,N_5749);
nor U10741 (N_10741,N_9952,N_6045);
and U10742 (N_10742,N_9110,N_5812);
or U10743 (N_10743,N_8018,N_8553);
or U10744 (N_10744,N_5719,N_7239);
and U10745 (N_10745,N_6942,N_5199);
and U10746 (N_10746,N_8132,N_5076);
and U10747 (N_10747,N_8700,N_6459);
or U10748 (N_10748,N_5656,N_6617);
or U10749 (N_10749,N_6783,N_7668);
or U10750 (N_10750,N_6637,N_8411);
and U10751 (N_10751,N_5539,N_7804);
nor U10752 (N_10752,N_5554,N_5214);
or U10753 (N_10753,N_5439,N_5515);
or U10754 (N_10754,N_7640,N_6931);
or U10755 (N_10755,N_6622,N_7684);
nand U10756 (N_10756,N_9668,N_6549);
or U10757 (N_10757,N_9868,N_7485);
nand U10758 (N_10758,N_7830,N_8232);
nand U10759 (N_10759,N_5570,N_9067);
or U10760 (N_10760,N_9969,N_8243);
nand U10761 (N_10761,N_5339,N_8238);
and U10762 (N_10762,N_8604,N_9670);
nor U10763 (N_10763,N_8235,N_6387);
xnor U10764 (N_10764,N_9292,N_8032);
and U10765 (N_10765,N_7915,N_9152);
nor U10766 (N_10766,N_7945,N_5894);
nand U10767 (N_10767,N_7040,N_8897);
nand U10768 (N_10768,N_6109,N_9097);
or U10769 (N_10769,N_9188,N_7826);
nor U10770 (N_10770,N_9826,N_7506);
nor U10771 (N_10771,N_8179,N_7822);
and U10772 (N_10772,N_8147,N_8558);
nor U10773 (N_10773,N_9086,N_5437);
or U10774 (N_10774,N_8594,N_7843);
nor U10775 (N_10775,N_6173,N_7589);
nor U10776 (N_10776,N_6866,N_7686);
nor U10777 (N_10777,N_5802,N_9973);
nand U10778 (N_10778,N_5068,N_6155);
nand U10779 (N_10779,N_9178,N_7321);
and U10780 (N_10780,N_8861,N_8796);
or U10781 (N_10781,N_7581,N_6034);
nor U10782 (N_10782,N_9013,N_7157);
or U10783 (N_10783,N_6314,N_9092);
nor U10784 (N_10784,N_8626,N_6324);
nor U10785 (N_10785,N_9640,N_8027);
and U10786 (N_10786,N_9094,N_6921);
nor U10787 (N_10787,N_6876,N_5498);
nor U10788 (N_10788,N_5677,N_5166);
and U10789 (N_10789,N_5982,N_7518);
nand U10790 (N_10790,N_6167,N_8706);
nand U10791 (N_10791,N_5406,N_5596);
nand U10792 (N_10792,N_6610,N_9757);
nand U10793 (N_10793,N_8278,N_5567);
nor U10794 (N_10794,N_5123,N_7878);
or U10795 (N_10795,N_9851,N_9796);
nor U10796 (N_10796,N_5947,N_8102);
nor U10797 (N_10797,N_7566,N_9716);
nor U10798 (N_10798,N_7738,N_6941);
or U10799 (N_10799,N_7647,N_8815);
nand U10800 (N_10800,N_8981,N_8702);
nand U10801 (N_10801,N_5281,N_7335);
and U10802 (N_10802,N_6701,N_9980);
or U10803 (N_10803,N_9597,N_8287);
nand U10804 (N_10804,N_7730,N_8395);
and U10805 (N_10805,N_9637,N_7462);
nand U10806 (N_10806,N_8420,N_5627);
nand U10807 (N_10807,N_6665,N_7665);
nand U10808 (N_10808,N_9599,N_9054);
nand U10809 (N_10809,N_9002,N_6300);
or U10810 (N_10810,N_9030,N_9044);
or U10811 (N_10811,N_9090,N_8364);
nor U10812 (N_10812,N_6975,N_6265);
or U10813 (N_10813,N_5178,N_6234);
nor U10814 (N_10814,N_9765,N_8820);
and U10815 (N_10815,N_6504,N_6062);
or U10816 (N_10816,N_8312,N_8222);
and U10817 (N_10817,N_7366,N_7693);
nor U10818 (N_10818,N_9908,N_7310);
nand U10819 (N_10819,N_6943,N_8044);
or U10820 (N_10820,N_7977,N_5613);
nand U10821 (N_10821,N_5962,N_7397);
nand U10822 (N_10822,N_6953,N_8841);
and U10823 (N_10823,N_6350,N_9840);
nand U10824 (N_10824,N_7702,N_6238);
nand U10825 (N_10825,N_5424,N_5133);
and U10826 (N_10826,N_9150,N_5000);
nor U10827 (N_10827,N_7026,N_8168);
or U10828 (N_10828,N_7340,N_8575);
nand U10829 (N_10829,N_7225,N_9836);
nor U10830 (N_10830,N_9368,N_8542);
or U10831 (N_10831,N_5747,N_7549);
or U10832 (N_10832,N_9808,N_8859);
nor U10833 (N_10833,N_6724,N_5354);
nor U10834 (N_10834,N_8299,N_8862);
and U10835 (N_10835,N_8035,N_5632);
nand U10836 (N_10836,N_6044,N_8611);
nor U10837 (N_10837,N_8247,N_6348);
nor U10838 (N_10838,N_9672,N_8746);
and U10839 (N_10839,N_9209,N_5922);
nand U10840 (N_10840,N_7995,N_6386);
nand U10841 (N_10841,N_8468,N_9163);
or U10842 (N_10842,N_5119,N_6078);
or U10843 (N_10843,N_6812,N_7384);
nor U10844 (N_10844,N_6856,N_6570);
and U10845 (N_10845,N_9823,N_7880);
or U10846 (N_10846,N_7277,N_6813);
nand U10847 (N_10847,N_8582,N_9718);
nor U10848 (N_10848,N_8494,N_6365);
and U10849 (N_10849,N_8878,N_5967);
and U10850 (N_10850,N_7300,N_5325);
nand U10851 (N_10851,N_7303,N_9197);
or U10852 (N_10852,N_9654,N_5081);
and U10853 (N_10853,N_6679,N_8456);
and U10854 (N_10854,N_5265,N_6154);
and U10855 (N_10855,N_8501,N_7734);
and U10856 (N_10856,N_8376,N_5844);
or U10857 (N_10857,N_7032,N_6241);
and U10858 (N_10858,N_8905,N_8550);
nand U10859 (N_10859,N_9551,N_6111);
or U10860 (N_10860,N_9083,N_8113);
nor U10861 (N_10861,N_9141,N_9231);
nor U10862 (N_10862,N_9589,N_8360);
and U10863 (N_10863,N_6715,N_6500);
and U10864 (N_10864,N_5673,N_9219);
nor U10865 (N_10865,N_7569,N_7573);
or U10866 (N_10866,N_9814,N_5940);
nor U10867 (N_10867,N_8256,N_5994);
nor U10868 (N_10868,N_8321,N_7325);
nor U10869 (N_10869,N_8990,N_7951);
nor U10870 (N_10870,N_8166,N_8387);
and U10871 (N_10871,N_6497,N_7148);
nor U10872 (N_10872,N_6506,N_7410);
nor U10873 (N_10873,N_9353,N_7936);
and U10874 (N_10874,N_6469,N_8663);
and U10875 (N_10875,N_6996,N_6016);
nor U10876 (N_10876,N_5551,N_8602);
and U10877 (N_10877,N_7687,N_9101);
or U10878 (N_10878,N_6161,N_7598);
or U10879 (N_10879,N_8249,N_6825);
nand U10880 (N_10880,N_5695,N_8757);
nand U10881 (N_10881,N_6702,N_6548);
nand U10882 (N_10882,N_5220,N_8641);
or U10883 (N_10883,N_6805,N_8733);
nand U10884 (N_10884,N_5320,N_8866);
nand U10885 (N_10885,N_5868,N_7257);
nor U10886 (N_10886,N_7701,N_8540);
nand U10887 (N_10887,N_7203,N_9548);
and U10888 (N_10888,N_9311,N_7240);
or U10889 (N_10889,N_9949,N_9006);
nor U10890 (N_10890,N_5853,N_7634);
nand U10891 (N_10891,N_9133,N_7137);
nor U10892 (N_10892,N_8493,N_9176);
and U10893 (N_10893,N_6609,N_6875);
and U10894 (N_10894,N_8810,N_6517);
and U10895 (N_10895,N_8769,N_8025);
and U10896 (N_10896,N_5528,N_8766);
and U10897 (N_10897,N_6833,N_9992);
nor U10898 (N_10898,N_6176,N_7177);
nand U10899 (N_10899,N_8041,N_9869);
or U10900 (N_10900,N_8063,N_6734);
nand U10901 (N_10901,N_9831,N_6017);
nor U10902 (N_10902,N_8400,N_8484);
or U10903 (N_10903,N_7752,N_6505);
or U10904 (N_10904,N_8050,N_8961);
nand U10905 (N_10905,N_7333,N_5644);
nor U10906 (N_10906,N_5902,N_6961);
or U10907 (N_10907,N_6992,N_6804);
nand U10908 (N_10908,N_7590,N_7788);
nand U10909 (N_10909,N_8785,N_5249);
nor U10910 (N_10910,N_9681,N_8633);
or U10911 (N_10911,N_9507,N_8385);
and U10912 (N_10912,N_7331,N_8358);
nand U10913 (N_10913,N_6367,N_7762);
or U10914 (N_10914,N_7482,N_6421);
and U10915 (N_10915,N_9933,N_9469);
and U10916 (N_10916,N_5652,N_6584);
or U10917 (N_10917,N_7898,N_9809);
or U10918 (N_10918,N_6933,N_9562);
nor U10919 (N_10919,N_9380,N_6697);
nand U10920 (N_10920,N_5650,N_6647);
xor U10921 (N_10921,N_9144,N_9136);
or U10922 (N_10922,N_9166,N_9699);
or U10923 (N_10923,N_6611,N_6717);
nor U10924 (N_10924,N_9497,N_8957);
or U10925 (N_10925,N_6289,N_9017);
or U10926 (N_10926,N_8927,N_9232);
and U10927 (N_10927,N_7487,N_9381);
nand U10928 (N_10928,N_7523,N_5306);
nor U10929 (N_10929,N_6052,N_6684);
or U10930 (N_10930,N_8691,N_7510);
nor U10931 (N_10931,N_7209,N_8843);
and U10932 (N_10932,N_5630,N_7856);
nand U10933 (N_10933,N_9046,N_6245);
nor U10934 (N_10934,N_8382,N_7127);
or U10935 (N_10935,N_7389,N_5827);
and U10936 (N_10936,N_9616,N_6327);
nor U10937 (N_10937,N_6473,N_6147);
or U10938 (N_10938,N_9060,N_6079);
or U10939 (N_10939,N_9256,N_9098);
nor U10940 (N_10940,N_9828,N_5446);
nor U10941 (N_10941,N_9413,N_7882);
or U10942 (N_10942,N_5344,N_9410);
nor U10943 (N_10943,N_9822,N_5351);
nor U10944 (N_10944,N_7165,N_9468);
or U10945 (N_10945,N_9175,N_9817);
and U10946 (N_10946,N_5300,N_6626);
xor U10947 (N_10947,N_6464,N_5895);
or U10948 (N_10948,N_7588,N_9014);
nor U10949 (N_10949,N_8930,N_8827);
and U10950 (N_10950,N_9114,N_5851);
or U10951 (N_10951,N_7110,N_8965);
or U10952 (N_10952,N_6755,N_9491);
nor U10953 (N_10953,N_7198,N_9055);
or U10954 (N_10954,N_5565,N_6557);
nor U10955 (N_10955,N_7242,N_6306);
or U10956 (N_10956,N_8178,N_8681);
or U10957 (N_10957,N_7400,N_5725);
nand U10958 (N_10958,N_5044,N_8664);
and U10959 (N_10959,N_7078,N_6085);
nand U10960 (N_10960,N_8972,N_9195);
nor U10961 (N_10961,N_9623,N_8982);
nand U10962 (N_10962,N_6404,N_6870);
and U10963 (N_10963,N_9888,N_6336);
or U10964 (N_10964,N_9248,N_5759);
nor U10965 (N_10965,N_5775,N_8020);
nor U10966 (N_10966,N_8209,N_6251);
nand U10967 (N_10967,N_5273,N_8750);
or U10968 (N_10968,N_5874,N_5819);
nand U10969 (N_10969,N_5961,N_9860);
and U10970 (N_10970,N_5824,N_8437);
nand U10971 (N_10971,N_6510,N_5764);
and U10972 (N_10972,N_5560,N_8823);
nand U10973 (N_10973,N_9124,N_5722);
nand U10974 (N_10974,N_5717,N_5384);
nand U10975 (N_10975,N_7599,N_8061);
nor U10976 (N_10976,N_9154,N_8658);
nand U10977 (N_10977,N_9773,N_9566);
and U10978 (N_10978,N_7108,N_5906);
and U10979 (N_10979,N_7405,N_8485);
nor U10980 (N_10980,N_7807,N_9960);
or U10981 (N_10981,N_9508,N_5488);
and U10982 (N_10982,N_5907,N_6526);
nor U10983 (N_10983,N_8780,N_7781);
and U10984 (N_10984,N_5140,N_8947);
and U10985 (N_10985,N_5169,N_6248);
or U10986 (N_10986,N_6509,N_5710);
nand U10987 (N_10987,N_9034,N_8565);
or U10988 (N_10988,N_7498,N_8194);
and U10989 (N_10989,N_9505,N_5871);
nand U10990 (N_10990,N_7367,N_8344);
nor U10991 (N_10991,N_8642,N_5376);
and U10992 (N_10992,N_8595,N_6839);
nor U10993 (N_10993,N_5990,N_8251);
and U10994 (N_10994,N_6529,N_6714);
nand U10995 (N_10995,N_5866,N_5520);
or U10996 (N_10996,N_7596,N_7782);
and U10997 (N_10997,N_7801,N_9971);
nor U10998 (N_10998,N_8955,N_5319);
and U10999 (N_10999,N_8433,N_5075);
or U11000 (N_11000,N_8762,N_9427);
nand U11001 (N_11001,N_5608,N_5468);
or U11002 (N_11002,N_8078,N_5280);
nand U11003 (N_11003,N_7540,N_6623);
and U11004 (N_11004,N_9569,N_7450);
or U11005 (N_11005,N_7954,N_7561);
nor U11006 (N_11006,N_8236,N_8505);
nand U11007 (N_11007,N_9471,N_8454);
nor U11008 (N_11008,N_8821,N_7611);
nor U11009 (N_11009,N_5524,N_5198);
nand U11010 (N_11010,N_6950,N_5586);
and U11011 (N_11011,N_7963,N_9089);
and U11012 (N_11012,N_7900,N_7837);
nand U11013 (N_11013,N_8478,N_7786);
nor U11014 (N_11014,N_9198,N_8834);
and U11015 (N_11015,N_6460,N_5549);
or U11016 (N_11016,N_9458,N_5660);
and U11017 (N_11017,N_7509,N_5796);
nor U11018 (N_11018,N_7299,N_6249);
or U11019 (N_11019,N_9898,N_5175);
nor U11020 (N_11020,N_8666,N_8759);
and U11021 (N_11021,N_6356,N_8819);
and U11022 (N_11022,N_7307,N_6148);
nor U11023 (N_11023,N_6447,N_5242);
and U11024 (N_11024,N_7997,N_7775);
nand U11025 (N_11025,N_7377,N_8465);
nor U11026 (N_11026,N_7937,N_5408);
nor U11027 (N_11027,N_5744,N_9821);
or U11028 (N_11028,N_5035,N_9003);
or U11029 (N_11029,N_9161,N_9258);
or U11030 (N_11030,N_9356,N_6131);
nand U11031 (N_11031,N_7473,N_6005);
nor U11032 (N_11032,N_7088,N_6971);
nand U11033 (N_11033,N_7058,N_7477);
or U11034 (N_11034,N_5066,N_8802);
nor U11035 (N_11035,N_8564,N_5986);
nand U11036 (N_11036,N_5566,N_5955);
nor U11037 (N_11037,N_7342,N_7721);
nor U11038 (N_11038,N_8292,N_7873);
and U11039 (N_11039,N_6650,N_9620);
nand U11040 (N_11040,N_6384,N_7252);
nor U11041 (N_11041,N_6310,N_9557);
or U11042 (N_11042,N_7336,N_8596);
or U11043 (N_11043,N_7776,N_9946);
and U11044 (N_11044,N_6105,N_7107);
nand U11045 (N_11045,N_5059,N_5750);
nand U11046 (N_11046,N_7324,N_9382);
nor U11047 (N_11047,N_8338,N_9667);
nor U11048 (N_11048,N_7126,N_9572);
nand U11049 (N_11049,N_6130,N_6534);
nand U11050 (N_11050,N_6067,N_5295);
or U11051 (N_11051,N_8083,N_6318);
nand U11052 (N_11052,N_6817,N_7445);
and U11053 (N_11053,N_5552,N_6727);
and U11054 (N_11054,N_5451,N_9900);
nor U11055 (N_11055,N_7539,N_8717);
and U11056 (N_11056,N_8089,N_8148);
nand U11057 (N_11057,N_6196,N_8938);
or U11058 (N_11058,N_8997,N_8877);
and U11059 (N_11059,N_8998,N_9416);
or U11060 (N_11060,N_6162,N_8614);
or U11061 (N_11061,N_9304,N_9193);
nand U11062 (N_11062,N_5849,N_9352);
and U11063 (N_11063,N_6305,N_5670);
nor U11064 (N_11064,N_9517,N_5721);
nor U11065 (N_11065,N_8670,N_7700);
or U11066 (N_11066,N_8239,N_6750);
or U11067 (N_11067,N_5736,N_6949);
or U11068 (N_11068,N_9657,N_8098);
nor U11069 (N_11069,N_6142,N_8177);
and U11070 (N_11070,N_5056,N_9648);
or U11071 (N_11071,N_9639,N_8648);
or U11072 (N_11072,N_7232,N_8217);
xnor U11073 (N_11073,N_8872,N_8645);
and U11074 (N_11074,N_6431,N_5078);
or U11075 (N_11075,N_7534,N_7208);
nor U11076 (N_11076,N_9490,N_5113);
and U11077 (N_11077,N_6232,N_7314);
nor U11078 (N_11078,N_6475,N_7757);
or U11079 (N_11079,N_6224,N_7152);
nand U11080 (N_11080,N_7517,N_6277);
or U11081 (N_11081,N_8839,N_6347);
nor U11082 (N_11082,N_8983,N_8443);
and U11083 (N_11083,N_7966,N_6097);
nor U11084 (N_11084,N_5489,N_9721);
and U11085 (N_11085,N_9139,N_5120);
and U11086 (N_11086,N_9157,N_9682);
and U11087 (N_11087,N_7174,N_9601);
and U11088 (N_11088,N_9035,N_8734);
and U11089 (N_11089,N_7481,N_6994);
nor U11090 (N_11090,N_6778,N_6390);
nand U11091 (N_11091,N_6673,N_6071);
or U11092 (N_11092,N_6836,N_6223);
nand U11093 (N_11093,N_6262,N_9185);
nand U11094 (N_11094,N_6579,N_5774);
nor U11095 (N_11095,N_7984,N_8009);
nand U11096 (N_11096,N_7245,N_8434);
or U11097 (N_11097,N_5789,N_7841);
nor U11098 (N_11098,N_9253,N_7759);
nand U11099 (N_11099,N_5218,N_7131);
and U11100 (N_11100,N_8324,N_8921);
nand U11101 (N_11101,N_5753,N_5862);
xnor U11102 (N_11102,N_9028,N_6121);
nor U11103 (N_11103,N_9709,N_9233);
or U11104 (N_11104,N_5599,N_9422);
nand U11105 (N_11105,N_6736,N_5128);
or U11106 (N_11106,N_5727,N_5779);
and U11107 (N_11107,N_9730,N_9211);
nand U11108 (N_11108,N_6025,N_7244);
nor U11109 (N_11109,N_5101,N_5788);
nand U11110 (N_11110,N_6180,N_9451);
and U11111 (N_11111,N_5358,N_9762);
and U11112 (N_11112,N_8290,N_5334);
or U11113 (N_11113,N_7705,N_8778);
nand U11114 (N_11114,N_7188,N_9996);
and U11115 (N_11115,N_6102,N_9521);
nor U11116 (N_11116,N_8074,N_8002);
and U11117 (N_11117,N_7416,N_8985);
nor U11118 (N_11118,N_7537,N_8926);
nand U11119 (N_11119,N_8416,N_9694);
and U11120 (N_11120,N_6371,N_6257);
nor U11121 (N_11121,N_7883,N_7376);
nor U11122 (N_11122,N_9515,N_7711);
or U11123 (N_11123,N_5031,N_8699);
and U11124 (N_11124,N_7607,N_9355);
nand U11125 (N_11125,N_5008,N_5327);
or U11126 (N_11126,N_6198,N_6560);
nand U11127 (N_11127,N_6021,N_7917);
and U11128 (N_11128,N_9241,N_9924);
xnor U11129 (N_11129,N_8019,N_8458);
and U11130 (N_11130,N_7238,N_5192);
and U11131 (N_11131,N_7633,N_5705);
nand U11132 (N_11132,N_7204,N_7346);
nor U11133 (N_11133,N_6807,N_8518);
nor U11134 (N_11134,N_7877,N_6728);
and U11135 (N_11135,N_8679,N_7971);
nor U11136 (N_11136,N_6363,N_9036);
or U11137 (N_11137,N_6424,N_5533);
and U11138 (N_11138,N_8913,N_5785);
or U11139 (N_11139,N_6201,N_9845);
or U11140 (N_11140,N_9272,N_9619);
and U11141 (N_11141,N_6657,N_6048);
nand U11142 (N_11142,N_9603,N_7429);
nor U11143 (N_11143,N_6853,N_6857);
and U11144 (N_11144,N_8367,N_9435);
nand U11145 (N_11145,N_7938,N_7187);
or U11146 (N_11146,N_8451,N_9174);
nand U11147 (N_11147,N_9479,N_6656);
nand U11148 (N_11148,N_9839,N_9289);
nor U11149 (N_11149,N_7283,N_5182);
and U11150 (N_11150,N_9608,N_9751);
nand U11151 (N_11151,N_7390,N_7112);
and U11152 (N_11152,N_8795,N_6929);
or U11153 (N_11153,N_9588,N_9473);
nand U11154 (N_11154,N_7932,N_9935);
and U11155 (N_11155,N_7564,N_7816);
and U11156 (N_11156,N_6049,N_6020);
and U11157 (N_11157,N_9630,N_9600);
or U11158 (N_11158,N_7042,N_6392);
or U11159 (N_11159,N_7755,N_5365);
or U11160 (N_11160,N_9558,N_9214);
nand U11161 (N_11161,N_6658,N_9771);
and U11162 (N_11162,N_6991,N_6352);
and U11163 (N_11163,N_6225,N_7978);
or U11164 (N_11164,N_9404,N_7249);
and U11165 (N_11165,N_5206,N_6004);
or U11166 (N_11166,N_7434,N_8693);
nor U11167 (N_11167,N_5784,N_5825);
nand U11168 (N_11168,N_6938,N_8886);
and U11169 (N_11169,N_8086,N_6389);
or U11170 (N_11170,N_6125,N_6686);
and U11171 (N_11171,N_5841,N_5538);
nand U11172 (N_11172,N_8284,N_5912);
nor U11173 (N_11173,N_6171,N_8580);
and U11174 (N_11174,N_7006,N_6295);
nand U11175 (N_11175,N_9301,N_6722);
nand U11176 (N_11176,N_7316,N_6311);
or U11177 (N_11177,N_9286,N_7353);
nor U11178 (N_11178,N_9883,N_7176);
or U11179 (N_11179,N_5142,N_9991);
or U11180 (N_11180,N_7472,N_8234);
xor U11181 (N_11181,N_6370,N_6601);
and U11182 (N_11182,N_5476,N_5525);
nor U11183 (N_11183,N_6537,N_6104);
and U11184 (N_11184,N_8805,N_6503);
nand U11185 (N_11185,N_6157,N_9555);
or U11186 (N_11186,N_8160,N_7853);
and U11187 (N_11187,N_7423,N_8634);
nor U11188 (N_11188,N_8714,N_5236);
nor U11189 (N_11189,N_6572,N_7285);
and U11190 (N_11190,N_8230,N_8474);
nand U11191 (N_11191,N_5797,N_6683);
or U11192 (N_11192,N_5235,N_5651);
and U11193 (N_11193,N_5681,N_6707);
nor U11194 (N_11194,N_7910,N_5256);
xor U11195 (N_11195,N_9644,N_9327);
nand U11196 (N_11196,N_6434,N_5572);
and U11197 (N_11197,N_5693,N_8574);
or U11198 (N_11198,N_9020,N_7370);
nand U11199 (N_11199,N_7067,N_6801);
and U11200 (N_11200,N_7621,N_8563);
nor U11201 (N_11201,N_5569,N_6671);
nand U11202 (N_11202,N_8138,N_9274);
or U11203 (N_11203,N_5260,N_8840);
and U11204 (N_11204,N_7210,N_8967);
or U11205 (N_11205,N_8781,N_9243);
and U11206 (N_11206,N_8669,N_7334);
or U11207 (N_11207,N_5811,N_9283);
nand U11208 (N_11208,N_5699,N_7544);
nand U11209 (N_11209,N_7379,N_5276);
or U11210 (N_11210,N_8071,N_8047);
and U11211 (N_11211,N_6040,N_7170);
and U11212 (N_11212,N_6988,N_6195);
nand U11213 (N_11213,N_5935,N_7034);
or U11214 (N_11214,N_8342,N_5591);
nand U11215 (N_11215,N_5854,N_5829);
and U11216 (N_11216,N_7039,N_5223);
and U11217 (N_11217,N_8414,N_7223);
nor U11218 (N_11218,N_9378,N_8662);
and U11219 (N_11219,N_9578,N_6200);
nor U11220 (N_11220,N_5502,N_8758);
nand U11221 (N_11221,N_6956,N_6705);
nand U11222 (N_11222,N_6213,N_9587);
nor U11223 (N_11223,N_9923,N_5027);
xnor U11224 (N_11224,N_6328,N_5314);
and U11225 (N_11225,N_8369,N_6508);
nand U11226 (N_11226,N_7597,N_9963);
and U11227 (N_11227,N_9115,N_6862);
nor U11228 (N_11228,N_6646,N_8381);
or U11229 (N_11229,N_7767,N_7454);
nor U11230 (N_11230,N_7976,N_5702);
nor U11231 (N_11231,N_6140,N_6743);
or U11232 (N_11232,N_5036,N_9962);
or U11233 (N_11233,N_8076,N_6708);
nor U11234 (N_11234,N_6719,N_9951);
and U11235 (N_11235,N_5978,N_7872);
and U11236 (N_11236,N_5316,N_7466);
nor U11237 (N_11237,N_6425,N_6253);
or U11238 (N_11238,N_9570,N_8644);
nand U11239 (N_11239,N_8302,N_9444);
or U11240 (N_11240,N_5672,N_9604);
nand U11241 (N_11241,N_9148,N_5976);
or U11242 (N_11242,N_5177,N_8901);
nand U11243 (N_11243,N_7724,N_5304);
and U11244 (N_11244,N_9595,N_7093);
nor U11245 (N_11245,N_8764,N_6826);
nand U11246 (N_11246,N_9659,N_5152);
and U11247 (N_11247,N_5429,N_6299);
nand U11248 (N_11248,N_7745,N_6235);
and U11249 (N_11249,N_6141,N_7638);
or U11250 (N_11250,N_5640,N_8765);
nor U11251 (N_11251,N_6547,N_9786);
nand U11252 (N_11252,N_8616,N_8943);
nand U11253 (N_11253,N_6628,N_5817);
or U11254 (N_11254,N_5001,N_7432);
and U11255 (N_11255,N_9591,N_9164);
and U11256 (N_11256,N_6518,N_5229);
and U11257 (N_11257,N_5945,N_9140);
or U11258 (N_11258,N_7975,N_5418);
and U11259 (N_11259,N_6768,N_5180);
nor U11260 (N_11260,N_7772,N_7351);
or U11261 (N_11261,N_5070,N_7374);
or U11262 (N_11262,N_7422,N_5159);
or U11263 (N_11263,N_8870,N_9224);
and U11264 (N_11264,N_8874,N_9800);
nand U11265 (N_11265,N_6592,N_5441);
and U11266 (N_11266,N_8554,N_9915);
nand U11267 (N_11267,N_9008,N_7819);
and U11268 (N_11268,N_7812,N_9437);
or U11269 (N_11269,N_9785,N_7998);
nor U11270 (N_11270,N_8603,N_7521);
nor U11271 (N_11271,N_6591,N_6317);
or U11272 (N_11272,N_7543,N_5998);
or U11273 (N_11273,N_5798,N_6713);
nor U11274 (N_11274,N_9737,N_9349);
and U11275 (N_11275,N_9012,N_7991);
nor U11276 (N_11276,N_7622,N_5951);
and U11277 (N_11277,N_5541,N_6369);
or U11278 (N_11278,N_5882,N_5296);
nand U11279 (N_11279,N_5509,N_7095);
and U11280 (N_11280,N_8798,N_7284);
or U11281 (N_11281,N_9196,N_9221);
and U11282 (N_11282,N_7262,N_7832);
or U11283 (N_11283,N_9778,N_8271);
nor U11284 (N_11284,N_9590,N_6912);
nor U11285 (N_11285,N_8797,N_7349);
nand U11286 (N_11286,N_6582,N_6634);
nand U11287 (N_11287,N_7286,N_6842);
or U11288 (N_11288,N_8557,N_5609);
nand U11289 (N_11289,N_8500,N_5741);
or U11290 (N_11290,N_6255,N_6764);
or U11291 (N_11291,N_9707,N_7312);
nor U11292 (N_11292,N_7315,N_8282);
and U11293 (N_11293,N_5919,N_5760);
and U11294 (N_11294,N_7409,N_6319);
or U11295 (N_11295,N_5347,N_7090);
nand U11296 (N_11296,N_5023,N_7503);
nor U11297 (N_11297,N_7251,N_9537);
and U11298 (N_11298,N_5987,N_7909);
nand U11299 (N_11299,N_6050,N_9455);
or U11300 (N_11300,N_9586,N_8127);
or U11301 (N_11301,N_9793,N_6760);
or U11302 (N_11302,N_6022,N_6824);
or U11303 (N_11303,N_5461,N_6828);
and U11304 (N_11304,N_9135,N_6237);
nand U11305 (N_11305,N_7455,N_9004);
or U11306 (N_11306,N_6165,N_9890);
nor U11307 (N_11307,N_6800,N_8472);
nand U11308 (N_11308,N_7005,N_5504);
nor U11309 (N_11309,N_5193,N_9419);
and U11310 (N_11310,N_9612,N_6461);
or U11311 (N_11311,N_7584,N_6226);
and U11312 (N_11312,N_8065,N_8261);
nor U11313 (N_11313,N_5843,N_6720);
or U11314 (N_11314,N_6641,N_6845);
and U11315 (N_11315,N_6939,N_5312);
nand U11316 (N_11316,N_5149,N_5246);
nor U11317 (N_11317,N_9244,N_6852);
nor U11318 (N_11318,N_6041,N_9275);
nand U11319 (N_11319,N_7448,N_6420);
nand U11320 (N_11320,N_6436,N_8293);
or U11321 (N_11321,N_6753,N_5861);
and U11322 (N_11322,N_5792,N_8635);
or U11323 (N_11323,N_7673,N_5653);
nand U11324 (N_11324,N_5857,N_7806);
or U11325 (N_11325,N_6482,N_9863);
nand U11326 (N_11326,N_9613,N_7387);
and U11327 (N_11327,N_8077,N_7406);
and U11328 (N_11328,N_6915,N_7623);
and U11329 (N_11329,N_6769,N_9117);
nand U11330 (N_11330,N_9541,N_5864);
nand U11331 (N_11331,N_9571,N_6086);
or U11332 (N_11332,N_9710,N_6084);
nand U11333 (N_11333,N_5191,N_5631);
or U11334 (N_11334,N_7274,N_8971);
nor U11335 (N_11335,N_5991,N_7398);
or U11336 (N_11336,N_5359,N_5615);
nand U11337 (N_11337,N_9780,N_5731);
and U11338 (N_11338,N_8551,N_5372);
and U11339 (N_11339,N_5706,N_5675);
nor U11340 (N_11340,N_5014,N_7582);
nand U11341 (N_11341,N_8791,N_5257);
nor U11342 (N_11342,N_7282,N_6410);
nand U11343 (N_11343,N_7615,N_8118);
nor U11344 (N_11344,N_9099,N_6476);
nand U11345 (N_11345,N_5678,N_5767);
and U11346 (N_11346,N_8711,N_6729);
nor U11347 (N_11347,N_8891,N_9626);
and U11348 (N_11348,N_6288,N_7495);
nor U11349 (N_11349,N_6146,N_6541);
and U11350 (N_11350,N_6107,N_8600);
and U11351 (N_11351,N_5542,N_6627);
or U11352 (N_11352,N_7565,N_7874);
and U11353 (N_11353,N_8636,N_8610);
or U11354 (N_11354,N_9964,N_7030);
nor U11355 (N_11355,N_9834,N_8305);
nor U11356 (N_11356,N_9057,N_9711);
xnor U11357 (N_11357,N_7741,N_8825);
and U11358 (N_11358,N_6927,N_9294);
nor U11359 (N_11359,N_5174,N_7430);
nor U11360 (N_11360,N_7190,N_8535);
nand U11361 (N_11361,N_6844,N_9986);
nand U11362 (N_11362,N_9143,N_5102);
nor U11363 (N_11363,N_5029,N_6662);
nor U11364 (N_11364,N_8182,N_7008);
and U11365 (N_11365,N_7707,N_9235);
nand U11366 (N_11366,N_5151,N_8285);
and U11367 (N_11367,N_5146,N_6907);
nor U11368 (N_11368,N_5886,N_9799);
and U11369 (N_11369,N_9593,N_9025);
and U11370 (N_11370,N_6869,N_8736);
nand U11371 (N_11371,N_5571,N_6691);
nand U11372 (N_11372,N_9683,N_6485);
and U11373 (N_11373,N_9267,N_9250);
or U11374 (N_11374,N_5282,N_7396);
or U11375 (N_11375,N_5002,N_7142);
or U11376 (N_11376,N_5400,N_5293);
or U11377 (N_11377,N_5328,N_7178);
or U11378 (N_11378,N_8640,N_8153);
nor U11379 (N_11379,N_5949,N_6069);
or U11380 (N_11380,N_6358,N_7120);
nor U11381 (N_11381,N_9819,N_5637);
nor U11382 (N_11382,N_6761,N_8362);
nor U11383 (N_11383,N_7736,N_9000);
or U11384 (N_11384,N_6184,N_7691);
nand U11385 (N_11385,N_7697,N_8375);
nand U11386 (N_11386,N_8470,N_9331);
nand U11387 (N_11387,N_6655,N_6645);
nand U11388 (N_11388,N_6762,N_6353);
nand U11389 (N_11389,N_9246,N_8198);
nor U11390 (N_11390,N_9848,N_9519);
and U11391 (N_11391,N_7022,N_6924);
nor U11392 (N_11392,N_5355,N_6695);
nand U11393 (N_11393,N_5239,N_9023);
nand U11394 (N_11394,N_8743,N_9120);
or U11395 (N_11395,N_5674,N_5272);
nor U11396 (N_11396,N_7357,N_9467);
or U11397 (N_11397,N_8390,N_8201);
and U11398 (N_11398,N_5720,N_5464);
nor U11399 (N_11399,N_7047,N_6360);
nand U11400 (N_11400,N_5593,N_8272);
nor U11401 (N_11401,N_9546,N_7881);
nor U11402 (N_11402,N_5603,N_9685);
nor U11403 (N_11403,N_5885,N_7919);
nand U11404 (N_11404,N_9950,N_5427);
or U11405 (N_11405,N_8008,N_7600);
nand U11406 (N_11406,N_8617,N_7546);
and U11407 (N_11407,N_7901,N_7964);
and U11408 (N_11408,N_8237,N_8388);
nand U11409 (N_11409,N_5916,N_7195);
xor U11410 (N_11410,N_5501,N_9351);
and U11411 (N_11411,N_8879,N_8205);
nand U11412 (N_11412,N_8749,N_7879);
nor U11413 (N_11413,N_6580,N_6143);
and U11414 (N_11414,N_8742,N_5646);
and U11415 (N_11415,N_8374,N_9134);
nor U11416 (N_11416,N_5340,N_6969);
and U11417 (N_11417,N_5692,N_7571);
or U11418 (N_11418,N_8094,N_5633);
nor U11419 (N_11419,N_9953,N_9690);
nand U11420 (N_11420,N_6979,N_8315);
or U11421 (N_11421,N_7028,N_7268);
or U11422 (N_11422,N_8242,N_7083);
and U11423 (N_11423,N_7275,N_9594);
xor U11424 (N_11424,N_9187,N_5469);
nor U11425 (N_11425,N_7102,N_9204);
and U11426 (N_11426,N_9483,N_7236);
or U11427 (N_11427,N_9810,N_9212);
or U11428 (N_11428,N_5160,N_9927);
or U11429 (N_11429,N_8356,N_9742);
nor U11430 (N_11430,N_9944,N_6922);
nand U11431 (N_11431,N_7713,N_9287);
nand U11432 (N_11432,N_8933,N_9449);
nand U11433 (N_11433,N_8218,N_5209);
nand U11434 (N_11434,N_7891,N_7636);
nand U11435 (N_11435,N_6990,N_8732);
nor U11436 (N_11436,N_6699,N_6136);
or U11437 (N_11437,N_8197,N_5395);
nor U11438 (N_11438,N_7595,N_6023);
nor U11439 (N_11439,N_6733,N_9565);
or U11440 (N_11440,N_5013,N_9424);
or U11441 (N_11441,N_6794,N_6449);
nor U11442 (N_11442,N_7514,N_6909);
nor U11443 (N_11443,N_6351,N_6700);
or U11444 (N_11444,N_5253,N_5307);
or U11445 (N_11445,N_9596,N_6888);
or U11446 (N_11446,N_7465,N_7682);
and U11447 (N_11447,N_5980,N_8729);
and U11448 (N_11448,N_7769,N_7007);
and U11449 (N_11449,N_7044,N_8531);
nor U11450 (N_11450,N_8818,N_8993);
nor U11451 (N_11451,N_5617,N_5112);
nand U11452 (N_11452,N_8829,N_7483);
nand U11453 (N_11453,N_7531,N_7031);
and U11454 (N_11454,N_5311,N_5374);
nand U11455 (N_11455,N_6494,N_6731);
and U11456 (N_11456,N_6716,N_7743);
or U11457 (N_11457,N_7644,N_7886);
nand U11458 (N_11458,N_9540,N_7360);
nor U11459 (N_11459,N_9547,N_8310);
nand U11460 (N_11460,N_6936,N_6550);
nand U11461 (N_11461,N_6406,N_6680);
or U11462 (N_11462,N_9835,N_7192);
nor U11463 (N_11463,N_9705,N_7023);
nand U11464 (N_11464,N_6341,N_9531);
nor U11465 (N_11465,N_9414,N_8322);
nor U11466 (N_11466,N_8833,N_5597);
or U11467 (N_11467,N_6563,N_8335);
nand U11468 (N_11468,N_5518,N_8850);
nand U11469 (N_11469,N_6139,N_7446);
nand U11470 (N_11470,N_9723,N_8665);
and U11471 (N_11471,N_6189,N_6654);
and U11472 (N_11472,N_5208,N_9056);
and U11473 (N_11473,N_7447,N_9239);
and U11474 (N_11474,N_9031,N_6168);
xor U11475 (N_11475,N_7580,N_8192);
nand U11476 (N_11476,N_7281,N_8070);
nand U11477 (N_11477,N_6799,N_5536);
or U11478 (N_11478,N_8904,N_7664);
nor U11479 (N_11479,N_6042,N_8112);
and U11480 (N_11480,N_8948,N_9855);
and U11481 (N_11481,N_8730,N_5286);
nor U11482 (N_11482,N_5873,N_9858);
and U11483 (N_11483,N_5039,N_9932);
nand U11484 (N_11484,N_5598,N_7320);
and U11485 (N_11485,N_8379,N_5292);
or U11486 (N_11486,N_9516,N_6577);
or U11487 (N_11487,N_7592,N_8692);
and U11488 (N_11488,N_8566,N_6018);
nor U11489 (N_11489,N_6177,N_6297);
nand U11490 (N_11490,N_8885,N_5350);
and U11491 (N_11491,N_5684,N_8026);
or U11492 (N_11492,N_6443,N_5975);
nand U11493 (N_11493,N_5914,N_6536);
nand U11494 (N_11494,N_5781,N_5131);
nor U11495 (N_11495,N_7264,N_8004);
nand U11496 (N_11496,N_7237,N_7612);
and U11497 (N_11497,N_9893,N_7011);
nor U11498 (N_11498,N_6521,N_8854);
nor U11499 (N_11499,N_5834,N_5318);
nor U11500 (N_11500,N_6615,N_9184);
nor U11501 (N_11501,N_8296,N_9217);
and U11502 (N_11502,N_7222,N_7354);
or U11503 (N_11503,N_9371,N_7586);
or U11504 (N_11504,N_8404,N_6281);
and U11505 (N_11505,N_8130,N_8895);
or U11506 (N_11506,N_6831,N_7685);
nand U11507 (N_11507,N_5668,N_6642);
nand U11508 (N_11508,N_5492,N_7922);
or U11509 (N_11509,N_7169,N_9007);
nand U11510 (N_11510,N_8513,N_8081);
and U11511 (N_11511,N_5346,N_6321);
and U11512 (N_11512,N_8619,N_6193);
and U11513 (N_11513,N_8038,N_5932);
or U11514 (N_11514,N_8298,N_9713);
or U11515 (N_11515,N_8245,N_6395);
or U11516 (N_11516,N_7563,N_5100);
nand U11517 (N_11517,N_6966,N_9666);
and U11518 (N_11518,N_6891,N_7754);
or U11519 (N_11519,N_8908,N_7217);
and U11520 (N_11520,N_5924,N_8154);
nand U11521 (N_11521,N_8066,N_9489);
nor U11522 (N_11522,N_5337,N_7863);
nand U11523 (N_11523,N_6145,N_5197);
nor U11524 (N_11524,N_7403,N_7929);
nand U11525 (N_11525,N_5777,N_5362);
nand U11526 (N_11526,N_5645,N_8773);
nand U11527 (N_11527,N_8010,N_9585);
and U11528 (N_11528,N_8646,N_7363);
nand U11529 (N_11529,N_7328,N_6774);
xnor U11530 (N_11530,N_8150,N_7247);
nand U11531 (N_11531,N_9956,N_6668);
and U11532 (N_11532,N_9813,N_5782);
and U11533 (N_11533,N_6940,N_7894);
nor U11534 (N_11534,N_9506,N_6430);
and U11535 (N_11535,N_7512,N_7548);
nand U11536 (N_11536,N_8583,N_5845);
or U11537 (N_11537,N_6567,N_7362);
and U11538 (N_11538,N_5718,N_7016);
nor U11539 (N_11539,N_6057,N_6597);
or U11540 (N_11540,N_8495,N_5363);
and U11541 (N_11541,N_5881,N_6378);
nor U11542 (N_11542,N_7787,N_9618);
and U11543 (N_11543,N_8067,N_9728);
nor U11544 (N_11544,N_8317,N_6259);
or U11545 (N_11545,N_7166,N_9421);
nor U11546 (N_11546,N_7452,N_7436);
nor U11547 (N_11547,N_7025,N_7999);
xnor U11548 (N_11548,N_5888,N_5589);
and U11549 (N_11549,N_5959,N_5278);
nor U11550 (N_11550,N_5444,N_7567);
nor U11551 (N_11551,N_7985,N_8873);
nand U11552 (N_11552,N_8530,N_7182);
nor U11553 (N_11553,N_9553,N_6925);
and U11554 (N_11554,N_5279,N_5288);
nor U11555 (N_11555,N_5153,N_5255);
and U11556 (N_11556,N_7803,N_6216);
or U11557 (N_11557,N_5137,N_6968);
nand U11558 (N_11558,N_7542,N_6094);
and U11559 (N_11559,N_7556,N_9925);
nand U11560 (N_11560,N_7440,N_6499);
nand U11561 (N_11561,N_9897,N_8532);
or U11562 (N_11562,N_5595,N_5165);
and U11563 (N_11563,N_9978,N_9307);
or U11564 (N_11564,N_8498,N_9333);
and U11565 (N_11565,N_6918,N_9528);
nor U11566 (N_11566,N_5244,N_8966);
or U11567 (N_11567,N_7570,N_5833);
and U11568 (N_11568,N_7866,N_7557);
or U11569 (N_11569,N_9102,N_9321);
or U11570 (N_11570,N_8893,N_7073);
and U11571 (N_11571,N_6423,N_8040);
and U11572 (N_11572,N_5641,N_7831);
nor U11573 (N_11573,N_6093,N_9129);
nor U11574 (N_11574,N_8627,N_8625);
and U11575 (N_11575,N_6551,N_6540);
or U11576 (N_11576,N_8731,N_8608);
and U11577 (N_11577,N_7206,N_6820);
or U11578 (N_11578,N_5121,N_8722);
xor U11579 (N_11579,N_5122,N_9263);
nor U11580 (N_11580,N_9202,N_6908);
or U11581 (N_11581,N_6863,N_9220);
xnor U11582 (N_11582,N_6230,N_9132);
or U11583 (N_11583,N_5333,N_9325);
and U11584 (N_11584,N_6077,N_6954);
nor U11585 (N_11585,N_9965,N_5867);
and U11586 (N_11586,N_6445,N_9290);
nand U11587 (N_11587,N_7808,N_8459);
or U11588 (N_11588,N_7468,N_6746);
or U11589 (N_11589,N_9567,N_5585);
nand U11590 (N_11590,N_5086,N_8361);
nor U11591 (N_11591,N_9717,N_9266);
nand U11592 (N_11592,N_6542,N_6156);
or U11593 (N_11593,N_5755,N_5405);
or U11594 (N_11594,N_7260,N_9615);
or U11595 (N_11595,N_6873,N_6882);
and U11596 (N_11596,N_6376,N_5428);
nor U11597 (N_11597,N_5269,N_5740);
nand U11598 (N_11598,N_5201,N_5115);
xnor U11599 (N_11599,N_8216,N_7193);
and U11600 (N_11600,N_8808,N_5850);
or U11601 (N_11601,N_8682,N_9062);
nand U11602 (N_11602,N_6466,N_8092);
nor U11603 (N_11603,N_9480,N_5024);
nand U11604 (N_11604,N_9194,N_5022);
or U11605 (N_11605,N_6614,N_6847);
nand U11606 (N_11606,N_5411,N_7292);
and U11607 (N_11607,N_5649,N_6046);
and U11608 (N_11608,N_7990,N_6502);
nand U11609 (N_11609,N_6688,N_6911);
nand U11610 (N_11610,N_9191,N_9638);
or U11611 (N_11611,N_9446,N_5923);
nand U11612 (N_11612,N_5776,N_6191);
nor U11613 (N_11613,N_8405,N_5665);
or U11614 (N_11614,N_5046,N_6519);
and U11615 (N_11615,N_9330,N_8486);
nor U11616 (N_11616,N_7024,N_6511);
nor U11617 (N_11617,N_9797,N_6242);
nor U11618 (N_11618,N_9782,N_9806);
nor U11619 (N_11619,N_9627,N_5238);
or U11620 (N_11620,N_6590,N_8223);
or U11621 (N_11621,N_8613,N_8940);
nor U11622 (N_11622,N_7861,N_5723);
nor U11623 (N_11623,N_9385,N_9005);
nand U11624 (N_11624,N_8620,N_7258);
or U11625 (N_11625,N_5041,N_8430);
nand U11626 (N_11626,N_9732,N_6393);
nor U11627 (N_11627,N_7967,N_8014);
and U11628 (N_11628,N_8195,N_9750);
nor U11629 (N_11629,N_7833,N_9983);
nand U11630 (N_11630,N_7811,N_8984);
nor U11631 (N_11631,N_9525,N_7124);
and U11632 (N_11632,N_8880,N_5547);
and U11633 (N_11633,N_7004,N_9549);
or U11634 (N_11634,N_8655,N_9877);
and U11635 (N_11635,N_8075,N_6112);
or U11636 (N_11636,N_8171,N_7940);
or U11637 (N_11637,N_8537,N_8962);
nor U11638 (N_11638,N_6399,N_7660);
nor U11639 (N_11639,N_7479,N_8445);
and U11640 (N_11640,N_6205,N_6031);
and U11641 (N_11641,N_5034,N_8483);
or U11642 (N_11642,N_8186,N_9167);
and U11643 (N_11643,N_5537,N_8093);
nor U11644 (N_11644,N_5508,N_6470);
or U11645 (N_11645,N_9411,N_8143);
or U11646 (N_11646,N_8300,N_9001);
and U11647 (N_11647,N_8497,N_6861);
or U11648 (N_11648,N_8755,N_5482);
or U11649 (N_11649,N_5391,N_5003);
and U11650 (N_11650,N_7717,N_7710);
and U11651 (N_11651,N_5138,N_9543);
or U11652 (N_11652,N_8950,N_7749);
nor U11653 (N_11653,N_5440,N_9069);
or U11654 (N_11654,N_5299,N_7988);
or U11655 (N_11655,N_7269,N_5545);
nor U11656 (N_11656,N_8776,N_9047);
or U11657 (N_11657,N_6669,N_5189);
nand U11658 (N_11658,N_7154,N_5680);
nand U11659 (N_11659,N_7175,N_5527);
xor U11660 (N_11660,N_6151,N_7048);
nor U11661 (N_11661,N_8012,N_6015);
or U11662 (N_11662,N_5018,N_8215);
or U11663 (N_11663,N_6488,N_8865);
nand U11664 (N_11664,N_5402,N_7758);
or U11665 (N_11665,N_6439,N_7778);
nor U11666 (N_11666,N_5960,N_5051);
and U11667 (N_11667,N_7918,N_9402);
nor U11668 (N_11668,N_9719,N_6188);
or U11669 (N_11669,N_9842,N_7019);
or U11670 (N_11670,N_9614,N_9015);
and U11671 (N_11671,N_9354,N_9039);
nor U11672 (N_11672,N_6672,N_9664);
nand U11673 (N_11673,N_8979,N_8704);
nand U11674 (N_11674,N_5040,N_5981);
nor U11675 (N_11675,N_8308,N_9319);
nand U11676 (N_11676,N_6745,N_6640);
and U11677 (N_11677,N_7368,N_9313);
nor U11678 (N_11678,N_5729,N_6561);
and U11679 (N_11679,N_7461,N_9545);
nand U11680 (N_11680,N_5968,N_8912);
nand U11681 (N_11681,N_9734,N_5423);
or U11682 (N_11682,N_9119,N_9384);
or U11683 (N_11683,N_9794,N_5389);
nor U11684 (N_11684,N_5163,N_5634);
nand U11685 (N_11685,N_8489,N_5080);
and U11686 (N_11686,N_8145,N_6910);
or U11687 (N_11687,N_6090,N_8259);
nand U11688 (N_11688,N_5187,N_8206);
and U11689 (N_11689,N_7934,N_8719);
and U11690 (N_11690,N_7579,N_5709);
nor U11691 (N_11691,N_5462,N_6490);
xnor U11692 (N_11692,N_7655,N_8572);
and U11693 (N_11693,N_7106,N_8318);
or U11694 (N_11694,N_7610,N_5648);
nand U11695 (N_11695,N_5847,N_5514);
nand U11696 (N_11696,N_9254,N_6903);
nor U11697 (N_11697,N_6725,N_6578);
or U11698 (N_11698,N_6368,N_5763);
nor U11699 (N_11699,N_7550,N_9605);
or U11700 (N_11700,N_9874,N_6935);
or U11701 (N_11701,N_8678,N_7259);
nor U11702 (N_11702,N_6589,N_9180);
nand U11703 (N_11703,N_8685,N_8705);
nor U11704 (N_11704,N_5421,N_9492);
nor U11705 (N_11705,N_7068,N_9691);
or U11706 (N_11706,N_5262,N_8787);
and U11707 (N_11707,N_9760,N_9142);
and U11708 (N_11708,N_6292,N_8816);
nand U11709 (N_11709,N_5019,N_7747);
or U11710 (N_11710,N_5179,N_6970);
nand U11711 (N_11711,N_7844,N_5064);
nand U11712 (N_11712,N_6834,N_8107);
or U11713 (N_11713,N_8849,N_7161);
or U11714 (N_11714,N_8403,N_9328);
and U11715 (N_11715,N_5188,N_5103);
and U11716 (N_11716,N_8831,N_7796);
and U11717 (N_11717,N_5992,N_5918);
nor U11718 (N_11718,N_8286,N_8522);
and U11719 (N_11719,N_5085,N_7606);
nor U11720 (N_11720,N_8103,N_9255);
and U11721 (N_11721,N_6246,N_9145);
nor U11722 (N_11722,N_7233,N_7792);
nor U11723 (N_11723,N_8448,N_6674);
or U11724 (N_11724,N_5207,N_9789);
nor U11725 (N_11725,N_7947,N_6349);
or U11726 (N_11726,N_6984,N_5573);
nor U11727 (N_11727,N_7092,N_9736);
or U11728 (N_11728,N_5315,N_9853);
or U11729 (N_11729,N_8227,N_9470);
nand U11730 (N_11730,N_6076,N_7791);
nand U11731 (N_11731,N_8452,N_6282);
nand U11732 (N_11732,N_5701,N_9609);
or U11733 (N_11733,N_6635,N_6796);
nand U11734 (N_11734,N_5473,N_8124);
and U11735 (N_11735,N_6272,N_6427);
nor U11736 (N_11736,N_6599,N_8330);
xor U11737 (N_11737,N_7562,N_9684);
nand U11738 (N_11738,N_5463,N_6624);
nand U11739 (N_11739,N_5712,N_6072);
nand U11740 (N_11740,N_6982,N_7972);
or U11741 (N_11741,N_7805,N_8502);
or U11742 (N_11742,N_8939,N_7577);
or U11743 (N_11743,N_7293,N_6838);
and U11744 (N_11744,N_5413,N_6885);
nor U11745 (N_11745,N_5984,N_7905);
or U11746 (N_11746,N_5099,N_8233);
nor U11747 (N_11747,N_7449,N_5908);
nor U11748 (N_11748,N_5915,N_7641);
and U11749 (N_11749,N_9079,N_5050);
and U11750 (N_11750,N_7035,N_7070);
nand U11751 (N_11751,N_6357,N_6790);
or U11752 (N_11752,N_9403,N_6228);
or U11753 (N_11753,N_5715,N_9201);
nor U11754 (N_11754,N_7373,N_6600);
nand U11755 (N_11755,N_7764,N_9818);
or U11756 (N_11756,N_9078,N_8937);
or U11757 (N_11757,N_9857,N_9859);
and U11758 (N_11758,N_5531,N_8254);
or U11759 (N_11759,N_8651,N_6832);
or U11760 (N_11760,N_9066,N_8212);
or U11761 (N_11761,N_7197,N_7653);
or U11762 (N_11762,N_9300,N_7074);
and U11763 (N_11763,N_8432,N_9577);
and U11764 (N_11764,N_5814,N_9643);
and U11765 (N_11765,N_9938,N_5126);
nor U11766 (N_11766,N_5093,N_7296);
xor U11767 (N_11767,N_8191,N_8476);
nand U11768 (N_11768,N_9738,N_5465);
nand U11769 (N_11769,N_5830,N_8151);
nand U11770 (N_11770,N_9805,N_8161);
nor U11771 (N_11771,N_6066,N_8165);
and U11772 (N_11772,N_7235,N_9937);
nor U11773 (N_11773,N_5228,N_5517);
and U11774 (N_11774,N_8341,N_5452);
or U11775 (N_11775,N_6895,N_6070);
nand U11776 (N_11776,N_8156,N_7491);
nand U11777 (N_11777,N_9169,N_9522);
nand U11778 (N_11778,N_8657,N_5484);
nand U11779 (N_11779,N_8325,N_6115);
nor U11780 (N_11780,N_9021,N_8431);
nor U11781 (N_11781,N_9884,N_5069);
or U11782 (N_11782,N_7470,N_9775);
or U11783 (N_11783,N_5828,N_8695);
or U11784 (N_11784,N_5497,N_5342);
nor U11785 (N_11785,N_7552,N_8126);
and U11786 (N_11786,N_9628,N_5963);
nand U11787 (N_11787,N_9303,N_8062);
nor U11788 (N_11788,N_9875,N_5147);
nor U11789 (N_11789,N_7224,N_5226);
or U11790 (N_11790,N_9207,N_7802);
or U11791 (N_11791,N_6980,N_9846);
or U11792 (N_11792,N_6119,N_5910);
and U11793 (N_11793,N_5390,N_5232);
and U11794 (N_11794,N_6901,N_8534);
nand U11795 (N_11795,N_9259,N_6693);
nor U11796 (N_11796,N_9579,N_5267);
or U11797 (N_11797,N_7994,N_7780);
nand U11798 (N_11798,N_9406,N_9484);
or U11799 (N_11799,N_5820,N_7973);
nor U11800 (N_11800,N_6809,N_7138);
nand U11801 (N_11801,N_5732,N_8085);
or U11802 (N_11802,N_8457,N_8059);
and U11803 (N_11803,N_9696,N_5432);
and U11804 (N_11804,N_8509,N_7840);
or U11805 (N_11805,N_6786,N_7912);
nor U11806 (N_11806,N_5616,N_8826);
nand U11807 (N_11807,N_9554,N_5890);
and U11808 (N_11808,N_9636,N_7322);
nor U11809 (N_11809,N_8994,N_6664);
nor U11810 (N_11810,N_9767,N_6897);
and U11811 (N_11811,N_6585,N_8407);
or U11812 (N_11812,N_5079,N_6362);
and U11813 (N_11813,N_6192,N_5522);
nor U11814 (N_11814,N_8162,N_7876);
nand U11815 (N_11815,N_8587,N_5092);
nand U11816 (N_11816,N_7834,N_8579);
or U11817 (N_11817,N_9162,N_5420);
and U11818 (N_11818,N_6276,N_9038);
nor U11819 (N_11819,N_7444,N_8852);
and U11820 (N_11820,N_8738,N_8270);
or U11821 (N_11821,N_9216,N_8853);
nor U11822 (N_11822,N_5116,N_5948);
and U11823 (N_11823,N_5495,N_6456);
nor U11824 (N_11824,N_8311,N_8351);
or U11825 (N_11825,N_5216,N_7185);
and U11826 (N_11826,N_7652,N_5135);
nand U11827 (N_11827,N_6043,N_8688);
or U11828 (N_11828,N_9149,N_5758);
nand U11829 (N_11829,N_6014,N_9237);
and U11830 (N_11830,N_5196,N_8005);
or U11831 (N_11831,N_9867,N_9081);
and U11832 (N_11832,N_7629,N_8423);
and U11833 (N_11833,N_8593,N_8916);
nand U11834 (N_11834,N_7828,N_6326);
nor U11835 (N_11835,N_8056,N_8869);
and U11836 (N_11836,N_5364,N_5448);
nand U11837 (N_11837,N_9316,N_9617);
nand U11838 (N_11838,N_8276,N_6258);
nand U11839 (N_11839,N_5694,N_7719);
xor U11840 (N_11840,N_6401,N_8329);
and U11841 (N_11841,N_9939,N_6780);
nand U11842 (N_11842,N_9856,N_6340);
xor U11843 (N_11843,N_8868,N_5143);
nand U11844 (N_11844,N_6172,N_9306);
and U11845 (N_11845,N_7578,N_6726);
and U11846 (N_11846,N_6920,N_9118);
nand U11847 (N_11847,N_9726,N_9336);
nor U11848 (N_11848,N_7760,N_7402);
and U11849 (N_11849,N_7753,N_8813);
nand U11850 (N_11850,N_6816,N_5869);
and U11851 (N_11851,N_5966,N_9990);
or U11852 (N_11852,N_7854,N_8116);
or U11853 (N_11853,N_6477,N_6986);
nor U11854 (N_11854,N_9343,N_7017);
and U11855 (N_11855,N_7359,N_9909);
or U11856 (N_11856,N_7100,N_8119);
or U11857 (N_11857,N_8945,N_8586);
and U11858 (N_11858,N_7810,N_8519);
nand U11859 (N_11859,N_9447,N_8017);
nor U11860 (N_11860,N_8568,N_9741);
nand U11861 (N_11861,N_9277,N_6028);
nand U11862 (N_11862,N_9523,N_6493);
nor U11863 (N_11863,N_9346,N_7979);
or U11864 (N_11864,N_7199,N_8898);
nand U11865 (N_11865,N_7002,N_6012);
nand U11866 (N_11866,N_8105,N_7896);
and U11867 (N_11867,N_6035,N_8464);
nand U11868 (N_11868,N_6663,N_6217);
or U11869 (N_11869,N_6878,N_9885);
and U11870 (N_11870,N_5011,N_6718);
nor U11871 (N_11871,N_9697,N_5017);
or U11872 (N_11872,N_9332,N_9478);
nor U11873 (N_11873,N_9390,N_6703);
nor U11874 (N_11874,N_5356,N_9442);
or U11875 (N_11875,N_6837,N_8964);
or U11876 (N_11876,N_7467,N_7339);
nor U11877 (N_11877,N_6446,N_8180);
nand U11878 (N_11878,N_6787,N_6366);
and U11879 (N_11879,N_8429,N_7365);
nand U11880 (N_11880,N_6758,N_9564);
nand U11881 (N_11881,N_8783,N_9389);
and U11882 (N_11882,N_9358,N_5425);
nor U11883 (N_11883,N_9369,N_8352);
or U11884 (N_11884,N_8894,N_6659);
nand U11885 (N_11885,N_5856,N_7341);
nor U11886 (N_11886,N_9159,N_8545);
or U11887 (N_11887,N_6038,N_5939);
and U11888 (N_11888,N_8248,N_9881);
nor U11889 (N_11889,N_8989,N_6462);
nand U11890 (N_11890,N_9999,N_8929);
and U11891 (N_11891,N_7263,N_7194);
nor U11892 (N_11892,N_8946,N_8372);
or U11893 (N_11893,N_6525,N_7924);
nor U11894 (N_11894,N_5240,N_5730);
nand U11895 (N_11895,N_8618,N_6457);
or U11896 (N_11896,N_6053,N_5049);
nand U11897 (N_11897,N_7167,N_6287);
or U11898 (N_11898,N_9445,N_7415);
nand U11899 (N_11899,N_6183,N_8708);
nand U11900 (N_11900,N_5450,N_9727);
nand U11901 (N_11901,N_9179,N_9671);
or U11902 (N_11902,N_8741,N_8569);
nor U11903 (N_11903,N_6065,N_6886);
and U11904 (N_11904,N_9542,N_9847);
nor U11905 (N_11905,N_9486,N_7164);
or U11906 (N_11906,N_7018,N_6538);
and U11907 (N_11907,N_9043,N_9104);
or U11908 (N_11908,N_8134,N_9911);
or U11909 (N_11909,N_7818,N_7956);
or U11910 (N_11910,N_6313,N_9692);
nor U11911 (N_11911,N_6247,N_7009);
and U11912 (N_11912,N_5676,N_5329);
nor U11913 (N_11913,N_5025,N_8621);
nor U11914 (N_11914,N_6892,N_8649);
nand U11915 (N_11915,N_9854,N_6377);
nor U11916 (N_11916,N_6906,N_9318);
nor U11917 (N_11917,N_7382,N_8560);
nand U11918 (N_11918,N_6394,N_9647);
xor U11919 (N_11919,N_5691,N_9920);
and U11920 (N_11920,N_9724,N_8504);
nand U11921 (N_11921,N_7862,N_7196);
nor U11922 (N_11922,N_5490,N_8920);
or U11923 (N_11923,N_7948,N_9774);
nor U11924 (N_11924,N_8789,N_6723);
or U11925 (N_11925,N_6342,N_9536);
and U11926 (N_11926,N_7372,N_9689);
nand U11927 (N_11927,N_7064,N_7459);
nand U11928 (N_11928,N_8007,N_5129);
nor U11929 (N_11929,N_9393,N_7243);
and U11930 (N_11930,N_7575,N_8629);
xnor U11931 (N_11931,N_6602,N_6904);
or U11932 (N_11932,N_7513,N_7475);
nor U11933 (N_11933,N_6080,N_8121);
or U11934 (N_11934,N_8419,N_9985);
and U11935 (N_11935,N_8170,N_9879);
and U11936 (N_11936,N_5756,N_9128);
and U11937 (N_11937,N_9731,N_9138);
or U11938 (N_11938,N_9257,N_9894);
xnor U11939 (N_11939,N_6739,N_7086);
or U11940 (N_11940,N_6706,N_5324);
nand U11941 (N_11941,N_6952,N_7737);
or U11942 (N_11942,N_7520,N_7708);
xor U11943 (N_11943,N_6418,N_5512);
and U11944 (N_11944,N_9748,N_6391);
nand U11945 (N_11945,N_7201,N_9456);
and U11946 (N_11946,N_5625,N_8900);
xnor U11947 (N_11947,N_7926,N_9702);
and U11948 (N_11948,N_5543,N_7530);
nand U11949 (N_11949,N_6815,N_9704);
and U11950 (N_11950,N_7981,N_9386);
nor U11951 (N_11951,N_9629,N_5559);
or U11952 (N_11952,N_9182,N_7227);
or U11953 (N_11953,N_8753,N_7089);
and U11954 (N_11954,N_9866,N_7168);
nor U11955 (N_11955,N_8354,N_7779);
nor U11956 (N_11956,N_5472,N_7241);
or U11957 (N_11957,N_8931,N_6690);
nor U11958 (N_11958,N_5601,N_8045);
or U11959 (N_11959,N_9320,N_7134);
nor U11960 (N_11960,N_5006,N_9961);
and U11961 (N_11961,N_8080,N_6355);
nand U11962 (N_11962,N_6024,N_9607);
nor U11963 (N_11963,N_6643,N_9803);
nor U11964 (N_11964,N_6312,N_7191);
nand U11965 (N_11965,N_9701,N_6330);
nand U11966 (N_11966,N_8975,N_9075);
or U11967 (N_11967,N_8133,N_9610);
nor U11968 (N_11968,N_8694,N_5105);
or U11969 (N_11969,N_9749,N_8023);
or U11970 (N_11970,N_6532,N_7675);
nor U11971 (N_11971,N_5619,N_8609);
and U11972 (N_11972,N_9899,N_8033);
xor U11973 (N_11973,N_7618,N_9107);
nor U11974 (N_11974,N_7783,N_6766);
and U11975 (N_11975,N_7330,N_7765);
and U11976 (N_11976,N_8412,N_6932);
nor U11977 (N_11977,N_9966,N_9229);
nor U11978 (N_11978,N_5535,N_5393);
nor U11979 (N_11979,N_7378,N_8099);
and U11980 (N_11980,N_8487,N_5285);
nand U11981 (N_11981,N_8226,N_8482);
or U11982 (N_11982,N_7347,N_8928);
and U11983 (N_11983,N_5392,N_5751);
nand U11984 (N_11984,N_5909,N_5663);
nor U11985 (N_11985,N_8221,N_8355);
nand U11986 (N_11986,N_5422,N_8914);
nand U11987 (N_11987,N_7645,N_6163);
or U11988 (N_11988,N_5793,N_5842);
or U11989 (N_11989,N_6523,N_7054);
and U11990 (N_11990,N_5768,N_9024);
nand U11991 (N_11991,N_6851,N_8883);
nand U11992 (N_11992,N_5973,N_7519);
and U11993 (N_11993,N_8393,N_6417);
or U11994 (N_11994,N_7709,N_5274);
and U11995 (N_11995,N_7094,N_5394);
xnor U11996 (N_11996,N_6308,N_9345);
nand U11997 (N_11997,N_5398,N_6110);
nor U11998 (N_11998,N_9477,N_8320);
nand U11999 (N_11999,N_5477,N_5332);
or U12000 (N_12000,N_8111,N_5370);
nor U12001 (N_12001,N_7533,N_6871);
nand U12002 (N_12002,N_5417,N_7572);
nor U12003 (N_12003,N_5800,N_8169);
and U12004 (N_12004,N_5905,N_8523);
or U12005 (N_12005,N_6359,N_8701);
nor U12006 (N_12006,N_5430,N_8309);
or U12007 (N_12007,N_8737,N_9338);
and U12008 (N_12008,N_9037,N_6605);
nor U12009 (N_12009,N_6670,N_5671);
and U12010 (N_12010,N_7728,N_7906);
and U12011 (N_12011,N_6294,N_8088);
nor U12012 (N_12012,N_5925,N_5832);
nand U12013 (N_12013,N_6989,N_5704);
nand U12014 (N_12014,N_5804,N_7953);
nand U12015 (N_12015,N_7139,N_9131);
nand U12016 (N_12016,N_7085,N_5222);
nor U12017 (N_12017,N_8450,N_7825);
nor U12018 (N_12018,N_8417,N_6581);
and U12019 (N_12019,N_6426,N_5977);
and U12020 (N_12020,N_6185,N_8347);
and U12021 (N_12021,N_6458,N_7650);
nor U12022 (N_12022,N_5284,N_5173);
nand U12023 (N_12023,N_7041,N_6027);
or U12024 (N_12024,N_6240,N_9532);
or U12025 (N_12025,N_5983,N_8036);
and U12026 (N_12026,N_9606,N_9904);
nand U12027 (N_12027,N_6451,N_6822);
nand U12028 (N_12028,N_9708,N_8571);
and U12029 (N_12029,N_7696,N_8527);
nand U12030 (N_12030,N_8240,N_6285);
or U12031 (N_12031,N_7027,N_8684);
nand U12032 (N_12032,N_6829,N_7871);
and U12033 (N_12033,N_6323,N_7790);
nor U12034 (N_12034,N_7642,N_6254);
and U12035 (N_12035,N_8830,N_9759);
nor U12036 (N_12036,N_6088,N_9400);
and U12037 (N_12037,N_9688,N_9575);
and U12038 (N_12038,N_6867,N_6621);
and U12039 (N_12039,N_6978,N_8740);
xor U12040 (N_12040,N_7541,N_7212);
or U12041 (N_12041,N_7635,N_6948);
or U12042 (N_12042,N_9493,N_8999);
nor U12043 (N_12043,N_8763,N_6612);
or U12044 (N_12044,N_7695,N_6564);
nor U12045 (N_12045,N_8110,N_7267);
or U12046 (N_12046,N_9048,N_5513);
nand U12047 (N_12047,N_7418,N_6098);
or U12048 (N_12048,N_6868,N_7601);
nand U12049 (N_12049,N_8289,N_7055);
or U12050 (N_12050,N_7231,N_8492);
or U12051 (N_12051,N_6329,N_9625);
nor U12052 (N_12052,N_5091,N_7690);
and U12053 (N_12053,N_7136,N_7486);
nand U12054 (N_12054,N_6164,N_7428);
and U12055 (N_12055,N_5043,N_8422);
and U12056 (N_12056,N_6987,N_6818);
nand U12057 (N_12057,N_5283,N_5577);
and U12058 (N_12058,N_6995,N_8924);
xnor U12059 (N_12059,N_6416,N_5614);
nor U12060 (N_12060,N_7740,N_7460);
nor U12061 (N_12061,N_6919,N_9170);
nor U12062 (N_12062,N_7553,N_6202);
and U12063 (N_12063,N_5996,N_6233);
and U12064 (N_12064,N_8204,N_7949);
or U12065 (N_12065,N_9297,N_7680);
nand U12066 (N_12066,N_9829,N_7674);
or U12067 (N_12067,N_5309,N_8142);
or U12068 (N_12068,N_8125,N_5054);
nor U12069 (N_12069,N_9087,N_8053);
and U12070 (N_12070,N_9498,N_6413);
and U12071 (N_12071,N_5298,N_7489);
nand U12072 (N_12072,N_5021,N_7554);
nand U12073 (N_12073,N_5806,N_7369);
or U12074 (N_12074,N_9945,N_7858);
and U12075 (N_12075,N_7375,N_8190);
nand U12076 (N_12076,N_9864,N_7939);
and U12077 (N_12077,N_8804,N_9679);
nand U12078 (N_12078,N_7855,N_6946);
nor U12079 (N_12079,N_7982,N_6361);
nor U12080 (N_12080,N_7774,N_6898);
nand U12081 (N_12081,N_8444,N_6039);
and U12082 (N_12082,N_5799,N_6150);
or U12083 (N_12083,N_9245,N_8413);
and U12084 (N_12084,N_9948,N_7115);
or U12085 (N_12085,N_7842,N_9171);
and U12086 (N_12086,N_5584,N_6738);
and U12087 (N_12087,N_6271,N_6256);
or U12088 (N_12088,N_9112,N_7712);
and U12089 (N_12089,N_7658,N_6266);
or U12090 (N_12090,N_8231,N_5746);
nor U12091 (N_12091,N_9461,N_7560);
or U12092 (N_12092,N_8506,N_8229);
or U12093 (N_12093,N_6916,N_9474);
nand U12094 (N_12094,N_9496,N_9592);
or U12095 (N_12095,N_7628,N_7494);
or U12096 (N_12096,N_6118,N_6797);
or U12097 (N_12097,N_7248,N_6129);
nor U12098 (N_12098,N_8115,N_6749);
or U12099 (N_12099,N_5127,N_7962);
and U12100 (N_12100,N_9954,N_9880);
nand U12101 (N_12101,N_7870,N_7128);
and U12102 (N_12102,N_9225,N_5063);
and U12103 (N_12103,N_8631,N_7735);
and U12104 (N_12104,N_5892,N_6096);
nor U12105 (N_12105,N_7824,N_5762);
nand U12106 (N_12106,N_9972,N_9982);
and U12107 (N_12107,N_6467,N_8343);
or U12108 (N_12108,N_7098,N_7725);
and U12109 (N_12109,N_7942,N_8015);
or U12110 (N_12110,N_7348,N_6428);
or U12111 (N_12111,N_8048,N_6127);
xnor U12112 (N_12112,N_6122,N_5875);
nand U12113 (N_12113,N_9249,N_8262);
or U12114 (N_12114,N_8273,N_7394);
or U12115 (N_12115,N_6073,N_8524);
nor U12116 (N_12116,N_8446,N_5264);
or U12117 (N_12117,N_6415,N_9611);
nand U12118 (N_12118,N_8001,N_5225);
nor U12119 (N_12119,N_5481,N_8887);
and U12120 (N_12120,N_9070,N_8345);
and U12121 (N_12121,N_5058,N_6667);
nand U12122 (N_12122,N_8397,N_9655);
nand U12123 (N_12123,N_6487,N_5383);
nand U12124 (N_12124,N_8418,N_5321);
and U12125 (N_12125,N_8922,N_7229);
nor U12126 (N_12126,N_5602,N_8323);
nor U12127 (N_12127,N_8959,N_7226);
nor U12128 (N_12128,N_5348,N_8072);
and U12129 (N_12129,N_8453,N_7651);
and U12130 (N_12130,N_9210,N_9454);
nand U12131 (N_12131,N_8174,N_6074);
or U12132 (N_12132,N_9852,N_8510);
nor U12133 (N_12133,N_8263,N_6219);
and U12134 (N_12134,N_9293,N_9669);
and U12135 (N_12135,N_8690,N_6089);
nor U12136 (N_12136,N_8980,N_5500);
nor U12137 (N_12137,N_6239,N_5953);
nor U12138 (N_12138,N_5136,N_7104);
or U12139 (N_12139,N_9423,N_9916);
nand U12140 (N_12140,N_6279,N_7545);
or U12141 (N_12141,N_6877,N_6696);
nand U12142 (N_12142,N_9399,N_6166);
and U12143 (N_12143,N_7386,N_5964);
nor U12144 (N_12144,N_7777,N_6181);
nor U12145 (N_12145,N_6414,N_9634);
or U12146 (N_12146,N_8313,N_9735);
nand U12147 (N_12147,N_5865,N_6091);
nor U12148 (N_12148,N_8728,N_5679);
nor U12149 (N_12149,N_8057,N_7959);
nand U12150 (N_12150,N_7323,N_8562);
and U12151 (N_12151,N_7555,N_8546);
nand U12152 (N_12152,N_6675,N_8760);
nand U12153 (N_12153,N_5737,N_8337);
nand U12154 (N_12154,N_6468,N_8585);
or U12155 (N_12155,N_7706,N_6174);
nand U12156 (N_12156,N_8867,N_8297);
and U12157 (N_12157,N_9296,N_7205);
or U12158 (N_12158,N_5211,N_7332);
nor U12159 (N_12159,N_5837,N_6530);
or U12160 (N_12160,N_6113,N_8969);
nor U12161 (N_12161,N_9844,N_8331);
or U12162 (N_12162,N_6397,N_7761);
or U12163 (N_12163,N_8268,N_8756);
and U12164 (N_12164,N_7069,N_9651);
nand U12165 (N_12165,N_6616,N_6763);
xnor U12166 (N_12166,N_9100,N_6565);
nand U12167 (N_12167,N_9462,N_8120);
nand U12168 (N_12168,N_9921,N_8172);
nand U12169 (N_12169,N_5397,N_8136);
and U12170 (N_12170,N_5470,N_5224);
nor U12171 (N_12171,N_8521,N_9076);
or U12172 (N_12172,N_5190,N_7729);
nand U12173 (N_12173,N_7391,N_6827);
nand U12174 (N_12174,N_8888,N_5487);
nand U12175 (N_12175,N_7836,N_5212);
nor U12176 (N_12176,N_6747,N_9929);
nor U12177 (N_12177,N_5783,N_7215);
nor U12178 (N_12178,N_9582,N_5954);
nor U12179 (N_12179,N_5442,N_6440);
nand U12180 (N_12180,N_9886,N_5241);
nor U12181 (N_12181,N_7681,N_8654);
and U12182 (N_12182,N_7153,N_9205);
nand U12183 (N_12183,N_5658,N_5416);
or U12184 (N_12184,N_7511,N_5664);
nand U12185 (N_12185,N_6595,N_9529);
or U12186 (N_12186,N_6694,N_5233);
nand U12187 (N_12187,N_7925,N_9261);
nor U12188 (N_12188,N_6608,N_9218);
nor U12189 (N_12189,N_7253,N_7532);
and U12190 (N_12190,N_5999,N_6594);
or U12191 (N_12191,N_8529,N_7504);
and U12192 (N_12192,N_5772,N_9213);
and U12193 (N_12193,N_5846,N_6252);
nor U12194 (N_12194,N_9556,N_9016);
nand U12195 (N_12195,N_6850,N_7033);
nor U12196 (N_12196,N_7214,N_9661);
nand U12197 (N_12197,N_7852,N_7147);
xor U12198 (N_12198,N_5711,N_9192);
nand U12199 (N_12199,N_5104,N_8748);
and U12200 (N_12200,N_6026,N_8183);
and U12201 (N_12201,N_5818,N_9387);
nand U12202 (N_12202,N_6879,N_5771);
nor U12203 (N_12203,N_5438,N_5532);
nor U12204 (N_12204,N_5605,N_7983);
and U12205 (N_12205,N_6776,N_5194);
nor U12206 (N_12206,N_9993,N_5157);
nor U12207 (N_12207,N_7123,N_7413);
nand U12208 (N_12208,N_8101,N_6636);
or U12209 (N_12209,N_6830,N_7059);
nand U12210 (N_12210,N_8277,N_6545);
nand U12211 (N_12211,N_9776,N_8193);
or U12212 (N_12212,N_7742,N_5988);
nor U12213 (N_12213,N_9485,N_7667);
and U12214 (N_12214,N_7079,N_5623);
or U12215 (N_12215,N_8283,N_7289);
nor U12216 (N_12216,N_9106,N_5415);
or U12217 (N_12217,N_5726,N_9281);
and U12218 (N_12218,N_6302,N_9260);
or U12219 (N_12219,N_7000,N_5289);
nand U12220 (N_12220,N_8996,N_9339);
nor U12221 (N_12221,N_6575,N_9362);
nor U12222 (N_12222,N_8176,N_6374);
nand U12223 (N_12223,N_5231,N_5366);
or U12224 (N_12224,N_6544,N_9095);
and U12225 (N_12225,N_9807,N_8225);
and U12226 (N_12226,N_5689,N_7887);
nor U12227 (N_12227,N_8561,N_8339);
and U12228 (N_12228,N_5618,N_8096);
and U12229 (N_12229,N_8473,N_8832);
and U12230 (N_12230,N_8544,N_5243);
and U12231 (N_12231,N_9156,N_9230);
nor U12232 (N_12232,N_6652,N_9027);
nand U12233 (N_12233,N_6379,N_9108);
nand U12234 (N_12234,N_5859,N_6059);
and U12235 (N_12235,N_5899,N_8164);
and U12236 (N_12236,N_9761,N_6874);
xor U12237 (N_12237,N_6692,N_9302);
or U12238 (N_12238,N_7158,N_5927);
and U12239 (N_12239,N_9552,N_6765);
and U12240 (N_12240,N_9383,N_9830);
or U12241 (N_12241,N_8909,N_8525);
nand U12242 (N_12242,N_9825,N_6552);
nor U12243 (N_12243,N_6598,N_9337);
nand U12244 (N_12244,N_9706,N_7813);
nor U12245 (N_12245,N_8392,N_5860);
xor U12246 (N_12246,N_7276,N_7488);
and U12247 (N_12247,N_7431,N_9714);
and U12248 (N_12248,N_8095,N_7817);
nand U12249 (N_12249,N_7986,N_5592);
and U12250 (N_12250,N_7613,N_5997);
nand U12251 (N_12251,N_9466,N_7508);
nor U12252 (N_12252,N_7114,N_5062);
nand U12253 (N_12253,N_5606,N_6483);
or U12254 (N_12254,N_5700,N_5661);
or U12255 (N_12255,N_6973,N_9173);
nand U12256 (N_12256,N_7895,N_8220);
and U12257 (N_12257,N_8469,N_7980);
nor U12258 (N_12258,N_8163,N_8304);
nand U12259 (N_12259,N_7731,N_5752);
or U12260 (N_12260,N_8941,N_5386);
nand U12261 (N_12261,N_6381,N_6058);
and U12262 (N_12262,N_9539,N_6682);
nor U12263 (N_12263,N_5901,N_8881);
or U12264 (N_12264,N_7528,N_5941);
nand U12265 (N_12265,N_5610,N_7631);
or U12266 (N_12266,N_8774,N_7218);
or U12267 (N_12267,N_6055,N_9745);
or U12268 (N_12268,N_6914,N_8207);
or U12269 (N_12269,N_6754,N_6889);
and U12270 (N_12270,N_6569,N_8661);
and U12271 (N_12271,N_9622,N_9093);
and U12272 (N_12272,N_5073,N_9452);
nor U12273 (N_12273,N_8715,N_7228);
or U12274 (N_12274,N_9889,N_7385);
and U12275 (N_12275,N_8265,N_5769);
nand U12276 (N_12276,N_5942,N_7720);
or U12277 (N_12277,N_5858,N_5956);
and U12278 (N_12278,N_9559,N_9137);
and U12279 (N_12279,N_6354,N_7515);
nand U12280 (N_12280,N_8398,N_5148);
nand U12281 (N_12281,N_5038,N_5639);
or U12282 (N_12282,N_6478,N_9440);
or U12283 (N_12283,N_6344,N_7326);
nor U12284 (N_12284,N_8031,N_8173);
nor U12285 (N_12285,N_9827,N_8624);
nor U12286 (N_12286,N_6757,N_6864);
nand U12287 (N_12287,N_7045,N_9500);
and U12288 (N_12288,N_6814,N_9022);
and U12289 (N_12289,N_5735,N_5176);
and U12290 (N_12290,N_7313,N_5946);
and U12291 (N_12291,N_9907,N_9926);
and U12292 (N_12292,N_6899,N_6207);
nand U12293 (N_12293,N_7864,N_7437);
nand U12294 (N_12294,N_7603,N_7931);
nor U12295 (N_12295,N_5302,N_5690);
or U12296 (N_12296,N_7768,N_7051);
nand U12297 (N_12297,N_5004,N_9631);
and U12298 (N_12298,N_6945,N_5042);
nand U12299 (N_12299,N_7392,N_7427);
nor U12300 (N_12300,N_5060,N_6859);
nor U12301 (N_12301,N_8281,N_6751);
or U12302 (N_12302,N_5754,N_6117);
and U12303 (N_12303,N_7290,N_6137);
and U12304 (N_12304,N_9725,N_9918);
nor U12305 (N_12305,N_6759,N_9560);
nand U12306 (N_12306,N_7750,N_7624);
and U12307 (N_12307,N_5564,N_7525);
nand U12308 (N_12308,N_6677,N_6767);
nand U12309 (N_12309,N_8157,N_8402);
nor U12310 (N_12310,N_6206,N_9418);
and U12311 (N_12311,N_5433,N_7490);
nor U12312 (N_12312,N_6472,N_8963);
or U12313 (N_12313,N_6533,N_7773);
or U12314 (N_12314,N_8386,N_5326);
and U12315 (N_12315,N_5089,N_8782);
nor U12316 (N_12316,N_6553,N_5144);
or U12317 (N_12317,N_8806,N_6454);
or U12318 (N_12318,N_6587,N_9397);
or U12319 (N_12319,N_5361,N_7604);
or U12320 (N_12320,N_9802,N_6651);
and U12321 (N_12321,N_6008,N_9703);
or U12322 (N_12322,N_7278,N_9441);
nand U12323 (N_12323,N_6032,N_7061);
nor U12324 (N_12324,N_9792,N_9512);
and U12325 (N_12325,N_8366,N_8817);
nand U12326 (N_12326,N_8725,N_7605);
nand U12327 (N_12327,N_7358,N_9434);
nand U12328 (N_12328,N_6781,N_5629);
nor U12329 (N_12329,N_8812,N_9123);
nor U12330 (N_12330,N_6231,N_5110);
nand U12331 (N_12331,N_9677,N_8754);
or U12332 (N_12332,N_5965,N_8526);
or U12333 (N_12333,N_8114,N_8051);
nor U12334 (N_12334,N_9242,N_6450);
nand U12335 (N_12335,N_5620,N_7659);
nor U12336 (N_12336,N_5467,N_6962);
nor U12337 (N_12337,N_7920,N_6630);
and U12338 (N_12338,N_9887,N_7897);
nand U12339 (N_12339,N_7075,N_6802);
or U12340 (N_12340,N_8158,N_6382);
and U12341 (N_12341,N_8303,N_5636);
or U12342 (N_12342,N_5277,N_8552);
nand U12343 (N_12343,N_9645,N_7255);
nand U12344 (N_12344,N_5738,N_9919);
nor U12345 (N_12345,N_9524,N_5510);
or U12346 (N_12346,N_7080,N_6402);
nor U12347 (N_12347,N_9234,N_9906);
and U12348 (N_12348,N_8006,N_7704);
or U12349 (N_12349,N_7458,N_7371);
and U12350 (N_12350,N_6793,N_9649);
nand U12351 (N_12351,N_9970,N_7671);
nor U12352 (N_12352,N_9633,N_9329);
nor U12353 (N_12353,N_6571,N_8391);
and U12354 (N_12354,N_9396,N_8460);
and U12355 (N_12355,N_6346,N_9153);
nor U12356 (N_12356,N_7950,N_7672);
and U12357 (N_12357,N_5270,N_5310);
and U12358 (N_12358,N_9049,N_7109);
and U12359 (N_12359,N_6343,N_5373);
and U12360 (N_12360,N_7839,N_6883);
and U12361 (N_12361,N_8589,N_8716);
nor U12362 (N_12362,N_7943,N_5090);
or U12363 (N_12363,N_7800,N_8747);
nor U12364 (N_12364,N_5088,N_6083);
or U12365 (N_12365,N_8479,N_8973);
or U12366 (N_12366,N_7608,N_7893);
and U12367 (N_12367,N_6917,N_7594);
nor U12368 (N_12368,N_8721,N_7933);
and U12369 (N_12369,N_5352,N_6890);
or U12370 (N_12370,N_8274,N_7968);
nor U12371 (N_12371,N_6784,N_7160);
nand U12372 (N_12372,N_9509,N_6396);
nor U12373 (N_12373,N_6260,N_6132);
xnor U12374 (N_12374,N_8858,N_6661);
nand U12375 (N_12375,N_9460,N_9495);
and U12376 (N_12376,N_8837,N_5485);
nor U12377 (N_12377,N_6531,N_7180);
nand U12378 (N_12378,N_7099,N_9146);
and U12379 (N_12379,N_5252,N_9463);
and U12380 (N_12380,N_7273,N_7012);
nand U12381 (N_12381,N_7211,N_9074);
nand U12382 (N_12382,N_5134,N_7439);
and U12383 (N_12383,N_5378,N_8890);
nand U12384 (N_12384,N_6455,N_7457);
nor U12385 (N_12385,N_8064,N_6712);
nor U12386 (N_12386,N_9186,N_9190);
or U12387 (N_12387,N_6835,N_5170);
nor U12388 (N_12388,N_8652,N_9096);
and U12389 (N_12389,N_6730,N_9488);
nor U12390 (N_12390,N_5626,N_6965);
nor U12391 (N_12391,N_9862,N_8488);
nand U12392 (N_12392,N_6186,N_7649);
and U12393 (N_12393,N_6593,N_5445);
nor U12394 (N_12394,N_6993,N_5548);
or U12395 (N_12395,N_8428,N_6092);
and U12396 (N_12396,N_7096,N_6267);
nand U12397 (N_12397,N_6709,N_8334);
and U12398 (N_12398,N_9084,N_6515);
and U12399 (N_12399,N_5893,N_5823);
nand U12400 (N_12400,N_8674,N_6559);
nand U12401 (N_12401,N_5480,N_7763);
and U12402 (N_12402,N_6010,N_6400);
nand U12403 (N_12403,N_8368,N_7848);
nand U12404 (N_12404,N_7144,N_5540);
or U12405 (N_12405,N_8415,N_6222);
nor U12406 (N_12406,N_6128,N_8672);
nor U12407 (N_12407,N_7130,N_5553);
and U12408 (N_12408,N_5387,N_8954);
nor U12409 (N_12409,N_9535,N_5341);
nand U12410 (N_12410,N_5247,N_9361);
nand U12411 (N_12411,N_5125,N_5544);
nand U12412 (N_12412,N_9464,N_6159);
nand U12413 (N_12413,N_6625,N_5479);
or U12414 (N_12414,N_6527,N_7916);
nor U12415 (N_12415,N_7049,N_7189);
or U12416 (N_12416,N_6855,N_8477);
nor U12417 (N_12417,N_8410,N_9841);
nand U12418 (N_12418,N_8801,N_6576);
nand U12419 (N_12419,N_7865,N_5379);
and U12420 (N_12420,N_5369,N_5950);
nor U12421 (N_12421,N_9913,N_5124);
nand U12422 (N_12422,N_7756,N_8258);
and U12423 (N_12423,N_8576,N_7678);
and U12424 (N_12424,N_9849,N_6756);
xor U12425 (N_12425,N_6124,N_8567);
and U12426 (N_12426,N_5530,N_6149);
and U12427 (N_12427,N_9584,N_9058);
or U12428 (N_12428,N_5154,N_9550);
or U12429 (N_12429,N_7084,N_6187);
and U12430 (N_12430,N_6619,N_7551);
nand U12431 (N_12431,N_6681,N_6486);
and U12432 (N_12432,N_5757,N_9527);
nor U12433 (N_12433,N_8555,N_9967);
and U12434 (N_12434,N_5258,N_8911);
or U12435 (N_12435,N_8668,N_9376);
nor U12436 (N_12436,N_7654,N_6660);
and U12437 (N_12437,N_9271,N_5933);
and U12438 (N_12438,N_8707,N_5210);
and U12439 (N_12439,N_8461,N_6325);
nor U12440 (N_12440,N_8396,N_6977);
nor U12441 (N_12441,N_6923,N_5047);
nor U12442 (N_12442,N_5203,N_6064);
nor U12443 (N_12443,N_8275,N_8129);
xnor U12444 (N_12444,N_6422,N_8889);
nand U12445 (N_12445,N_5118,N_6100);
or U12446 (N_12446,N_7593,N_7911);
and U12447 (N_12447,N_8547,N_7559);
and U12448 (N_12448,N_8726,N_6632);
nor U12449 (N_12449,N_8842,N_8847);
and U12450 (N_12450,N_6964,N_8653);
nand U12451 (N_12451,N_8543,N_6268);
and U12452 (N_12452,N_5496,N_5158);
and U12453 (N_12453,N_5926,N_9305);
and U12454 (N_12454,N_7254,N_9781);
nand U12455 (N_12455,N_9975,N_7789);
nor U12456 (N_12456,N_6631,N_6009);
or U12457 (N_12457,N_5453,N_6983);
and U12458 (N_12458,N_9526,N_8638);
nand U12459 (N_12459,N_6286,N_6250);
nand U12460 (N_12460,N_6644,N_6789);
or U12461 (N_12461,N_7535,N_6364);
nor U12462 (N_12462,N_9896,N_8424);
and U12463 (N_12463,N_6555,N_8189);
xor U12464 (N_12464,N_9481,N_9063);
nor U12465 (N_12465,N_6471,N_7036);
nor U12466 (N_12466,N_5172,N_9360);
nand U12467 (N_12467,N_6522,N_5993);
or U12468 (N_12468,N_7261,N_5414);
and U12469 (N_12469,N_8581,N_6618);
nor U12470 (N_12470,N_7726,N_9502);
or U12471 (N_12471,N_8013,N_6721);
xor U12472 (N_12472,N_9865,N_7464);
nor U12473 (N_12473,N_8340,N_5367);
or U12474 (N_12474,N_9783,N_6013);
nor U12475 (N_12475,N_5338,N_5254);
or U12476 (N_12476,N_9268,N_9676);
or U12477 (N_12477,N_7478,N_5815);
nand U12478 (N_12478,N_9308,N_8951);
nand U12479 (N_12479,N_6748,N_7173);
nor U12480 (N_12480,N_9367,N_9870);
nor U12481 (N_12481,N_6574,N_7732);
nor U12482 (N_12482,N_8246,N_9602);
nor U12483 (N_12483,N_5219,N_7692);
nand U12484 (N_12484,N_8919,N_7643);
nand U12485 (N_12485,N_9653,N_5558);
and U12486 (N_12486,N_8517,N_7141);
nand U12487 (N_12487,N_8377,N_8667);
nor U12488 (N_12488,N_5161,N_7380);
and U12489 (N_12489,N_6033,N_6218);
nor U12490 (N_12490,N_9861,N_9236);
nand U12491 (N_12491,N_5458,N_5891);
or U12492 (N_12492,N_6963,N_8788);
and U12493 (N_12493,N_8350,N_7103);
nor U12494 (N_12494,N_9199,N_7395);
and U12495 (N_12495,N_9443,N_5447);
or U12496 (N_12496,N_5574,N_7003);
nand U12497 (N_12497,N_9335,N_9976);
and U12498 (N_12498,N_9680,N_5563);
nor U12499 (N_12499,N_9746,N_8090);
and U12500 (N_12500,N_9837,N_6823);
nand U12501 (N_12501,N_7153,N_5335);
nor U12502 (N_12502,N_6922,N_7356);
or U12503 (N_12503,N_7302,N_9673);
nand U12504 (N_12504,N_9196,N_7101);
and U12505 (N_12505,N_7400,N_7036);
and U12506 (N_12506,N_5639,N_7286);
or U12507 (N_12507,N_5225,N_6369);
or U12508 (N_12508,N_7971,N_8546);
and U12509 (N_12509,N_9468,N_7089);
nor U12510 (N_12510,N_5306,N_9957);
nor U12511 (N_12511,N_6692,N_8258);
nor U12512 (N_12512,N_7436,N_7428);
nand U12513 (N_12513,N_7666,N_7793);
or U12514 (N_12514,N_8048,N_9454);
nor U12515 (N_12515,N_6866,N_5931);
nor U12516 (N_12516,N_5564,N_9399);
nand U12517 (N_12517,N_9998,N_8806);
nor U12518 (N_12518,N_5122,N_6280);
and U12519 (N_12519,N_7993,N_9548);
nor U12520 (N_12520,N_7731,N_7584);
nor U12521 (N_12521,N_5587,N_6482);
and U12522 (N_12522,N_9527,N_9690);
and U12523 (N_12523,N_6445,N_6514);
nand U12524 (N_12524,N_8831,N_5918);
and U12525 (N_12525,N_9556,N_6275);
or U12526 (N_12526,N_9903,N_5496);
nor U12527 (N_12527,N_8934,N_5547);
and U12528 (N_12528,N_6476,N_5078);
and U12529 (N_12529,N_9605,N_7822);
nand U12530 (N_12530,N_5936,N_8720);
nand U12531 (N_12531,N_6770,N_7266);
and U12532 (N_12532,N_9339,N_5724);
nor U12533 (N_12533,N_5143,N_6694);
nand U12534 (N_12534,N_9232,N_5655);
or U12535 (N_12535,N_7537,N_9561);
or U12536 (N_12536,N_9775,N_7731);
nand U12537 (N_12537,N_7495,N_7789);
or U12538 (N_12538,N_6507,N_8217);
and U12539 (N_12539,N_9336,N_6333);
and U12540 (N_12540,N_7830,N_6063);
or U12541 (N_12541,N_7802,N_8454);
nand U12542 (N_12542,N_5798,N_9679);
nor U12543 (N_12543,N_5127,N_8621);
or U12544 (N_12544,N_9256,N_8035);
or U12545 (N_12545,N_9951,N_7304);
nand U12546 (N_12546,N_7323,N_9079);
and U12547 (N_12547,N_6910,N_8441);
nand U12548 (N_12548,N_8291,N_5570);
nand U12549 (N_12549,N_6981,N_7440);
nand U12550 (N_12550,N_9397,N_7596);
nand U12551 (N_12551,N_8988,N_9347);
nor U12552 (N_12552,N_5142,N_9685);
or U12553 (N_12553,N_9157,N_7590);
and U12554 (N_12554,N_8983,N_6696);
or U12555 (N_12555,N_7145,N_8715);
nor U12556 (N_12556,N_5235,N_9251);
nand U12557 (N_12557,N_6381,N_6581);
xnor U12558 (N_12558,N_7222,N_8272);
or U12559 (N_12559,N_7338,N_8241);
and U12560 (N_12560,N_5269,N_9066);
and U12561 (N_12561,N_9322,N_8181);
and U12562 (N_12562,N_6711,N_8544);
or U12563 (N_12563,N_8606,N_9576);
nor U12564 (N_12564,N_9901,N_5656);
nand U12565 (N_12565,N_5722,N_8300);
and U12566 (N_12566,N_6375,N_6487);
and U12567 (N_12567,N_8411,N_7304);
nand U12568 (N_12568,N_9276,N_8712);
nor U12569 (N_12569,N_5079,N_8261);
nor U12570 (N_12570,N_9918,N_8151);
nor U12571 (N_12571,N_9705,N_9116);
nor U12572 (N_12572,N_5440,N_7896);
nand U12573 (N_12573,N_5889,N_5471);
or U12574 (N_12574,N_6149,N_8750);
nand U12575 (N_12575,N_6767,N_8445);
or U12576 (N_12576,N_5323,N_7030);
nand U12577 (N_12577,N_7347,N_5906);
nand U12578 (N_12578,N_6591,N_6502);
nand U12579 (N_12579,N_8421,N_9609);
nand U12580 (N_12580,N_8462,N_9553);
or U12581 (N_12581,N_6947,N_7877);
and U12582 (N_12582,N_7779,N_8556);
nor U12583 (N_12583,N_6822,N_9417);
or U12584 (N_12584,N_9042,N_7068);
nor U12585 (N_12585,N_5752,N_9732);
nand U12586 (N_12586,N_5923,N_7610);
or U12587 (N_12587,N_8063,N_5080);
or U12588 (N_12588,N_9011,N_6560);
nand U12589 (N_12589,N_8947,N_6797);
and U12590 (N_12590,N_9225,N_6810);
and U12591 (N_12591,N_7600,N_9670);
or U12592 (N_12592,N_7570,N_6704);
or U12593 (N_12593,N_9192,N_5249);
xor U12594 (N_12594,N_5611,N_6040);
and U12595 (N_12595,N_9815,N_7353);
and U12596 (N_12596,N_9431,N_5633);
or U12597 (N_12597,N_5832,N_5862);
and U12598 (N_12598,N_5712,N_9913);
nand U12599 (N_12599,N_8451,N_9818);
nand U12600 (N_12600,N_6573,N_5918);
nand U12601 (N_12601,N_8373,N_6811);
and U12602 (N_12602,N_9302,N_6161);
nor U12603 (N_12603,N_8514,N_6637);
nor U12604 (N_12604,N_8413,N_7490);
nor U12605 (N_12605,N_7083,N_9104);
nor U12606 (N_12606,N_9565,N_9861);
nor U12607 (N_12607,N_9809,N_8391);
and U12608 (N_12608,N_5117,N_5912);
and U12609 (N_12609,N_5435,N_6613);
and U12610 (N_12610,N_8975,N_8268);
nor U12611 (N_12611,N_9982,N_5443);
nor U12612 (N_12612,N_7925,N_7984);
and U12613 (N_12613,N_8870,N_5659);
and U12614 (N_12614,N_7695,N_9950);
or U12615 (N_12615,N_8856,N_9527);
nand U12616 (N_12616,N_7066,N_9566);
nor U12617 (N_12617,N_5340,N_7391);
or U12618 (N_12618,N_8423,N_9738);
or U12619 (N_12619,N_5626,N_8233);
nand U12620 (N_12620,N_5429,N_8237);
and U12621 (N_12621,N_6593,N_9446);
or U12622 (N_12622,N_6141,N_6667);
and U12623 (N_12623,N_6313,N_9472);
nor U12624 (N_12624,N_9504,N_6662);
xor U12625 (N_12625,N_9560,N_6510);
or U12626 (N_12626,N_6601,N_9570);
and U12627 (N_12627,N_8666,N_9882);
nor U12628 (N_12628,N_8069,N_5088);
and U12629 (N_12629,N_5628,N_7927);
nand U12630 (N_12630,N_7147,N_5007);
nand U12631 (N_12631,N_6679,N_9789);
nand U12632 (N_12632,N_5454,N_6671);
and U12633 (N_12633,N_7177,N_5115);
and U12634 (N_12634,N_8430,N_5397);
nand U12635 (N_12635,N_5287,N_7662);
or U12636 (N_12636,N_7220,N_8562);
and U12637 (N_12637,N_8286,N_7376);
and U12638 (N_12638,N_9616,N_6465);
xor U12639 (N_12639,N_5777,N_7793);
nand U12640 (N_12640,N_8981,N_6752);
nand U12641 (N_12641,N_6403,N_7255);
nor U12642 (N_12642,N_8111,N_6226);
nor U12643 (N_12643,N_7722,N_5011);
and U12644 (N_12644,N_8981,N_6139);
and U12645 (N_12645,N_8586,N_8259);
nand U12646 (N_12646,N_5922,N_6455);
and U12647 (N_12647,N_8241,N_6535);
and U12648 (N_12648,N_7516,N_8404);
nand U12649 (N_12649,N_9002,N_6115);
nand U12650 (N_12650,N_6825,N_8989);
and U12651 (N_12651,N_8287,N_9171);
nor U12652 (N_12652,N_9084,N_6767);
nor U12653 (N_12653,N_8660,N_6147);
nor U12654 (N_12654,N_7112,N_6836);
or U12655 (N_12655,N_5378,N_7807);
or U12656 (N_12656,N_5305,N_7586);
and U12657 (N_12657,N_6112,N_7215);
nor U12658 (N_12658,N_9135,N_5202);
nor U12659 (N_12659,N_6245,N_6197);
or U12660 (N_12660,N_7983,N_6149);
nor U12661 (N_12661,N_6321,N_5512);
nand U12662 (N_12662,N_8974,N_9565);
or U12663 (N_12663,N_7609,N_7381);
and U12664 (N_12664,N_7160,N_5962);
nand U12665 (N_12665,N_9535,N_8046);
nand U12666 (N_12666,N_5952,N_6024);
nand U12667 (N_12667,N_8924,N_5878);
or U12668 (N_12668,N_7829,N_7218);
and U12669 (N_12669,N_5361,N_6810);
or U12670 (N_12670,N_7300,N_5596);
or U12671 (N_12671,N_5494,N_7083);
or U12672 (N_12672,N_5671,N_7453);
or U12673 (N_12673,N_5426,N_8540);
and U12674 (N_12674,N_7425,N_9664);
nand U12675 (N_12675,N_5494,N_7823);
nor U12676 (N_12676,N_5112,N_8967);
and U12677 (N_12677,N_9830,N_7322);
and U12678 (N_12678,N_7028,N_6729);
and U12679 (N_12679,N_7643,N_7895);
nor U12680 (N_12680,N_7928,N_6562);
nor U12681 (N_12681,N_8093,N_9381);
or U12682 (N_12682,N_7666,N_6548);
and U12683 (N_12683,N_8702,N_8728);
and U12684 (N_12684,N_9368,N_9662);
and U12685 (N_12685,N_7799,N_9391);
nor U12686 (N_12686,N_8484,N_5142);
or U12687 (N_12687,N_9393,N_9508);
nand U12688 (N_12688,N_6864,N_7562);
nor U12689 (N_12689,N_5744,N_6264);
nand U12690 (N_12690,N_9642,N_8938);
nand U12691 (N_12691,N_7921,N_7655);
or U12692 (N_12692,N_9676,N_6934);
nor U12693 (N_12693,N_7657,N_7577);
and U12694 (N_12694,N_6412,N_9023);
nor U12695 (N_12695,N_6504,N_8317);
and U12696 (N_12696,N_9824,N_5672);
or U12697 (N_12697,N_8819,N_9123);
and U12698 (N_12698,N_5491,N_5583);
nor U12699 (N_12699,N_6977,N_8731);
nand U12700 (N_12700,N_5516,N_8966);
nand U12701 (N_12701,N_9170,N_7019);
or U12702 (N_12702,N_6191,N_8870);
xor U12703 (N_12703,N_6521,N_5179);
nor U12704 (N_12704,N_9155,N_7304);
or U12705 (N_12705,N_8808,N_8039);
nor U12706 (N_12706,N_9113,N_7128);
nand U12707 (N_12707,N_5914,N_9918);
and U12708 (N_12708,N_8434,N_8914);
nand U12709 (N_12709,N_5275,N_5489);
or U12710 (N_12710,N_7591,N_6463);
or U12711 (N_12711,N_7749,N_9485);
nor U12712 (N_12712,N_6473,N_6120);
nor U12713 (N_12713,N_5183,N_7960);
and U12714 (N_12714,N_8311,N_9499);
and U12715 (N_12715,N_8616,N_7107);
and U12716 (N_12716,N_9548,N_6080);
nor U12717 (N_12717,N_6087,N_7157);
nand U12718 (N_12718,N_5605,N_9819);
and U12719 (N_12719,N_5490,N_7191);
nor U12720 (N_12720,N_5088,N_6589);
and U12721 (N_12721,N_7143,N_8922);
nor U12722 (N_12722,N_6521,N_9119);
or U12723 (N_12723,N_7765,N_5389);
or U12724 (N_12724,N_6666,N_6964);
and U12725 (N_12725,N_7022,N_7584);
and U12726 (N_12726,N_8889,N_7025);
nor U12727 (N_12727,N_7792,N_7279);
and U12728 (N_12728,N_9556,N_6612);
or U12729 (N_12729,N_6202,N_8119);
nand U12730 (N_12730,N_8867,N_7892);
nand U12731 (N_12731,N_8434,N_8174);
or U12732 (N_12732,N_7486,N_6480);
and U12733 (N_12733,N_8426,N_9608);
nand U12734 (N_12734,N_9531,N_6219);
nand U12735 (N_12735,N_7286,N_9485);
nor U12736 (N_12736,N_8061,N_9689);
nand U12737 (N_12737,N_7103,N_6809);
or U12738 (N_12738,N_5242,N_7667);
nand U12739 (N_12739,N_6890,N_9344);
or U12740 (N_12740,N_7610,N_8874);
nor U12741 (N_12741,N_9117,N_6141);
nand U12742 (N_12742,N_7224,N_7212);
nor U12743 (N_12743,N_6042,N_5829);
nor U12744 (N_12744,N_8490,N_9539);
xnor U12745 (N_12745,N_7215,N_9208);
nand U12746 (N_12746,N_7119,N_7130);
nor U12747 (N_12747,N_9661,N_9948);
or U12748 (N_12748,N_9735,N_5745);
xnor U12749 (N_12749,N_9280,N_7578);
or U12750 (N_12750,N_7713,N_8995);
nor U12751 (N_12751,N_9920,N_9403);
nand U12752 (N_12752,N_7250,N_8634);
nand U12753 (N_12753,N_9852,N_5418);
nor U12754 (N_12754,N_5361,N_7147);
or U12755 (N_12755,N_9460,N_5822);
or U12756 (N_12756,N_5843,N_8166);
nor U12757 (N_12757,N_7280,N_7338);
nor U12758 (N_12758,N_9790,N_6718);
nand U12759 (N_12759,N_8099,N_9358);
and U12760 (N_12760,N_7868,N_5074);
nor U12761 (N_12761,N_5186,N_9964);
or U12762 (N_12762,N_7974,N_6024);
nor U12763 (N_12763,N_7159,N_8788);
and U12764 (N_12764,N_9211,N_7746);
nand U12765 (N_12765,N_6722,N_7464);
and U12766 (N_12766,N_9645,N_6444);
and U12767 (N_12767,N_5866,N_8170);
or U12768 (N_12768,N_5429,N_5403);
or U12769 (N_12769,N_5299,N_9588);
xnor U12770 (N_12770,N_8163,N_5735);
nand U12771 (N_12771,N_7840,N_5806);
nor U12772 (N_12772,N_8150,N_5602);
nand U12773 (N_12773,N_8928,N_5441);
nor U12774 (N_12774,N_9639,N_8160);
or U12775 (N_12775,N_8977,N_9997);
nor U12776 (N_12776,N_7919,N_5985);
or U12777 (N_12777,N_8226,N_7721);
or U12778 (N_12778,N_7507,N_5872);
and U12779 (N_12779,N_6117,N_8407);
nor U12780 (N_12780,N_5703,N_5117);
nand U12781 (N_12781,N_8794,N_8739);
nand U12782 (N_12782,N_5176,N_9704);
nand U12783 (N_12783,N_8555,N_9258);
nor U12784 (N_12784,N_7555,N_8722);
or U12785 (N_12785,N_7717,N_7788);
and U12786 (N_12786,N_6412,N_7720);
or U12787 (N_12787,N_7252,N_7438);
xnor U12788 (N_12788,N_7278,N_5650);
or U12789 (N_12789,N_8956,N_5976);
and U12790 (N_12790,N_7657,N_5844);
or U12791 (N_12791,N_8538,N_5478);
and U12792 (N_12792,N_7838,N_5354);
nor U12793 (N_12793,N_5564,N_8634);
and U12794 (N_12794,N_6022,N_8787);
and U12795 (N_12795,N_8935,N_5880);
or U12796 (N_12796,N_7946,N_5373);
nand U12797 (N_12797,N_8411,N_5658);
or U12798 (N_12798,N_7516,N_8221);
and U12799 (N_12799,N_5872,N_6211);
nor U12800 (N_12800,N_8528,N_7501);
nand U12801 (N_12801,N_6985,N_7245);
nand U12802 (N_12802,N_6985,N_9214);
nand U12803 (N_12803,N_5329,N_6016);
xor U12804 (N_12804,N_8248,N_8019);
or U12805 (N_12805,N_7047,N_6407);
and U12806 (N_12806,N_7309,N_9890);
nor U12807 (N_12807,N_5644,N_6838);
nor U12808 (N_12808,N_9491,N_5381);
nand U12809 (N_12809,N_8195,N_5490);
nor U12810 (N_12810,N_9351,N_7387);
nand U12811 (N_12811,N_5499,N_6943);
nand U12812 (N_12812,N_6582,N_6105);
or U12813 (N_12813,N_8932,N_7806);
or U12814 (N_12814,N_7617,N_9215);
nor U12815 (N_12815,N_5659,N_7026);
or U12816 (N_12816,N_5496,N_7785);
xnor U12817 (N_12817,N_7218,N_7211);
or U12818 (N_12818,N_5727,N_8048);
and U12819 (N_12819,N_9509,N_8048);
and U12820 (N_12820,N_7938,N_6816);
and U12821 (N_12821,N_9100,N_6154);
nor U12822 (N_12822,N_8538,N_7904);
nand U12823 (N_12823,N_8292,N_9967);
nor U12824 (N_12824,N_9916,N_7892);
nor U12825 (N_12825,N_7309,N_5382);
nand U12826 (N_12826,N_8364,N_7075);
nor U12827 (N_12827,N_5866,N_8015);
or U12828 (N_12828,N_5666,N_6967);
nand U12829 (N_12829,N_8113,N_7865);
or U12830 (N_12830,N_9232,N_6037);
nand U12831 (N_12831,N_5389,N_9124);
nand U12832 (N_12832,N_7352,N_7524);
nor U12833 (N_12833,N_5259,N_8758);
nand U12834 (N_12834,N_5687,N_9390);
and U12835 (N_12835,N_5427,N_5508);
or U12836 (N_12836,N_7601,N_7086);
or U12837 (N_12837,N_5914,N_6292);
nor U12838 (N_12838,N_9634,N_5419);
nor U12839 (N_12839,N_8321,N_8410);
nor U12840 (N_12840,N_8525,N_6376);
or U12841 (N_12841,N_6496,N_5516);
and U12842 (N_12842,N_9038,N_8505);
nand U12843 (N_12843,N_7281,N_7593);
and U12844 (N_12844,N_9620,N_7108);
and U12845 (N_12845,N_5403,N_9769);
nor U12846 (N_12846,N_7974,N_5112);
nand U12847 (N_12847,N_5649,N_5587);
and U12848 (N_12848,N_5638,N_5369);
or U12849 (N_12849,N_8705,N_9367);
or U12850 (N_12850,N_9428,N_6177);
nor U12851 (N_12851,N_7146,N_7955);
nor U12852 (N_12852,N_8078,N_9512);
and U12853 (N_12853,N_6129,N_7197);
or U12854 (N_12854,N_9516,N_9380);
and U12855 (N_12855,N_8209,N_6370);
or U12856 (N_12856,N_5312,N_8033);
and U12857 (N_12857,N_5923,N_9257);
nand U12858 (N_12858,N_9098,N_8256);
nand U12859 (N_12859,N_8777,N_5132);
nand U12860 (N_12860,N_8870,N_6311);
nor U12861 (N_12861,N_7573,N_6067);
nand U12862 (N_12862,N_8065,N_7352);
nand U12863 (N_12863,N_5080,N_7802);
nand U12864 (N_12864,N_8865,N_5513);
and U12865 (N_12865,N_9689,N_6344);
and U12866 (N_12866,N_9312,N_8597);
nor U12867 (N_12867,N_7713,N_6551);
nor U12868 (N_12868,N_6659,N_6234);
nor U12869 (N_12869,N_8810,N_8223);
or U12870 (N_12870,N_9791,N_7755);
nor U12871 (N_12871,N_9700,N_8373);
nor U12872 (N_12872,N_9774,N_6089);
nand U12873 (N_12873,N_5873,N_7837);
nand U12874 (N_12874,N_9884,N_7486);
nor U12875 (N_12875,N_9479,N_6138);
nand U12876 (N_12876,N_9904,N_8334);
and U12877 (N_12877,N_9605,N_5243);
nor U12878 (N_12878,N_6143,N_8246);
or U12879 (N_12879,N_6588,N_8452);
and U12880 (N_12880,N_6627,N_9025);
nand U12881 (N_12881,N_7657,N_8797);
or U12882 (N_12882,N_5424,N_7626);
or U12883 (N_12883,N_7105,N_9804);
or U12884 (N_12884,N_8036,N_8251);
and U12885 (N_12885,N_5939,N_7710);
nand U12886 (N_12886,N_8813,N_8347);
nand U12887 (N_12887,N_7751,N_9238);
or U12888 (N_12888,N_7077,N_5609);
or U12889 (N_12889,N_8210,N_8660);
nor U12890 (N_12890,N_8561,N_9317);
nand U12891 (N_12891,N_7550,N_6182);
and U12892 (N_12892,N_8314,N_7979);
nand U12893 (N_12893,N_6799,N_9167);
nand U12894 (N_12894,N_7289,N_6939);
and U12895 (N_12895,N_5290,N_7271);
nand U12896 (N_12896,N_7521,N_7631);
nor U12897 (N_12897,N_9758,N_6732);
nand U12898 (N_12898,N_9374,N_7509);
nand U12899 (N_12899,N_8902,N_5965);
nand U12900 (N_12900,N_6521,N_9337);
and U12901 (N_12901,N_7925,N_6740);
or U12902 (N_12902,N_6245,N_6750);
nand U12903 (N_12903,N_7311,N_7922);
nor U12904 (N_12904,N_5659,N_8873);
and U12905 (N_12905,N_8120,N_6061);
nand U12906 (N_12906,N_6456,N_7140);
and U12907 (N_12907,N_6972,N_6011);
nand U12908 (N_12908,N_9356,N_6199);
and U12909 (N_12909,N_6737,N_6971);
nand U12910 (N_12910,N_9610,N_5098);
xnor U12911 (N_12911,N_8726,N_7553);
nand U12912 (N_12912,N_9818,N_6832);
or U12913 (N_12913,N_6661,N_7372);
or U12914 (N_12914,N_6563,N_9133);
or U12915 (N_12915,N_6114,N_9300);
or U12916 (N_12916,N_8851,N_8490);
nor U12917 (N_12917,N_5895,N_7284);
nand U12918 (N_12918,N_6722,N_8118);
nand U12919 (N_12919,N_9295,N_7815);
or U12920 (N_12920,N_7942,N_8247);
and U12921 (N_12921,N_5633,N_9776);
or U12922 (N_12922,N_6678,N_7944);
nor U12923 (N_12923,N_7058,N_5410);
nand U12924 (N_12924,N_6995,N_6864);
and U12925 (N_12925,N_7041,N_9720);
nand U12926 (N_12926,N_8958,N_7128);
xnor U12927 (N_12927,N_7558,N_6057);
nand U12928 (N_12928,N_9505,N_9348);
and U12929 (N_12929,N_7337,N_7406);
or U12930 (N_12930,N_6623,N_6127);
nand U12931 (N_12931,N_7345,N_6512);
nor U12932 (N_12932,N_5308,N_9737);
and U12933 (N_12933,N_5651,N_5829);
and U12934 (N_12934,N_6492,N_7311);
nand U12935 (N_12935,N_7240,N_9811);
nand U12936 (N_12936,N_9447,N_5670);
and U12937 (N_12937,N_5767,N_6410);
and U12938 (N_12938,N_8908,N_7286);
or U12939 (N_12939,N_5592,N_6641);
nor U12940 (N_12940,N_9742,N_8244);
or U12941 (N_12941,N_5092,N_9405);
and U12942 (N_12942,N_7290,N_8150);
or U12943 (N_12943,N_5528,N_9557);
nor U12944 (N_12944,N_8022,N_6284);
nor U12945 (N_12945,N_5219,N_5842);
and U12946 (N_12946,N_9256,N_8421);
and U12947 (N_12947,N_7555,N_6528);
nor U12948 (N_12948,N_5743,N_8332);
and U12949 (N_12949,N_7692,N_7087);
nand U12950 (N_12950,N_9465,N_8546);
nor U12951 (N_12951,N_9230,N_9416);
or U12952 (N_12952,N_6063,N_9112);
nor U12953 (N_12953,N_8268,N_6910);
and U12954 (N_12954,N_8134,N_6235);
or U12955 (N_12955,N_8887,N_9348);
nor U12956 (N_12956,N_8429,N_6291);
and U12957 (N_12957,N_6741,N_7771);
nor U12958 (N_12958,N_5412,N_8476);
nor U12959 (N_12959,N_8336,N_9530);
and U12960 (N_12960,N_7656,N_8572);
and U12961 (N_12961,N_7126,N_9035);
and U12962 (N_12962,N_9363,N_7353);
and U12963 (N_12963,N_8754,N_6800);
nor U12964 (N_12964,N_9823,N_7268);
or U12965 (N_12965,N_7416,N_8733);
or U12966 (N_12966,N_8426,N_7479);
nand U12967 (N_12967,N_9671,N_6657);
nor U12968 (N_12968,N_7467,N_5287);
nand U12969 (N_12969,N_5847,N_9283);
or U12970 (N_12970,N_6788,N_5536);
nor U12971 (N_12971,N_5935,N_9434);
nor U12972 (N_12972,N_6639,N_8125);
or U12973 (N_12973,N_9610,N_6112);
nand U12974 (N_12974,N_8428,N_6315);
nor U12975 (N_12975,N_8911,N_8113);
or U12976 (N_12976,N_9940,N_5105);
nor U12977 (N_12977,N_9210,N_5254);
or U12978 (N_12978,N_7332,N_7830);
nor U12979 (N_12979,N_5420,N_6267);
or U12980 (N_12980,N_5351,N_8396);
nor U12981 (N_12981,N_6455,N_8072);
nand U12982 (N_12982,N_8373,N_7030);
nor U12983 (N_12983,N_9991,N_7454);
nor U12984 (N_12984,N_5909,N_8861);
nand U12985 (N_12985,N_8920,N_8699);
nand U12986 (N_12986,N_7846,N_9813);
and U12987 (N_12987,N_7232,N_7096);
nor U12988 (N_12988,N_5211,N_5405);
and U12989 (N_12989,N_9488,N_7769);
or U12990 (N_12990,N_7469,N_9102);
nand U12991 (N_12991,N_7015,N_6699);
or U12992 (N_12992,N_9098,N_5861);
or U12993 (N_12993,N_8604,N_6034);
or U12994 (N_12994,N_6108,N_9595);
and U12995 (N_12995,N_6096,N_7803);
nand U12996 (N_12996,N_9288,N_7248);
nor U12997 (N_12997,N_8191,N_6032);
and U12998 (N_12998,N_6261,N_7192);
nor U12999 (N_12999,N_7973,N_7585);
or U13000 (N_13000,N_5973,N_8598);
nand U13001 (N_13001,N_9243,N_8709);
or U13002 (N_13002,N_6828,N_5693);
nor U13003 (N_13003,N_8468,N_7420);
nand U13004 (N_13004,N_6171,N_6492);
nand U13005 (N_13005,N_8236,N_6590);
and U13006 (N_13006,N_8143,N_5822);
nor U13007 (N_13007,N_8732,N_6046);
nor U13008 (N_13008,N_5786,N_9627);
nand U13009 (N_13009,N_7429,N_5935);
nand U13010 (N_13010,N_5405,N_6012);
and U13011 (N_13011,N_5574,N_9967);
or U13012 (N_13012,N_8737,N_5549);
nand U13013 (N_13013,N_7684,N_5792);
and U13014 (N_13014,N_6032,N_7654);
nor U13015 (N_13015,N_6834,N_5299);
or U13016 (N_13016,N_5014,N_6332);
nand U13017 (N_13017,N_8533,N_7324);
nor U13018 (N_13018,N_6866,N_7849);
and U13019 (N_13019,N_8372,N_8472);
nand U13020 (N_13020,N_5740,N_7906);
or U13021 (N_13021,N_8070,N_8286);
nand U13022 (N_13022,N_8163,N_6725);
and U13023 (N_13023,N_8974,N_8382);
or U13024 (N_13024,N_9721,N_9795);
nor U13025 (N_13025,N_6816,N_5440);
nand U13026 (N_13026,N_9012,N_7017);
nand U13027 (N_13027,N_5787,N_8387);
nor U13028 (N_13028,N_6805,N_6844);
nor U13029 (N_13029,N_8857,N_8588);
nor U13030 (N_13030,N_8496,N_5873);
nand U13031 (N_13031,N_5461,N_8199);
nand U13032 (N_13032,N_9607,N_7039);
or U13033 (N_13033,N_7903,N_5578);
nor U13034 (N_13034,N_9007,N_9219);
nand U13035 (N_13035,N_7097,N_8012);
nor U13036 (N_13036,N_8342,N_8205);
or U13037 (N_13037,N_7208,N_9677);
nor U13038 (N_13038,N_7749,N_5133);
nor U13039 (N_13039,N_7719,N_5986);
and U13040 (N_13040,N_7670,N_9447);
nor U13041 (N_13041,N_9891,N_6067);
and U13042 (N_13042,N_7171,N_6605);
or U13043 (N_13043,N_6052,N_6013);
nor U13044 (N_13044,N_6008,N_6114);
nand U13045 (N_13045,N_7359,N_5757);
and U13046 (N_13046,N_9725,N_7268);
nor U13047 (N_13047,N_5993,N_8413);
or U13048 (N_13048,N_9524,N_8559);
or U13049 (N_13049,N_8798,N_7507);
or U13050 (N_13050,N_5092,N_6879);
nand U13051 (N_13051,N_9652,N_8341);
and U13052 (N_13052,N_6943,N_6951);
nor U13053 (N_13053,N_6986,N_5536);
and U13054 (N_13054,N_6865,N_9166);
nor U13055 (N_13055,N_9824,N_7267);
nor U13056 (N_13056,N_5789,N_7673);
and U13057 (N_13057,N_6833,N_5641);
nand U13058 (N_13058,N_6862,N_9455);
nand U13059 (N_13059,N_7050,N_8188);
nand U13060 (N_13060,N_9921,N_6465);
and U13061 (N_13061,N_6320,N_9146);
and U13062 (N_13062,N_8701,N_6749);
nor U13063 (N_13063,N_6664,N_5875);
or U13064 (N_13064,N_7339,N_5813);
nand U13065 (N_13065,N_5424,N_7270);
or U13066 (N_13066,N_6209,N_8432);
nor U13067 (N_13067,N_7462,N_7169);
or U13068 (N_13068,N_7448,N_9915);
or U13069 (N_13069,N_5721,N_9474);
or U13070 (N_13070,N_9047,N_7681);
nand U13071 (N_13071,N_9743,N_6089);
nor U13072 (N_13072,N_6342,N_8021);
and U13073 (N_13073,N_7546,N_5372);
and U13074 (N_13074,N_6379,N_7472);
nand U13075 (N_13075,N_9665,N_9619);
nand U13076 (N_13076,N_5431,N_7590);
or U13077 (N_13077,N_8645,N_8543);
and U13078 (N_13078,N_8063,N_8430);
nand U13079 (N_13079,N_8095,N_5480);
and U13080 (N_13080,N_5838,N_8333);
and U13081 (N_13081,N_5365,N_6278);
and U13082 (N_13082,N_6005,N_7245);
nand U13083 (N_13083,N_7250,N_9497);
or U13084 (N_13084,N_9586,N_7981);
nor U13085 (N_13085,N_6034,N_6155);
and U13086 (N_13086,N_9138,N_9955);
nor U13087 (N_13087,N_6593,N_7536);
or U13088 (N_13088,N_8269,N_8307);
or U13089 (N_13089,N_5671,N_6454);
or U13090 (N_13090,N_8180,N_9852);
or U13091 (N_13091,N_8649,N_8926);
nor U13092 (N_13092,N_6715,N_8632);
or U13093 (N_13093,N_8262,N_5927);
or U13094 (N_13094,N_7471,N_5633);
or U13095 (N_13095,N_5967,N_8287);
nor U13096 (N_13096,N_8781,N_8444);
nor U13097 (N_13097,N_5901,N_6431);
or U13098 (N_13098,N_9637,N_6970);
xor U13099 (N_13099,N_6684,N_8569);
nand U13100 (N_13100,N_6981,N_6314);
nor U13101 (N_13101,N_8830,N_7605);
nor U13102 (N_13102,N_6970,N_8606);
or U13103 (N_13103,N_8280,N_6287);
nor U13104 (N_13104,N_8882,N_5320);
nor U13105 (N_13105,N_8704,N_5045);
and U13106 (N_13106,N_6973,N_8332);
and U13107 (N_13107,N_8324,N_8499);
nor U13108 (N_13108,N_5857,N_9433);
and U13109 (N_13109,N_6931,N_7959);
or U13110 (N_13110,N_5537,N_6327);
and U13111 (N_13111,N_7971,N_6549);
nand U13112 (N_13112,N_7113,N_6012);
or U13113 (N_13113,N_5283,N_9738);
nand U13114 (N_13114,N_8862,N_9757);
or U13115 (N_13115,N_6432,N_6019);
and U13116 (N_13116,N_7391,N_8285);
and U13117 (N_13117,N_7935,N_5924);
nor U13118 (N_13118,N_5792,N_8590);
and U13119 (N_13119,N_5849,N_7709);
or U13120 (N_13120,N_8405,N_6995);
or U13121 (N_13121,N_8054,N_5341);
nor U13122 (N_13122,N_9884,N_5516);
nor U13123 (N_13123,N_8299,N_5013);
nor U13124 (N_13124,N_9599,N_7766);
nor U13125 (N_13125,N_7332,N_9334);
nand U13126 (N_13126,N_6199,N_5079);
nor U13127 (N_13127,N_9060,N_6928);
nand U13128 (N_13128,N_8979,N_6083);
and U13129 (N_13129,N_7299,N_7091);
and U13130 (N_13130,N_6930,N_7461);
nor U13131 (N_13131,N_6895,N_9439);
and U13132 (N_13132,N_6946,N_5752);
xor U13133 (N_13133,N_7091,N_7456);
nor U13134 (N_13134,N_6935,N_8091);
nand U13135 (N_13135,N_9249,N_6346);
and U13136 (N_13136,N_8703,N_6961);
nor U13137 (N_13137,N_8455,N_8135);
nand U13138 (N_13138,N_7021,N_9693);
or U13139 (N_13139,N_6885,N_8305);
nand U13140 (N_13140,N_5501,N_9144);
and U13141 (N_13141,N_7816,N_6425);
nand U13142 (N_13142,N_6172,N_6655);
nand U13143 (N_13143,N_9723,N_8328);
or U13144 (N_13144,N_8447,N_8617);
nor U13145 (N_13145,N_9023,N_9967);
or U13146 (N_13146,N_6353,N_9478);
and U13147 (N_13147,N_7220,N_8203);
nor U13148 (N_13148,N_7142,N_6394);
or U13149 (N_13149,N_7555,N_6353);
nor U13150 (N_13150,N_8555,N_6066);
nor U13151 (N_13151,N_6390,N_6890);
or U13152 (N_13152,N_8040,N_9142);
or U13153 (N_13153,N_5875,N_7396);
nand U13154 (N_13154,N_6037,N_9783);
nor U13155 (N_13155,N_6026,N_5168);
and U13156 (N_13156,N_8998,N_8002);
or U13157 (N_13157,N_5111,N_5514);
nand U13158 (N_13158,N_7426,N_5154);
and U13159 (N_13159,N_9431,N_9237);
and U13160 (N_13160,N_6766,N_8448);
and U13161 (N_13161,N_5933,N_5222);
nand U13162 (N_13162,N_5028,N_9684);
or U13163 (N_13163,N_8625,N_8524);
or U13164 (N_13164,N_9094,N_8642);
nor U13165 (N_13165,N_6809,N_9140);
nand U13166 (N_13166,N_9440,N_5432);
nand U13167 (N_13167,N_8026,N_8716);
and U13168 (N_13168,N_5771,N_8669);
nor U13169 (N_13169,N_5537,N_6230);
nor U13170 (N_13170,N_7854,N_6653);
nor U13171 (N_13171,N_7602,N_5741);
nor U13172 (N_13172,N_6861,N_9810);
nand U13173 (N_13173,N_8580,N_6424);
and U13174 (N_13174,N_9209,N_8526);
nor U13175 (N_13175,N_8335,N_7803);
or U13176 (N_13176,N_9334,N_9655);
nand U13177 (N_13177,N_5548,N_5238);
nand U13178 (N_13178,N_8457,N_9853);
or U13179 (N_13179,N_8748,N_7988);
nand U13180 (N_13180,N_5803,N_9690);
and U13181 (N_13181,N_9189,N_9629);
and U13182 (N_13182,N_9365,N_7999);
xor U13183 (N_13183,N_7126,N_7352);
or U13184 (N_13184,N_7445,N_9228);
nand U13185 (N_13185,N_9107,N_9173);
nor U13186 (N_13186,N_9639,N_6243);
nand U13187 (N_13187,N_6885,N_8550);
nor U13188 (N_13188,N_8636,N_8389);
or U13189 (N_13189,N_9622,N_7652);
nand U13190 (N_13190,N_7812,N_8180);
nand U13191 (N_13191,N_6174,N_8460);
nor U13192 (N_13192,N_8548,N_6943);
nor U13193 (N_13193,N_7906,N_9412);
nor U13194 (N_13194,N_7092,N_7987);
nand U13195 (N_13195,N_9911,N_9624);
or U13196 (N_13196,N_9454,N_5396);
and U13197 (N_13197,N_5246,N_5261);
nor U13198 (N_13198,N_8135,N_5845);
nand U13199 (N_13199,N_5518,N_8540);
nor U13200 (N_13200,N_9067,N_7561);
and U13201 (N_13201,N_6394,N_7795);
nor U13202 (N_13202,N_8440,N_9723);
and U13203 (N_13203,N_8999,N_8311);
nand U13204 (N_13204,N_7148,N_9647);
nand U13205 (N_13205,N_9772,N_9756);
nor U13206 (N_13206,N_6194,N_5977);
or U13207 (N_13207,N_6169,N_7157);
nor U13208 (N_13208,N_8332,N_8432);
nand U13209 (N_13209,N_9754,N_6852);
and U13210 (N_13210,N_9251,N_9413);
xnor U13211 (N_13211,N_9470,N_9468);
or U13212 (N_13212,N_9260,N_7656);
nand U13213 (N_13213,N_8093,N_8552);
nand U13214 (N_13214,N_6419,N_9812);
nand U13215 (N_13215,N_7155,N_8664);
nand U13216 (N_13216,N_8520,N_8263);
or U13217 (N_13217,N_8596,N_7907);
nor U13218 (N_13218,N_7488,N_5514);
nor U13219 (N_13219,N_8473,N_7455);
nand U13220 (N_13220,N_6663,N_6193);
and U13221 (N_13221,N_5527,N_7800);
or U13222 (N_13222,N_7315,N_9169);
and U13223 (N_13223,N_5701,N_9303);
or U13224 (N_13224,N_8813,N_7310);
and U13225 (N_13225,N_9491,N_5036);
or U13226 (N_13226,N_7946,N_9273);
nand U13227 (N_13227,N_8154,N_9454);
and U13228 (N_13228,N_5873,N_9445);
or U13229 (N_13229,N_8658,N_7183);
or U13230 (N_13230,N_6355,N_7767);
or U13231 (N_13231,N_9194,N_7640);
nand U13232 (N_13232,N_9723,N_7939);
or U13233 (N_13233,N_8081,N_6458);
nor U13234 (N_13234,N_9965,N_9897);
nor U13235 (N_13235,N_5746,N_8515);
nand U13236 (N_13236,N_6242,N_7335);
nor U13237 (N_13237,N_6609,N_9776);
nand U13238 (N_13238,N_9667,N_7796);
nor U13239 (N_13239,N_5479,N_6195);
or U13240 (N_13240,N_7940,N_8967);
and U13241 (N_13241,N_7438,N_8464);
xnor U13242 (N_13242,N_5245,N_6332);
or U13243 (N_13243,N_5797,N_6736);
nand U13244 (N_13244,N_8455,N_6656);
nor U13245 (N_13245,N_8885,N_8309);
nand U13246 (N_13246,N_7710,N_5727);
or U13247 (N_13247,N_9263,N_8725);
nor U13248 (N_13248,N_8077,N_7458);
nor U13249 (N_13249,N_8784,N_9463);
and U13250 (N_13250,N_5945,N_8332);
nand U13251 (N_13251,N_7479,N_7418);
or U13252 (N_13252,N_7080,N_6163);
and U13253 (N_13253,N_9661,N_7752);
or U13254 (N_13254,N_6993,N_5327);
nor U13255 (N_13255,N_8178,N_6700);
or U13256 (N_13256,N_8269,N_9980);
nand U13257 (N_13257,N_6370,N_6139);
nand U13258 (N_13258,N_7391,N_6428);
or U13259 (N_13259,N_7322,N_5234);
and U13260 (N_13260,N_5997,N_8457);
nand U13261 (N_13261,N_8106,N_8367);
or U13262 (N_13262,N_9324,N_6226);
nand U13263 (N_13263,N_9696,N_8129);
or U13264 (N_13264,N_8212,N_6215);
and U13265 (N_13265,N_8469,N_6342);
nand U13266 (N_13266,N_7430,N_9998);
nor U13267 (N_13267,N_5788,N_8177);
nor U13268 (N_13268,N_5446,N_8353);
nand U13269 (N_13269,N_5645,N_5711);
and U13270 (N_13270,N_8908,N_7627);
and U13271 (N_13271,N_5883,N_9833);
or U13272 (N_13272,N_5421,N_6477);
or U13273 (N_13273,N_8617,N_7430);
nor U13274 (N_13274,N_9283,N_7880);
or U13275 (N_13275,N_9460,N_5837);
nor U13276 (N_13276,N_6622,N_9832);
nor U13277 (N_13277,N_8074,N_5743);
and U13278 (N_13278,N_6069,N_8678);
xnor U13279 (N_13279,N_6234,N_5374);
nor U13280 (N_13280,N_8838,N_7985);
nor U13281 (N_13281,N_8746,N_6454);
nor U13282 (N_13282,N_7328,N_5548);
nor U13283 (N_13283,N_7381,N_8901);
nor U13284 (N_13284,N_8483,N_5992);
nor U13285 (N_13285,N_8983,N_5287);
nor U13286 (N_13286,N_6997,N_8484);
and U13287 (N_13287,N_5032,N_5886);
nand U13288 (N_13288,N_5346,N_7950);
or U13289 (N_13289,N_6848,N_9045);
nand U13290 (N_13290,N_7610,N_5133);
nand U13291 (N_13291,N_7237,N_9130);
and U13292 (N_13292,N_6876,N_6086);
xnor U13293 (N_13293,N_6682,N_9717);
nor U13294 (N_13294,N_6922,N_6283);
and U13295 (N_13295,N_5306,N_9458);
or U13296 (N_13296,N_5489,N_7517);
and U13297 (N_13297,N_8075,N_8405);
or U13298 (N_13298,N_9864,N_7446);
and U13299 (N_13299,N_8593,N_6850);
and U13300 (N_13300,N_8415,N_7242);
nor U13301 (N_13301,N_7310,N_7362);
or U13302 (N_13302,N_7310,N_5177);
and U13303 (N_13303,N_5718,N_5912);
nor U13304 (N_13304,N_5307,N_6045);
nor U13305 (N_13305,N_8814,N_6557);
nor U13306 (N_13306,N_7045,N_7331);
nand U13307 (N_13307,N_9739,N_5214);
nand U13308 (N_13308,N_8532,N_9228);
nor U13309 (N_13309,N_6720,N_7054);
or U13310 (N_13310,N_7645,N_5873);
or U13311 (N_13311,N_7315,N_9528);
nand U13312 (N_13312,N_7413,N_5899);
or U13313 (N_13313,N_5169,N_6230);
and U13314 (N_13314,N_7683,N_6603);
nor U13315 (N_13315,N_9722,N_9846);
nand U13316 (N_13316,N_7456,N_5125);
nor U13317 (N_13317,N_8547,N_5444);
or U13318 (N_13318,N_5382,N_9736);
or U13319 (N_13319,N_6853,N_9220);
and U13320 (N_13320,N_5540,N_7313);
or U13321 (N_13321,N_9280,N_8459);
and U13322 (N_13322,N_8565,N_7576);
nand U13323 (N_13323,N_5028,N_6968);
or U13324 (N_13324,N_8177,N_7954);
nand U13325 (N_13325,N_7918,N_8267);
nand U13326 (N_13326,N_5720,N_5098);
nand U13327 (N_13327,N_8770,N_5112);
nand U13328 (N_13328,N_8293,N_7282);
nor U13329 (N_13329,N_8716,N_5434);
nand U13330 (N_13330,N_5770,N_7364);
nor U13331 (N_13331,N_6309,N_7809);
nor U13332 (N_13332,N_7573,N_5620);
nand U13333 (N_13333,N_6533,N_5749);
and U13334 (N_13334,N_5969,N_7686);
nor U13335 (N_13335,N_9391,N_6359);
or U13336 (N_13336,N_9059,N_9667);
or U13337 (N_13337,N_5221,N_8955);
nor U13338 (N_13338,N_5606,N_9049);
and U13339 (N_13339,N_7553,N_9624);
nand U13340 (N_13340,N_9131,N_8891);
and U13341 (N_13341,N_5743,N_8318);
nor U13342 (N_13342,N_6611,N_9271);
nor U13343 (N_13343,N_6094,N_9728);
nand U13344 (N_13344,N_5399,N_9562);
and U13345 (N_13345,N_5250,N_7210);
and U13346 (N_13346,N_6376,N_6587);
nor U13347 (N_13347,N_6432,N_5200);
nor U13348 (N_13348,N_8102,N_6146);
and U13349 (N_13349,N_5760,N_5293);
nor U13350 (N_13350,N_8677,N_8678);
nand U13351 (N_13351,N_6921,N_8915);
nor U13352 (N_13352,N_7328,N_9121);
nand U13353 (N_13353,N_9331,N_9338);
nand U13354 (N_13354,N_7148,N_6553);
or U13355 (N_13355,N_9593,N_5178);
nor U13356 (N_13356,N_6617,N_6128);
and U13357 (N_13357,N_9273,N_7083);
nand U13358 (N_13358,N_8046,N_5579);
or U13359 (N_13359,N_6955,N_9131);
nor U13360 (N_13360,N_6701,N_8602);
or U13361 (N_13361,N_6129,N_7913);
nor U13362 (N_13362,N_8719,N_7604);
nor U13363 (N_13363,N_6060,N_8771);
and U13364 (N_13364,N_9495,N_8065);
nand U13365 (N_13365,N_5565,N_5818);
and U13366 (N_13366,N_8532,N_8145);
or U13367 (N_13367,N_6775,N_6638);
or U13368 (N_13368,N_6905,N_6245);
nor U13369 (N_13369,N_5473,N_5953);
nand U13370 (N_13370,N_8615,N_5146);
nand U13371 (N_13371,N_5213,N_7490);
or U13372 (N_13372,N_7198,N_7605);
nor U13373 (N_13373,N_7540,N_8429);
nand U13374 (N_13374,N_9594,N_6698);
nand U13375 (N_13375,N_8797,N_8276);
and U13376 (N_13376,N_5053,N_6843);
xor U13377 (N_13377,N_7176,N_7310);
nor U13378 (N_13378,N_8456,N_8636);
and U13379 (N_13379,N_9069,N_7877);
and U13380 (N_13380,N_5116,N_9416);
nor U13381 (N_13381,N_7716,N_6828);
nand U13382 (N_13382,N_6404,N_7417);
nor U13383 (N_13383,N_6383,N_5890);
and U13384 (N_13384,N_7457,N_5695);
nand U13385 (N_13385,N_7833,N_5865);
nor U13386 (N_13386,N_7195,N_6797);
or U13387 (N_13387,N_5780,N_8449);
nor U13388 (N_13388,N_5547,N_8865);
nand U13389 (N_13389,N_6354,N_7788);
nand U13390 (N_13390,N_9292,N_5967);
and U13391 (N_13391,N_6989,N_8509);
nor U13392 (N_13392,N_6698,N_5151);
or U13393 (N_13393,N_8705,N_9553);
nand U13394 (N_13394,N_8770,N_6355);
nor U13395 (N_13395,N_9169,N_5175);
nor U13396 (N_13396,N_6117,N_6108);
nand U13397 (N_13397,N_8842,N_6884);
nor U13398 (N_13398,N_6418,N_8607);
and U13399 (N_13399,N_8469,N_5186);
or U13400 (N_13400,N_6162,N_7044);
nor U13401 (N_13401,N_9344,N_8204);
nor U13402 (N_13402,N_5887,N_8240);
and U13403 (N_13403,N_5452,N_7138);
nand U13404 (N_13404,N_6837,N_8881);
and U13405 (N_13405,N_9808,N_7122);
nand U13406 (N_13406,N_7387,N_7252);
nor U13407 (N_13407,N_8990,N_9106);
and U13408 (N_13408,N_6328,N_7940);
nor U13409 (N_13409,N_6854,N_5752);
nand U13410 (N_13410,N_8578,N_7652);
and U13411 (N_13411,N_7737,N_8014);
and U13412 (N_13412,N_7960,N_9069);
and U13413 (N_13413,N_6868,N_8816);
and U13414 (N_13414,N_8634,N_5727);
or U13415 (N_13415,N_5461,N_7242);
nor U13416 (N_13416,N_6631,N_8928);
and U13417 (N_13417,N_8610,N_5728);
or U13418 (N_13418,N_9483,N_5548);
xor U13419 (N_13419,N_8946,N_8730);
nor U13420 (N_13420,N_6399,N_6814);
or U13421 (N_13421,N_5622,N_9260);
nor U13422 (N_13422,N_7289,N_7236);
and U13423 (N_13423,N_8617,N_9785);
nor U13424 (N_13424,N_8916,N_5454);
nor U13425 (N_13425,N_9654,N_9061);
nor U13426 (N_13426,N_8092,N_9233);
nor U13427 (N_13427,N_7838,N_6532);
nand U13428 (N_13428,N_9557,N_8792);
nand U13429 (N_13429,N_8134,N_9959);
nand U13430 (N_13430,N_7810,N_7058);
nand U13431 (N_13431,N_8126,N_7121);
nand U13432 (N_13432,N_9288,N_9708);
and U13433 (N_13433,N_7084,N_5482);
nand U13434 (N_13434,N_7940,N_6644);
and U13435 (N_13435,N_9783,N_5634);
and U13436 (N_13436,N_8527,N_9325);
nand U13437 (N_13437,N_8831,N_9096);
and U13438 (N_13438,N_8673,N_7006);
nor U13439 (N_13439,N_8595,N_5742);
and U13440 (N_13440,N_7203,N_6251);
or U13441 (N_13441,N_5948,N_8485);
nor U13442 (N_13442,N_7094,N_7675);
or U13443 (N_13443,N_8322,N_5002);
or U13444 (N_13444,N_5975,N_6158);
nand U13445 (N_13445,N_5373,N_9437);
nand U13446 (N_13446,N_7643,N_8083);
nand U13447 (N_13447,N_5859,N_9648);
nor U13448 (N_13448,N_5272,N_9233);
and U13449 (N_13449,N_7723,N_8938);
or U13450 (N_13450,N_5842,N_6061);
or U13451 (N_13451,N_5858,N_6516);
nor U13452 (N_13452,N_8419,N_5377);
nand U13453 (N_13453,N_7369,N_7245);
nand U13454 (N_13454,N_8119,N_7170);
nand U13455 (N_13455,N_8267,N_6147);
or U13456 (N_13456,N_7691,N_7496);
nor U13457 (N_13457,N_7165,N_7659);
and U13458 (N_13458,N_8441,N_8524);
and U13459 (N_13459,N_8979,N_6318);
nand U13460 (N_13460,N_5837,N_9694);
nor U13461 (N_13461,N_8027,N_7427);
nor U13462 (N_13462,N_9878,N_6107);
and U13463 (N_13463,N_8855,N_9166);
nand U13464 (N_13464,N_7517,N_6631);
nor U13465 (N_13465,N_6478,N_5217);
nand U13466 (N_13466,N_8940,N_5197);
nor U13467 (N_13467,N_7784,N_5807);
nand U13468 (N_13468,N_8694,N_9078);
nor U13469 (N_13469,N_5981,N_9302);
and U13470 (N_13470,N_9985,N_6543);
or U13471 (N_13471,N_7764,N_8024);
or U13472 (N_13472,N_9189,N_8243);
nor U13473 (N_13473,N_5373,N_5262);
and U13474 (N_13474,N_9602,N_8108);
nand U13475 (N_13475,N_5591,N_8983);
and U13476 (N_13476,N_6862,N_9033);
nand U13477 (N_13477,N_8443,N_9430);
nor U13478 (N_13478,N_6246,N_7374);
nor U13479 (N_13479,N_9712,N_5463);
and U13480 (N_13480,N_8182,N_7977);
and U13481 (N_13481,N_9316,N_8761);
nand U13482 (N_13482,N_9465,N_7288);
nand U13483 (N_13483,N_6966,N_6205);
nand U13484 (N_13484,N_8254,N_8688);
or U13485 (N_13485,N_8132,N_6795);
and U13486 (N_13486,N_9551,N_7627);
and U13487 (N_13487,N_6146,N_5721);
or U13488 (N_13488,N_7832,N_9092);
and U13489 (N_13489,N_8686,N_6715);
nor U13490 (N_13490,N_7375,N_8849);
nor U13491 (N_13491,N_9950,N_8966);
and U13492 (N_13492,N_6336,N_5011);
nor U13493 (N_13493,N_8637,N_8028);
and U13494 (N_13494,N_7888,N_7711);
and U13495 (N_13495,N_6207,N_8270);
nand U13496 (N_13496,N_9406,N_5717);
or U13497 (N_13497,N_9633,N_7984);
nand U13498 (N_13498,N_5582,N_8437);
nor U13499 (N_13499,N_5125,N_6779);
and U13500 (N_13500,N_8065,N_9812);
or U13501 (N_13501,N_7917,N_9035);
or U13502 (N_13502,N_6361,N_9827);
nor U13503 (N_13503,N_5934,N_5132);
or U13504 (N_13504,N_5811,N_5406);
or U13505 (N_13505,N_5774,N_9478);
or U13506 (N_13506,N_7722,N_9420);
nor U13507 (N_13507,N_8887,N_7850);
and U13508 (N_13508,N_7004,N_5200);
and U13509 (N_13509,N_6694,N_5609);
or U13510 (N_13510,N_6986,N_6111);
or U13511 (N_13511,N_6651,N_6033);
nor U13512 (N_13512,N_8847,N_8127);
or U13513 (N_13513,N_9058,N_5878);
nand U13514 (N_13514,N_7985,N_8149);
nand U13515 (N_13515,N_8201,N_8310);
or U13516 (N_13516,N_9969,N_5413);
or U13517 (N_13517,N_9546,N_9739);
or U13518 (N_13518,N_6547,N_5451);
nand U13519 (N_13519,N_8331,N_7336);
and U13520 (N_13520,N_6352,N_5020);
and U13521 (N_13521,N_6091,N_9199);
or U13522 (N_13522,N_5832,N_6258);
or U13523 (N_13523,N_5756,N_5627);
and U13524 (N_13524,N_6862,N_7969);
and U13525 (N_13525,N_8740,N_5753);
or U13526 (N_13526,N_5774,N_6028);
nor U13527 (N_13527,N_9268,N_5860);
or U13528 (N_13528,N_5919,N_5055);
nand U13529 (N_13529,N_5891,N_8808);
or U13530 (N_13530,N_9219,N_8115);
or U13531 (N_13531,N_7794,N_8958);
nand U13532 (N_13532,N_9611,N_9975);
or U13533 (N_13533,N_9896,N_6998);
and U13534 (N_13534,N_6639,N_8545);
nand U13535 (N_13535,N_5861,N_6572);
nor U13536 (N_13536,N_7496,N_7169);
xor U13537 (N_13537,N_6321,N_7112);
nor U13538 (N_13538,N_7506,N_6533);
nor U13539 (N_13539,N_7968,N_5486);
nand U13540 (N_13540,N_9109,N_7539);
xor U13541 (N_13541,N_5951,N_6360);
and U13542 (N_13542,N_5787,N_9822);
and U13543 (N_13543,N_5177,N_5868);
nand U13544 (N_13544,N_9572,N_5337);
nor U13545 (N_13545,N_5442,N_5332);
nor U13546 (N_13546,N_8496,N_5021);
and U13547 (N_13547,N_9332,N_8469);
nand U13548 (N_13548,N_8783,N_8768);
nor U13549 (N_13549,N_5772,N_8265);
nor U13550 (N_13550,N_7040,N_9872);
nor U13551 (N_13551,N_5237,N_6871);
nand U13552 (N_13552,N_7353,N_9251);
nor U13553 (N_13553,N_5470,N_7718);
and U13554 (N_13554,N_7036,N_8949);
nor U13555 (N_13555,N_8132,N_9282);
nand U13556 (N_13556,N_8806,N_5299);
and U13557 (N_13557,N_9156,N_5976);
and U13558 (N_13558,N_7705,N_8775);
nor U13559 (N_13559,N_6115,N_9135);
or U13560 (N_13560,N_8191,N_6064);
xnor U13561 (N_13561,N_7207,N_7292);
and U13562 (N_13562,N_6342,N_6276);
and U13563 (N_13563,N_6943,N_7723);
nand U13564 (N_13564,N_7298,N_7132);
and U13565 (N_13565,N_7257,N_6967);
or U13566 (N_13566,N_7501,N_6247);
and U13567 (N_13567,N_6821,N_8698);
nand U13568 (N_13568,N_9984,N_5499);
nand U13569 (N_13569,N_9111,N_8841);
and U13570 (N_13570,N_8655,N_5933);
nand U13571 (N_13571,N_7683,N_7389);
and U13572 (N_13572,N_9677,N_5937);
nand U13573 (N_13573,N_5234,N_7195);
nand U13574 (N_13574,N_7586,N_8078);
nand U13575 (N_13575,N_9405,N_9802);
and U13576 (N_13576,N_5159,N_7001);
and U13577 (N_13577,N_7734,N_9727);
nor U13578 (N_13578,N_9713,N_6247);
and U13579 (N_13579,N_7913,N_6983);
or U13580 (N_13580,N_7498,N_7537);
or U13581 (N_13581,N_8790,N_9975);
nand U13582 (N_13582,N_7265,N_7789);
or U13583 (N_13583,N_5185,N_5291);
nand U13584 (N_13584,N_7400,N_8525);
nand U13585 (N_13585,N_8871,N_9154);
and U13586 (N_13586,N_7581,N_5544);
nor U13587 (N_13587,N_7359,N_7732);
and U13588 (N_13588,N_8171,N_6838);
or U13589 (N_13589,N_9653,N_6495);
nand U13590 (N_13590,N_7326,N_8639);
or U13591 (N_13591,N_5087,N_6942);
nand U13592 (N_13592,N_8535,N_5792);
and U13593 (N_13593,N_9137,N_9696);
or U13594 (N_13594,N_5048,N_5263);
nand U13595 (N_13595,N_6799,N_7714);
nand U13596 (N_13596,N_9676,N_6024);
nand U13597 (N_13597,N_8603,N_7058);
nor U13598 (N_13598,N_5038,N_7541);
or U13599 (N_13599,N_5919,N_8652);
nor U13600 (N_13600,N_8453,N_9242);
xor U13601 (N_13601,N_9251,N_9114);
and U13602 (N_13602,N_7586,N_8441);
or U13603 (N_13603,N_6733,N_9100);
nor U13604 (N_13604,N_7584,N_5949);
and U13605 (N_13605,N_8669,N_8610);
or U13606 (N_13606,N_9675,N_9238);
and U13607 (N_13607,N_9065,N_9530);
and U13608 (N_13608,N_5198,N_9229);
nand U13609 (N_13609,N_7795,N_9581);
nor U13610 (N_13610,N_9575,N_5046);
and U13611 (N_13611,N_7905,N_7449);
or U13612 (N_13612,N_7331,N_6314);
nand U13613 (N_13613,N_6072,N_8796);
and U13614 (N_13614,N_7066,N_7726);
nor U13615 (N_13615,N_5666,N_6032);
nor U13616 (N_13616,N_5208,N_9792);
nand U13617 (N_13617,N_5926,N_8419);
or U13618 (N_13618,N_7308,N_6802);
or U13619 (N_13619,N_5083,N_6165);
nor U13620 (N_13620,N_6969,N_5265);
or U13621 (N_13621,N_8476,N_5294);
and U13622 (N_13622,N_9271,N_6576);
and U13623 (N_13623,N_6544,N_8119);
or U13624 (N_13624,N_9096,N_7663);
nand U13625 (N_13625,N_7834,N_9204);
or U13626 (N_13626,N_7052,N_6423);
nand U13627 (N_13627,N_6735,N_6690);
or U13628 (N_13628,N_7347,N_7134);
or U13629 (N_13629,N_6777,N_9373);
nand U13630 (N_13630,N_5221,N_5675);
and U13631 (N_13631,N_5177,N_7069);
nor U13632 (N_13632,N_9277,N_9107);
nor U13633 (N_13633,N_8427,N_8076);
or U13634 (N_13634,N_8734,N_6896);
nand U13635 (N_13635,N_8299,N_8896);
and U13636 (N_13636,N_9941,N_5498);
and U13637 (N_13637,N_9281,N_5348);
nor U13638 (N_13638,N_6167,N_9856);
nor U13639 (N_13639,N_6635,N_9349);
nand U13640 (N_13640,N_8911,N_7586);
and U13641 (N_13641,N_6164,N_5043);
nand U13642 (N_13642,N_5529,N_5980);
or U13643 (N_13643,N_8780,N_9393);
or U13644 (N_13644,N_9720,N_5824);
nor U13645 (N_13645,N_7797,N_7169);
and U13646 (N_13646,N_7340,N_7540);
nand U13647 (N_13647,N_8583,N_6558);
nor U13648 (N_13648,N_7093,N_5734);
or U13649 (N_13649,N_7092,N_6463);
nand U13650 (N_13650,N_5522,N_5616);
and U13651 (N_13651,N_6260,N_8237);
and U13652 (N_13652,N_6269,N_8814);
xor U13653 (N_13653,N_8140,N_7615);
or U13654 (N_13654,N_7816,N_8860);
and U13655 (N_13655,N_7121,N_8521);
nand U13656 (N_13656,N_8686,N_7302);
nand U13657 (N_13657,N_8786,N_6066);
or U13658 (N_13658,N_8156,N_9010);
and U13659 (N_13659,N_8009,N_5015);
or U13660 (N_13660,N_8109,N_5034);
and U13661 (N_13661,N_8298,N_9700);
and U13662 (N_13662,N_7830,N_5741);
or U13663 (N_13663,N_6603,N_5636);
nor U13664 (N_13664,N_5742,N_6521);
nand U13665 (N_13665,N_5085,N_8813);
nor U13666 (N_13666,N_9263,N_8778);
and U13667 (N_13667,N_5997,N_9525);
nor U13668 (N_13668,N_6370,N_9898);
nand U13669 (N_13669,N_6769,N_8646);
or U13670 (N_13670,N_8574,N_9992);
or U13671 (N_13671,N_9115,N_5584);
nor U13672 (N_13672,N_8496,N_8283);
nor U13673 (N_13673,N_7314,N_7204);
nand U13674 (N_13674,N_6546,N_6627);
or U13675 (N_13675,N_6446,N_5674);
nand U13676 (N_13676,N_6996,N_8331);
nand U13677 (N_13677,N_7535,N_5990);
nor U13678 (N_13678,N_5004,N_6499);
nor U13679 (N_13679,N_6369,N_9339);
nor U13680 (N_13680,N_5605,N_7766);
or U13681 (N_13681,N_7861,N_9322);
or U13682 (N_13682,N_8802,N_5127);
nor U13683 (N_13683,N_5857,N_8432);
or U13684 (N_13684,N_6494,N_7039);
nand U13685 (N_13685,N_9996,N_7720);
or U13686 (N_13686,N_5497,N_5576);
and U13687 (N_13687,N_9362,N_6694);
nand U13688 (N_13688,N_7130,N_9491);
nor U13689 (N_13689,N_5909,N_5044);
nand U13690 (N_13690,N_8226,N_6472);
or U13691 (N_13691,N_6395,N_9718);
or U13692 (N_13692,N_6092,N_8083);
nor U13693 (N_13693,N_7716,N_6026);
and U13694 (N_13694,N_7228,N_7374);
nor U13695 (N_13695,N_6267,N_7174);
and U13696 (N_13696,N_8735,N_5489);
nand U13697 (N_13697,N_8130,N_7307);
nor U13698 (N_13698,N_6217,N_5182);
or U13699 (N_13699,N_6408,N_8981);
nor U13700 (N_13700,N_8554,N_8228);
nand U13701 (N_13701,N_5791,N_8872);
and U13702 (N_13702,N_6306,N_6682);
or U13703 (N_13703,N_7612,N_6110);
and U13704 (N_13704,N_7713,N_6415);
nand U13705 (N_13705,N_8826,N_7903);
and U13706 (N_13706,N_5227,N_8635);
and U13707 (N_13707,N_5327,N_9199);
nor U13708 (N_13708,N_8130,N_9246);
nor U13709 (N_13709,N_5761,N_7623);
and U13710 (N_13710,N_8774,N_8258);
and U13711 (N_13711,N_8960,N_5125);
and U13712 (N_13712,N_5946,N_8580);
nor U13713 (N_13713,N_8167,N_6955);
and U13714 (N_13714,N_5561,N_9722);
nand U13715 (N_13715,N_5156,N_8980);
nor U13716 (N_13716,N_5601,N_5585);
nand U13717 (N_13717,N_6161,N_8211);
and U13718 (N_13718,N_9496,N_5249);
and U13719 (N_13719,N_9119,N_7580);
or U13720 (N_13720,N_9770,N_9985);
xnor U13721 (N_13721,N_6860,N_8271);
nand U13722 (N_13722,N_6752,N_8083);
and U13723 (N_13723,N_5993,N_7275);
and U13724 (N_13724,N_8684,N_5246);
and U13725 (N_13725,N_8033,N_9345);
or U13726 (N_13726,N_6132,N_9999);
or U13727 (N_13727,N_9133,N_5676);
nand U13728 (N_13728,N_8264,N_7821);
and U13729 (N_13729,N_7470,N_7684);
nand U13730 (N_13730,N_6144,N_9041);
nand U13731 (N_13731,N_5876,N_7672);
and U13732 (N_13732,N_6046,N_8395);
and U13733 (N_13733,N_9656,N_6149);
nor U13734 (N_13734,N_6419,N_8091);
or U13735 (N_13735,N_5351,N_9722);
or U13736 (N_13736,N_5618,N_6380);
nand U13737 (N_13737,N_7910,N_6333);
and U13738 (N_13738,N_9017,N_8912);
or U13739 (N_13739,N_9059,N_9844);
or U13740 (N_13740,N_8023,N_7701);
nor U13741 (N_13741,N_5966,N_7316);
or U13742 (N_13742,N_5981,N_5507);
nand U13743 (N_13743,N_8537,N_6636);
or U13744 (N_13744,N_5103,N_6168);
and U13745 (N_13745,N_6379,N_6184);
nand U13746 (N_13746,N_7524,N_7134);
nor U13747 (N_13747,N_9530,N_6169);
or U13748 (N_13748,N_5985,N_9183);
or U13749 (N_13749,N_6482,N_6875);
nand U13750 (N_13750,N_7352,N_6797);
nand U13751 (N_13751,N_6673,N_8695);
nand U13752 (N_13752,N_9605,N_8617);
nor U13753 (N_13753,N_8037,N_8867);
or U13754 (N_13754,N_6682,N_9089);
or U13755 (N_13755,N_8273,N_5621);
or U13756 (N_13756,N_7157,N_7393);
nor U13757 (N_13757,N_7514,N_6762);
and U13758 (N_13758,N_7668,N_5734);
nor U13759 (N_13759,N_8299,N_5993);
nand U13760 (N_13760,N_5365,N_9086);
nor U13761 (N_13761,N_9056,N_8941);
or U13762 (N_13762,N_6213,N_9798);
nor U13763 (N_13763,N_5884,N_9276);
nor U13764 (N_13764,N_7007,N_9912);
nor U13765 (N_13765,N_6339,N_6158);
or U13766 (N_13766,N_8740,N_9043);
and U13767 (N_13767,N_9113,N_7429);
or U13768 (N_13768,N_5489,N_6439);
or U13769 (N_13769,N_9969,N_6112);
nor U13770 (N_13770,N_6319,N_5808);
and U13771 (N_13771,N_6574,N_7249);
nand U13772 (N_13772,N_9343,N_6060);
nand U13773 (N_13773,N_8069,N_8965);
or U13774 (N_13774,N_9177,N_8441);
and U13775 (N_13775,N_9212,N_9413);
or U13776 (N_13776,N_6395,N_6785);
and U13777 (N_13777,N_7919,N_7072);
nand U13778 (N_13778,N_9331,N_8666);
or U13779 (N_13779,N_9614,N_8570);
nand U13780 (N_13780,N_8276,N_7714);
nand U13781 (N_13781,N_5850,N_8882);
or U13782 (N_13782,N_9641,N_7484);
nor U13783 (N_13783,N_6275,N_7074);
nor U13784 (N_13784,N_8757,N_5103);
or U13785 (N_13785,N_8044,N_6473);
nand U13786 (N_13786,N_7198,N_6283);
or U13787 (N_13787,N_8650,N_6455);
nand U13788 (N_13788,N_5174,N_5340);
nor U13789 (N_13789,N_9373,N_7612);
and U13790 (N_13790,N_7122,N_5755);
and U13791 (N_13791,N_6773,N_7703);
nor U13792 (N_13792,N_5234,N_7031);
and U13793 (N_13793,N_8518,N_7033);
nand U13794 (N_13794,N_9003,N_8565);
or U13795 (N_13795,N_6127,N_8229);
nand U13796 (N_13796,N_5480,N_5068);
or U13797 (N_13797,N_8899,N_8223);
nand U13798 (N_13798,N_7031,N_5085);
or U13799 (N_13799,N_6928,N_6914);
nand U13800 (N_13800,N_7892,N_9509);
nor U13801 (N_13801,N_8054,N_5171);
and U13802 (N_13802,N_6400,N_6498);
or U13803 (N_13803,N_6168,N_8627);
or U13804 (N_13804,N_8667,N_8619);
nand U13805 (N_13805,N_6406,N_8037);
and U13806 (N_13806,N_5114,N_5260);
and U13807 (N_13807,N_6728,N_7287);
nor U13808 (N_13808,N_7642,N_5930);
or U13809 (N_13809,N_6043,N_7584);
nor U13810 (N_13810,N_6731,N_6112);
and U13811 (N_13811,N_9291,N_6589);
or U13812 (N_13812,N_5751,N_9487);
and U13813 (N_13813,N_8462,N_6096);
nor U13814 (N_13814,N_5296,N_6229);
nand U13815 (N_13815,N_7925,N_7037);
or U13816 (N_13816,N_6270,N_6044);
and U13817 (N_13817,N_8871,N_7620);
nand U13818 (N_13818,N_8586,N_9102);
and U13819 (N_13819,N_6539,N_7393);
nor U13820 (N_13820,N_9213,N_9665);
and U13821 (N_13821,N_5073,N_8886);
nor U13822 (N_13822,N_7319,N_7039);
nor U13823 (N_13823,N_7029,N_7534);
nor U13824 (N_13824,N_6302,N_6775);
nor U13825 (N_13825,N_7798,N_9546);
and U13826 (N_13826,N_9563,N_8411);
nand U13827 (N_13827,N_8806,N_9827);
nor U13828 (N_13828,N_8581,N_9157);
and U13829 (N_13829,N_8645,N_7298);
nor U13830 (N_13830,N_8147,N_9289);
nand U13831 (N_13831,N_6813,N_5104);
or U13832 (N_13832,N_8343,N_6118);
or U13833 (N_13833,N_7287,N_7718);
nand U13834 (N_13834,N_6616,N_5656);
and U13835 (N_13835,N_6366,N_8857);
and U13836 (N_13836,N_8116,N_9534);
nor U13837 (N_13837,N_8694,N_5189);
nor U13838 (N_13838,N_8004,N_6855);
and U13839 (N_13839,N_5418,N_7643);
nor U13840 (N_13840,N_8865,N_5663);
nand U13841 (N_13841,N_5292,N_6943);
nor U13842 (N_13842,N_9968,N_5725);
nor U13843 (N_13843,N_7472,N_6758);
nor U13844 (N_13844,N_8155,N_5487);
or U13845 (N_13845,N_9130,N_5815);
nand U13846 (N_13846,N_5252,N_9807);
nand U13847 (N_13847,N_5302,N_8586);
nor U13848 (N_13848,N_7125,N_6666);
and U13849 (N_13849,N_6133,N_7456);
xnor U13850 (N_13850,N_9349,N_8000);
and U13851 (N_13851,N_8671,N_8565);
and U13852 (N_13852,N_6639,N_8473);
nand U13853 (N_13853,N_7819,N_8089);
nand U13854 (N_13854,N_7838,N_6014);
nor U13855 (N_13855,N_8698,N_8281);
or U13856 (N_13856,N_7308,N_9059);
and U13857 (N_13857,N_6749,N_9421);
or U13858 (N_13858,N_6088,N_5127);
nand U13859 (N_13859,N_6239,N_7188);
or U13860 (N_13860,N_9706,N_8457);
and U13861 (N_13861,N_9109,N_9222);
and U13862 (N_13862,N_5657,N_6765);
nor U13863 (N_13863,N_6087,N_7531);
nand U13864 (N_13864,N_5716,N_7785);
nor U13865 (N_13865,N_6263,N_6146);
and U13866 (N_13866,N_7169,N_9600);
nand U13867 (N_13867,N_7763,N_5819);
or U13868 (N_13868,N_6113,N_6550);
and U13869 (N_13869,N_5366,N_7918);
and U13870 (N_13870,N_9236,N_7693);
or U13871 (N_13871,N_6698,N_5372);
or U13872 (N_13872,N_8084,N_7157);
nand U13873 (N_13873,N_6993,N_7323);
nor U13874 (N_13874,N_9404,N_5095);
xor U13875 (N_13875,N_8045,N_9548);
nor U13876 (N_13876,N_5717,N_8685);
and U13877 (N_13877,N_8263,N_6699);
nand U13878 (N_13878,N_5064,N_9789);
nor U13879 (N_13879,N_6774,N_8122);
nor U13880 (N_13880,N_8758,N_7390);
nand U13881 (N_13881,N_8569,N_7045);
or U13882 (N_13882,N_7776,N_5189);
nand U13883 (N_13883,N_8205,N_6323);
and U13884 (N_13884,N_8431,N_9488);
or U13885 (N_13885,N_8293,N_5926);
and U13886 (N_13886,N_9155,N_7389);
nor U13887 (N_13887,N_7239,N_7937);
and U13888 (N_13888,N_8271,N_9535);
or U13889 (N_13889,N_8646,N_7169);
and U13890 (N_13890,N_6204,N_5903);
or U13891 (N_13891,N_9859,N_5615);
nor U13892 (N_13892,N_6875,N_7144);
or U13893 (N_13893,N_7279,N_7164);
nand U13894 (N_13894,N_9446,N_7395);
or U13895 (N_13895,N_5851,N_6665);
and U13896 (N_13896,N_5247,N_8821);
and U13897 (N_13897,N_9588,N_7267);
nand U13898 (N_13898,N_8359,N_5261);
or U13899 (N_13899,N_5273,N_9742);
nand U13900 (N_13900,N_5362,N_5981);
nor U13901 (N_13901,N_8885,N_7021);
nor U13902 (N_13902,N_5758,N_7246);
nor U13903 (N_13903,N_6241,N_5858);
and U13904 (N_13904,N_8539,N_7265);
or U13905 (N_13905,N_9357,N_7579);
nor U13906 (N_13906,N_8834,N_9801);
nor U13907 (N_13907,N_7780,N_5080);
nor U13908 (N_13908,N_9327,N_5726);
and U13909 (N_13909,N_5367,N_6639);
nor U13910 (N_13910,N_7529,N_5064);
and U13911 (N_13911,N_8824,N_6742);
nand U13912 (N_13912,N_7040,N_6237);
and U13913 (N_13913,N_7197,N_6496);
or U13914 (N_13914,N_8256,N_6285);
and U13915 (N_13915,N_6896,N_8974);
nand U13916 (N_13916,N_9754,N_5918);
nand U13917 (N_13917,N_9777,N_9938);
nand U13918 (N_13918,N_5088,N_9602);
nor U13919 (N_13919,N_9310,N_5789);
or U13920 (N_13920,N_8523,N_6617);
or U13921 (N_13921,N_5715,N_6519);
or U13922 (N_13922,N_7594,N_9681);
or U13923 (N_13923,N_5583,N_9165);
nor U13924 (N_13924,N_7263,N_5220);
and U13925 (N_13925,N_7162,N_9126);
nand U13926 (N_13926,N_9025,N_6238);
and U13927 (N_13927,N_5960,N_7478);
and U13928 (N_13928,N_5572,N_7075);
or U13929 (N_13929,N_8780,N_7094);
and U13930 (N_13930,N_7619,N_9460);
or U13931 (N_13931,N_6787,N_7110);
nor U13932 (N_13932,N_5587,N_5178);
nor U13933 (N_13933,N_8041,N_9708);
nor U13934 (N_13934,N_5056,N_6047);
nor U13935 (N_13935,N_7119,N_8668);
or U13936 (N_13936,N_5169,N_5851);
and U13937 (N_13937,N_6299,N_6235);
or U13938 (N_13938,N_9457,N_8628);
and U13939 (N_13939,N_7064,N_5452);
nor U13940 (N_13940,N_5137,N_9597);
nor U13941 (N_13941,N_8915,N_6709);
nand U13942 (N_13942,N_8428,N_5680);
and U13943 (N_13943,N_8508,N_5217);
nor U13944 (N_13944,N_8416,N_8558);
nand U13945 (N_13945,N_9058,N_7637);
nand U13946 (N_13946,N_7000,N_5270);
nand U13947 (N_13947,N_9852,N_8909);
nand U13948 (N_13948,N_5898,N_6846);
nor U13949 (N_13949,N_9313,N_8193);
nor U13950 (N_13950,N_7327,N_9236);
nand U13951 (N_13951,N_9372,N_7982);
and U13952 (N_13952,N_5392,N_9104);
nor U13953 (N_13953,N_5933,N_8138);
nand U13954 (N_13954,N_7236,N_6609);
nor U13955 (N_13955,N_7178,N_9165);
or U13956 (N_13956,N_6870,N_6510);
nor U13957 (N_13957,N_6435,N_6677);
nor U13958 (N_13958,N_5624,N_7019);
nor U13959 (N_13959,N_9949,N_8732);
and U13960 (N_13960,N_9932,N_7648);
and U13961 (N_13961,N_8467,N_7502);
nor U13962 (N_13962,N_6872,N_9079);
nand U13963 (N_13963,N_6259,N_7053);
or U13964 (N_13964,N_6791,N_8223);
nand U13965 (N_13965,N_6556,N_7258);
nand U13966 (N_13966,N_8911,N_7689);
and U13967 (N_13967,N_5163,N_9508);
nand U13968 (N_13968,N_8805,N_9832);
nor U13969 (N_13969,N_6205,N_6721);
nor U13970 (N_13970,N_5391,N_8768);
or U13971 (N_13971,N_5498,N_9698);
nor U13972 (N_13972,N_5000,N_5958);
and U13973 (N_13973,N_5392,N_9365);
nand U13974 (N_13974,N_8830,N_5548);
and U13975 (N_13975,N_9876,N_9306);
nand U13976 (N_13976,N_7034,N_9822);
or U13977 (N_13977,N_8911,N_8507);
nor U13978 (N_13978,N_8584,N_9086);
or U13979 (N_13979,N_7724,N_7722);
or U13980 (N_13980,N_9831,N_8496);
and U13981 (N_13981,N_8974,N_8426);
or U13982 (N_13982,N_6287,N_6892);
nor U13983 (N_13983,N_6602,N_8591);
nor U13984 (N_13984,N_6190,N_7000);
nor U13985 (N_13985,N_9290,N_9049);
and U13986 (N_13986,N_8349,N_5802);
nor U13987 (N_13987,N_9687,N_7345);
or U13988 (N_13988,N_5646,N_7131);
nand U13989 (N_13989,N_5700,N_6261);
or U13990 (N_13990,N_5019,N_8195);
nor U13991 (N_13991,N_9128,N_6648);
or U13992 (N_13992,N_5925,N_6038);
and U13993 (N_13993,N_8415,N_6768);
or U13994 (N_13994,N_8924,N_7827);
and U13995 (N_13995,N_6726,N_5948);
or U13996 (N_13996,N_6586,N_9394);
nand U13997 (N_13997,N_9305,N_7179);
nand U13998 (N_13998,N_8611,N_8178);
nor U13999 (N_13999,N_9384,N_7904);
and U14000 (N_14000,N_8173,N_6219);
and U14001 (N_14001,N_6430,N_8812);
nor U14002 (N_14002,N_7784,N_8125);
or U14003 (N_14003,N_8852,N_7650);
or U14004 (N_14004,N_8837,N_5180);
and U14005 (N_14005,N_6807,N_6870);
and U14006 (N_14006,N_8790,N_8753);
and U14007 (N_14007,N_9285,N_6705);
nand U14008 (N_14008,N_6034,N_6445);
and U14009 (N_14009,N_8956,N_5208);
or U14010 (N_14010,N_7765,N_5710);
or U14011 (N_14011,N_5429,N_8309);
or U14012 (N_14012,N_6242,N_6512);
nor U14013 (N_14013,N_8215,N_9917);
nand U14014 (N_14014,N_5727,N_9203);
and U14015 (N_14015,N_8148,N_7943);
and U14016 (N_14016,N_9798,N_6235);
nand U14017 (N_14017,N_7741,N_8812);
or U14018 (N_14018,N_6954,N_6028);
and U14019 (N_14019,N_8517,N_8472);
nor U14020 (N_14020,N_6651,N_5286);
and U14021 (N_14021,N_8590,N_9567);
nor U14022 (N_14022,N_5706,N_9049);
or U14023 (N_14023,N_9224,N_8820);
nand U14024 (N_14024,N_5108,N_8002);
xnor U14025 (N_14025,N_6201,N_5368);
nor U14026 (N_14026,N_7639,N_9867);
or U14027 (N_14027,N_6622,N_8978);
nor U14028 (N_14028,N_9840,N_6062);
and U14029 (N_14029,N_7757,N_9517);
and U14030 (N_14030,N_6160,N_5941);
nor U14031 (N_14031,N_9207,N_9513);
or U14032 (N_14032,N_7551,N_8479);
nor U14033 (N_14033,N_7927,N_6464);
nand U14034 (N_14034,N_8755,N_9495);
or U14035 (N_14035,N_9502,N_8261);
nand U14036 (N_14036,N_9301,N_5643);
nor U14037 (N_14037,N_9502,N_9139);
nand U14038 (N_14038,N_9839,N_8349);
nand U14039 (N_14039,N_7963,N_9152);
or U14040 (N_14040,N_8901,N_7565);
or U14041 (N_14041,N_9752,N_6901);
nor U14042 (N_14042,N_9486,N_8752);
nand U14043 (N_14043,N_8788,N_6830);
nor U14044 (N_14044,N_7603,N_9141);
and U14045 (N_14045,N_5551,N_7596);
and U14046 (N_14046,N_6126,N_9677);
and U14047 (N_14047,N_8557,N_8305);
or U14048 (N_14048,N_5134,N_8931);
nor U14049 (N_14049,N_7707,N_9954);
nor U14050 (N_14050,N_7411,N_7598);
or U14051 (N_14051,N_5454,N_9742);
or U14052 (N_14052,N_5722,N_5992);
nor U14053 (N_14053,N_9302,N_6900);
or U14054 (N_14054,N_9645,N_5001);
nand U14055 (N_14055,N_6577,N_7257);
and U14056 (N_14056,N_6614,N_5854);
or U14057 (N_14057,N_8546,N_7742);
nor U14058 (N_14058,N_9168,N_5676);
or U14059 (N_14059,N_5249,N_9275);
nand U14060 (N_14060,N_7999,N_9452);
nand U14061 (N_14061,N_7929,N_7111);
or U14062 (N_14062,N_6785,N_7794);
nand U14063 (N_14063,N_8470,N_6296);
nand U14064 (N_14064,N_8036,N_8250);
or U14065 (N_14065,N_8996,N_7778);
nor U14066 (N_14066,N_5762,N_9055);
nand U14067 (N_14067,N_9361,N_5956);
nor U14068 (N_14068,N_7626,N_6371);
nor U14069 (N_14069,N_7748,N_8505);
or U14070 (N_14070,N_8539,N_8999);
or U14071 (N_14071,N_8563,N_9847);
or U14072 (N_14072,N_8111,N_5958);
nand U14073 (N_14073,N_8244,N_6597);
nor U14074 (N_14074,N_9288,N_7826);
and U14075 (N_14075,N_7627,N_8981);
nor U14076 (N_14076,N_6098,N_6613);
and U14077 (N_14077,N_7265,N_8470);
and U14078 (N_14078,N_6715,N_6725);
nand U14079 (N_14079,N_6547,N_5050);
nor U14080 (N_14080,N_7035,N_8931);
and U14081 (N_14081,N_9494,N_6472);
nand U14082 (N_14082,N_7117,N_9477);
and U14083 (N_14083,N_9294,N_8816);
and U14084 (N_14084,N_5811,N_9813);
nor U14085 (N_14085,N_9681,N_9674);
or U14086 (N_14086,N_7825,N_6726);
or U14087 (N_14087,N_9101,N_5527);
or U14088 (N_14088,N_7026,N_8436);
or U14089 (N_14089,N_7479,N_5618);
nor U14090 (N_14090,N_7693,N_7338);
or U14091 (N_14091,N_8715,N_5465);
and U14092 (N_14092,N_5421,N_8319);
nand U14093 (N_14093,N_9291,N_5845);
nor U14094 (N_14094,N_8118,N_9853);
xnor U14095 (N_14095,N_7150,N_5086);
nor U14096 (N_14096,N_9721,N_6379);
and U14097 (N_14097,N_8220,N_8328);
nand U14098 (N_14098,N_7205,N_6106);
nand U14099 (N_14099,N_9684,N_9948);
nor U14100 (N_14100,N_9681,N_8622);
nand U14101 (N_14101,N_8225,N_7709);
nor U14102 (N_14102,N_9949,N_6485);
nand U14103 (N_14103,N_7183,N_6643);
nor U14104 (N_14104,N_7164,N_9908);
or U14105 (N_14105,N_5882,N_6024);
and U14106 (N_14106,N_7493,N_8773);
nand U14107 (N_14107,N_8919,N_8246);
and U14108 (N_14108,N_7536,N_8684);
or U14109 (N_14109,N_6658,N_8387);
nand U14110 (N_14110,N_5311,N_9811);
and U14111 (N_14111,N_7631,N_5639);
or U14112 (N_14112,N_6477,N_9843);
nor U14113 (N_14113,N_6789,N_6248);
nand U14114 (N_14114,N_6393,N_9900);
or U14115 (N_14115,N_6507,N_5121);
and U14116 (N_14116,N_7853,N_6908);
and U14117 (N_14117,N_6768,N_6291);
nand U14118 (N_14118,N_8110,N_9462);
nor U14119 (N_14119,N_9845,N_7864);
nand U14120 (N_14120,N_6556,N_9034);
and U14121 (N_14121,N_7529,N_5235);
or U14122 (N_14122,N_9562,N_9201);
nor U14123 (N_14123,N_5258,N_5131);
and U14124 (N_14124,N_5726,N_5674);
nor U14125 (N_14125,N_5993,N_8846);
and U14126 (N_14126,N_7902,N_9850);
nand U14127 (N_14127,N_5944,N_9813);
or U14128 (N_14128,N_8462,N_7422);
and U14129 (N_14129,N_5370,N_8687);
nand U14130 (N_14130,N_9793,N_6097);
nand U14131 (N_14131,N_9834,N_7467);
and U14132 (N_14132,N_6264,N_9491);
nand U14133 (N_14133,N_7261,N_6923);
and U14134 (N_14134,N_8508,N_7912);
or U14135 (N_14135,N_6277,N_9432);
nor U14136 (N_14136,N_9943,N_5894);
and U14137 (N_14137,N_7111,N_6157);
nand U14138 (N_14138,N_7279,N_8187);
nand U14139 (N_14139,N_9501,N_7428);
nor U14140 (N_14140,N_9623,N_5610);
nor U14141 (N_14141,N_5745,N_8558);
and U14142 (N_14142,N_8043,N_6563);
and U14143 (N_14143,N_9187,N_9007);
and U14144 (N_14144,N_8247,N_8316);
or U14145 (N_14145,N_7075,N_9802);
nor U14146 (N_14146,N_9224,N_8077);
and U14147 (N_14147,N_9684,N_6980);
nand U14148 (N_14148,N_9371,N_6409);
and U14149 (N_14149,N_6706,N_5158);
nand U14150 (N_14150,N_6549,N_8826);
nor U14151 (N_14151,N_8081,N_7332);
or U14152 (N_14152,N_9770,N_6274);
nand U14153 (N_14153,N_8939,N_8523);
nand U14154 (N_14154,N_5941,N_5962);
and U14155 (N_14155,N_8257,N_9812);
nor U14156 (N_14156,N_8037,N_7931);
nand U14157 (N_14157,N_9033,N_8764);
or U14158 (N_14158,N_5959,N_7031);
nor U14159 (N_14159,N_6620,N_8901);
nand U14160 (N_14160,N_8380,N_6719);
or U14161 (N_14161,N_6976,N_9972);
nor U14162 (N_14162,N_9538,N_6489);
or U14163 (N_14163,N_6709,N_8757);
or U14164 (N_14164,N_7781,N_7617);
nor U14165 (N_14165,N_7918,N_6640);
or U14166 (N_14166,N_9711,N_6905);
nor U14167 (N_14167,N_7690,N_9095);
nor U14168 (N_14168,N_9336,N_6798);
nor U14169 (N_14169,N_5984,N_7240);
or U14170 (N_14170,N_5625,N_6434);
and U14171 (N_14171,N_7591,N_9603);
nand U14172 (N_14172,N_7786,N_9301);
and U14173 (N_14173,N_8336,N_8327);
nor U14174 (N_14174,N_6900,N_7844);
and U14175 (N_14175,N_8838,N_5701);
and U14176 (N_14176,N_9237,N_8688);
and U14177 (N_14177,N_6417,N_8435);
or U14178 (N_14178,N_6548,N_5318);
nand U14179 (N_14179,N_7113,N_6167);
nor U14180 (N_14180,N_7566,N_5020);
nand U14181 (N_14181,N_6799,N_9224);
and U14182 (N_14182,N_9415,N_5998);
and U14183 (N_14183,N_7655,N_8239);
nand U14184 (N_14184,N_5779,N_9114);
nand U14185 (N_14185,N_7420,N_8079);
nor U14186 (N_14186,N_6705,N_8482);
nor U14187 (N_14187,N_6332,N_8365);
or U14188 (N_14188,N_9374,N_7156);
nand U14189 (N_14189,N_6623,N_8587);
or U14190 (N_14190,N_9334,N_9434);
and U14191 (N_14191,N_5639,N_7608);
and U14192 (N_14192,N_5997,N_9880);
xnor U14193 (N_14193,N_6926,N_6286);
or U14194 (N_14194,N_5501,N_7406);
nand U14195 (N_14195,N_5166,N_9519);
nand U14196 (N_14196,N_7139,N_9833);
or U14197 (N_14197,N_6824,N_6625);
nand U14198 (N_14198,N_7873,N_9005);
nand U14199 (N_14199,N_5093,N_7521);
and U14200 (N_14200,N_8157,N_9995);
nand U14201 (N_14201,N_8632,N_6218);
and U14202 (N_14202,N_8368,N_8868);
nor U14203 (N_14203,N_7996,N_7398);
or U14204 (N_14204,N_8517,N_6627);
nor U14205 (N_14205,N_5804,N_6429);
nor U14206 (N_14206,N_5513,N_5889);
nor U14207 (N_14207,N_9560,N_5171);
and U14208 (N_14208,N_9262,N_7680);
or U14209 (N_14209,N_9123,N_7417);
nor U14210 (N_14210,N_9308,N_6717);
nor U14211 (N_14211,N_9187,N_9805);
nand U14212 (N_14212,N_5519,N_6730);
and U14213 (N_14213,N_9513,N_6494);
nor U14214 (N_14214,N_6726,N_6460);
nand U14215 (N_14215,N_6090,N_6880);
nand U14216 (N_14216,N_7018,N_8961);
nand U14217 (N_14217,N_8325,N_9647);
nand U14218 (N_14218,N_8210,N_6600);
nor U14219 (N_14219,N_8628,N_8222);
nand U14220 (N_14220,N_8255,N_5389);
or U14221 (N_14221,N_5019,N_7862);
nand U14222 (N_14222,N_5254,N_6605);
nor U14223 (N_14223,N_5423,N_8441);
and U14224 (N_14224,N_6887,N_5945);
nand U14225 (N_14225,N_8780,N_6397);
nand U14226 (N_14226,N_9740,N_8774);
nand U14227 (N_14227,N_5409,N_9254);
nand U14228 (N_14228,N_8589,N_9592);
nor U14229 (N_14229,N_6833,N_5449);
nand U14230 (N_14230,N_8088,N_9152);
nor U14231 (N_14231,N_9131,N_7174);
nand U14232 (N_14232,N_6391,N_6584);
and U14233 (N_14233,N_8022,N_9377);
nor U14234 (N_14234,N_8886,N_7657);
nand U14235 (N_14235,N_7283,N_7708);
and U14236 (N_14236,N_5305,N_5909);
nand U14237 (N_14237,N_6684,N_6121);
and U14238 (N_14238,N_6172,N_5548);
nor U14239 (N_14239,N_5412,N_9101);
nand U14240 (N_14240,N_9367,N_9994);
nor U14241 (N_14241,N_6371,N_7310);
nor U14242 (N_14242,N_8381,N_5468);
and U14243 (N_14243,N_8313,N_6676);
or U14244 (N_14244,N_8186,N_7505);
or U14245 (N_14245,N_7575,N_8803);
or U14246 (N_14246,N_7748,N_9641);
nand U14247 (N_14247,N_8768,N_8602);
nor U14248 (N_14248,N_7371,N_6864);
and U14249 (N_14249,N_5587,N_8481);
and U14250 (N_14250,N_6997,N_6705);
nand U14251 (N_14251,N_8356,N_8246);
and U14252 (N_14252,N_9359,N_9730);
or U14253 (N_14253,N_7670,N_7284);
nor U14254 (N_14254,N_6286,N_7565);
nor U14255 (N_14255,N_8242,N_7344);
nor U14256 (N_14256,N_8745,N_8757);
nand U14257 (N_14257,N_8043,N_7000);
and U14258 (N_14258,N_5014,N_8409);
nor U14259 (N_14259,N_6597,N_9989);
nand U14260 (N_14260,N_6520,N_9744);
and U14261 (N_14261,N_9820,N_9342);
and U14262 (N_14262,N_7030,N_5994);
nand U14263 (N_14263,N_5412,N_7625);
or U14264 (N_14264,N_6343,N_9864);
or U14265 (N_14265,N_5453,N_9261);
nor U14266 (N_14266,N_8352,N_5670);
or U14267 (N_14267,N_7307,N_8399);
nand U14268 (N_14268,N_9281,N_5373);
and U14269 (N_14269,N_9561,N_5138);
nand U14270 (N_14270,N_8053,N_9412);
or U14271 (N_14271,N_5305,N_5715);
nand U14272 (N_14272,N_5468,N_6742);
nor U14273 (N_14273,N_7121,N_9594);
or U14274 (N_14274,N_5796,N_8817);
or U14275 (N_14275,N_6560,N_9880);
nand U14276 (N_14276,N_9997,N_7128);
and U14277 (N_14277,N_8369,N_6325);
or U14278 (N_14278,N_9246,N_6372);
and U14279 (N_14279,N_7665,N_6642);
nand U14280 (N_14280,N_8071,N_7495);
and U14281 (N_14281,N_8916,N_6090);
nand U14282 (N_14282,N_9380,N_9522);
or U14283 (N_14283,N_5268,N_6418);
nor U14284 (N_14284,N_8529,N_6069);
or U14285 (N_14285,N_6259,N_6412);
nand U14286 (N_14286,N_7114,N_6495);
nand U14287 (N_14287,N_6775,N_5322);
or U14288 (N_14288,N_8801,N_6011);
nor U14289 (N_14289,N_5839,N_9406);
xnor U14290 (N_14290,N_6732,N_8668);
and U14291 (N_14291,N_5289,N_5287);
nand U14292 (N_14292,N_5016,N_5118);
nor U14293 (N_14293,N_5769,N_7809);
or U14294 (N_14294,N_8655,N_6088);
nor U14295 (N_14295,N_9644,N_6037);
or U14296 (N_14296,N_6574,N_5992);
nor U14297 (N_14297,N_5016,N_6944);
nor U14298 (N_14298,N_6848,N_5970);
or U14299 (N_14299,N_6326,N_5333);
nor U14300 (N_14300,N_7461,N_9104);
or U14301 (N_14301,N_6450,N_8450);
or U14302 (N_14302,N_6539,N_5953);
nand U14303 (N_14303,N_5954,N_6362);
nand U14304 (N_14304,N_5731,N_5875);
and U14305 (N_14305,N_8374,N_6484);
or U14306 (N_14306,N_7145,N_6697);
nor U14307 (N_14307,N_9036,N_7953);
or U14308 (N_14308,N_9617,N_5138);
and U14309 (N_14309,N_7599,N_5226);
or U14310 (N_14310,N_5844,N_5659);
nor U14311 (N_14311,N_9549,N_5773);
and U14312 (N_14312,N_8254,N_6722);
nand U14313 (N_14313,N_5310,N_8934);
or U14314 (N_14314,N_9560,N_9588);
or U14315 (N_14315,N_7614,N_6193);
nand U14316 (N_14316,N_5119,N_5653);
nand U14317 (N_14317,N_5114,N_8195);
or U14318 (N_14318,N_9337,N_8929);
nand U14319 (N_14319,N_7733,N_5829);
nor U14320 (N_14320,N_6130,N_8819);
xnor U14321 (N_14321,N_7526,N_7762);
nand U14322 (N_14322,N_5464,N_7752);
nand U14323 (N_14323,N_9025,N_6429);
and U14324 (N_14324,N_6556,N_6937);
or U14325 (N_14325,N_7299,N_8278);
and U14326 (N_14326,N_5832,N_5000);
and U14327 (N_14327,N_6799,N_7695);
nor U14328 (N_14328,N_7576,N_9021);
and U14329 (N_14329,N_5480,N_8194);
nor U14330 (N_14330,N_8452,N_6078);
and U14331 (N_14331,N_6799,N_7040);
or U14332 (N_14332,N_5753,N_9613);
or U14333 (N_14333,N_9499,N_8149);
nor U14334 (N_14334,N_5059,N_5483);
or U14335 (N_14335,N_6701,N_6269);
nand U14336 (N_14336,N_7162,N_6032);
and U14337 (N_14337,N_5288,N_5592);
or U14338 (N_14338,N_9432,N_6860);
nor U14339 (N_14339,N_7266,N_5144);
nor U14340 (N_14340,N_8751,N_5661);
or U14341 (N_14341,N_5133,N_5131);
nor U14342 (N_14342,N_8373,N_6336);
nor U14343 (N_14343,N_8237,N_8419);
nor U14344 (N_14344,N_7253,N_8944);
or U14345 (N_14345,N_5216,N_5717);
and U14346 (N_14346,N_8479,N_6729);
nor U14347 (N_14347,N_6056,N_6581);
or U14348 (N_14348,N_6709,N_5442);
nor U14349 (N_14349,N_7604,N_8791);
and U14350 (N_14350,N_8110,N_8106);
nand U14351 (N_14351,N_6828,N_5840);
nand U14352 (N_14352,N_5364,N_7335);
nand U14353 (N_14353,N_7762,N_6244);
and U14354 (N_14354,N_6016,N_8979);
or U14355 (N_14355,N_6041,N_8344);
or U14356 (N_14356,N_6172,N_5877);
nor U14357 (N_14357,N_7960,N_5925);
nand U14358 (N_14358,N_7018,N_7741);
or U14359 (N_14359,N_8000,N_6860);
and U14360 (N_14360,N_6288,N_8516);
nand U14361 (N_14361,N_6443,N_8274);
or U14362 (N_14362,N_5764,N_5963);
nor U14363 (N_14363,N_6367,N_8335);
or U14364 (N_14364,N_5211,N_6792);
nand U14365 (N_14365,N_5487,N_8624);
nand U14366 (N_14366,N_6978,N_7524);
and U14367 (N_14367,N_9446,N_6640);
nor U14368 (N_14368,N_8641,N_9179);
and U14369 (N_14369,N_8024,N_7015);
and U14370 (N_14370,N_9885,N_6316);
nor U14371 (N_14371,N_7155,N_6891);
nand U14372 (N_14372,N_7318,N_7342);
nor U14373 (N_14373,N_8352,N_6178);
nand U14374 (N_14374,N_5061,N_5222);
and U14375 (N_14375,N_7544,N_9335);
or U14376 (N_14376,N_9556,N_9296);
or U14377 (N_14377,N_6725,N_7068);
nand U14378 (N_14378,N_9529,N_5930);
or U14379 (N_14379,N_9071,N_8783);
nand U14380 (N_14380,N_7304,N_9756);
or U14381 (N_14381,N_9525,N_8609);
or U14382 (N_14382,N_5621,N_7090);
nand U14383 (N_14383,N_7773,N_5309);
or U14384 (N_14384,N_8914,N_8007);
nor U14385 (N_14385,N_7990,N_7470);
or U14386 (N_14386,N_9831,N_5776);
nand U14387 (N_14387,N_9893,N_7411);
nor U14388 (N_14388,N_5338,N_7601);
nor U14389 (N_14389,N_8329,N_7330);
nand U14390 (N_14390,N_5309,N_5487);
nand U14391 (N_14391,N_6194,N_9631);
or U14392 (N_14392,N_5084,N_5024);
nand U14393 (N_14393,N_8330,N_9121);
or U14394 (N_14394,N_7334,N_9086);
nor U14395 (N_14395,N_7124,N_6153);
and U14396 (N_14396,N_6344,N_6007);
nand U14397 (N_14397,N_9833,N_5055);
nand U14398 (N_14398,N_5157,N_5999);
or U14399 (N_14399,N_9691,N_5514);
or U14400 (N_14400,N_9804,N_6492);
and U14401 (N_14401,N_9166,N_8690);
or U14402 (N_14402,N_6943,N_6537);
nor U14403 (N_14403,N_9387,N_5439);
nand U14404 (N_14404,N_7803,N_9073);
nor U14405 (N_14405,N_9442,N_6688);
and U14406 (N_14406,N_5264,N_6568);
or U14407 (N_14407,N_9293,N_8071);
and U14408 (N_14408,N_5232,N_9351);
and U14409 (N_14409,N_9551,N_5064);
nor U14410 (N_14410,N_7219,N_8829);
nor U14411 (N_14411,N_7792,N_7891);
nor U14412 (N_14412,N_8987,N_8575);
or U14413 (N_14413,N_8811,N_6549);
and U14414 (N_14414,N_6901,N_6538);
nor U14415 (N_14415,N_8535,N_8234);
and U14416 (N_14416,N_6197,N_7607);
or U14417 (N_14417,N_9816,N_7876);
or U14418 (N_14418,N_8481,N_9608);
nand U14419 (N_14419,N_6079,N_6704);
nor U14420 (N_14420,N_9218,N_8166);
and U14421 (N_14421,N_5499,N_7109);
nand U14422 (N_14422,N_7859,N_9757);
or U14423 (N_14423,N_7102,N_7980);
xor U14424 (N_14424,N_9738,N_6943);
nand U14425 (N_14425,N_7200,N_7851);
nor U14426 (N_14426,N_6110,N_5091);
and U14427 (N_14427,N_5338,N_7849);
or U14428 (N_14428,N_5122,N_7830);
nor U14429 (N_14429,N_5885,N_7058);
nor U14430 (N_14430,N_9559,N_5171);
nand U14431 (N_14431,N_5065,N_8597);
xnor U14432 (N_14432,N_7627,N_9545);
nand U14433 (N_14433,N_8252,N_7339);
nor U14434 (N_14434,N_7536,N_6251);
or U14435 (N_14435,N_5744,N_8475);
nand U14436 (N_14436,N_9182,N_8248);
nor U14437 (N_14437,N_5111,N_7784);
nor U14438 (N_14438,N_6264,N_6260);
nor U14439 (N_14439,N_6796,N_5392);
xnor U14440 (N_14440,N_6295,N_7518);
or U14441 (N_14441,N_8820,N_8129);
or U14442 (N_14442,N_6739,N_8182);
or U14443 (N_14443,N_5663,N_9948);
nor U14444 (N_14444,N_6476,N_7320);
nand U14445 (N_14445,N_9818,N_9759);
nor U14446 (N_14446,N_6201,N_7074);
nor U14447 (N_14447,N_6639,N_5671);
nor U14448 (N_14448,N_6867,N_6306);
nor U14449 (N_14449,N_6214,N_5743);
or U14450 (N_14450,N_7716,N_7175);
and U14451 (N_14451,N_6673,N_9133);
nor U14452 (N_14452,N_8305,N_6044);
or U14453 (N_14453,N_6461,N_9045);
or U14454 (N_14454,N_5692,N_7998);
nand U14455 (N_14455,N_5572,N_6133);
nand U14456 (N_14456,N_5195,N_9610);
or U14457 (N_14457,N_8148,N_6232);
nand U14458 (N_14458,N_7320,N_7560);
or U14459 (N_14459,N_5214,N_7133);
nor U14460 (N_14460,N_7436,N_8721);
nor U14461 (N_14461,N_5230,N_7005);
nor U14462 (N_14462,N_7194,N_8253);
or U14463 (N_14463,N_5357,N_6397);
nor U14464 (N_14464,N_7248,N_7594);
and U14465 (N_14465,N_8142,N_9477);
nand U14466 (N_14466,N_6808,N_6228);
nand U14467 (N_14467,N_7291,N_9272);
nand U14468 (N_14468,N_8529,N_8668);
nor U14469 (N_14469,N_6534,N_7379);
nand U14470 (N_14470,N_7396,N_8480);
and U14471 (N_14471,N_7618,N_7905);
or U14472 (N_14472,N_9370,N_5515);
or U14473 (N_14473,N_8645,N_7401);
nand U14474 (N_14474,N_6916,N_7181);
nor U14475 (N_14475,N_5309,N_8414);
nor U14476 (N_14476,N_7161,N_6872);
and U14477 (N_14477,N_7041,N_6236);
nand U14478 (N_14478,N_8358,N_5441);
nor U14479 (N_14479,N_9043,N_9818);
or U14480 (N_14480,N_8595,N_5198);
nand U14481 (N_14481,N_9989,N_6368);
and U14482 (N_14482,N_6489,N_8231);
nor U14483 (N_14483,N_6193,N_7885);
xor U14484 (N_14484,N_5829,N_8137);
nor U14485 (N_14485,N_5115,N_8010);
and U14486 (N_14486,N_5492,N_7648);
nor U14487 (N_14487,N_8911,N_8664);
nor U14488 (N_14488,N_6538,N_9803);
and U14489 (N_14489,N_6282,N_9844);
and U14490 (N_14490,N_6631,N_8706);
and U14491 (N_14491,N_5929,N_8571);
and U14492 (N_14492,N_8645,N_5634);
nand U14493 (N_14493,N_6096,N_5691);
and U14494 (N_14494,N_9012,N_5215);
nand U14495 (N_14495,N_8976,N_6618);
or U14496 (N_14496,N_6969,N_7690);
or U14497 (N_14497,N_9839,N_8918);
nand U14498 (N_14498,N_9361,N_5054);
nor U14499 (N_14499,N_7048,N_8462);
nor U14500 (N_14500,N_6181,N_6592);
nor U14501 (N_14501,N_9823,N_8463);
nor U14502 (N_14502,N_9055,N_9028);
nor U14503 (N_14503,N_8459,N_6872);
nor U14504 (N_14504,N_5827,N_5433);
and U14505 (N_14505,N_7264,N_9796);
nand U14506 (N_14506,N_9465,N_8401);
nor U14507 (N_14507,N_6390,N_9496);
nor U14508 (N_14508,N_9591,N_6005);
nor U14509 (N_14509,N_5059,N_5247);
nand U14510 (N_14510,N_5927,N_9193);
nor U14511 (N_14511,N_9978,N_7405);
nor U14512 (N_14512,N_8092,N_8750);
or U14513 (N_14513,N_9454,N_7438);
nand U14514 (N_14514,N_9697,N_7462);
nor U14515 (N_14515,N_6719,N_9102);
nor U14516 (N_14516,N_6577,N_7152);
nand U14517 (N_14517,N_5638,N_6070);
or U14518 (N_14518,N_9554,N_7537);
nand U14519 (N_14519,N_5157,N_7114);
and U14520 (N_14520,N_8731,N_8199);
and U14521 (N_14521,N_7069,N_7257);
nor U14522 (N_14522,N_5857,N_8621);
or U14523 (N_14523,N_7776,N_6651);
or U14524 (N_14524,N_9197,N_5491);
nor U14525 (N_14525,N_6095,N_8674);
nand U14526 (N_14526,N_9685,N_5748);
nand U14527 (N_14527,N_9060,N_5026);
nor U14528 (N_14528,N_7470,N_9152);
nand U14529 (N_14529,N_7098,N_9090);
and U14530 (N_14530,N_5058,N_6922);
or U14531 (N_14531,N_5215,N_9073);
nand U14532 (N_14532,N_7382,N_7769);
and U14533 (N_14533,N_8885,N_8044);
nand U14534 (N_14534,N_8687,N_8298);
nor U14535 (N_14535,N_6074,N_9144);
or U14536 (N_14536,N_9860,N_7030);
or U14537 (N_14537,N_5844,N_9810);
and U14538 (N_14538,N_8597,N_6205);
nand U14539 (N_14539,N_6003,N_9389);
nand U14540 (N_14540,N_7702,N_9357);
or U14541 (N_14541,N_9512,N_6241);
and U14542 (N_14542,N_8248,N_6246);
nand U14543 (N_14543,N_6427,N_9953);
and U14544 (N_14544,N_7053,N_7504);
and U14545 (N_14545,N_5975,N_6322);
nand U14546 (N_14546,N_8554,N_9283);
or U14547 (N_14547,N_6673,N_6356);
nand U14548 (N_14548,N_6009,N_6865);
and U14549 (N_14549,N_7628,N_6416);
and U14550 (N_14550,N_9653,N_6330);
and U14551 (N_14551,N_8651,N_5582);
or U14552 (N_14552,N_6118,N_8033);
nand U14553 (N_14553,N_9421,N_6600);
nor U14554 (N_14554,N_8253,N_8097);
nor U14555 (N_14555,N_8541,N_7785);
nand U14556 (N_14556,N_6886,N_5417);
and U14557 (N_14557,N_9153,N_7494);
nand U14558 (N_14558,N_9384,N_8451);
nor U14559 (N_14559,N_6080,N_5724);
nand U14560 (N_14560,N_8653,N_5312);
xor U14561 (N_14561,N_5280,N_5220);
or U14562 (N_14562,N_9094,N_9457);
and U14563 (N_14563,N_7253,N_6778);
nor U14564 (N_14564,N_6088,N_6995);
and U14565 (N_14565,N_8210,N_9742);
or U14566 (N_14566,N_7419,N_7782);
or U14567 (N_14567,N_8366,N_5207);
nand U14568 (N_14568,N_7385,N_5034);
or U14569 (N_14569,N_9744,N_8054);
nand U14570 (N_14570,N_6960,N_6082);
or U14571 (N_14571,N_5754,N_8747);
xnor U14572 (N_14572,N_5836,N_8294);
nand U14573 (N_14573,N_5250,N_7654);
or U14574 (N_14574,N_5655,N_8978);
or U14575 (N_14575,N_6035,N_5531);
nand U14576 (N_14576,N_6902,N_8864);
and U14577 (N_14577,N_7366,N_8453);
or U14578 (N_14578,N_6613,N_5726);
nand U14579 (N_14579,N_5344,N_9475);
nor U14580 (N_14580,N_7717,N_7646);
or U14581 (N_14581,N_6582,N_5357);
and U14582 (N_14582,N_9550,N_9812);
nand U14583 (N_14583,N_7506,N_9436);
and U14584 (N_14584,N_7749,N_8612);
or U14585 (N_14585,N_7846,N_6923);
nor U14586 (N_14586,N_9401,N_7378);
and U14587 (N_14587,N_8056,N_8643);
and U14588 (N_14588,N_7852,N_5136);
or U14589 (N_14589,N_9288,N_5021);
and U14590 (N_14590,N_5997,N_8612);
nor U14591 (N_14591,N_6346,N_7632);
nand U14592 (N_14592,N_8153,N_7310);
or U14593 (N_14593,N_6539,N_7565);
nand U14594 (N_14594,N_8843,N_7256);
nand U14595 (N_14595,N_8768,N_5797);
and U14596 (N_14596,N_9638,N_8634);
nor U14597 (N_14597,N_7485,N_7795);
and U14598 (N_14598,N_8134,N_9240);
nand U14599 (N_14599,N_6563,N_7721);
or U14600 (N_14600,N_5085,N_6217);
nand U14601 (N_14601,N_9273,N_9035);
nor U14602 (N_14602,N_6344,N_7037);
or U14603 (N_14603,N_7351,N_6257);
nor U14604 (N_14604,N_7801,N_6090);
or U14605 (N_14605,N_8166,N_5795);
nand U14606 (N_14606,N_8843,N_8860);
nor U14607 (N_14607,N_6800,N_7740);
and U14608 (N_14608,N_7830,N_5135);
or U14609 (N_14609,N_7487,N_8316);
nor U14610 (N_14610,N_7526,N_6508);
or U14611 (N_14611,N_5316,N_5645);
and U14612 (N_14612,N_9233,N_6546);
or U14613 (N_14613,N_9808,N_6855);
and U14614 (N_14614,N_9920,N_7804);
nand U14615 (N_14615,N_5240,N_5565);
nor U14616 (N_14616,N_7179,N_7397);
nand U14617 (N_14617,N_5087,N_5547);
and U14618 (N_14618,N_6203,N_7419);
or U14619 (N_14619,N_5406,N_6170);
nand U14620 (N_14620,N_8510,N_8466);
nand U14621 (N_14621,N_7102,N_7025);
nor U14622 (N_14622,N_9017,N_7489);
nand U14623 (N_14623,N_9880,N_7365);
and U14624 (N_14624,N_8862,N_5865);
or U14625 (N_14625,N_7098,N_7090);
xnor U14626 (N_14626,N_6252,N_6012);
and U14627 (N_14627,N_6694,N_8060);
or U14628 (N_14628,N_9541,N_8529);
and U14629 (N_14629,N_8335,N_5363);
or U14630 (N_14630,N_9761,N_8479);
nand U14631 (N_14631,N_8062,N_6007);
nor U14632 (N_14632,N_8787,N_9024);
or U14633 (N_14633,N_9833,N_8241);
nor U14634 (N_14634,N_6363,N_5084);
and U14635 (N_14635,N_5586,N_9794);
nor U14636 (N_14636,N_5299,N_7198);
and U14637 (N_14637,N_6719,N_7446);
nor U14638 (N_14638,N_8551,N_9610);
or U14639 (N_14639,N_7139,N_5622);
xor U14640 (N_14640,N_6908,N_8148);
and U14641 (N_14641,N_6975,N_7265);
or U14642 (N_14642,N_7293,N_9156);
or U14643 (N_14643,N_6785,N_8348);
or U14644 (N_14644,N_6418,N_9361);
and U14645 (N_14645,N_6562,N_9159);
or U14646 (N_14646,N_5866,N_6331);
or U14647 (N_14647,N_5744,N_5165);
nand U14648 (N_14648,N_7134,N_6065);
or U14649 (N_14649,N_8914,N_5374);
and U14650 (N_14650,N_7971,N_9998);
and U14651 (N_14651,N_6257,N_8118);
or U14652 (N_14652,N_6298,N_5256);
or U14653 (N_14653,N_7840,N_9531);
nand U14654 (N_14654,N_9545,N_8871);
and U14655 (N_14655,N_9618,N_9475);
nor U14656 (N_14656,N_9773,N_6171);
and U14657 (N_14657,N_5857,N_9832);
nand U14658 (N_14658,N_7857,N_7381);
nand U14659 (N_14659,N_8690,N_9652);
or U14660 (N_14660,N_5743,N_7805);
nor U14661 (N_14661,N_9265,N_8882);
and U14662 (N_14662,N_7203,N_7923);
nand U14663 (N_14663,N_6817,N_7713);
nand U14664 (N_14664,N_9928,N_8701);
or U14665 (N_14665,N_7659,N_8683);
or U14666 (N_14666,N_7651,N_6817);
or U14667 (N_14667,N_6490,N_8922);
or U14668 (N_14668,N_6583,N_9484);
and U14669 (N_14669,N_7369,N_7232);
and U14670 (N_14670,N_6285,N_6060);
or U14671 (N_14671,N_5342,N_7563);
or U14672 (N_14672,N_6117,N_8963);
or U14673 (N_14673,N_7309,N_7003);
or U14674 (N_14674,N_6313,N_5054);
nor U14675 (N_14675,N_7830,N_9106);
nand U14676 (N_14676,N_9224,N_8725);
nand U14677 (N_14677,N_8997,N_7581);
and U14678 (N_14678,N_5505,N_6410);
and U14679 (N_14679,N_8180,N_7396);
nand U14680 (N_14680,N_5597,N_6628);
and U14681 (N_14681,N_9735,N_8177);
or U14682 (N_14682,N_5796,N_9678);
nand U14683 (N_14683,N_5667,N_9656);
nor U14684 (N_14684,N_7419,N_5587);
and U14685 (N_14685,N_7493,N_7789);
or U14686 (N_14686,N_7892,N_9354);
nand U14687 (N_14687,N_5245,N_7400);
nor U14688 (N_14688,N_5850,N_9647);
nand U14689 (N_14689,N_7552,N_7071);
nand U14690 (N_14690,N_6948,N_9173);
nor U14691 (N_14691,N_7350,N_9604);
nand U14692 (N_14692,N_5054,N_5876);
and U14693 (N_14693,N_5998,N_6915);
or U14694 (N_14694,N_5930,N_9061);
nand U14695 (N_14695,N_8416,N_5862);
nor U14696 (N_14696,N_6710,N_5954);
and U14697 (N_14697,N_9888,N_5779);
nor U14698 (N_14698,N_8638,N_8799);
nor U14699 (N_14699,N_6317,N_8027);
and U14700 (N_14700,N_8785,N_6370);
and U14701 (N_14701,N_7111,N_9080);
and U14702 (N_14702,N_7137,N_7918);
nand U14703 (N_14703,N_8515,N_5007);
and U14704 (N_14704,N_9386,N_9672);
nand U14705 (N_14705,N_8225,N_8083);
nand U14706 (N_14706,N_5835,N_9193);
or U14707 (N_14707,N_7433,N_5577);
or U14708 (N_14708,N_8982,N_9620);
or U14709 (N_14709,N_5440,N_5197);
or U14710 (N_14710,N_7614,N_9451);
or U14711 (N_14711,N_5916,N_9479);
nand U14712 (N_14712,N_9354,N_5494);
and U14713 (N_14713,N_5921,N_6025);
and U14714 (N_14714,N_5248,N_7261);
and U14715 (N_14715,N_8091,N_5196);
and U14716 (N_14716,N_7925,N_5411);
nor U14717 (N_14717,N_7967,N_9388);
xnor U14718 (N_14718,N_7343,N_8772);
nand U14719 (N_14719,N_5352,N_6589);
and U14720 (N_14720,N_8626,N_5755);
and U14721 (N_14721,N_5896,N_5760);
and U14722 (N_14722,N_5282,N_9879);
and U14723 (N_14723,N_5293,N_7839);
nand U14724 (N_14724,N_9455,N_6247);
or U14725 (N_14725,N_6077,N_5510);
or U14726 (N_14726,N_9747,N_8903);
nor U14727 (N_14727,N_7711,N_7121);
nor U14728 (N_14728,N_9284,N_5986);
or U14729 (N_14729,N_7654,N_8500);
or U14730 (N_14730,N_8276,N_6616);
nor U14731 (N_14731,N_8205,N_8179);
nor U14732 (N_14732,N_8265,N_6955);
or U14733 (N_14733,N_5900,N_9009);
nor U14734 (N_14734,N_6761,N_6459);
or U14735 (N_14735,N_5636,N_8357);
nor U14736 (N_14736,N_9181,N_8781);
and U14737 (N_14737,N_8762,N_8088);
and U14738 (N_14738,N_8863,N_8716);
nor U14739 (N_14739,N_5171,N_5429);
nand U14740 (N_14740,N_7149,N_8558);
nor U14741 (N_14741,N_9457,N_7551);
nor U14742 (N_14742,N_5107,N_7730);
nor U14743 (N_14743,N_8571,N_8654);
or U14744 (N_14744,N_8679,N_9941);
and U14745 (N_14745,N_7835,N_9247);
or U14746 (N_14746,N_8919,N_9212);
and U14747 (N_14747,N_5916,N_8259);
or U14748 (N_14748,N_9674,N_8059);
xnor U14749 (N_14749,N_8282,N_5691);
nand U14750 (N_14750,N_5665,N_7064);
or U14751 (N_14751,N_6090,N_5290);
nand U14752 (N_14752,N_8663,N_7407);
nand U14753 (N_14753,N_5195,N_8299);
nand U14754 (N_14754,N_9025,N_7712);
and U14755 (N_14755,N_5320,N_8947);
and U14756 (N_14756,N_6189,N_7527);
and U14757 (N_14757,N_7894,N_9097);
nor U14758 (N_14758,N_9218,N_8445);
nor U14759 (N_14759,N_8575,N_5996);
or U14760 (N_14760,N_5357,N_7664);
nand U14761 (N_14761,N_8098,N_6693);
nand U14762 (N_14762,N_7555,N_5363);
or U14763 (N_14763,N_9496,N_7618);
nor U14764 (N_14764,N_7635,N_5320);
nor U14765 (N_14765,N_6416,N_9245);
nand U14766 (N_14766,N_6049,N_5585);
or U14767 (N_14767,N_7901,N_9877);
or U14768 (N_14768,N_6193,N_5609);
and U14769 (N_14769,N_7613,N_8802);
nand U14770 (N_14770,N_9240,N_7545);
nand U14771 (N_14771,N_7604,N_6875);
or U14772 (N_14772,N_8710,N_5950);
nor U14773 (N_14773,N_6223,N_6875);
nor U14774 (N_14774,N_7637,N_5370);
nand U14775 (N_14775,N_5619,N_5922);
and U14776 (N_14776,N_5113,N_5038);
nor U14777 (N_14777,N_6926,N_9662);
xnor U14778 (N_14778,N_6337,N_6108);
and U14779 (N_14779,N_5570,N_9138);
and U14780 (N_14780,N_5774,N_5102);
or U14781 (N_14781,N_9018,N_9517);
nand U14782 (N_14782,N_9717,N_7164);
and U14783 (N_14783,N_8695,N_7253);
and U14784 (N_14784,N_6227,N_9356);
nand U14785 (N_14785,N_5905,N_9748);
and U14786 (N_14786,N_6609,N_7083);
or U14787 (N_14787,N_7847,N_5302);
nor U14788 (N_14788,N_7255,N_6303);
nand U14789 (N_14789,N_8471,N_5221);
or U14790 (N_14790,N_8319,N_8919);
nand U14791 (N_14791,N_8428,N_5815);
or U14792 (N_14792,N_7537,N_9968);
or U14793 (N_14793,N_5891,N_8620);
nor U14794 (N_14794,N_6716,N_5315);
and U14795 (N_14795,N_6360,N_6035);
and U14796 (N_14796,N_6350,N_9277);
and U14797 (N_14797,N_6971,N_7562);
and U14798 (N_14798,N_6588,N_7201);
nand U14799 (N_14799,N_9868,N_6042);
and U14800 (N_14800,N_6145,N_5633);
nor U14801 (N_14801,N_6437,N_9233);
nor U14802 (N_14802,N_5162,N_9798);
nor U14803 (N_14803,N_9311,N_7702);
nand U14804 (N_14804,N_7222,N_9651);
or U14805 (N_14805,N_8450,N_5839);
nand U14806 (N_14806,N_9731,N_5026);
and U14807 (N_14807,N_8803,N_7345);
nor U14808 (N_14808,N_9350,N_9720);
or U14809 (N_14809,N_6412,N_7917);
or U14810 (N_14810,N_7769,N_9690);
nor U14811 (N_14811,N_7607,N_8191);
nand U14812 (N_14812,N_9369,N_6751);
nand U14813 (N_14813,N_6030,N_7248);
and U14814 (N_14814,N_9310,N_6308);
or U14815 (N_14815,N_6563,N_6599);
nor U14816 (N_14816,N_8325,N_5380);
or U14817 (N_14817,N_9983,N_6857);
or U14818 (N_14818,N_7060,N_9204);
or U14819 (N_14819,N_5256,N_8225);
or U14820 (N_14820,N_7231,N_8373);
nand U14821 (N_14821,N_5914,N_8455);
xor U14822 (N_14822,N_6070,N_9546);
nor U14823 (N_14823,N_7631,N_8108);
nor U14824 (N_14824,N_9347,N_7430);
or U14825 (N_14825,N_9135,N_8083);
nand U14826 (N_14826,N_7592,N_6644);
and U14827 (N_14827,N_8251,N_6067);
and U14828 (N_14828,N_5982,N_6704);
or U14829 (N_14829,N_8161,N_6671);
or U14830 (N_14830,N_8579,N_8127);
and U14831 (N_14831,N_7002,N_7045);
nand U14832 (N_14832,N_5942,N_9530);
nand U14833 (N_14833,N_8943,N_5261);
nor U14834 (N_14834,N_7853,N_9350);
nand U14835 (N_14835,N_7927,N_8821);
nand U14836 (N_14836,N_5890,N_7091);
or U14837 (N_14837,N_6969,N_6057);
and U14838 (N_14838,N_7374,N_8125);
nor U14839 (N_14839,N_7388,N_8254);
nand U14840 (N_14840,N_6525,N_6046);
nor U14841 (N_14841,N_7161,N_5667);
nand U14842 (N_14842,N_8266,N_8558);
or U14843 (N_14843,N_5389,N_5542);
or U14844 (N_14844,N_6314,N_9686);
nand U14845 (N_14845,N_5383,N_9897);
or U14846 (N_14846,N_6097,N_7444);
nand U14847 (N_14847,N_6573,N_9765);
or U14848 (N_14848,N_6211,N_8755);
nor U14849 (N_14849,N_7020,N_8249);
nor U14850 (N_14850,N_6072,N_5677);
and U14851 (N_14851,N_7688,N_9159);
nand U14852 (N_14852,N_6430,N_8712);
nor U14853 (N_14853,N_5650,N_7785);
or U14854 (N_14854,N_9866,N_7031);
nor U14855 (N_14855,N_7717,N_5504);
nor U14856 (N_14856,N_5146,N_5984);
and U14857 (N_14857,N_5876,N_9492);
and U14858 (N_14858,N_9339,N_7157);
or U14859 (N_14859,N_7207,N_9092);
nand U14860 (N_14860,N_9804,N_8531);
and U14861 (N_14861,N_7128,N_7097);
or U14862 (N_14862,N_8280,N_5462);
nor U14863 (N_14863,N_5068,N_9740);
nand U14864 (N_14864,N_6884,N_8664);
nor U14865 (N_14865,N_7776,N_9821);
or U14866 (N_14866,N_5537,N_5862);
nor U14867 (N_14867,N_7095,N_5434);
or U14868 (N_14868,N_7674,N_7191);
or U14869 (N_14869,N_7095,N_8006);
nand U14870 (N_14870,N_8212,N_6774);
nand U14871 (N_14871,N_9442,N_6372);
nor U14872 (N_14872,N_5022,N_9439);
nand U14873 (N_14873,N_8846,N_5727);
nand U14874 (N_14874,N_9910,N_9327);
nor U14875 (N_14875,N_9706,N_8889);
nor U14876 (N_14876,N_8080,N_7515);
or U14877 (N_14877,N_9523,N_5564);
nand U14878 (N_14878,N_7399,N_7341);
and U14879 (N_14879,N_7536,N_8750);
nand U14880 (N_14880,N_8421,N_5333);
or U14881 (N_14881,N_8966,N_6462);
nor U14882 (N_14882,N_6011,N_8572);
nand U14883 (N_14883,N_7009,N_5511);
nand U14884 (N_14884,N_9061,N_8331);
nand U14885 (N_14885,N_8548,N_9556);
nand U14886 (N_14886,N_9647,N_6779);
nor U14887 (N_14887,N_9714,N_6510);
nand U14888 (N_14888,N_5709,N_8601);
nand U14889 (N_14889,N_9447,N_7209);
nor U14890 (N_14890,N_8812,N_5497);
or U14891 (N_14891,N_8089,N_5936);
nand U14892 (N_14892,N_7954,N_6605);
nand U14893 (N_14893,N_6914,N_8020);
and U14894 (N_14894,N_8978,N_9809);
nor U14895 (N_14895,N_5593,N_9712);
or U14896 (N_14896,N_7585,N_6712);
or U14897 (N_14897,N_5779,N_6086);
nand U14898 (N_14898,N_9884,N_5182);
nor U14899 (N_14899,N_9182,N_5376);
nor U14900 (N_14900,N_7491,N_7480);
and U14901 (N_14901,N_8252,N_8146);
nand U14902 (N_14902,N_6149,N_5043);
nand U14903 (N_14903,N_8910,N_5566);
and U14904 (N_14904,N_6117,N_9408);
nand U14905 (N_14905,N_7140,N_7697);
nor U14906 (N_14906,N_9587,N_7207);
nand U14907 (N_14907,N_9759,N_7130);
nand U14908 (N_14908,N_9467,N_9802);
nand U14909 (N_14909,N_6144,N_5472);
nor U14910 (N_14910,N_5089,N_5506);
or U14911 (N_14911,N_7905,N_5374);
and U14912 (N_14912,N_8041,N_5944);
or U14913 (N_14913,N_5494,N_7538);
nor U14914 (N_14914,N_6073,N_5392);
or U14915 (N_14915,N_8624,N_7855);
nand U14916 (N_14916,N_6622,N_9019);
nor U14917 (N_14917,N_7772,N_9516);
nand U14918 (N_14918,N_6186,N_5546);
xnor U14919 (N_14919,N_8899,N_9723);
nor U14920 (N_14920,N_9459,N_6617);
nor U14921 (N_14921,N_7948,N_7684);
nor U14922 (N_14922,N_6828,N_9048);
and U14923 (N_14923,N_5198,N_5347);
and U14924 (N_14924,N_5354,N_7307);
nor U14925 (N_14925,N_9264,N_8273);
nor U14926 (N_14926,N_7956,N_8240);
nand U14927 (N_14927,N_5457,N_9482);
nand U14928 (N_14928,N_8373,N_5122);
or U14929 (N_14929,N_6579,N_8257);
nor U14930 (N_14930,N_6097,N_8771);
nor U14931 (N_14931,N_6462,N_5327);
and U14932 (N_14932,N_6557,N_9444);
nor U14933 (N_14933,N_6760,N_6427);
nand U14934 (N_14934,N_7600,N_9617);
and U14935 (N_14935,N_5207,N_6945);
or U14936 (N_14936,N_5673,N_5674);
nand U14937 (N_14937,N_8452,N_5485);
nor U14938 (N_14938,N_8020,N_9097);
or U14939 (N_14939,N_5796,N_6432);
or U14940 (N_14940,N_8978,N_6725);
nor U14941 (N_14941,N_5974,N_6665);
and U14942 (N_14942,N_9599,N_7094);
nand U14943 (N_14943,N_8715,N_9232);
nor U14944 (N_14944,N_9497,N_7349);
nor U14945 (N_14945,N_8682,N_8210);
nand U14946 (N_14946,N_9425,N_9103);
nand U14947 (N_14947,N_6707,N_8552);
nor U14948 (N_14948,N_9807,N_9193);
nor U14949 (N_14949,N_7225,N_8926);
and U14950 (N_14950,N_7904,N_5970);
nand U14951 (N_14951,N_7490,N_5584);
xnor U14952 (N_14952,N_8439,N_7266);
and U14953 (N_14953,N_7859,N_5011);
or U14954 (N_14954,N_9336,N_9116);
and U14955 (N_14955,N_9648,N_7681);
nand U14956 (N_14956,N_5744,N_8435);
nand U14957 (N_14957,N_7996,N_6851);
and U14958 (N_14958,N_9290,N_6317);
and U14959 (N_14959,N_7006,N_5343);
xor U14960 (N_14960,N_5100,N_5715);
or U14961 (N_14961,N_8165,N_5150);
nand U14962 (N_14962,N_7454,N_6105);
or U14963 (N_14963,N_7387,N_8670);
nand U14964 (N_14964,N_9031,N_5019);
and U14965 (N_14965,N_9729,N_9114);
nand U14966 (N_14966,N_5322,N_5935);
nor U14967 (N_14967,N_5840,N_7578);
nor U14968 (N_14968,N_5747,N_7614);
nor U14969 (N_14969,N_5378,N_5644);
nand U14970 (N_14970,N_8156,N_8384);
or U14971 (N_14971,N_9278,N_8870);
nand U14972 (N_14972,N_8177,N_7905);
nand U14973 (N_14973,N_9565,N_9211);
and U14974 (N_14974,N_7660,N_9201);
or U14975 (N_14975,N_6713,N_5829);
nand U14976 (N_14976,N_7126,N_8929);
nor U14977 (N_14977,N_6392,N_5345);
nand U14978 (N_14978,N_8228,N_7144);
or U14979 (N_14979,N_8357,N_7880);
nor U14980 (N_14980,N_8772,N_9032);
and U14981 (N_14981,N_7552,N_9747);
and U14982 (N_14982,N_6854,N_5841);
and U14983 (N_14983,N_6468,N_6173);
or U14984 (N_14984,N_7916,N_9876);
nor U14985 (N_14985,N_8347,N_8816);
and U14986 (N_14986,N_7499,N_7413);
nor U14987 (N_14987,N_8436,N_8354);
and U14988 (N_14988,N_7577,N_6553);
or U14989 (N_14989,N_8341,N_5614);
or U14990 (N_14990,N_8274,N_9875);
nor U14991 (N_14991,N_6131,N_5812);
nor U14992 (N_14992,N_6222,N_7722);
nand U14993 (N_14993,N_6490,N_8896);
nand U14994 (N_14994,N_9773,N_7803);
and U14995 (N_14995,N_6558,N_8751);
or U14996 (N_14996,N_7586,N_7105);
and U14997 (N_14997,N_6574,N_8993);
nor U14998 (N_14998,N_6620,N_9722);
nor U14999 (N_14999,N_5429,N_8866);
or UO_0 (O_0,N_11720,N_13277);
nor UO_1 (O_1,N_12091,N_13011);
or UO_2 (O_2,N_14325,N_13216);
or UO_3 (O_3,N_13284,N_10495);
nor UO_4 (O_4,N_13671,N_13678);
nand UO_5 (O_5,N_13474,N_10344);
nand UO_6 (O_6,N_14732,N_13456);
and UO_7 (O_7,N_10094,N_14003);
nor UO_8 (O_8,N_11955,N_13365);
nor UO_9 (O_9,N_14263,N_10521);
and UO_10 (O_10,N_13281,N_11047);
and UO_11 (O_11,N_11007,N_12674);
nand UO_12 (O_12,N_14835,N_14246);
nor UO_13 (O_13,N_14944,N_13394);
and UO_14 (O_14,N_11609,N_13217);
nor UO_15 (O_15,N_11029,N_12843);
nor UO_16 (O_16,N_10171,N_11094);
nor UO_17 (O_17,N_11156,N_12805);
nand UO_18 (O_18,N_12334,N_12149);
nand UO_19 (O_19,N_12501,N_11719);
and UO_20 (O_20,N_11906,N_10505);
or UO_21 (O_21,N_14032,N_13135);
nor UO_22 (O_22,N_10480,N_12868);
and UO_23 (O_23,N_11469,N_10439);
nand UO_24 (O_24,N_11359,N_11220);
or UO_25 (O_25,N_14783,N_11916);
or UO_26 (O_26,N_13165,N_10782);
or UO_27 (O_27,N_10602,N_11848);
or UO_28 (O_28,N_12835,N_12598);
and UO_29 (O_29,N_14213,N_14753);
and UO_30 (O_30,N_13734,N_11541);
and UO_31 (O_31,N_14361,N_13212);
nor UO_32 (O_32,N_11880,N_13289);
and UO_33 (O_33,N_11276,N_10147);
and UO_34 (O_34,N_11624,N_12148);
and UO_35 (O_35,N_10246,N_12790);
nand UO_36 (O_36,N_10283,N_11074);
or UO_37 (O_37,N_13654,N_10691);
nor UO_38 (O_38,N_13798,N_13552);
or UO_39 (O_39,N_11213,N_11451);
or UO_40 (O_40,N_10962,N_14181);
nand UO_41 (O_41,N_11164,N_14646);
nor UO_42 (O_42,N_11499,N_13684);
and UO_43 (O_43,N_14049,N_12888);
nand UO_44 (O_44,N_11344,N_10012);
and UO_45 (O_45,N_10506,N_13746);
and UO_46 (O_46,N_10587,N_10637);
nor UO_47 (O_47,N_14566,N_12647);
nor UO_48 (O_48,N_11377,N_11999);
nor UO_49 (O_49,N_13717,N_13962);
xnor UO_50 (O_50,N_13451,N_11982);
and UO_51 (O_51,N_10225,N_13816);
and UO_52 (O_52,N_12352,N_13703);
nand UO_53 (O_53,N_11885,N_14296);
or UO_54 (O_54,N_13527,N_13181);
and UO_55 (O_55,N_11518,N_14083);
nand UO_56 (O_56,N_10211,N_11010);
or UO_57 (O_57,N_14828,N_13749);
or UO_58 (O_58,N_14184,N_12948);
nor UO_59 (O_59,N_12739,N_12183);
nor UO_60 (O_60,N_13543,N_13064);
nand UO_61 (O_61,N_13015,N_12241);
and UO_62 (O_62,N_10957,N_13042);
or UO_63 (O_63,N_14793,N_13959);
or UO_64 (O_64,N_10747,N_13120);
or UO_65 (O_65,N_10373,N_14444);
and UO_66 (O_66,N_14358,N_13292);
and UO_67 (O_67,N_10054,N_14587);
or UO_68 (O_68,N_13305,N_13248);
and UO_69 (O_69,N_14250,N_14654);
nand UO_70 (O_70,N_11846,N_12252);
nand UO_71 (O_71,N_13779,N_14157);
and UO_72 (O_72,N_10825,N_14661);
and UO_73 (O_73,N_14995,N_14599);
nor UO_74 (O_74,N_14681,N_10323);
or UO_75 (O_75,N_14096,N_13311);
nor UO_76 (O_76,N_14253,N_14387);
nor UO_77 (O_77,N_11328,N_10628);
or UO_78 (O_78,N_11819,N_11153);
and UO_79 (O_79,N_14969,N_13761);
nor UO_80 (O_80,N_11909,N_11943);
and UO_81 (O_81,N_12399,N_10905);
nand UO_82 (O_82,N_10207,N_12066);
nor UO_83 (O_83,N_13274,N_11605);
and UO_84 (O_84,N_10220,N_13435);
or UO_85 (O_85,N_12933,N_11250);
and UO_86 (O_86,N_11653,N_13742);
nor UO_87 (O_87,N_14231,N_13252);
or UO_88 (O_88,N_13355,N_10697);
nor UO_89 (O_89,N_11867,N_14019);
nand UO_90 (O_90,N_11808,N_14927);
nand UO_91 (O_91,N_11496,N_10787);
nand UO_92 (O_92,N_11107,N_13743);
or UO_93 (O_93,N_14173,N_13698);
nand UO_94 (O_94,N_10789,N_13740);
and UO_95 (O_95,N_12500,N_13434);
and UO_96 (O_96,N_14490,N_10202);
nand UO_97 (O_97,N_10315,N_12829);
nor UO_98 (O_98,N_10101,N_14576);
nand UO_99 (O_99,N_14151,N_12012);
nand UO_100 (O_100,N_11455,N_13868);
and UO_101 (O_101,N_12119,N_13668);
nand UO_102 (O_102,N_12759,N_13834);
nor UO_103 (O_103,N_10167,N_14028);
or UO_104 (O_104,N_14419,N_14024);
and UO_105 (O_105,N_12086,N_12258);
nand UO_106 (O_106,N_14354,N_10862);
nor UO_107 (O_107,N_13149,N_13446);
nand UO_108 (O_108,N_11505,N_13488);
and UO_109 (O_109,N_13636,N_10792);
nand UO_110 (O_110,N_14116,N_12416);
nand UO_111 (O_111,N_14824,N_10332);
and UO_112 (O_112,N_13041,N_12643);
or UO_113 (O_113,N_13310,N_14657);
nand UO_114 (O_114,N_10065,N_13610);
and UO_115 (O_115,N_13321,N_12980);
or UO_116 (O_116,N_14457,N_13117);
or UO_117 (O_117,N_10208,N_12010);
nand UO_118 (O_118,N_11835,N_11268);
or UO_119 (O_119,N_14477,N_11594);
or UO_120 (O_120,N_12410,N_12295);
nand UO_121 (O_121,N_11474,N_14653);
or UO_122 (O_122,N_14284,N_11773);
nand UO_123 (O_123,N_10509,N_11516);
and UO_124 (O_124,N_12540,N_12931);
and UO_125 (O_125,N_12532,N_13713);
and UO_126 (O_126,N_11475,N_12880);
nand UO_127 (O_127,N_14016,N_10817);
or UO_128 (O_128,N_11569,N_10514);
or UO_129 (O_129,N_10530,N_12428);
and UO_130 (O_130,N_14478,N_14560);
nor UO_131 (O_131,N_10286,N_11882);
or UO_132 (O_132,N_13964,N_11187);
and UO_133 (O_133,N_10939,N_10206);
and UO_134 (O_134,N_10491,N_12026);
or UO_135 (O_135,N_11812,N_11096);
and UO_136 (O_136,N_10646,N_12212);
nand UO_137 (O_137,N_13098,N_13634);
nand UO_138 (O_138,N_12798,N_11067);
nand UO_139 (O_139,N_11162,N_13087);
or UO_140 (O_140,N_11315,N_10417);
or UO_141 (O_141,N_14752,N_14971);
nor UO_142 (O_142,N_10562,N_14264);
nor UO_143 (O_143,N_14497,N_12042);
and UO_144 (O_144,N_14711,N_14171);
nand UO_145 (O_145,N_10176,N_10608);
nand UO_146 (O_146,N_11218,N_12577);
nor UO_147 (O_147,N_13264,N_10650);
nor UO_148 (O_148,N_11995,N_14225);
nand UO_149 (O_149,N_11224,N_12648);
nand UO_150 (O_150,N_11945,N_14312);
nor UO_151 (O_151,N_10821,N_12713);
and UO_152 (O_152,N_13092,N_11211);
and UO_153 (O_153,N_12693,N_14965);
and UO_154 (O_154,N_10857,N_14866);
and UO_155 (O_155,N_11381,N_10039);
nor UO_156 (O_156,N_10927,N_10112);
nor UO_157 (O_157,N_10104,N_13839);
or UO_158 (O_158,N_12411,N_10268);
and UO_159 (O_159,N_10199,N_10959);
and UO_160 (O_160,N_10129,N_10389);
nand UO_161 (O_161,N_12811,N_11969);
nand UO_162 (O_162,N_11019,N_14289);
or UO_163 (O_163,N_14622,N_13119);
or UO_164 (O_164,N_14105,N_14122);
or UO_165 (O_165,N_13697,N_13232);
and UO_166 (O_166,N_12355,N_12579);
nand UO_167 (O_167,N_14875,N_13626);
and UO_168 (O_168,N_13757,N_11749);
or UO_169 (O_169,N_14124,N_10056);
and UO_170 (O_170,N_10791,N_13835);
nand UO_171 (O_171,N_14704,N_12907);
nand UO_172 (O_172,N_14235,N_12682);
and UO_173 (O_173,N_14913,N_14287);
nor UO_174 (O_174,N_12310,N_12903);
or UO_175 (O_175,N_12595,N_11763);
nor UO_176 (O_176,N_11484,N_12237);
nor UO_177 (O_177,N_14099,N_11636);
and UO_178 (O_178,N_13763,N_12286);
nand UO_179 (O_179,N_14210,N_13578);
and UO_180 (O_180,N_14574,N_10696);
and UO_181 (O_181,N_10615,N_14161);
nand UO_182 (O_182,N_11361,N_13551);
nor UO_183 (O_183,N_14418,N_14816);
nor UO_184 (O_184,N_11266,N_11168);
or UO_185 (O_185,N_14836,N_13526);
and UO_186 (O_186,N_14484,N_14042);
nand UO_187 (O_187,N_14953,N_14773);
or UO_188 (O_188,N_14685,N_11581);
nand UO_189 (O_189,N_12626,N_12074);
and UO_190 (O_190,N_10617,N_11369);
and UO_191 (O_191,N_12225,N_12642);
and UO_192 (O_192,N_14807,N_13785);
or UO_193 (O_193,N_13937,N_12944);
nand UO_194 (O_194,N_11396,N_14515);
and UO_195 (O_195,N_13114,N_13439);
nand UO_196 (O_196,N_13519,N_14277);
nor UO_197 (O_197,N_10422,N_14226);
and UO_198 (O_198,N_11037,N_14201);
and UO_199 (O_199,N_13948,N_10543);
or UO_200 (O_200,N_13029,N_13662);
nor UO_201 (O_201,N_11273,N_10548);
or UO_202 (O_202,N_11589,N_14898);
nor UO_203 (O_203,N_11663,N_10731);
and UO_204 (O_204,N_12985,N_11558);
nor UO_205 (O_205,N_11537,N_11648);
or UO_206 (O_206,N_13554,N_12180);
nand UO_207 (O_207,N_13141,N_12618);
nand UO_208 (O_208,N_12262,N_11005);
nor UO_209 (O_209,N_11545,N_14809);
and UO_210 (O_210,N_14382,N_12883);
and UO_211 (O_211,N_10024,N_14797);
nor UO_212 (O_212,N_10403,N_13807);
or UO_213 (O_213,N_11504,N_10970);
nand UO_214 (O_214,N_11843,N_14544);
nor UO_215 (O_215,N_14819,N_12623);
nor UO_216 (O_216,N_12530,N_13424);
or UO_217 (O_217,N_10964,N_13857);
or UO_218 (O_218,N_10410,N_12794);
nor UO_219 (O_219,N_10236,N_11802);
nand UO_220 (O_220,N_12476,N_10979);
nor UO_221 (O_221,N_14785,N_13334);
or UO_222 (O_222,N_14984,N_11336);
nand UO_223 (O_223,N_10191,N_11950);
or UO_224 (O_224,N_12005,N_14430);
nor UO_225 (O_225,N_13251,N_10856);
nor UO_226 (O_226,N_13235,N_11294);
or UO_227 (O_227,N_14321,N_10799);
nand UO_228 (O_228,N_13214,N_12502);
and UO_229 (O_229,N_10183,N_11927);
nor UO_230 (O_230,N_14505,N_14053);
nand UO_231 (O_231,N_14108,N_11065);
and UO_232 (O_232,N_14391,N_11866);
or UO_233 (O_233,N_13129,N_10255);
or UO_234 (O_234,N_14278,N_10145);
or UO_235 (O_235,N_14949,N_14005);
and UO_236 (O_236,N_10128,N_10513);
nand UO_237 (O_237,N_10947,N_14687);
or UO_238 (O_238,N_11741,N_13190);
nand UO_239 (O_239,N_11136,N_11321);
or UO_240 (O_240,N_13912,N_12049);
and UO_241 (O_241,N_14460,N_10461);
nand UO_242 (O_242,N_13019,N_14413);
and UO_243 (O_243,N_13416,N_11728);
nor UO_244 (O_244,N_11761,N_14182);
or UO_245 (O_245,N_10658,N_11608);
nand UO_246 (O_246,N_10418,N_13445);
nor UO_247 (O_247,N_14102,N_13316);
or UO_248 (O_248,N_11743,N_10861);
or UO_249 (O_249,N_10911,N_13601);
nand UO_250 (O_250,N_12079,N_14852);
or UO_251 (O_251,N_11422,N_10758);
or UO_252 (O_252,N_13187,N_12402);
nand UO_253 (O_253,N_14390,N_10574);
nor UO_254 (O_254,N_10975,N_12124);
or UO_255 (O_255,N_10355,N_12337);
and UO_256 (O_256,N_10638,N_12503);
and UO_257 (O_257,N_12118,N_10692);
and UO_258 (O_258,N_11473,N_12218);
or UO_259 (O_259,N_11772,N_11132);
or UO_260 (O_260,N_13861,N_10898);
nor UO_261 (O_261,N_14468,N_10441);
nand UO_262 (O_262,N_14609,N_10262);
or UO_263 (O_263,N_10035,N_12413);
and UO_264 (O_264,N_11888,N_13370);
nand UO_265 (O_265,N_14344,N_12731);
and UO_266 (O_266,N_12475,N_11941);
and UO_267 (O_267,N_13173,N_14485);
and UO_268 (O_268,N_13025,N_12612);
xor UO_269 (O_269,N_11073,N_12709);
nor UO_270 (O_270,N_14690,N_11724);
nand UO_271 (O_271,N_13920,N_11851);
and UO_272 (O_272,N_12009,N_11873);
nand UO_273 (O_273,N_12667,N_13775);
or UO_274 (O_274,N_11394,N_12581);
nand UO_275 (O_275,N_14536,N_14650);
or UO_276 (O_276,N_12832,N_11402);
or UO_277 (O_277,N_10775,N_14856);
or UO_278 (O_278,N_13317,N_10840);
nor UO_279 (O_279,N_14061,N_14466);
nor UO_280 (O_280,N_11138,N_10729);
nor UO_281 (O_281,N_14345,N_11899);
nor UO_282 (O_282,N_13977,N_12436);
or UO_283 (O_283,N_10477,N_11350);
and UO_284 (O_284,N_12704,N_14802);
or UO_285 (O_285,N_13598,N_13517);
or UO_286 (O_286,N_11521,N_10143);
or UO_287 (O_287,N_14189,N_13633);
nand UO_288 (O_288,N_11553,N_13627);
and UO_289 (O_289,N_11531,N_14327);
nor UO_290 (O_290,N_10594,N_13909);
nor UO_291 (O_291,N_11988,N_12940);
nor UO_292 (O_292,N_11022,N_11607);
nor UO_293 (O_293,N_12403,N_12011);
nand UO_294 (O_294,N_14366,N_12488);
nand UO_295 (O_295,N_13819,N_13147);
nand UO_296 (O_296,N_10958,N_10843);
or UO_297 (O_297,N_10778,N_12962);
or UO_298 (O_298,N_12353,N_12523);
or UO_299 (O_299,N_10592,N_10468);
and UO_300 (O_300,N_11011,N_11118);
nand UO_301 (O_301,N_12784,N_14672);
nor UO_302 (O_302,N_12472,N_10447);
nor UO_303 (O_303,N_13789,N_14668);
or UO_304 (O_304,N_12250,N_10013);
nand UO_305 (O_305,N_10100,N_14332);
or UO_306 (O_306,N_13006,N_11041);
nand UO_307 (O_307,N_14219,N_14050);
nand UO_308 (O_308,N_10230,N_10070);
or UO_309 (O_309,N_12307,N_13108);
and UO_310 (O_310,N_13840,N_14873);
and UO_311 (O_311,N_10448,N_14352);
nand UO_312 (O_312,N_14946,N_13282);
nor UO_313 (O_313,N_11014,N_11303);
and UO_314 (O_314,N_11254,N_10405);
or UO_315 (O_315,N_13781,N_10260);
or UO_316 (O_316,N_13796,N_12344);
nand UO_317 (O_317,N_13271,N_13470);
nor UO_318 (O_318,N_10660,N_12208);
nand UO_319 (O_319,N_13701,N_13245);
and UO_320 (O_320,N_11380,N_14805);
nand UO_321 (O_321,N_11706,N_10163);
nor UO_322 (O_322,N_13965,N_12849);
and UO_323 (O_323,N_10281,N_12157);
and UO_324 (O_324,N_12186,N_10348);
and UO_325 (O_325,N_13824,N_14166);
nor UO_326 (O_326,N_14133,N_14733);
nor UO_327 (O_327,N_10576,N_14494);
nor UO_328 (O_328,N_12806,N_14769);
or UO_329 (O_329,N_12365,N_13609);
or UO_330 (O_330,N_13299,N_12946);
or UO_331 (O_331,N_14818,N_13947);
nand UO_332 (O_332,N_14339,N_13385);
or UO_333 (O_333,N_10105,N_11676);
or UO_334 (O_334,N_12022,N_14156);
xor UO_335 (O_335,N_13125,N_13453);
nor UO_336 (O_336,N_12763,N_11967);
nand UO_337 (O_337,N_12261,N_13597);
nand UO_338 (O_338,N_11353,N_10838);
nand UO_339 (O_339,N_13345,N_11280);
and UO_340 (O_340,N_14942,N_12951);
nand UO_341 (O_341,N_10215,N_10426);
or UO_342 (O_342,N_14320,N_10115);
and UO_343 (O_343,N_14677,N_11201);
nand UO_344 (O_344,N_11340,N_10526);
nand UO_345 (O_345,N_13501,N_10783);
nand UO_346 (O_346,N_10231,N_11371);
or UO_347 (O_347,N_10198,N_14996);
nor UO_348 (O_348,N_12434,N_10107);
nor UO_349 (O_349,N_10682,N_14578);
nand UO_350 (O_350,N_13706,N_12167);
nand UO_351 (O_351,N_12377,N_12840);
and UO_352 (O_352,N_12382,N_14861);
nand UO_353 (O_353,N_12553,N_10307);
nand UO_354 (O_354,N_12514,N_14710);
and UO_355 (O_355,N_13624,N_13686);
nand UO_356 (O_356,N_11751,N_13710);
nand UO_357 (O_357,N_13258,N_11021);
and UO_358 (O_358,N_14409,N_11234);
or UO_359 (O_359,N_10459,N_10681);
and UO_360 (O_360,N_12546,N_13685);
nand UO_361 (O_361,N_12121,N_10093);
and UO_362 (O_362,N_14090,N_10683);
nor UO_363 (O_363,N_11035,N_12904);
and UO_364 (O_364,N_14867,N_10925);
nand UO_365 (O_365,N_11642,N_14735);
and UO_366 (O_366,N_10040,N_10566);
nor UO_367 (O_367,N_13016,N_10294);
nand UO_368 (O_368,N_14338,N_14465);
nor UO_369 (O_369,N_13646,N_12802);
and UO_370 (O_370,N_13239,N_12653);
or UO_371 (O_371,N_10282,N_13148);
nand UO_372 (O_372,N_12447,N_11680);
nor UO_373 (O_373,N_10641,N_12740);
nand UO_374 (O_374,N_11869,N_13081);
nand UO_375 (O_375,N_10913,N_13536);
nor UO_376 (O_376,N_12699,N_10695);
and UO_377 (O_377,N_10714,N_13290);
or UO_378 (O_378,N_11855,N_14665);
and UO_379 (O_379,N_11739,N_14127);
or UO_380 (O_380,N_13233,N_11199);
or UO_381 (O_381,N_13509,N_10451);
and UO_382 (O_382,N_14731,N_14741);
and UO_383 (O_383,N_11833,N_12779);
or UO_384 (O_384,N_10270,N_14571);
nor UO_385 (O_385,N_10014,N_14307);
nand UO_386 (O_386,N_12110,N_14489);
nand UO_387 (O_387,N_13047,N_12383);
or UO_388 (O_388,N_10337,N_14521);
and UO_389 (O_389,N_14087,N_13930);
or UO_390 (O_390,N_13485,N_13707);
and UO_391 (O_391,N_14216,N_10705);
and UO_392 (O_392,N_11388,N_14736);
nor UO_393 (O_393,N_13452,N_14383);
nand UO_394 (O_394,N_12204,N_12677);
or UO_395 (O_395,N_13102,N_14720);
and UO_396 (O_396,N_12267,N_10730);
and UO_397 (O_397,N_14977,N_10341);
nor UO_398 (O_398,N_12467,N_11032);
nand UO_399 (O_399,N_14832,N_13990);
or UO_400 (O_400,N_12926,N_12321);
nand UO_401 (O_401,N_12977,N_12730);
nor UO_402 (O_402,N_14041,N_10693);
and UO_403 (O_403,N_12151,N_13872);
nand UO_404 (O_404,N_11183,N_13926);
or UO_405 (O_405,N_13998,N_12238);
nor UO_406 (O_406,N_11818,N_14459);
or UO_407 (O_407,N_13658,N_13441);
nand UO_408 (O_408,N_12761,N_12804);
or UO_409 (O_409,N_14365,N_13814);
and UO_410 (O_410,N_12785,N_11111);
nor UO_411 (O_411,N_10607,N_11391);
and UO_412 (O_412,N_14186,N_14367);
and UO_413 (O_413,N_14956,N_10431);
and UO_414 (O_414,N_10485,N_12879);
nand UO_415 (O_415,N_10442,N_11288);
nor UO_416 (O_416,N_12441,N_10849);
and UO_417 (O_417,N_11914,N_12629);
or UO_418 (O_418,N_13225,N_13167);
nand UO_419 (O_419,N_14118,N_10896);
nor UO_420 (O_420,N_10452,N_13155);
nand UO_421 (O_421,N_14180,N_10175);
nor UO_422 (O_422,N_14568,N_13419);
nor UO_423 (O_423,N_14857,N_12437);
nand UO_424 (O_424,N_10233,N_11229);
nand UO_425 (O_425,N_14359,N_10584);
and UO_426 (O_426,N_13637,N_12300);
and UO_427 (O_427,N_13644,N_11244);
or UO_428 (O_428,N_12791,N_11495);
nor UO_429 (O_429,N_11262,N_12768);
or UO_430 (O_430,N_14052,N_13862);
nand UO_431 (O_431,N_11954,N_14017);
or UO_432 (O_432,N_14285,N_10921);
or UO_433 (O_433,N_12935,N_12795);
and UO_434 (O_434,N_11717,N_12526);
or UO_435 (O_435,N_14146,N_14663);
and UO_436 (O_436,N_11490,N_12178);
and UO_437 (O_437,N_11650,N_10284);
and UO_438 (O_438,N_10570,N_12673);
or UO_439 (O_439,N_11614,N_11146);
nor UO_440 (O_440,N_11860,N_12493);
or UO_441 (O_441,N_12645,N_12260);
nand UO_442 (O_442,N_10733,N_11951);
or UO_443 (O_443,N_11633,N_10771);
nor UO_444 (O_444,N_10713,N_10750);
nor UO_445 (O_445,N_10850,N_12095);
and UO_446 (O_446,N_13306,N_13246);
and UO_447 (O_447,N_13238,N_11998);
and UO_448 (O_448,N_12810,N_14316);
or UO_449 (O_449,N_10810,N_10325);
and UO_450 (O_450,N_12210,N_12229);
nand UO_451 (O_451,N_11471,N_14794);
nand UO_452 (O_452,N_11815,N_14271);
or UO_453 (O_453,N_10865,N_13675);
or UO_454 (O_454,N_12752,N_12996);
and UO_455 (O_455,N_14728,N_14762);
or UO_456 (O_456,N_12519,N_14559);
or UO_457 (O_457,N_14274,N_11528);
or UO_458 (O_458,N_10851,N_13894);
nand UO_459 (O_459,N_11030,N_11525);
nor UO_460 (O_460,N_10989,N_13567);
nand UO_461 (O_461,N_13161,N_12296);
nand UO_462 (O_462,N_12615,N_10580);
nor UO_463 (O_463,N_12253,N_10425);
nand UO_464 (O_464,N_12717,N_11345);
and UO_465 (O_465,N_12187,N_11522);
or UO_466 (O_466,N_14636,N_13145);
and UO_467 (O_467,N_13066,N_14426);
or UO_468 (O_468,N_10358,N_10872);
and UO_469 (O_469,N_10803,N_13454);
nand UO_470 (O_470,N_12886,N_14813);
nand UO_471 (O_471,N_12316,N_11444);
nor UO_472 (O_472,N_12734,N_13974);
nor UO_473 (O_473,N_12608,N_11735);
or UO_474 (O_474,N_12590,N_12562);
or UO_475 (O_475,N_13262,N_13286);
nand UO_476 (O_476,N_13309,N_12989);
or UO_477 (O_477,N_13681,N_12409);
and UO_478 (O_478,N_14695,N_11367);
or UO_479 (O_479,N_11063,N_11202);
nor UO_480 (O_480,N_10305,N_12000);
and UO_481 (O_481,N_13587,N_13897);
or UO_482 (O_482,N_10854,N_14167);
or UO_483 (O_483,N_11448,N_13495);
nand UO_484 (O_484,N_13139,N_11348);
nor UO_485 (O_485,N_10518,N_14493);
and UO_486 (O_486,N_10438,N_12830);
nor UO_487 (O_487,N_13287,N_13090);
xor UO_488 (O_488,N_14230,N_13660);
and UO_489 (O_489,N_14084,N_10372);
or UO_490 (O_490,N_13194,N_14770);
and UO_491 (O_491,N_11920,N_12376);
nor UO_492 (O_492,N_10642,N_13157);
nor UO_493 (O_493,N_13344,N_14011);
nor UO_494 (O_494,N_11316,N_10906);
nor UO_495 (O_495,N_13350,N_12299);
or UO_496 (O_496,N_12508,N_10460);
and UO_497 (O_497,N_12446,N_10336);
and UO_498 (O_498,N_14619,N_12451);
and UO_499 (O_499,N_14691,N_12465);
nand UO_500 (O_500,N_12536,N_14403);
nand UO_501 (O_501,N_13091,N_11631);
and UO_502 (O_502,N_14254,N_12466);
or UO_503 (O_503,N_11274,N_12702);
or UO_504 (O_504,N_12837,N_12181);
or UO_505 (O_505,N_11887,N_12978);
or UO_506 (O_506,N_14744,N_13753);
nor UO_507 (O_507,N_13576,N_13705);
nand UO_508 (O_508,N_14834,N_12057);
nor UO_509 (O_509,N_14565,N_12970);
nor UO_510 (O_510,N_13423,N_13017);
and UO_511 (O_511,N_10918,N_13691);
nor UO_512 (O_512,N_12567,N_11436);
nand UO_513 (O_513,N_13569,N_11894);
nor UO_514 (O_514,N_11686,N_10313);
nor UO_515 (O_515,N_13522,N_13422);
nor UO_516 (O_516,N_10836,N_11807);
and UO_517 (O_517,N_14340,N_11926);
and UO_518 (O_518,N_12272,N_10572);
or UO_519 (O_519,N_12587,N_11181);
nand UO_520 (O_520,N_11755,N_14803);
or UO_521 (O_521,N_13295,N_10804);
and UO_522 (O_522,N_12325,N_11442);
and UO_523 (O_523,N_14266,N_13390);
and UO_524 (O_524,N_13179,N_13563);
nand UO_525 (O_525,N_14393,N_10021);
or UO_526 (O_526,N_12930,N_11520);
and UO_527 (O_527,N_12478,N_12559);
nor UO_528 (O_528,N_12782,N_13213);
or UO_529 (O_529,N_13766,N_11679);
nor UO_530 (O_530,N_12848,N_12314);
and UO_531 (O_531,N_12264,N_13402);
nand UO_532 (O_532,N_10735,N_10569);
nor UO_533 (O_533,N_10251,N_10721);
and UO_534 (O_534,N_11568,N_11102);
nor UO_535 (O_535,N_10819,N_10604);
nand UO_536 (O_536,N_12177,N_13860);
and UO_537 (O_537,N_11801,N_14002);
nor UO_538 (O_538,N_14280,N_12720);
or UO_539 (O_539,N_13810,N_10719);
or UO_540 (O_540,N_12239,N_10203);
nand UO_541 (O_541,N_13459,N_12958);
and UO_542 (O_542,N_12006,N_12571);
nand UO_543 (O_543,N_12769,N_12408);
or UO_544 (O_544,N_14886,N_12471);
nand UO_545 (O_545,N_13648,N_11659);
nor UO_546 (O_546,N_11125,N_14326);
and UO_547 (O_547,N_10928,N_12669);
or UO_548 (O_548,N_11506,N_12834);
or UO_549 (O_549,N_11810,N_11934);
nor UO_550 (O_550,N_11456,N_10492);
nand UO_551 (O_551,N_10444,N_11570);
or UO_552 (O_552,N_11189,N_11269);
nor UO_553 (O_553,N_10583,N_13399);
or UO_554 (O_554,N_12351,N_10739);
nor UO_555 (O_555,N_13116,N_14742);
and UO_556 (O_556,N_14772,N_14778);
and UO_557 (O_557,N_10603,N_10412);
and UO_558 (O_558,N_11298,N_13778);
or UO_559 (O_559,N_14006,N_11373);
and UO_560 (O_560,N_13996,N_11806);
nand UO_561 (O_561,N_12135,N_14217);
and UO_562 (O_562,N_11123,N_13342);
and UO_563 (O_563,N_13566,N_12509);
and UO_564 (O_564,N_14979,N_10727);
and UO_565 (O_565,N_12067,N_11251);
nor UO_566 (O_566,N_11064,N_13191);
nand UO_567 (O_567,N_14992,N_10924);
and UO_568 (O_568,N_13969,N_11072);
and UO_569 (O_569,N_11657,N_14651);
nor UO_570 (O_570,N_11879,N_11709);
nor UO_571 (O_571,N_13588,N_11219);
and UO_572 (O_572,N_13592,N_14104);
and UO_573 (O_573,N_14228,N_10036);
nand UO_574 (O_574,N_13794,N_14652);
or UO_575 (O_575,N_10776,N_13069);
or UO_576 (O_576,N_13103,N_11771);
xnor UO_577 (O_577,N_10591,N_12282);
nor UO_578 (O_578,N_11492,N_12141);
or UO_579 (O_579,N_11864,N_11645);
nand UO_580 (O_580,N_10349,N_10279);
nor UO_581 (O_581,N_12914,N_11134);
nand UO_582 (O_582,N_14829,N_13620);
nor UO_583 (O_583,N_11939,N_12788);
nor UO_584 (O_584,N_14222,N_13606);
nor UO_585 (O_585,N_13944,N_12694);
and UO_586 (O_586,N_11237,N_14131);
or UO_587 (O_587,N_14922,N_13546);
and UO_588 (O_588,N_12481,N_14594);
nand UO_589 (O_589,N_14738,N_13099);
nor UO_590 (O_590,N_14799,N_13097);
or UO_591 (O_591,N_11296,N_10133);
nand UO_592 (O_592,N_12202,N_12222);
nor UO_593 (O_593,N_11382,N_13655);
and UO_594 (O_594,N_11309,N_14943);
nand UO_595 (O_595,N_11640,N_14072);
or UO_596 (O_596,N_11983,N_13226);
nor UO_597 (O_597,N_12456,N_10728);
and UO_598 (O_598,N_10968,N_12963);
and UO_599 (O_599,N_14048,N_14139);
nor UO_600 (O_600,N_12288,N_10159);
nand UO_601 (O_601,N_12214,N_12331);
and UO_602 (O_602,N_14684,N_12976);
nand UO_603 (O_603,N_10200,N_14449);
and UO_604 (O_604,N_12518,N_11300);
nor UO_605 (O_605,N_10032,N_10984);
nor UO_606 (O_606,N_13545,N_11793);
nand UO_607 (O_607,N_14404,N_11750);
and UO_608 (O_608,N_10829,N_13267);
nor UO_609 (O_609,N_12381,N_10503);
nand UO_610 (O_610,N_11364,N_10618);
or UO_611 (O_611,N_11690,N_11721);
and UO_612 (O_612,N_14331,N_14939);
or UO_613 (O_613,N_10007,N_14585);
and UO_614 (O_614,N_10867,N_12171);
nand UO_615 (O_615,N_10529,N_13672);
or UO_616 (O_616,N_13003,N_12027);
and UO_617 (O_617,N_14840,N_12248);
or UO_618 (O_618,N_12609,N_10309);
nor UO_619 (O_619,N_11868,N_13244);
nand UO_620 (O_620,N_10746,N_13542);
nand UO_621 (O_621,N_10184,N_12550);
and UO_622 (O_622,N_10394,N_11637);
or UO_623 (O_623,N_12343,N_13038);
nor UO_624 (O_624,N_13367,N_13673);
nand UO_625 (O_625,N_13797,N_11515);
or UO_626 (O_626,N_12658,N_11891);
nor UO_627 (O_627,N_10037,N_12913);
or UO_628 (O_628,N_12706,N_14158);
or UO_629 (O_629,N_14305,N_14877);
nor UO_630 (O_630,N_14434,N_13549);
nand UO_631 (O_631,N_13219,N_12736);
nor UO_632 (O_632,N_10333,N_13348);
nor UO_633 (O_633,N_14060,N_10816);
nor UO_634 (O_634,N_14592,N_14103);
nor UO_635 (O_635,N_14441,N_12226);
nor UO_636 (O_636,N_11355,N_14392);
or UO_637 (O_637,N_13884,N_13095);
and UO_638 (O_638,N_11536,N_11874);
or UO_639 (O_639,N_12039,N_12290);
and UO_640 (O_640,N_12711,N_10868);
and UO_641 (O_641,N_11433,N_13484);
nor UO_642 (O_642,N_12748,N_13085);
nor UO_643 (O_643,N_10297,N_10455);
or UO_644 (O_644,N_10076,N_14420);
or UO_645 (O_645,N_11859,N_12861);
and UO_646 (O_646,N_11768,N_13525);
nor UO_647 (O_647,N_11223,N_12610);
nor UO_648 (O_648,N_14207,N_14514);
and UO_649 (O_649,N_11649,N_13083);
and UO_650 (O_650,N_12230,N_11781);
or UO_651 (O_651,N_11928,N_10470);
nor UO_652 (O_652,N_12722,N_10437);
xor UO_653 (O_653,N_10549,N_14190);
nand UO_654 (O_654,N_12084,N_10474);
nand UO_655 (O_655,N_14513,N_13487);
nor UO_656 (O_656,N_14934,N_12139);
nor UO_657 (O_657,N_10339,N_12999);
or UO_658 (O_658,N_11068,N_14518);
nand UO_659 (O_659,N_10568,N_12863);
nor UO_660 (O_660,N_12644,N_13323);
or UO_661 (O_661,N_12961,N_11236);
or UO_662 (O_662,N_14267,N_11503);
nor UO_663 (O_663,N_13450,N_11311);
nand UO_664 (O_664,N_14147,N_12496);
nor UO_665 (O_665,N_11795,N_13531);
nor UO_666 (O_666,N_14265,N_12942);
or UO_667 (O_667,N_10579,N_13851);
and UO_668 (O_668,N_14906,N_13031);
nand UO_669 (O_669,N_10963,N_11104);
and UO_670 (O_670,N_10222,N_11994);
and UO_671 (O_671,N_14531,N_10933);
nand UO_672 (O_672,N_14261,N_11427);
nand UO_673 (O_673,N_12034,N_10280);
nand UO_674 (O_674,N_12822,N_10807);
and UO_675 (O_675,N_10930,N_12812);
nor UO_676 (O_676,N_13584,N_11840);
or UO_677 (O_677,N_10929,N_10125);
nand UO_678 (O_678,N_13720,N_11870);
nand UO_679 (O_679,N_10015,N_14701);
and UO_680 (O_680,N_12982,N_14273);
or UO_681 (O_681,N_10106,N_10234);
and UO_682 (O_682,N_11404,N_12729);
and UO_683 (O_683,N_10310,N_11040);
or UO_684 (O_684,N_11500,N_14454);
nand UO_685 (O_685,N_12168,N_13725);
nor UO_686 (O_686,N_12104,N_10919);
nand UO_687 (O_687,N_10082,N_13918);
or UO_688 (O_688,N_13140,N_11200);
and UO_689 (O_689,N_10150,N_10986);
and UO_690 (O_690,N_14980,N_13372);
nand UO_691 (O_691,N_14232,N_14908);
nand UO_692 (O_692,N_12522,N_13301);
or UO_693 (O_693,N_11465,N_11789);
or UO_694 (O_694,N_10009,N_11667);
or UO_695 (O_695,N_14159,N_14512);
nand UO_696 (O_696,N_11039,N_13844);
or UO_697 (O_697,N_12125,N_10702);
or UO_698 (O_698,N_11100,N_11527);
nand UO_699 (O_699,N_10457,N_10764);
and UO_700 (O_700,N_11192,N_11434);
nor UO_701 (O_701,N_13493,N_11968);
or UO_702 (O_702,N_10419,N_10050);
or UO_703 (O_703,N_11924,N_13958);
nor UO_704 (O_704,N_14496,N_10060);
and UO_705 (O_705,N_13168,N_13056);
nand UO_706 (O_706,N_14725,N_11082);
nor UO_707 (O_707,N_13967,N_12555);
nand UO_708 (O_708,N_11263,N_12342);
or UO_709 (O_709,N_11261,N_11413);
nand UO_710 (O_710,N_13783,N_14279);
nor UO_711 (O_711,N_10146,N_12712);
nand UO_712 (O_712,N_10088,N_12727);
nor UO_713 (O_713,N_12263,N_12224);
or UO_714 (O_714,N_11576,N_10665);
nand UO_715 (O_715,N_12162,N_10811);
or UO_716 (O_716,N_10823,N_11150);
nand UO_717 (O_717,N_13621,N_11126);
nand UO_718 (O_718,N_11108,N_12454);
nor UO_719 (O_719,N_14903,N_11152);
nor UO_720 (O_720,N_11331,N_12341);
nand UO_721 (O_721,N_13680,N_10052);
nand UO_722 (O_722,N_14329,N_14739);
and UO_723 (O_723,N_12771,N_14581);
nor UO_724 (O_724,N_12070,N_14086);
and UO_725 (O_725,N_10551,N_13300);
nor UO_726 (O_726,N_11259,N_12543);
or UO_727 (O_727,N_13022,N_13315);
nor UO_728 (O_728,N_10774,N_12657);
nor UO_729 (O_729,N_14874,N_11900);
nand UO_730 (O_730,N_11131,N_12032);
nand UO_731 (O_731,N_11405,N_12199);
or UO_732 (O_732,N_14111,N_13960);
nor UO_733 (O_733,N_14808,N_14849);
nand UO_734 (O_734,N_10252,N_11343);
nand UO_735 (O_735,N_12979,N_14612);
nand UO_736 (O_736,N_10001,N_10785);
and UO_737 (O_737,N_10327,N_11519);
or UO_738 (O_738,N_12892,N_10780);
nand UO_739 (O_739,N_10654,N_14697);
and UO_740 (O_740,N_12469,N_11089);
or UO_741 (O_741,N_10272,N_13647);
or UO_742 (O_742,N_14437,N_13773);
or UO_743 (O_743,N_12796,N_11163);
or UO_744 (O_744,N_10732,N_11956);
nand UO_745 (O_745,N_12158,N_12767);
and UO_746 (O_746,N_11902,N_12495);
or UO_747 (O_747,N_14826,N_10894);
nand UO_748 (O_748,N_12603,N_14341);
nor UO_749 (O_749,N_10177,N_12015);
and UO_750 (O_750,N_10784,N_11711);
and UO_751 (O_751,N_11986,N_11790);
nor UO_752 (O_752,N_13336,N_13055);
nor UO_753 (O_753,N_11824,N_10224);
and UO_754 (O_754,N_14973,N_11905);
and UO_755 (O_755,N_13882,N_14200);
xor UO_756 (O_756,N_11003,N_13461);
nor UO_757 (O_757,N_13280,N_13302);
nand UO_758 (O_758,N_10723,N_11066);
nor UO_759 (O_759,N_11511,N_10322);
nand UO_760 (O_760,N_13210,N_14342);
or UO_761 (O_761,N_14895,N_10744);
or UO_762 (O_762,N_10258,N_10876);
nand UO_763 (O_763,N_10786,N_13380);
nand UO_764 (O_764,N_12714,N_13983);
nand UO_765 (O_765,N_13397,N_14885);
nor UO_766 (O_766,N_10320,N_12368);
or UO_767 (O_767,N_11559,N_12442);
or UO_768 (O_768,N_13723,N_10400);
nor UO_769 (O_769,N_13997,N_12990);
nand UO_770 (O_770,N_11601,N_14362);
nand UO_771 (O_771,N_13115,N_13028);
and UO_772 (O_772,N_14281,N_11682);
nor UO_773 (O_773,N_14112,N_11227);
nand UO_774 (O_774,N_10376,N_14486);
nor UO_775 (O_775,N_14747,N_11159);
nand UO_776 (O_776,N_14976,N_10891);
or UO_777 (O_777,N_11117,N_12678);
nor UO_778 (O_778,N_13358,N_11991);
nor UO_779 (O_779,N_13270,N_14858);
and UO_780 (O_780,N_10625,N_11430);
or UO_781 (O_781,N_12242,N_11171);
or UO_782 (O_782,N_14626,N_14789);
and UO_783 (O_783,N_13492,N_11360);
nand UO_784 (O_784,N_11352,N_12773);
nor UO_785 (O_785,N_11349,N_13486);
nand UO_786 (O_786,N_12405,N_13650);
nand UO_787 (O_787,N_14333,N_13975);
nor UO_788 (O_788,N_14179,N_10067);
or UO_789 (O_789,N_11036,N_14970);
nor UO_790 (O_790,N_12430,N_14206);
nor UO_791 (O_791,N_11307,N_12619);
or UO_792 (O_792,N_13935,N_13366);
nand UO_793 (O_793,N_10414,N_14297);
nand UO_794 (O_794,N_10915,N_10025);
nor UO_795 (O_795,N_13198,N_14034);
nand UO_796 (O_796,N_13068,N_13051);
nor UO_797 (O_797,N_14044,N_11612);
or UO_798 (O_798,N_10490,N_13639);
nand UO_799 (O_799,N_10762,N_10170);
or UO_800 (O_800,N_11792,N_11575);
or UO_801 (O_801,N_12542,N_13018);
nand UO_802 (O_802,N_13871,N_10293);
nand UO_803 (O_803,N_12576,N_11708);
nor UO_804 (O_804,N_13261,N_12313);
nor UO_805 (O_805,N_10656,N_14597);
nor UO_806 (O_806,N_14029,N_13611);
nand UO_807 (O_807,N_14351,N_11529);
nand UO_808 (O_808,N_14379,N_12431);
nor UO_809 (O_809,N_14255,N_10997);
nand UO_810 (O_810,N_10187,N_12504);
or UO_811 (O_811,N_13171,N_14948);
and UO_812 (O_812,N_11256,N_11464);
nand UO_813 (O_813,N_11912,N_13771);
nor UO_814 (O_814,N_14205,N_11441);
or UO_815 (O_815,N_13330,N_11195);
nor UO_816 (O_816,N_11713,N_14500);
or UO_817 (O_817,N_13482,N_12602);
nor UO_818 (O_818,N_13253,N_10196);
nand UO_819 (O_819,N_14456,N_11754);
nand UO_820 (O_820,N_11147,N_14696);
or UO_821 (O_821,N_14698,N_13273);
or UO_822 (O_822,N_10381,N_11615);
or UO_823 (O_823,N_14079,N_12176);
or UO_824 (O_824,N_10298,N_14945);
nand UO_825 (O_825,N_12556,N_11946);
or UO_826 (O_826,N_10113,N_11587);
and UO_827 (O_827,N_10842,N_10985);
and UO_828 (O_828,N_11319,N_14850);
or UO_829 (O_829,N_10064,N_10462);
nor UO_830 (O_830,N_11674,N_13714);
nor UO_831 (O_831,N_10680,N_10934);
nand UO_832 (O_832,N_14841,N_11557);
or UO_833 (O_833,N_10226,N_11257);
nor UO_834 (O_834,N_13278,N_14707);
nand UO_835 (O_835,N_10122,N_10398);
nor UO_836 (O_836,N_13952,N_13208);
and UO_837 (O_837,N_14119,N_10507);
nand UO_838 (O_838,N_14530,N_11155);
and UO_839 (O_839,N_10832,N_11206);
nand UO_840 (O_840,N_14990,N_13533);
or UO_841 (O_841,N_12746,N_13818);
and UO_842 (O_842,N_13847,N_10880);
or UO_843 (O_843,N_13946,N_11302);
and UO_844 (O_844,N_11597,N_14617);
nand UO_845 (O_845,N_13529,N_13747);
nor UO_846 (O_846,N_13298,N_12853);
nor UO_847 (O_847,N_11602,N_12628);
nor UO_848 (O_848,N_14046,N_11389);
nand UO_849 (O_849,N_12133,N_13793);
nor UO_850 (O_850,N_10338,N_10657);
nor UO_851 (O_851,N_10718,N_11744);
and UO_852 (O_852,N_10162,N_10845);
nand UO_853 (O_853,N_10289,N_12703);
nor UO_854 (O_854,N_10370,N_14998);
nand UO_855 (O_855,N_13436,N_12866);
and UO_856 (O_856,N_12081,N_13243);
nand UO_857 (O_857,N_13065,N_13513);
nor UO_858 (O_858,N_11463,N_10109);
nor UO_859 (O_859,N_13572,N_14925);
nand UO_860 (O_860,N_11826,N_12919);
or UO_861 (O_861,N_10292,N_12632);
and UO_862 (O_862,N_11318,N_10103);
nor UO_863 (O_863,N_14727,N_11952);
nor UO_864 (O_864,N_14384,N_12924);
and UO_865 (O_865,N_10770,N_13692);
or UO_866 (O_866,N_10519,N_13032);
nor UO_867 (O_867,N_12320,N_14155);
nand UO_868 (O_868,N_10369,N_14608);
and UO_869 (O_869,N_11705,N_12983);
and UO_870 (O_870,N_14153,N_14078);
and UO_871 (O_871,N_12132,N_11027);
nor UO_872 (O_872,N_10689,N_11446);
and UO_873 (O_873,N_13178,N_10554);
or UO_874 (O_874,N_14745,N_10777);
nor UO_875 (O_875,N_10471,N_10734);
nor UO_876 (O_876,N_13657,N_10741);
nand UO_877 (O_877,N_11411,N_14962);
or UO_878 (O_878,N_10449,N_13156);
xnor UO_879 (O_879,N_13448,N_13679);
and UO_880 (O_880,N_10110,N_10139);
nand UO_881 (O_881,N_13520,N_11876);
and UO_882 (O_882,N_11406,N_13727);
or UO_883 (O_883,N_11970,N_14959);
nor UO_884 (O_884,N_10424,N_11374);
nand UO_885 (O_885,N_13902,N_13084);
nor UO_886 (O_886,N_13458,N_12572);
and UO_887 (O_887,N_10329,N_13467);
nand UO_888 (O_888,N_13361,N_10890);
or UO_889 (O_889,N_13759,N_13622);
or UO_890 (O_890,N_12877,N_10144);
nand UO_891 (O_891,N_13376,N_13294);
or UO_892 (O_892,N_14251,N_13596);
nor UO_893 (O_893,N_10023,N_11012);
or UO_894 (O_894,N_10038,N_12064);
and UO_895 (O_895,N_12927,N_14678);
nor UO_896 (O_896,N_14757,N_10005);
nand UO_897 (O_897,N_11699,N_13923);
nor UO_898 (O_898,N_14313,N_13915);
nor UO_899 (O_899,N_12477,N_11090);
or UO_900 (O_900,N_10385,N_13184);
nor UO_901 (O_901,N_13729,N_11736);
and UO_902 (O_902,N_10326,N_14798);
nand UO_903 (O_903,N_11923,N_13349);
and UO_904 (O_904,N_13408,N_11683);
nand UO_905 (O_905,N_12107,N_14054);
or UO_906 (O_906,N_12048,N_13152);
and UO_907 (O_907,N_10084,N_13979);
and UO_908 (O_908,N_13221,N_14887);
and UO_909 (O_909,N_12474,N_10942);
or UO_910 (O_910,N_14963,N_10440);
or UO_911 (O_911,N_10879,N_12025);
and UO_912 (O_912,N_13266,N_11974);
and UO_913 (O_913,N_13971,N_12582);
or UO_914 (O_914,N_14713,N_13110);
or UO_915 (O_915,N_11337,N_13111);
nand UO_916 (O_916,N_12684,N_11861);
nand UO_917 (O_917,N_11672,N_14734);
and UO_918 (O_918,N_13508,N_13304);
and UO_919 (O_919,N_11813,N_12293);
nand UO_920 (O_920,N_13143,N_11731);
nand UO_921 (O_921,N_12386,N_11197);
nor UO_922 (O_922,N_11279,N_13437);
and UO_923 (O_923,N_11059,N_10154);
and UO_924 (O_924,N_14779,N_14822);
nor UO_925 (O_925,N_14007,N_13790);
and UO_926 (O_926,N_13712,N_14790);
and UO_927 (O_927,N_13269,N_13188);
and UO_928 (O_928,N_14800,N_10006);
nand UO_929 (O_929,N_11423,N_13573);
or UO_930 (O_930,N_11459,N_12599);
and UO_931 (O_931,N_12855,N_12449);
nand UO_932 (O_932,N_10610,N_11784);
or UO_933 (O_933,N_14106,N_13995);
nand UO_934 (O_934,N_12470,N_12560);
or UO_935 (O_935,N_14300,N_13322);
and UO_936 (O_936,N_13393,N_12586);
or UO_937 (O_937,N_12786,N_12511);
and UO_938 (O_938,N_11248,N_13715);
and UO_939 (O_939,N_11252,N_14142);
nor UO_940 (O_940,N_12373,N_13339);
nand UO_941 (O_941,N_13933,N_10875);
nor UO_942 (O_942,N_14396,N_14257);
and UO_943 (O_943,N_14252,N_13961);
nor UO_944 (O_944,N_13515,N_13821);
nor UO_945 (O_945,N_11742,N_12396);
and UO_946 (O_946,N_13815,N_11478);
nor UO_947 (O_947,N_12905,N_12219);
and UO_948 (O_948,N_13319,N_10627);
nor UO_949 (O_949,N_13758,N_11087);
nand UO_950 (O_950,N_12937,N_11493);
and UO_951 (O_951,N_11267,N_10267);
and UO_952 (O_952,N_11823,N_10528);
nand UO_953 (O_953,N_13966,N_11351);
or UO_954 (O_954,N_14328,N_12460);
or UO_955 (O_955,N_11099,N_11799);
and UO_956 (O_956,N_11762,N_12427);
nor UO_957 (O_957,N_14600,N_13968);
or UO_958 (O_958,N_14400,N_11175);
and UO_959 (O_959,N_13901,N_12043);
and UO_960 (O_960,N_13845,N_11368);
nand UO_961 (O_961,N_13182,N_14178);
nor UO_962 (O_962,N_12114,N_13938);
nand UO_963 (O_963,N_11573,N_10539);
or UO_964 (O_964,N_10779,N_12175);
nand UO_965 (O_965,N_14680,N_14020);
nor UO_966 (O_966,N_11854,N_12592);
xnor UO_967 (O_967,N_11978,N_11327);
xnor UO_968 (O_968,N_14545,N_10390);
and UO_969 (O_969,N_13333,N_13442);
or UO_970 (O_970,N_14033,N_13054);
or UO_971 (O_971,N_13885,N_14817);
and UO_972 (O_972,N_10002,N_13387);
nand UO_973 (O_973,N_14845,N_13548);
and UO_974 (O_974,N_11618,N_11655);
or UO_975 (O_975,N_14035,N_13291);
and UO_976 (O_976,N_12510,N_14491);
and UO_977 (O_977,N_11588,N_12021);
nor UO_978 (O_978,N_13303,N_11617);
or UO_979 (O_979,N_13656,N_14027);
nand UO_980 (O_980,N_14662,N_12285);
nand UO_981 (O_981,N_11688,N_13805);
and UO_982 (O_982,N_11188,N_10564);
nor UO_983 (O_983,N_11566,N_10228);
and UO_984 (O_984,N_10828,N_11910);
and UO_985 (O_985,N_13932,N_11556);
nor UO_986 (O_986,N_13558,N_13257);
and UO_987 (O_987,N_10489,N_12127);
nand UO_988 (O_988,N_10931,N_11872);
and UO_989 (O_989,N_10873,N_14981);
and UO_990 (O_990,N_14537,N_12008);
or UO_991 (O_991,N_13237,N_11215);
and UO_992 (O_992,N_13702,N_11565);
nand UO_993 (O_993,N_11692,N_14162);
or UO_994 (O_994,N_14294,N_14197);
and UO_995 (O_995,N_10126,N_12234);
and UO_996 (O_996,N_12281,N_12004);
nand UO_997 (O_997,N_14792,N_13724);
or UO_998 (O_998,N_12103,N_11695);
nand UO_999 (O_999,N_14242,N_13285);
and UO_1000 (O_1000,N_12040,N_11403);
nand UO_1001 (O_1001,N_11241,N_13591);
or UO_1002 (O_1002,N_13791,N_10415);
or UO_1003 (O_1003,N_14360,N_12498);
nand UO_1004 (O_1004,N_11948,N_10430);
and UO_1005 (O_1005,N_11783,N_11165);
nand UO_1006 (O_1006,N_14152,N_11277);
nand UO_1007 (O_1007,N_10402,N_10092);
nor UO_1008 (O_1008,N_11443,N_14896);
or UO_1009 (O_1009,N_11290,N_10029);
nand UO_1010 (O_1010,N_13313,N_10565);
nor UO_1011 (O_1011,N_12489,N_11638);
nand UO_1012 (O_1012,N_12774,N_12232);
or UO_1013 (O_1013,N_11347,N_10951);
nand UO_1014 (O_1014,N_10140,N_10500);
nand UO_1015 (O_1015,N_11417,N_13142);
and UO_1016 (O_1016,N_11509,N_10316);
nand UO_1017 (O_1017,N_10391,N_11386);
and UO_1018 (O_1018,N_12852,N_10022);
nand UO_1019 (O_1019,N_13823,N_10397);
or UO_1020 (O_1020,N_10668,N_12992);
or UO_1021 (O_1021,N_11222,N_14428);
nor UO_1022 (O_1022,N_11925,N_10809);
nor UO_1023 (O_1023,N_11884,N_14583);
and UO_1024 (O_1024,N_13838,N_14318);
and UO_1025 (O_1025,N_10609,N_11142);
and UO_1026 (O_1026,N_11561,N_10047);
and UO_1027 (O_1027,N_12326,N_13846);
or UO_1028 (O_1028,N_10749,N_10631);
nor UO_1029 (O_1029,N_11409,N_11748);
nand UO_1030 (O_1030,N_14185,N_10586);
nand UO_1031 (O_1031,N_10661,N_13193);
or UO_1032 (O_1032,N_11756,N_11775);
or UO_1033 (O_1033,N_11666,N_12591);
and UO_1034 (O_1034,N_12762,N_10945);
nor UO_1035 (O_1035,N_11458,N_14402);
or UO_1036 (O_1036,N_11524,N_13180);
nor UO_1037 (O_1037,N_10643,N_13381);
nor UO_1038 (O_1038,N_11727,N_13174);
and UO_1039 (O_1039,N_12742,N_11432);
nor UO_1040 (O_1040,N_11009,N_11834);
or UO_1041 (O_1041,N_13853,N_10102);
nor UO_1042 (O_1042,N_12792,N_14815);
nor UO_1043 (O_1043,N_14063,N_10956);
and UO_1044 (O_1044,N_11960,N_11769);
nor UO_1045 (O_1045,N_12613,N_11849);
xnor UO_1046 (O_1046,N_14830,N_10091);
or UO_1047 (O_1047,N_11154,N_14451);
or UO_1048 (O_1048,N_14075,N_13721);
nand UO_1049 (O_1049,N_10317,N_13052);
and UO_1050 (O_1050,N_10311,N_11028);
and UO_1051 (O_1051,N_10135,N_12634);
nor UO_1052 (O_1052,N_13831,N_14168);
and UO_1053 (O_1053,N_10217,N_12401);
or UO_1054 (O_1054,N_11317,N_12198);
and UO_1055 (O_1055,N_11161,N_14323);
nand UO_1056 (O_1056,N_14791,N_11383);
nor UO_1057 (O_1057,N_12680,N_13347);
and UO_1058 (O_1058,N_14863,N_14972);
nand UO_1059 (O_1059,N_11931,N_12654);
or UO_1060 (O_1060,N_12847,N_13795);
and UO_1061 (O_1061,N_11346,N_13616);
and UO_1062 (O_1062,N_13919,N_13708);
or UO_1063 (O_1063,N_13984,N_12770);
nand UO_1064 (O_1064,N_13020,N_11698);
or UO_1065 (O_1065,N_14525,N_10949);
and UO_1066 (O_1066,N_12338,N_13676);
and UO_1067 (O_1067,N_14929,N_12675);
and UO_1068 (O_1068,N_12685,N_11976);
and UO_1069 (O_1069,N_13629,N_14538);
nor UO_1070 (O_1070,N_14837,N_11746);
nor UO_1071 (O_1071,N_12231,N_12129);
nand UO_1072 (O_1072,N_14463,N_14502);
nor UO_1073 (O_1073,N_11740,N_10346);
and UO_1074 (O_1074,N_14893,N_13829);
or UO_1075 (O_1075,N_12424,N_13571);
nor UO_1076 (O_1076,N_14483,N_11580);
or UO_1077 (O_1077,N_10213,N_14135);
nand UO_1078 (O_1078,N_11964,N_10520);
nor UO_1079 (O_1079,N_13449,N_11467);
nand UO_1080 (O_1080,N_12981,N_11191);
nand UO_1081 (O_1081,N_10976,N_11042);
and UO_1082 (O_1082,N_14589,N_10142);
and UO_1083 (O_1083,N_14000,N_11634);
and UO_1084 (O_1084,N_14899,N_12020);
or UO_1085 (O_1085,N_10185,N_12433);
nor UO_1086 (O_1086,N_11639,N_11243);
nor UO_1087 (O_1087,N_10345,N_13976);
nand UO_1088 (O_1088,N_10864,N_11498);
nand UO_1089 (O_1089,N_12294,N_13279);
or UO_1090 (O_1090,N_13265,N_11270);
nand UO_1091 (O_1091,N_11949,N_12059);
or UO_1092 (O_1092,N_12301,N_11897);
nor UO_1093 (O_1093,N_11828,N_13945);
or UO_1094 (O_1094,N_11752,N_11562);
nand UO_1095 (O_1095,N_13888,N_12539);
nor UO_1096 (O_1096,N_12384,N_11543);
and UO_1097 (O_1097,N_12108,N_13730);
or UO_1098 (O_1098,N_12823,N_13128);
or UO_1099 (O_1099,N_13468,N_13539);
nand UO_1100 (O_1100,N_10965,N_12975);
or UO_1101 (O_1101,N_12764,N_13343);
or UO_1102 (O_1102,N_11992,N_13774);
nor UO_1103 (O_1103,N_11980,N_11730);
or UO_1104 (O_1104,N_13443,N_14699);
and UO_1105 (O_1105,N_14569,N_11774);
xor UO_1106 (O_1106,N_14136,N_13873);
and UO_1107 (O_1107,N_13170,N_11599);
and UO_1108 (O_1108,N_11817,N_10663);
and UO_1109 (O_1109,N_12220,N_11965);
nand UO_1110 (O_1110,N_10165,N_13159);
or UO_1111 (O_1111,N_11534,N_11714);
nand UO_1112 (O_1112,N_12607,N_10802);
and UO_1113 (O_1113,N_10003,N_13481);
nor UO_1114 (O_1114,N_10622,N_14314);
nand UO_1115 (O_1115,N_10511,N_11414);
nor UO_1116 (O_1116,N_12056,N_12797);
or UO_1117 (O_1117,N_14064,N_10678);
and UO_1118 (O_1118,N_13670,N_10754);
nand UO_1119 (O_1119,N_12035,N_12625);
or UO_1120 (O_1120,N_13483,N_10679);
nand UO_1121 (O_1121,N_14590,N_13096);
nor UO_1122 (O_1122,N_10190,N_11786);
nor UO_1123 (O_1123,N_14767,N_10766);
or UO_1124 (O_1124,N_12491,N_12458);
and UO_1125 (O_1125,N_10967,N_12826);
nor UO_1126 (O_1126,N_10844,N_10897);
nor UO_1127 (O_1127,N_11820,N_13630);
nand UO_1128 (O_1128,N_10285,N_14879);
nand UO_1129 (O_1129,N_11070,N_11084);
or UO_1130 (O_1130,N_14844,N_13378);
nand UO_1131 (O_1131,N_12101,N_11457);
nand UO_1132 (O_1132,N_13374,N_12878);
nand UO_1133 (O_1133,N_11567,N_13905);
nor UO_1134 (O_1134,N_10748,N_13556);
and UO_1135 (O_1135,N_11015,N_14095);
or UO_1136 (O_1136,N_13528,N_12429);
nand UO_1137 (O_1137,N_11357,N_14023);
or UO_1138 (O_1138,N_14260,N_12621);
and UO_1139 (O_1139,N_11632,N_14492);
or UO_1140 (O_1140,N_14693,N_10243);
nor UO_1141 (O_1141,N_12379,N_13695);
nor UO_1142 (O_1142,N_12029,N_11987);
and UO_1143 (O_1143,N_14275,N_10111);
nand UO_1144 (O_1144,N_13642,N_14974);
nor UO_1145 (O_1145,N_11616,N_12328);
and UO_1146 (O_1146,N_13075,N_13106);
and UO_1147 (O_1147,N_13559,N_10703);
and UO_1148 (O_1148,N_13391,N_13471);
or UO_1149 (O_1149,N_13619,N_12357);
nor UO_1150 (O_1150,N_14059,N_14422);
and UO_1151 (O_1151,N_13682,N_12359);
nor UO_1152 (O_1152,N_14407,N_12825);
and UO_1153 (O_1153,N_12069,N_10883);
nor UO_1154 (O_1154,N_10156,N_12611);
nor UO_1155 (O_1155,N_14353,N_11399);
or UO_1156 (O_1156,N_14012,N_10259);
nor UO_1157 (O_1157,N_14557,N_12637);
nor UO_1158 (O_1158,N_10446,N_14724);
and UO_1159 (O_1159,N_14902,N_14919);
nand UO_1160 (O_1160,N_13858,N_13241);
nor UO_1161 (O_1161,N_13940,N_12594);
nand UO_1162 (O_1162,N_11703,N_11054);
nor UO_1163 (O_1163,N_14203,N_13589);
or UO_1164 (O_1164,N_12687,N_10871);
nor UO_1165 (O_1165,N_12872,N_11702);
nor UO_1166 (O_1166,N_12223,N_12964);
nand UO_1167 (O_1167,N_10686,N_13535);
nand UO_1168 (O_1168,N_11930,N_11057);
nor UO_1169 (O_1169,N_12144,N_12865);
nand UO_1170 (O_1170,N_13754,N_11069);
nor UO_1171 (O_1171,N_14535,N_14509);
nand UO_1172 (O_1172,N_12705,N_10205);
nor UO_1173 (O_1173,N_14729,N_11513);
nand UO_1174 (O_1174,N_10651,N_11375);
and UO_1175 (O_1175,N_11001,N_13227);
and UO_1176 (O_1176,N_10363,N_14229);
nor UO_1177 (O_1177,N_12499,N_13560);
nor UO_1178 (O_1178,N_14511,N_14702);
nor UO_1179 (O_1179,N_14546,N_12700);
or UO_1180 (O_1180,N_12910,N_13623);
nand UO_1181 (O_1181,N_10710,N_11542);
nor UO_1182 (O_1182,N_13407,N_13507);
or UO_1183 (O_1183,N_10388,N_14337);
or UO_1184 (O_1184,N_14950,N_11190);
or UO_1185 (O_1185,N_13664,N_13689);
or UO_1186 (O_1186,N_12882,N_13878);
nand UO_1187 (O_1187,N_14975,N_10350);
nand UO_1188 (O_1188,N_13353,N_14833);
nor UO_1189 (O_1189,N_14021,N_14923);
or UO_1190 (O_1190,N_13201,N_14907);
nand UO_1191 (O_1191,N_12723,N_13079);
or UO_1192 (O_1192,N_10061,N_11660);
nor UO_1193 (O_1193,N_12420,N_12939);
nor UO_1194 (O_1194,N_13562,N_11759);
and UO_1195 (O_1195,N_10863,N_12123);
or UO_1196 (O_1196,N_13396,N_14638);
nor UO_1197 (O_1197,N_10193,N_12639);
and UO_1198 (O_1198,N_11652,N_11052);
nor UO_1199 (O_1199,N_12363,N_12757);
and UO_1200 (O_1200,N_14018,N_14564);
nand UO_1201 (O_1201,N_14633,N_12881);
nor UO_1202 (O_1202,N_11722,N_13073);
and UO_1203 (O_1203,N_14708,N_11081);
nor UO_1204 (O_1204,N_13674,N_13283);
nor UO_1205 (O_1205,N_11613,N_10377);
nand UO_1206 (O_1206,N_12335,N_10573);
or UO_1207 (O_1207,N_12336,N_14660);
nor UO_1208 (O_1208,N_10765,N_14480);
or UO_1209 (O_1209,N_10567,N_14584);
and UO_1210 (O_1210,N_11915,N_11415);
nand UO_1211 (O_1211,N_11517,N_13812);
nand UO_1212 (O_1212,N_11424,N_12052);
nor UO_1213 (O_1213,N_13822,N_11821);
or UO_1214 (O_1214,N_13440,N_10250);
nand UO_1215 (O_1215,N_14776,N_13700);
and UO_1216 (O_1216,N_11975,N_12112);
nand UO_1217 (O_1217,N_13893,N_13263);
or UO_1218 (O_1218,N_12589,N_11669);
or UO_1219 (O_1219,N_13476,N_10944);
or UO_1220 (O_1220,N_12959,N_10606);
or UO_1221 (O_1221,N_10711,N_10796);
and UO_1222 (O_1222,N_14909,N_10577);
nand UO_1223 (O_1223,N_14038,N_10257);
and UO_1224 (O_1224,N_11173,N_14172);
or UO_1225 (O_1225,N_13987,N_14115);
nor UO_1226 (O_1226,N_10808,N_11546);
nand UO_1227 (O_1227,N_14227,N_13544);
and UO_1228 (O_1228,N_13665,N_11918);
nor UO_1229 (O_1229,N_14134,N_14414);
nand UO_1230 (O_1230,N_14846,N_14472);
nor UO_1231 (O_1231,N_14716,N_12308);
nand UO_1232 (O_1232,N_14236,N_11611);
or UO_1233 (O_1233,N_10366,N_14175);
and UO_1234 (O_1234,N_11115,N_13503);
or UO_1235 (O_1235,N_10324,N_12036);
nor UO_1236 (O_1236,N_14801,N_14138);
or UO_1237 (O_1237,N_11677,N_13811);
nor UO_1238 (O_1238,N_11907,N_14239);
nor UO_1239 (O_1239,N_10992,N_13046);
and UO_1240 (O_1240,N_14637,N_11555);
nand UO_1241 (O_1241,N_10087,N_14070);
or UO_1242 (O_1242,N_12479,N_12869);
nand UO_1243 (O_1243,N_13134,N_12640);
nor UO_1244 (O_1244,N_10266,N_14220);
and UO_1245 (O_1245,N_10237,N_12333);
or UO_1246 (O_1246,N_13346,N_13428);
nor UO_1247 (O_1247,N_12406,N_11610);
nand UO_1248 (O_1248,N_14613,N_11582);
nand UO_1249 (O_1249,N_14291,N_10598);
nand UO_1250 (O_1250,N_11747,N_12649);
nor UO_1251 (O_1251,N_11306,N_10481);
or UO_1252 (O_1252,N_12159,N_11395);
nor UO_1253 (O_1253,N_10588,N_10995);
and UO_1254 (O_1254,N_11622,N_14448);
or UO_1255 (O_1255,N_12361,N_12063);
nand UO_1256 (O_1256,N_10593,N_10978);
nor UO_1257 (O_1257,N_13341,N_12776);
and UO_1258 (O_1258,N_10540,N_12099);
and UO_1259 (O_1259,N_12317,N_14089);
and UO_1260 (O_1260,N_12243,N_11538);
and UO_1261 (O_1261,N_14904,N_10134);
and UO_1262 (O_1262,N_12244,N_12857);
or UO_1263 (O_1263,N_11651,N_11079);
and UO_1264 (O_1264,N_10245,N_12743);
and UO_1265 (O_1265,N_10655,N_12534);
or UO_1266 (O_1266,N_13071,N_10062);
or UO_1267 (O_1267,N_13922,N_12309);
and UO_1268 (O_1268,N_13817,N_14869);
nor UO_1269 (O_1269,N_13259,N_10550);
nor UO_1270 (O_1270,N_11726,N_11858);
nor UO_1271 (O_1271,N_10045,N_11335);
or UO_1272 (O_1272,N_10794,N_13898);
and UO_1273 (O_1273,N_14377,N_12967);
and UO_1274 (O_1274,N_10450,N_11881);
or UO_1275 (O_1275,N_12093,N_10969);
nor UO_1276 (O_1276,N_10901,N_14160);
and UO_1277 (O_1277,N_14363,N_11619);
nor UO_1278 (O_1278,N_10432,N_13505);
and UO_1279 (O_1279,N_11051,N_14503);
nand UO_1280 (O_1280,N_12593,N_10303);
or UO_1281 (O_1281,N_13737,N_10707);
nor UO_1282 (O_1282,N_13058,N_13950);
or UO_1283 (O_1283,N_10961,N_11586);
nand UO_1284 (O_1284,N_12085,N_14504);
and UO_1285 (O_1285,N_11179,N_11076);
or UO_1286 (O_1286,N_12934,N_12662);
nor UO_1287 (O_1287,N_13328,N_10049);
nor UO_1288 (O_1288,N_10068,N_11418);
or UO_1289 (O_1289,N_11122,N_10484);
and UO_1290 (O_1290,N_10247,N_13988);
and UO_1291 (O_1291,N_13645,N_14634);
nand UO_1292 (O_1292,N_12439,N_12170);
nor UO_1293 (O_1293,N_11488,N_13750);
or UO_1294 (O_1294,N_13013,N_14968);
and UO_1295 (O_1295,N_11242,N_14306);
nor UO_1296 (O_1296,N_11026,N_12751);
or UO_1297 (O_1297,N_11701,N_12464);
nor UO_1298 (O_1298,N_11635,N_13082);
nor UO_1299 (O_1299,N_11620,N_14730);
nor UO_1300 (O_1300,N_14624,N_10396);
and UO_1301 (O_1301,N_12412,N_12116);
nand UO_1302 (O_1302,N_14916,N_10319);
and UO_1303 (O_1303,N_13880,N_14516);
nand UO_1304 (O_1304,N_10954,N_10522);
and UO_1305 (O_1305,N_14737,N_14026);
or UO_1306 (O_1306,N_10688,N_14811);
nor UO_1307 (O_1307,N_13359,N_14610);
nand UO_1308 (O_1308,N_12172,N_13683);
nor UO_1309 (O_1309,N_12908,N_13943);
nand UO_1310 (O_1310,N_11092,N_11539);
and UO_1311 (O_1311,N_13826,N_13895);
and UO_1312 (O_1312,N_12952,N_10633);
nand UO_1313 (O_1313,N_10219,N_14187);
nand UO_1314 (O_1314,N_12193,N_14582);
and UO_1315 (O_1315,N_11938,N_11675);
and UO_1316 (O_1316,N_12954,N_13568);
nand UO_1317 (O_1317,N_10235,N_14931);
nor UO_1318 (O_1318,N_13963,N_12695);
nor UO_1319 (O_1319,N_14442,N_14315);
nor UO_1320 (O_1320,N_13941,N_11485);
xnor UO_1321 (O_1321,N_12078,N_12265);
nand UO_1322 (O_1322,N_13044,N_14630);
nand UO_1323 (O_1323,N_13908,N_12909);
and UO_1324 (O_1324,N_13405,N_14523);
nand UO_1325 (O_1325,N_14982,N_11196);
and UO_1326 (O_1326,N_10684,N_14746);
nand UO_1327 (O_1327,N_14522,N_14398);
or UO_1328 (O_1328,N_11579,N_11145);
nand UO_1329 (O_1329,N_14346,N_14071);
and UO_1330 (O_1330,N_12568,N_14901);
and UO_1331 (O_1331,N_13392,N_13192);
or UO_1332 (O_1332,N_11363,N_14381);
xnor UO_1333 (O_1333,N_12164,N_10209);
or UO_1334 (O_1334,N_14921,N_11295);
and UO_1335 (O_1335,N_14416,N_13711);
and UO_1336 (O_1336,N_13109,N_11186);
xnor UO_1337 (O_1337,N_12033,N_13833);
and UO_1338 (O_1338,N_12280,N_14069);
nor UO_1339 (O_1339,N_11643,N_12283);
nand UO_1340 (O_1340,N_10083,N_11141);
or UO_1341 (O_1341,N_14411,N_11944);
and UO_1342 (O_1342,N_14202,N_10977);
and UO_1343 (O_1343,N_11563,N_13464);
nor UO_1344 (O_1344,N_13579,N_13957);
and UO_1345 (O_1345,N_12060,N_14475);
and UO_1346 (O_1346,N_10950,N_14595);
nor UO_1347 (O_1347,N_12683,N_10983);
nand UO_1348 (O_1348,N_12984,N_13690);
and UO_1349 (O_1349,N_11333,N_12138);
and UO_1350 (O_1350,N_14964,N_11210);
nand UO_1351 (O_1351,N_13491,N_13510);
and UO_1352 (O_1352,N_12324,N_12233);
nor UO_1353 (O_1353,N_11342,N_12163);
nor UO_1354 (O_1354,N_14714,N_14806);
or UO_1355 (O_1355,N_13832,N_11712);
nand UO_1356 (O_1356,N_13854,N_10848);
nand UO_1357 (O_1357,N_12912,N_14700);
and UO_1358 (O_1358,N_14259,N_12627);
nor UO_1359 (O_1359,N_12150,N_11289);
and UO_1360 (O_1360,N_12136,N_14369);
and UO_1361 (O_1361,N_10352,N_13236);
nor UO_1362 (O_1362,N_11002,N_12676);
nand UO_1363 (O_1363,N_12276,N_11963);
nor UO_1364 (O_1364,N_11979,N_11454);
nand UO_1365 (O_1365,N_11287,N_12092);
or UO_1366 (O_1366,N_14766,N_11101);
or UO_1367 (O_1367,N_10335,N_10180);
and UO_1368 (O_1368,N_10086,N_11048);
nor UO_1369 (O_1369,N_11665,N_14149);
and UO_1370 (O_1370,N_14796,N_10662);
nor UO_1371 (O_1371,N_11972,N_11322);
or UO_1372 (O_1372,N_11957,N_14195);
nand UO_1373 (O_1373,N_13635,N_10223);
or UO_1374 (O_1374,N_12566,N_10525);
nor UO_1375 (O_1375,N_12346,N_10544);
or UO_1376 (O_1376,N_10116,N_14567);
nor UO_1377 (O_1377,N_13577,N_13326);
or UO_1378 (O_1378,N_13164,N_10371);
or UO_1379 (O_1379,N_14628,N_12606);
nand UO_1380 (O_1380,N_10630,N_11438);
or UO_1381 (O_1381,N_14025,N_10434);
or UO_1382 (O_1382,N_14495,N_14288);
or UO_1383 (O_1383,N_12901,N_10497);
and UO_1384 (O_1384,N_14607,N_14208);
or UO_1385 (O_1385,N_11120,N_11572);
nor UO_1386 (O_1386,N_10935,N_12497);
or UO_1387 (O_1387,N_12065,N_14642);
xnor UO_1388 (O_1388,N_13154,N_12772);
and UO_1389 (O_1389,N_14188,N_13921);
nor UO_1390 (O_1390,N_13787,N_14825);
nand UO_1391 (O_1391,N_10153,N_12918);
nor UO_1392 (O_1392,N_12174,N_10515);
nand UO_1393 (O_1393,N_10334,N_10922);
nor UO_1394 (O_1394,N_11629,N_12391);
nand UO_1395 (O_1395,N_11551,N_13131);
or UO_1396 (O_1396,N_14659,N_11844);
or UO_1397 (O_1397,N_10304,N_10756);
nor UO_1398 (O_1398,N_12289,N_12385);
nor UO_1399 (O_1399,N_10535,N_12528);
or UO_1400 (O_1400,N_14141,N_14598);
and UO_1401 (O_1401,N_12780,N_10912);
nand UO_1402 (O_1402,N_10123,N_13413);
and UO_1403 (O_1403,N_13927,N_13939);
nor UO_1404 (O_1404,N_13615,N_13231);
nor UO_1405 (O_1405,N_14467,N_11839);
or UO_1406 (O_1406,N_11842,N_14091);
nor UO_1407 (O_1407,N_13113,N_14540);
nor UO_1408 (O_1408,N_11917,N_11124);
and UO_1409 (O_1409,N_10201,N_12256);
nand UO_1410 (O_1410,N_11060,N_13137);
and UO_1411 (O_1411,N_12873,N_10987);
and UO_1412 (O_1412,N_10990,N_12656);
nor UO_1413 (O_1413,N_12211,N_11554);
and UO_1414 (O_1414,N_13222,N_14709);
nand UO_1415 (O_1415,N_13913,N_12820);
and UO_1416 (O_1416,N_14507,N_13121);
nand UO_1417 (O_1417,N_11791,N_10328);
nand UO_1418 (O_1418,N_12195,N_13745);
and UO_1419 (O_1419,N_14248,N_14347);
or UO_1420 (O_1420,N_14286,N_11958);
or UO_1421 (O_1421,N_10501,N_10547);
or UO_1422 (O_1422,N_14040,N_12925);
nor UO_1423 (O_1423,N_13993,N_10026);
or UO_1424 (O_1424,N_10119,N_11853);
nand UO_1425 (O_1425,N_14795,N_12765);
and UO_1426 (O_1426,N_14774,N_10351);
and UO_1427 (O_1427,N_11627,N_13425);
or UO_1428 (O_1428,N_12370,N_10757);
nor UO_1429 (O_1429,N_13632,N_10290);
nor UO_1430 (O_1430,N_10465,N_11603);
nand UO_1431 (O_1431,N_14640,N_13506);
or UO_1432 (O_1432,N_14758,N_10639);
nor UO_1433 (O_1433,N_14851,N_13473);
nand UO_1434 (O_1434,N_11339,N_14999);
nor UO_1435 (O_1435,N_12051,N_12549);
nor UO_1436 (O_1436,N_10000,N_11113);
or UO_1437 (O_1437,N_10130,N_13254);
nand UO_1438 (O_1438,N_12340,N_10273);
nor UO_1439 (O_1439,N_14262,N_12329);
and UO_1440 (O_1440,N_14093,N_12841);
nand UO_1441 (O_1441,N_10619,N_13934);
nand UO_1442 (O_1442,N_11305,N_10561);
and UO_1443 (O_1443,N_12014,N_13377);
or UO_1444 (O_1444,N_14900,N_14244);
or UO_1445 (O_1445,N_14311,N_14883);
or UO_1446 (O_1446,N_10090,N_12760);
nand UO_1447 (O_1447,N_12941,N_10132);
nand UO_1448 (O_1448,N_14692,N_13410);
or UO_1449 (O_1449,N_14415,N_10354);
nand UO_1450 (O_1450,N_10614,N_14058);
and UO_1451 (O_1451,N_10330,N_14679);
nor UO_1452 (O_1452,N_10916,N_11985);
nand UO_1453 (O_1453,N_13039,N_14580);
nor UO_1454 (O_1454,N_11272,N_12659);
and UO_1455 (O_1455,N_14645,N_10938);
nor UO_1456 (O_1456,N_11625,N_13953);
nand UO_1457 (O_1457,N_13808,N_11033);
nand UO_1458 (O_1458,N_13403,N_14618);
nor UO_1459 (O_1459,N_14947,N_11420);
or UO_1460 (O_1460,N_12398,N_10907);
nor UO_1461 (O_1461,N_12630,N_10488);
and UO_1462 (O_1462,N_10464,N_12819);
and UO_1463 (O_1463,N_14649,N_11512);
and UO_1464 (O_1464,N_10063,N_11410);
nor UO_1465 (O_1465,N_12670,N_11540);
or UO_1466 (O_1466,N_12131,N_11788);
or UO_1467 (O_1467,N_12266,N_12524);
or UO_1468 (O_1468,N_14126,N_11691);
or UO_1469 (O_1469,N_13027,N_12808);
or UO_1470 (O_1470,N_13040,N_12453);
or UO_1471 (O_1471,N_13438,N_14719);
nor UO_1472 (O_1472,N_11407,N_13010);
or UO_1473 (O_1473,N_13499,N_11088);
nor UO_1474 (O_1474,N_12017,N_14814);
nand UO_1475 (O_1475,N_11185,N_11119);
or UO_1476 (O_1476,N_11308,N_14823);
and UO_1477 (O_1477,N_14827,N_13153);
or UO_1478 (O_1478,N_11392,N_14957);
nand UO_1479 (O_1479,N_14051,N_13479);
nand UO_1480 (O_1480,N_14871,N_13595);
or UO_1481 (O_1481,N_12884,N_13234);
and UO_1482 (O_1482,N_14408,N_10634);
and UO_1483 (O_1483,N_12897,N_10585);
or UO_1484 (O_1484,N_14031,N_14859);
xnor UO_1485 (O_1485,N_14097,N_10926);
or UO_1486 (O_1486,N_12287,N_11144);
or UO_1487 (O_1487,N_11668,N_12997);
or UO_1488 (O_1488,N_11372,N_10508);
nor UO_1489 (O_1489,N_11393,N_10795);
and UO_1490 (O_1490,N_11776,N_11647);
and UO_1491 (O_1491,N_14510,N_13852);
nor UO_1492 (O_1492,N_12671,N_13384);
and UO_1493 (O_1493,N_12605,N_11038);
nor UO_1494 (O_1494,N_13582,N_13514);
xnor UO_1495 (O_1495,N_11253,N_12097);
or UO_1496 (O_1496,N_13782,N_13466);
nand UO_1497 (O_1497,N_13200,N_13329);
or UO_1498 (O_1498,N_11850,N_11687);
and UO_1499 (O_1499,N_10952,N_11523);
nor UO_1500 (O_1500,N_12955,N_14722);
or UO_1501 (O_1501,N_13640,N_12444);
and UO_1502 (O_1502,N_14552,N_12077);
nor UO_1503 (O_1503,N_10423,N_14706);
and UO_1504 (O_1504,N_14292,N_10409);
and UO_1505 (O_1505,N_12426,N_10885);
nor UO_1506 (O_1506,N_14335,N_10458);
nor UO_1507 (O_1507,N_13314,N_12681);
nor UO_1508 (O_1508,N_12284,N_13666);
nor UO_1509 (O_1509,N_13421,N_11460);
or UO_1510 (O_1510,N_11425,N_12561);
xnor UO_1511 (O_1511,N_10149,N_11398);
or UO_1512 (O_1512,N_10051,N_14572);
nand UO_1513 (O_1513,N_10720,N_10466);
and UO_1514 (O_1514,N_13030,N_13776);
and UO_1515 (O_1515,N_14301,N_14364);
and UO_1516 (O_1516,N_12046,N_14555);
or UO_1517 (O_1517,N_13799,N_12949);
or UO_1518 (O_1518,N_11526,N_13447);
or UO_1519 (O_1519,N_11286,N_10670);
and UO_1520 (O_1520,N_12710,N_12080);
nor UO_1521 (O_1521,N_13792,N_14109);
and UO_1522 (O_1522,N_14298,N_12236);
nand UO_1523 (O_1523,N_10716,N_10300);
nor UO_1524 (O_1524,N_12102,N_12240);
and UO_1525 (O_1525,N_10046,N_10755);
and UO_1526 (O_1526,N_13489,N_11139);
or UO_1527 (O_1527,N_12716,N_12142);
or UO_1528 (O_1528,N_10124,N_10408);
nand UO_1529 (O_1529,N_14978,N_14055);
or UO_1530 (O_1530,N_11472,N_14788);
and UO_1531 (O_1531,N_13130,N_12686);
nand UO_1532 (O_1532,N_13325,N_11892);
and UO_1533 (O_1533,N_10240,N_13986);
and UO_1534 (O_1534,N_12915,N_13409);
and UO_1535 (O_1535,N_13911,N_10127);
and UO_1536 (O_1536,N_14986,N_10676);
and UO_1537 (O_1537,N_10478,N_13699);
nand UO_1538 (O_1538,N_10118,N_14994);
nand UO_1539 (O_1539,N_14013,N_11208);
or UO_1540 (O_1540,N_10726,N_13224);
and UO_1541 (O_1541,N_14030,N_11103);
and UO_1542 (O_1542,N_11942,N_10138);
nand UO_1543 (O_1543,N_14551,N_11590);
and UO_1544 (O_1544,N_14575,N_11707);
nor UO_1545 (O_1545,N_11544,N_10653);
nor UO_1546 (O_1546,N_14150,N_13431);
or UO_1547 (O_1547,N_10640,N_11255);
nor UO_1548 (O_1548,N_10261,N_12833);
nand UO_1549 (O_1549,N_10886,N_14164);
or UO_1550 (O_1550,N_13809,N_14417);
and UO_1551 (O_1551,N_10010,N_14370);
or UO_1552 (O_1552,N_13863,N_10988);
nand UO_1553 (O_1553,N_13523,N_14303);
and UO_1554 (O_1554,N_14751,N_12787);
nand UO_1555 (O_1555,N_12366,N_14639);
nor UO_1556 (O_1556,N_13230,N_11847);
or UO_1557 (O_1557,N_10852,N_12851);
xnor UO_1558 (O_1558,N_10081,N_12360);
or UO_1559 (O_1559,N_13900,N_10017);
and UO_1560 (O_1560,N_13767,N_12137);
nand UO_1561 (O_1561,N_13534,N_12516);
and UO_1562 (O_1562,N_11445,N_11510);
and UO_1563 (O_1563,N_11671,N_10685);
or UO_1564 (O_1564,N_12463,N_12443);
and UO_1565 (O_1565,N_11766,N_11297);
and UO_1566 (O_1566,N_12169,N_10623);
nor UO_1567 (O_1567,N_10179,N_13163);
and UO_1568 (O_1568,N_10900,N_10812);
or UO_1569 (O_1569,N_13185,N_10694);
nand UO_1570 (O_1570,N_11000,N_12173);
and UO_1571 (O_1571,N_12679,N_12120);
or UO_1572 (O_1572,N_14302,N_14558);
nand UO_1573 (O_1573,N_11129,N_12974);
and UO_1574 (O_1574,N_10814,N_12814);
and UO_1575 (O_1575,N_13813,N_14215);
nor UO_1576 (O_1576,N_10553,N_13726);
and UO_1577 (O_1577,N_13890,N_14648);
and UO_1578 (O_1578,N_12641,N_14591);
and UO_1579 (O_1579,N_13417,N_14935);
nand UO_1580 (O_1580,N_11973,N_10600);
nand UO_1581 (O_1581,N_14723,N_10704);
nor UO_1582 (O_1582,N_12152,N_11780);
and UO_1583 (O_1583,N_11400,N_11829);
and UO_1584 (O_1584,N_12856,N_13062);
and UO_1585 (O_1585,N_14596,N_12480);
nand UO_1586 (O_1586,N_14721,N_14717);
or UO_1587 (O_1587,N_14224,N_11889);
or UO_1588 (O_1588,N_14380,N_12274);
nand UO_1589 (O_1589,N_11301,N_13555);
or UO_1590 (O_1590,N_14110,N_10454);
and UO_1591 (O_1591,N_12906,N_13917);
or UO_1592 (O_1592,N_14199,N_12483);
and UO_1593 (O_1593,N_12744,N_14424);
nand UO_1594 (O_1594,N_14154,N_13427);
nand UO_1595 (O_1595,N_11664,N_10048);
nand UO_1596 (O_1596,N_14117,N_12201);
nor UO_1597 (O_1597,N_14718,N_10538);
nor UO_1598 (O_1598,N_12616,N_14937);
nand UO_1599 (O_1599,N_12358,N_14238);
and UO_1600 (O_1600,N_10899,N_12075);
nand UO_1601 (O_1601,N_12938,N_12354);
or UO_1602 (O_1602,N_12485,N_10089);
or UO_1603 (O_1603,N_13652,N_12374);
nand UO_1604 (O_1604,N_13035,N_10940);
or UO_1605 (O_1605,N_11693,N_13411);
or UO_1606 (O_1606,N_10181,N_10698);
and UO_1607 (O_1607,N_11452,N_13324);
or UO_1608 (O_1608,N_12545,N_11086);
nor UO_1609 (O_1609,N_10031,N_12207);
nand UO_1610 (O_1610,N_11098,N_12580);
or UO_1611 (O_1611,N_12758,N_11044);
or UO_1612 (O_1612,N_10847,N_11078);
or UO_1613 (O_1613,N_11816,N_14864);
nand UO_1614 (O_1614,N_11260,N_11971);
or UO_1615 (O_1615,N_11623,N_11794);
and UO_1616 (O_1616,N_14911,N_10699);
and UO_1617 (O_1617,N_11233,N_12024);
and UO_1618 (O_1618,N_14473,N_14905);
or UO_1619 (O_1619,N_12547,N_14009);
and UO_1620 (O_1620,N_13866,N_11329);
nand UO_1621 (O_1621,N_14882,N_13308);
or UO_1622 (O_1622,N_11809,N_12921);
and UO_1623 (O_1623,N_13538,N_14405);
or UO_1624 (O_1624,N_11993,N_12327);
and UO_1625 (O_1625,N_12473,N_13455);
nand UO_1626 (O_1626,N_10648,N_12697);
nor UO_1627 (O_1627,N_14958,N_12087);
nor UO_1628 (O_1628,N_10647,N_11489);
nand UO_1629 (O_1629,N_12859,N_10365);
nand UO_1630 (O_1630,N_12269,N_14223);
nand UO_1631 (O_1631,N_13189,N_12018);
nand UO_1632 (O_1632,N_10706,N_13126);
nand UO_1633 (O_1633,N_14547,N_14623);
nor UO_1634 (O_1634,N_13931,N_12045);
nand UO_1635 (O_1635,N_14435,N_12297);
nor UO_1636 (O_1636,N_14177,N_11049);
nor UO_1637 (O_1637,N_12235,N_11533);
or UO_1638 (O_1638,N_13828,N_13331);
and UO_1639 (O_1639,N_14062,N_11758);
nor UO_1640 (O_1640,N_11247,N_14376);
xnor UO_1641 (O_1641,N_12192,N_13537);
or UO_1642 (O_1642,N_11106,N_11935);
nor UO_1643 (O_1643,N_10318,N_13229);
and UO_1644 (O_1644,N_14388,N_12947);
nand UO_1645 (O_1645,N_13203,N_14412);
nor UO_1646 (O_1646,N_10189,N_12278);
nor UO_1647 (O_1647,N_10632,N_10443);
nor UO_1648 (O_1648,N_13078,N_14212);
and UO_1649 (O_1649,N_12923,N_10801);
and UO_1650 (O_1650,N_12389,N_12397);
nand UO_1651 (O_1651,N_11025,N_12548);
or UO_1652 (O_1652,N_14268,N_10357);
and UO_1653 (O_1653,N_12407,N_12870);
nor UO_1654 (O_1654,N_14563,N_10555);
nor UO_1655 (O_1655,N_10556,N_10674);
or UO_1656 (O_1656,N_12117,N_12505);
or UO_1657 (O_1657,N_12666,N_10937);
and UO_1658 (O_1658,N_12652,N_10364);
and UO_1659 (O_1659,N_10356,N_10331);
nor UO_1660 (O_1660,N_12512,N_12660);
nor UO_1661 (O_1661,N_13077,N_11779);
and UO_1662 (O_1662,N_14843,N_12076);
or UO_1663 (O_1663,N_12322,N_11334);
or UO_1664 (O_1664,N_10558,N_12100);
nand UO_1665 (O_1665,N_12251,N_10941);
nand UO_1666 (O_1666,N_11112,N_11095);
nand UO_1667 (O_1667,N_14641,N_12574);
xnor UO_1668 (O_1668,N_13612,N_10671);
or UO_1669 (O_1669,N_11550,N_14101);
nor UO_1670 (O_1670,N_12692,N_13457);
or UO_1671 (O_1671,N_10232,N_12781);
nor UO_1672 (O_1672,N_14755,N_11626);
and UO_1673 (O_1673,N_11379,N_10612);
or UO_1674 (O_1674,N_13891,N_14336);
or UO_1675 (O_1675,N_12725,N_14918);
nor UO_1676 (O_1676,N_11700,N_13240);
and UO_1677 (O_1677,N_11571,N_13012);
or UO_1678 (O_1678,N_10380,N_12874);
nand UO_1679 (O_1679,N_12090,N_12690);
and UO_1680 (O_1680,N_13788,N_12105);
nand UO_1681 (O_1681,N_12130,N_12525);
and UO_1682 (O_1682,N_12484,N_13296);
and UO_1683 (O_1683,N_13002,N_13956);
or UO_1684 (O_1684,N_10773,N_10878);
nor UO_1685 (O_1685,N_13924,N_11431);
or UO_1686 (O_1686,N_12190,N_14088);
or UO_1687 (O_1687,N_14625,N_13127);
nand UO_1688 (O_1688,N_11157,N_12019);
or UO_1689 (O_1689,N_11416,N_10971);
nand UO_1690 (O_1690,N_13756,N_12111);
nor UO_1691 (O_1691,N_11989,N_11354);
and UO_1692 (O_1692,N_11797,N_10456);
or UO_1693 (O_1693,N_14163,N_13360);
and UO_1694 (O_1694,N_10827,N_14194);
xnor UO_1695 (O_1695,N_11390,N_11841);
and UO_1696 (O_1696,N_11378,N_14839);
nor UO_1697 (O_1697,N_10435,N_14421);
nand UO_1698 (O_1698,N_12838,N_11228);
or UO_1699 (O_1699,N_13335,N_11583);
or UO_1700 (O_1700,N_10077,N_12228);
nand UO_1701 (O_1701,N_12664,N_11514);
nand UO_1702 (O_1702,N_11006,N_10624);
or UO_1703 (O_1703,N_13053,N_10108);
and UO_1704 (O_1704,N_14066,N_11412);
and UO_1705 (O_1705,N_14754,N_13600);
nor UO_1706 (O_1706,N_13255,N_11852);
or UO_1707 (O_1707,N_13197,N_14926);
nand UO_1708 (O_1708,N_13800,N_13004);
or UO_1709 (O_1709,N_11966,N_12850);
nand UO_1710 (O_1710,N_13613,N_11097);
or UO_1711 (O_1711,N_11265,N_12541);
or UO_1712 (O_1712,N_13617,N_13719);
or UO_1713 (O_1713,N_12620,N_14881);
and UO_1714 (O_1714,N_13000,N_11109);
nor UO_1715 (O_1715,N_10204,N_10483);
or UO_1716 (O_1716,N_13731,N_11600);
and UO_1717 (O_1717,N_11697,N_10428);
nor UO_1718 (O_1718,N_13049,N_12588);
and UO_1719 (O_1719,N_10302,N_13080);
nor UO_1720 (O_1720,N_13607,N_13883);
nand UO_1721 (O_1721,N_12221,N_13497);
nand UO_1722 (O_1722,N_14782,N_12754);
nor UO_1723 (O_1723,N_14556,N_10881);
nand UO_1724 (O_1724,N_11908,N_10932);
nor UO_1725 (O_1725,N_12636,N_13877);
or UO_1726 (O_1726,N_12896,N_14249);
nor UO_1727 (O_1727,N_12200,N_14243);
or UO_1728 (O_1728,N_11264,N_13429);
nor UO_1729 (O_1729,N_13223,N_13100);
nand UO_1730 (O_1730,N_11704,N_12440);
or UO_1731 (O_1731,N_11919,N_12887);
nand UO_1732 (O_1732,N_11282,N_12438);
nor UO_1733 (O_1733,N_10277,N_14211);
or UO_1734 (O_1734,N_11936,N_10581);
or UO_1735 (O_1735,N_13850,N_14553);
nor UO_1736 (O_1736,N_14247,N_10910);
or UO_1737 (O_1737,N_12987,N_14324);
or UO_1738 (O_1738,N_10767,N_11449);
nor UO_1739 (O_1739,N_12459,N_13651);
nor UO_1740 (O_1740,N_13169,N_12527);
or UO_1741 (O_1741,N_12038,N_11798);
or UO_1742 (O_1742,N_12651,N_10629);
or UO_1743 (O_1743,N_10155,N_13465);
nor UO_1744 (O_1744,N_14037,N_11685);
and UO_1745 (O_1745,N_12062,N_10645);
or UO_1746 (O_1746,N_13023,N_14269);
and UO_1747 (O_1747,N_13354,N_10709);
nor UO_1748 (O_1748,N_12415,N_14176);
nand UO_1749 (O_1749,N_12638,N_13570);
and UO_1750 (O_1750,N_14453,N_14355);
nand UO_1751 (O_1751,N_13837,N_13327);
nor UO_1752 (O_1752,N_10524,N_10874);
or UO_1753 (O_1753,N_13196,N_14533);
or UO_1754 (O_1754,N_12273,N_10841);
and UO_1755 (O_1755,N_11283,N_14123);
nor UO_1756 (O_1756,N_14784,N_13072);
and UO_1757 (O_1757,N_10229,N_14763);
nand UO_1758 (O_1758,N_11207,N_10936);
nand UO_1759 (O_1759,N_11913,N_13906);
and UO_1760 (O_1760,N_10532,N_10269);
or UO_1761 (O_1761,N_11016,N_13981);
and UO_1762 (O_1762,N_11249,N_13604);
nand UO_1763 (O_1763,N_14884,N_14036);
and UO_1764 (O_1764,N_14960,N_10276);
nor UO_1765 (O_1765,N_12858,N_13362);
or UO_1766 (O_1766,N_14357,N_12088);
or UO_1767 (O_1767,N_10362,N_12537);
and UO_1768 (O_1768,N_14295,N_13744);
nor UO_1769 (O_1769,N_14941,N_11172);
and UO_1770 (O_1770,N_10677,N_10395);
or UO_1771 (O_1771,N_12968,N_14045);
and UO_1772 (O_1772,N_12986,N_10659);
nand UO_1773 (O_1773,N_13970,N_13383);
nand UO_1774 (O_1774,N_10620,N_14860);
and UO_1775 (O_1775,N_13704,N_14092);
and UO_1776 (O_1776,N_11238,N_14330);
nor UO_1777 (O_1777,N_14427,N_13728);
and UO_1778 (O_1778,N_14894,N_10798);
nand UO_1779 (O_1779,N_13094,N_13060);
nor UO_1780 (O_1780,N_13843,N_13432);
nand UO_1781 (O_1781,N_14218,N_13942);
nand UO_1782 (O_1782,N_11385,N_12708);
nor UO_1783 (O_1783,N_14616,N_11814);
nor UO_1784 (O_1784,N_12414,N_12807);
nor UO_1785 (O_1785,N_14928,N_14065);
nand UO_1786 (O_1786,N_10822,N_11053);
or UO_1787 (O_1787,N_14954,N_14145);
nor UO_1788 (O_1788,N_11018,N_13859);
nor UO_1789 (O_1789,N_10264,N_14611);
nand UO_1790 (O_1790,N_13412,N_12013);
and UO_1791 (O_1791,N_13603,N_14245);
or UO_1792 (O_1792,N_13088,N_12691);
nand UO_1793 (O_1793,N_11447,N_10383);
nand UO_1794 (O_1794,N_12450,N_13123);
nor UO_1795 (O_1795,N_13496,N_11083);
or UO_1796 (O_1796,N_11678,N_12583);
and UO_1797 (O_1797,N_12364,N_12535);
nand UO_1798 (O_1798,N_11606,N_11246);
nand UO_1799 (O_1799,N_12507,N_13806);
and UO_1800 (O_1800,N_10413,N_11235);
nor UO_1801 (O_1801,N_11143,N_12422);
xnor UO_1802 (O_1802,N_12737,N_10981);
or UO_1803 (O_1803,N_14196,N_13999);
nand UO_1804 (O_1804,N_10429,N_10476);
or UO_1805 (O_1805,N_12348,N_14888);
nand UO_1806 (O_1806,N_13256,N_13166);
nand UO_1807 (O_1807,N_14452,N_14371);
or UO_1808 (O_1808,N_14865,N_10903);
and UO_1809 (O_1809,N_11320,N_13364);
nand UO_1810 (O_1810,N_14759,N_10173);
or UO_1811 (O_1811,N_14910,N_14520);
nand UO_1812 (O_1812,N_12793,N_10095);
and UO_1813 (O_1813,N_13849,N_13804);
nand UO_1814 (O_1814,N_12721,N_12513);
and UO_1815 (O_1815,N_10074,N_11871);
and UO_1816 (O_1816,N_10174,N_10752);
xor UO_1817 (O_1817,N_10839,N_12215);
or UO_1818 (O_1818,N_14740,N_12371);
nand UO_1819 (O_1819,N_12995,N_14272);
nand UO_1820 (O_1820,N_10537,N_13748);
nand UO_1821 (O_1821,N_11114,N_11091);
and UO_1822 (O_1822,N_13463,N_14543);
nor UO_1823 (O_1823,N_10160,N_12778);
nand UO_1824 (O_1824,N_11836,N_10420);
nor UO_1825 (O_1825,N_12098,N_10536);
nand UO_1826 (O_1826,N_13009,N_10993);
nand UO_1827 (O_1827,N_10141,N_13914);
nand UO_1828 (O_1828,N_12154,N_11656);
nor UO_1829 (O_1829,N_10469,N_14094);
nor UO_1830 (O_1830,N_13475,N_14658);
and UO_1831 (O_1831,N_12349,N_14425);
and UO_1832 (O_1832,N_12565,N_10920);
nand UO_1833 (O_1833,N_10073,N_13992);
and UO_1834 (O_1834,N_11831,N_11757);
nand UO_1835 (O_1835,N_11440,N_12001);
or UO_1836 (O_1836,N_12738,N_10837);
and UO_1837 (O_1837,N_14621,N_11901);
and UO_1838 (O_1838,N_10401,N_14077);
or UO_1839 (O_1839,N_13989,N_12552);
nor UO_1840 (O_1840,N_12894,N_12809);
nand UO_1841 (O_1841,N_11732,N_12813);
nor UO_1842 (O_1842,N_10096,N_11217);
and UO_1843 (O_1843,N_10761,N_12966);
nor UO_1844 (O_1844,N_13951,N_13460);
or UO_1845 (O_1845,N_12777,N_10475);
and UO_1846 (O_1846,N_14373,N_13780);
and UO_1847 (O_1847,N_10016,N_14487);
nand UO_1848 (O_1848,N_12246,N_14482);
and UO_1849 (O_1849,N_14304,N_14821);
nor UO_1850 (O_1850,N_14081,N_10131);
nor UO_1851 (O_1851,N_13357,N_10382);
and UO_1852 (O_1852,N_12418,N_12564);
nand UO_1853 (O_1853,N_12993,N_10546);
and UO_1854 (O_1854,N_10078,N_13400);
or UO_1855 (O_1855,N_10496,N_14812);
nor UO_1856 (O_1856,N_12165,N_10386);
nor UO_1857 (O_1857,N_12965,N_10172);
or UO_1858 (O_1858,N_14310,N_11437);
nand UO_1859 (O_1859,N_12179,N_14183);
and UO_1860 (O_1860,N_12622,N_11209);
or UO_1861 (O_1861,N_14670,N_10517);
nor UO_1862 (O_1862,N_13034,N_10374);
nand UO_1863 (O_1863,N_10393,N_14550);
nor UO_1864 (O_1864,N_11017,N_12971);
nor UO_1865 (O_1865,N_10806,N_11075);
nor UO_1866 (O_1866,N_12994,N_11832);
and UO_1867 (O_1867,N_14880,N_11856);
and UO_1868 (O_1868,N_14605,N_14787);
nand UO_1869 (O_1869,N_14057,N_13307);
or UO_1870 (O_1870,N_13070,N_11421);
nand UO_1871 (O_1871,N_11466,N_14113);
or UO_1872 (O_1872,N_10075,N_12305);
nor UO_1873 (O_1873,N_12247,N_10616);
nor UO_1874 (O_1874,N_12044,N_12733);
and UO_1875 (O_1875,N_12146,N_11684);
nand UO_1876 (O_1876,N_14855,N_10596);
nor UO_1877 (O_1877,N_14348,N_11178);
and UO_1878 (O_1878,N_11323,N_12390);
nor UO_1879 (O_1879,N_10436,N_10858);
and UO_1880 (O_1880,N_10948,N_12455);
nor UO_1881 (O_1881,N_14193,N_13512);
and UO_1882 (O_1882,N_13869,N_11630);
nor UO_1883 (O_1883,N_14671,N_11148);
or UO_1884 (O_1884,N_13910,N_11778);
nor UO_1885 (O_1885,N_13118,N_14433);
nor UO_1886 (O_1886,N_13207,N_11777);
nand UO_1887 (O_1887,N_13659,N_11299);
nor UO_1888 (O_1888,N_11584,N_11903);
and UO_1889 (O_1889,N_13892,N_11031);
or UO_1890 (O_1890,N_10743,N_14015);
nand UO_1891 (O_1891,N_13649,N_11494);
nor UO_1892 (O_1892,N_12554,N_13694);
and UO_1893 (O_1893,N_11376,N_11450);
nor UO_1894 (O_1894,N_13014,N_14308);
and UO_1895 (O_1895,N_12145,N_10826);
or UO_1896 (O_1896,N_11462,N_12213);
and UO_1897 (O_1897,N_12600,N_10712);
nor UO_1898 (O_1898,N_14987,N_10644);
nand UO_1899 (O_1899,N_12945,N_12696);
or UO_1900 (O_1900,N_11356,N_12929);
nor UO_1901 (O_1901,N_12998,N_11085);
nor UO_1902 (O_1902,N_14447,N_10973);
nor UO_1903 (O_1903,N_13389,N_12766);
or UO_1904 (O_1904,N_13836,N_11662);
nand UO_1905 (O_1905,N_10909,N_13480);
and UO_1906 (O_1906,N_11397,N_10182);
xnor UO_1907 (O_1907,N_14394,N_10137);
nor UO_1908 (O_1908,N_12665,N_13352);
and UO_1909 (O_1909,N_14952,N_11718);
and UO_1910 (O_1910,N_11962,N_11370);
and UO_1911 (O_1911,N_13593,N_14561);
nand UO_1912 (O_1912,N_10895,N_11332);
or UO_1913 (O_1913,N_10611,N_10321);
or UO_1914 (O_1914,N_12515,N_11461);
and UO_1915 (O_1915,N_10788,N_11644);
nand UO_1916 (O_1916,N_14319,N_13739);
nor UO_1917 (O_1917,N_13532,N_10813);
nand UO_1918 (O_1918,N_13043,N_10192);
and UO_1919 (O_1919,N_14374,N_11232);
and UO_1920 (O_1920,N_14445,N_14786);
nand UO_1921 (O_1921,N_11710,N_10242);
and UO_1922 (O_1922,N_11292,N_14528);
nor UO_1923 (O_1923,N_12380,N_11497);
nor UO_1924 (O_1924,N_11435,N_11689);
or UO_1925 (O_1925,N_10877,N_10534);
and UO_1926 (O_1926,N_14241,N_10999);
xor UO_1927 (O_1927,N_11180,N_10820);
or UO_1928 (O_1928,N_10361,N_13086);
nand UO_1929 (O_1929,N_11133,N_12185);
or UO_1930 (O_1930,N_11239,N_14988);
and UO_1931 (O_1931,N_12663,N_10221);
nand UO_1932 (O_1932,N_14132,N_13669);
nand UO_1933 (O_1933,N_13874,N_12312);
and UO_1934 (O_1934,N_10753,N_10502);
nor UO_1935 (O_1935,N_11149,N_12533);
and UO_1936 (O_1936,N_11177,N_10238);
nor UO_1937 (O_1937,N_10917,N_14951);
and UO_1938 (O_1938,N_13472,N_13379);
nor UO_1939 (O_1939,N_12672,N_14726);
and UO_1940 (O_1940,N_10499,N_10479);
nand UO_1941 (O_1941,N_14878,N_12161);
nand UO_1942 (O_1942,N_14299,N_10197);
xnor UO_1943 (O_1943,N_14527,N_13249);
or UO_1944 (O_1944,N_13985,N_11977);
and UO_1945 (O_1945,N_10392,N_11203);
nor UO_1946 (O_1946,N_10664,N_11811);
and UO_1947 (O_1947,N_12893,N_10288);
nand UO_1948 (O_1948,N_14462,N_10687);
or UO_1949 (O_1949,N_14082,N_10759);
or UO_1950 (O_1950,N_12388,N_10194);
nor UO_1951 (O_1951,N_13530,N_10853);
or UO_1952 (O_1952,N_14917,N_13498);
nor UO_1953 (O_1953,N_11468,N_12735);
nor UO_1954 (O_1954,N_12928,N_14666);
nand UO_1955 (O_1955,N_13418,N_14588);
and UO_1956 (O_1956,N_12041,N_12007);
and UO_1957 (O_1957,N_10740,N_10888);
and UO_1958 (O_1958,N_14570,N_11961);
and UO_1959 (O_1959,N_14043,N_10218);
nand UO_1960 (O_1960,N_13972,N_13772);
nor UO_1961 (O_1961,N_13211,N_14047);
or UO_1962 (O_1962,N_14632,N_13089);
nand UO_1963 (O_1963,N_10287,N_10152);
nor UO_1964 (O_1964,N_10980,N_13318);
or UO_1965 (O_1965,N_12404,N_11621);
or UO_1966 (O_1966,N_10760,N_14534);
nor UO_1967 (O_1967,N_10114,N_10751);
xor UO_1968 (O_1968,N_13586,N_11734);
or UO_1969 (O_1969,N_10552,N_12332);
and UO_1970 (O_1970,N_11715,N_12047);
and UO_1971 (O_1971,N_13733,N_14539);
nand UO_1972 (O_1972,N_14283,N_14056);
or UO_1973 (O_1973,N_12156,N_10169);
nor UO_1974 (O_1974,N_10055,N_13338);
nand UO_1975 (O_1975,N_12655,N_12836);
nor UO_1976 (O_1976,N_12028,N_14519);
nor UO_1977 (O_1977,N_10256,N_11723);
nand UO_1978 (O_1978,N_11174,N_11578);
nand UO_1979 (O_1979,N_13398,N_10527);
or UO_1980 (O_1980,N_11071,N_12520);
nor UO_1981 (O_1981,N_12827,N_13340);
and UO_1982 (O_1982,N_14450,N_13067);
nand UO_1983 (O_1983,N_12991,N_14603);
or UO_1984 (O_1984,N_12387,N_12203);
nor UO_1985 (O_1985,N_14389,N_10306);
nor UO_1986 (O_1986,N_13202,N_14756);
and UO_1987 (O_1987,N_14674,N_12058);
nand UO_1988 (O_1988,N_10406,N_14593);
and UO_1989 (O_1989,N_11929,N_12347);
or UO_1990 (O_1990,N_10531,N_13371);
and UO_1991 (O_1991,N_10831,N_10889);
nand UO_1992 (O_1992,N_10571,N_14204);
or UO_1993 (O_1993,N_10772,N_11061);
nand UO_1994 (O_1994,N_10158,N_14842);
nor UO_1995 (O_1995,N_14438,N_12707);
nor UO_1996 (O_1996,N_12775,N_13594);
and UO_1997 (O_1997,N_14395,N_10818);
or UO_1998 (O_1998,N_10960,N_10955);
and UO_1999 (O_1999,N_12249,N_10359);
endmodule