module basic_1000_10000_1500_5_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_731,In_22);
and U1 (N_1,In_428,In_880);
nand U2 (N_2,In_20,In_264);
and U3 (N_3,In_738,In_804);
or U4 (N_4,In_158,In_183);
or U5 (N_5,In_904,In_90);
or U6 (N_6,In_418,In_571);
nand U7 (N_7,In_956,In_859);
nor U8 (N_8,In_226,In_822);
and U9 (N_9,In_285,In_197);
nor U10 (N_10,In_11,In_792);
nor U11 (N_11,In_934,In_424);
and U12 (N_12,In_576,In_188);
or U13 (N_13,In_533,In_42);
nor U14 (N_14,In_797,In_714);
nand U15 (N_15,In_658,In_460);
and U16 (N_16,In_456,In_775);
or U17 (N_17,In_106,In_884);
nor U18 (N_18,In_132,In_139);
and U19 (N_19,In_899,In_490);
xor U20 (N_20,In_772,In_575);
nand U21 (N_21,In_830,In_19);
nor U22 (N_22,In_718,In_290);
or U23 (N_23,In_782,In_971);
or U24 (N_24,In_427,In_500);
and U25 (N_25,In_109,In_558);
nor U26 (N_26,In_610,In_778);
or U27 (N_27,In_431,In_279);
or U28 (N_28,In_31,In_517);
nor U29 (N_29,In_839,In_511);
and U30 (N_30,In_389,In_849);
or U31 (N_31,In_667,In_773);
or U32 (N_32,In_137,In_946);
and U33 (N_33,In_278,In_256);
and U34 (N_34,In_958,In_660);
nand U35 (N_35,In_873,In_524);
or U36 (N_36,In_84,In_855);
or U37 (N_37,In_259,In_229);
or U38 (N_38,In_730,In_846);
nand U39 (N_39,In_294,In_851);
nand U40 (N_40,In_193,In_916);
nand U41 (N_41,In_326,In_777);
and U42 (N_42,In_65,In_210);
or U43 (N_43,In_143,In_895);
or U44 (N_44,In_636,In_239);
nand U45 (N_45,In_66,In_888);
or U46 (N_46,In_759,In_117);
nor U47 (N_47,In_567,In_9);
nor U48 (N_48,In_268,In_453);
nor U49 (N_49,In_573,In_196);
nand U50 (N_50,In_876,In_982);
or U51 (N_51,In_754,In_497);
nor U52 (N_52,In_414,In_273);
or U53 (N_53,In_732,In_371);
nand U54 (N_54,In_920,In_905);
and U55 (N_55,In_823,In_409);
and U56 (N_56,In_26,In_421);
and U57 (N_57,In_400,In_875);
nor U58 (N_58,In_100,In_581);
and U59 (N_59,In_672,In_441);
or U60 (N_60,In_81,In_225);
or U61 (N_61,In_911,In_858);
nor U62 (N_62,In_391,In_551);
or U63 (N_63,In_108,In_646);
nor U64 (N_64,In_844,In_145);
or U65 (N_65,In_795,In_962);
and U66 (N_66,In_34,In_518);
or U67 (N_67,In_960,In_590);
nand U68 (N_68,In_640,In_645);
and U69 (N_69,In_36,In_944);
nor U70 (N_70,In_564,In_122);
or U71 (N_71,In_638,In_121);
nor U72 (N_72,In_639,In_127);
or U73 (N_73,In_402,In_311);
nor U74 (N_74,In_726,In_211);
and U75 (N_75,In_419,In_779);
nor U76 (N_76,In_396,In_350);
nand U77 (N_77,In_938,In_970);
or U78 (N_78,In_545,In_356);
nand U79 (N_79,In_522,In_801);
nor U80 (N_80,In_88,In_788);
and U81 (N_81,In_556,In_976);
or U82 (N_82,In_274,In_961);
nor U83 (N_83,In_159,In_783);
or U84 (N_84,In_458,In_119);
nand U85 (N_85,In_483,In_891);
or U86 (N_86,In_979,In_434);
nand U87 (N_87,In_77,In_463);
and U88 (N_88,In_711,In_998);
and U89 (N_89,In_848,In_198);
and U90 (N_90,In_530,In_491);
nand U91 (N_91,In_260,In_536);
nor U92 (N_92,In_896,In_351);
xor U93 (N_93,In_984,In_488);
or U94 (N_94,In_746,In_663);
and U95 (N_95,In_236,In_459);
and U96 (N_96,In_771,In_37);
or U97 (N_97,In_325,In_697);
nor U98 (N_98,In_552,In_887);
nor U99 (N_99,In_302,In_769);
nor U100 (N_100,In_366,In_446);
or U101 (N_101,In_331,In_316);
and U102 (N_102,In_923,In_681);
nor U103 (N_103,In_698,In_761);
nor U104 (N_104,In_76,In_883);
or U105 (N_105,In_364,In_49);
xnor U106 (N_106,In_149,In_69);
nor U107 (N_107,In_717,In_255);
and U108 (N_108,In_58,In_526);
nor U109 (N_109,In_954,In_622);
or U110 (N_110,In_104,In_365);
nor U111 (N_111,In_950,In_128);
or U112 (N_112,In_856,In_153);
nand U113 (N_113,In_678,In_355);
and U114 (N_114,In_941,In_444);
nor U115 (N_115,In_12,In_582);
nand U116 (N_116,In_919,In_955);
or U117 (N_117,In_560,In_947);
nand U118 (N_118,In_252,In_367);
and U119 (N_119,In_447,In_130);
and U120 (N_120,In_164,In_606);
and U121 (N_121,In_393,In_379);
nand U122 (N_122,In_872,In_413);
nand U123 (N_123,In_245,In_482);
and U124 (N_124,In_764,In_963);
nor U125 (N_125,In_965,In_794);
and U126 (N_126,In_468,In_123);
or U127 (N_127,In_257,In_177);
or U128 (N_128,In_643,In_83);
and U129 (N_129,In_692,In_803);
or U130 (N_130,In_319,In_230);
nand U131 (N_131,In_907,In_825);
nand U132 (N_132,In_261,In_175);
nand U133 (N_133,In_918,In_339);
and U134 (N_134,In_91,In_605);
and U135 (N_135,In_702,In_683);
nand U136 (N_136,In_641,In_470);
nand U137 (N_137,In_719,In_212);
nand U138 (N_138,In_398,In_99);
nor U139 (N_139,In_890,In_248);
or U140 (N_140,In_628,In_116);
or U141 (N_141,In_502,In_324);
nor U142 (N_142,In_345,In_834);
or U143 (N_143,In_996,In_602);
and U144 (N_144,In_332,In_360);
and U145 (N_145,In_922,In_29);
and U146 (N_146,In_190,In_312);
or U147 (N_147,In_288,In_748);
nand U148 (N_148,In_908,In_112);
and U149 (N_149,In_3,In_785);
nor U150 (N_150,In_675,In_724);
or U151 (N_151,In_43,In_301);
or U152 (N_152,In_320,In_654);
nand U153 (N_153,In_185,In_781);
or U154 (N_154,In_569,In_28);
or U155 (N_155,In_713,In_271);
or U156 (N_156,In_964,In_999);
and U157 (N_157,In_705,In_227);
nand U158 (N_158,In_725,In_932);
nor U159 (N_159,In_46,In_203);
nand U160 (N_160,In_747,In_587);
or U161 (N_161,In_852,In_498);
or U162 (N_162,In_160,In_712);
nand U163 (N_163,In_342,In_790);
or U164 (N_164,In_816,In_494);
nor U165 (N_165,In_977,In_2);
and U166 (N_166,In_450,In_72);
or U167 (N_167,In_579,In_512);
nor U168 (N_168,In_27,In_357);
or U169 (N_169,In_716,In_180);
nor U170 (N_170,In_352,In_611);
nor U171 (N_171,In_568,In_704);
and U172 (N_172,In_340,In_94);
nor U173 (N_173,In_809,In_666);
nand U174 (N_174,In_669,In_637);
nor U175 (N_175,In_644,In_687);
or U176 (N_176,In_63,In_559);
nand U177 (N_177,In_410,In_334);
nor U178 (N_178,In_975,In_862);
or U179 (N_179,In_519,In_457);
and U180 (N_180,In_59,In_565);
or U181 (N_181,In_737,In_169);
and U182 (N_182,In_251,In_656);
nor U183 (N_183,In_449,In_865);
and U184 (N_184,In_433,In_881);
or U185 (N_185,In_47,In_496);
nand U186 (N_186,In_609,In_394);
and U187 (N_187,In_987,In_86);
nor U188 (N_188,In_843,In_758);
nand U189 (N_189,In_613,In_89);
nand U190 (N_190,In_44,In_195);
and U191 (N_191,In_362,In_744);
and U192 (N_192,In_329,In_328);
and U193 (N_193,In_600,In_632);
nand U194 (N_194,In_743,In_485);
and U195 (N_195,In_313,In_385);
and U196 (N_196,In_115,In_201);
or U197 (N_197,In_405,In_280);
nand U198 (N_198,In_82,In_943);
nor U199 (N_199,In_240,In_793);
nor U200 (N_200,In_237,In_707);
nand U201 (N_201,In_384,In_307);
nand U202 (N_202,In_527,In_674);
or U203 (N_203,In_817,In_513);
or U204 (N_204,In_528,In_506);
or U205 (N_205,In_52,In_953);
and U206 (N_206,In_415,In_933);
nor U207 (N_207,In_734,In_436);
and U208 (N_208,In_550,In_157);
nand U209 (N_209,In_736,In_467);
and U210 (N_210,In_819,In_299);
or U211 (N_211,In_756,In_648);
or U212 (N_212,In_924,In_516);
nor U213 (N_213,In_995,In_75);
nor U214 (N_214,In_749,In_266);
nand U215 (N_215,In_780,In_570);
nor U216 (N_216,In_204,In_836);
and U217 (N_217,In_207,In_649);
and U218 (N_218,In_254,In_805);
nor U219 (N_219,In_623,In_18);
nor U220 (N_220,In_532,In_474);
nor U221 (N_221,In_304,In_912);
and U222 (N_222,In_8,In_306);
or U223 (N_223,In_437,In_466);
and U224 (N_224,In_471,In_287);
and U225 (N_225,In_105,In_189);
and U226 (N_226,In_231,In_464);
nor U227 (N_227,In_930,In_68);
nor U228 (N_228,In_727,In_79);
nand U229 (N_229,In_293,In_853);
nor U230 (N_230,In_765,In_200);
nor U231 (N_231,In_125,In_192);
nor U232 (N_232,In_298,In_915);
and U233 (N_233,In_92,In_499);
nand U234 (N_234,In_422,In_426);
nor U235 (N_235,In_465,In_53);
nand U236 (N_236,In_700,In_548);
and U237 (N_237,In_314,In_966);
nand U238 (N_238,In_289,In_165);
nor U239 (N_239,In_729,In_395);
nand U240 (N_240,In_489,In_676);
and U241 (N_241,In_776,In_163);
and U242 (N_242,In_509,In_878);
and U243 (N_243,In_343,In_662);
or U244 (N_244,In_32,In_625);
nor U245 (N_245,In_120,In_484);
nand U246 (N_246,In_828,In_507);
and U247 (N_247,In_572,In_135);
nor U248 (N_248,In_50,In_358);
or U249 (N_249,In_514,In_172);
or U250 (N_250,In_679,In_297);
or U251 (N_251,In_650,In_992);
and U252 (N_252,In_373,In_607);
nand U253 (N_253,In_603,In_96);
or U254 (N_254,In_857,In_860);
and U255 (N_255,In_715,In_430);
and U256 (N_256,In_906,In_741);
or U257 (N_257,In_6,In_978);
nand U258 (N_258,In_220,In_879);
nor U259 (N_259,In_0,In_337);
or U260 (N_260,In_840,In_118);
and U261 (N_261,In_346,In_814);
nor U262 (N_262,In_949,In_300);
or U263 (N_263,In_154,In_448);
and U264 (N_264,In_503,In_586);
or U265 (N_265,In_540,In_626);
nand U266 (N_266,In_721,In_208);
nor U267 (N_267,In_209,In_763);
nand U268 (N_268,In_847,In_408);
or U269 (N_269,In_330,In_945);
or U270 (N_270,In_936,In_802);
or U271 (N_271,In_336,In_595);
and U272 (N_272,In_940,In_553);
nor U273 (N_273,In_694,In_404);
nand U274 (N_274,In_495,In_686);
nor U275 (N_275,In_131,In_608);
nand U276 (N_276,In_796,In_25);
nor U277 (N_277,In_728,In_377);
or U278 (N_278,In_439,In_4);
or U279 (N_279,In_827,In_397);
nor U280 (N_280,In_191,In_866);
nand U281 (N_281,In_93,In_244);
nand U282 (N_282,In_253,In_126);
or U283 (N_283,In_826,In_344);
nor U284 (N_284,In_510,In_983);
nor U285 (N_285,In_146,In_411);
and U286 (N_286,In_291,In_753);
nand U287 (N_287,In_914,In_901);
or U288 (N_288,In_480,In_652);
and U289 (N_289,In_577,In_824);
nor U290 (N_290,In_486,In_869);
or U291 (N_291,In_263,In_21);
nand U292 (N_292,In_310,In_929);
nor U293 (N_293,In_994,In_752);
nand U294 (N_294,In_841,In_647);
nor U295 (N_295,In_113,In_17);
and U296 (N_296,In_655,In_243);
nor U297 (N_297,In_181,In_800);
and U298 (N_298,In_353,In_142);
or U299 (N_299,In_634,In_504);
nor U300 (N_300,In_720,In_443);
nor U301 (N_301,In_889,In_751);
and U302 (N_302,In_939,In_537);
or U303 (N_303,In_555,In_341);
nand U304 (N_304,In_452,In_845);
nand U305 (N_305,In_897,In_392);
nand U306 (N_306,In_696,In_680);
or U307 (N_307,In_205,In_733);
or U308 (N_308,In_766,In_653);
nand U309 (N_309,In_151,In_296);
nor U310 (N_310,In_219,In_78);
and U311 (N_311,In_39,In_442);
nor U312 (N_312,In_534,In_241);
nor U313 (N_313,In_184,In_61);
and U314 (N_314,In_767,In_178);
nand U315 (N_315,In_597,In_505);
and U316 (N_316,In_124,In_369);
or U317 (N_317,In_272,In_618);
nor U318 (N_318,In_593,In_258);
or U319 (N_319,In_703,In_806);
or U320 (N_320,In_454,In_171);
or U321 (N_321,In_850,In_152);
or U322 (N_322,In_308,In_882);
or U323 (N_323,In_584,In_832);
or U324 (N_324,In_829,In_740);
nor U325 (N_325,In_461,In_798);
nor U326 (N_326,In_276,In_903);
and U327 (N_327,In_492,In_627);
or U328 (N_328,In_682,In_57);
and U329 (N_329,In_842,In_213);
or U330 (N_330,In_403,In_224);
nand U331 (N_331,In_228,In_110);
or U332 (N_332,In_900,In_162);
and U333 (N_333,In_774,In_74);
nor U334 (N_334,In_921,In_927);
nor U335 (N_335,In_566,In_238);
or U336 (N_336,In_750,In_107);
nor U337 (N_337,In_969,In_863);
and U338 (N_338,In_815,In_1);
nor U339 (N_339,In_173,In_376);
nand U340 (N_340,In_67,In_784);
or U341 (N_341,In_665,In_813);
and U342 (N_342,In_981,In_138);
and U343 (N_343,In_885,In_60);
nor U344 (N_344,In_399,In_33);
nor U345 (N_345,In_166,In_51);
nor U346 (N_346,In_363,In_591);
nor U347 (N_347,In_554,In_38);
and U348 (N_348,In_48,In_902);
or U349 (N_349,In_598,In_925);
nor U350 (N_350,In_24,In_789);
and U351 (N_351,In_333,In_592);
nor U352 (N_352,In_194,In_547);
and U353 (N_353,In_580,In_242);
or U354 (N_354,In_635,In_386);
and U355 (N_355,In_133,In_420);
nor U356 (N_356,In_129,In_479);
nor U357 (N_357,In_926,In_161);
and U358 (N_358,In_501,In_382);
nand U359 (N_359,In_807,In_462);
nand U360 (N_360,In_735,In_630);
or U361 (N_361,In_657,In_561);
nand U362 (N_362,In_62,In_370);
and U363 (N_363,In_233,In_262);
or U364 (N_364,In_742,In_401);
or U365 (N_365,In_757,In_520);
nor U366 (N_366,In_85,In_283);
nand U367 (N_367,In_269,In_980);
nand U368 (N_368,In_15,In_838);
nand U369 (N_369,In_235,In_604);
nor U370 (N_370,In_664,In_282);
nor U371 (N_371,In_167,In_691);
nand U372 (N_372,In_810,In_378);
nor U373 (N_373,In_629,In_974);
and U374 (N_374,In_677,In_633);
or U375 (N_375,In_986,In_182);
or U376 (N_376,In_249,In_435);
and U377 (N_377,In_451,In_973);
nand U378 (N_378,In_372,In_689);
nor U379 (N_379,In_670,In_585);
or U380 (N_380,In_928,In_98);
nand U381 (N_381,In_596,In_438);
and U382 (N_382,In_892,In_621);
nand U383 (N_383,In_387,In_425);
and U384 (N_384,In_359,In_303);
nor U385 (N_385,In_327,In_948);
nand U386 (N_386,In_589,In_951);
nand U387 (N_387,In_972,In_854);
nand U388 (N_388,In_275,In_549);
and U389 (N_389,In_762,In_599);
nor U390 (N_390,In_745,In_232);
nand U391 (N_391,In_989,In_155);
and U392 (N_392,In_821,In_624);
or U393 (N_393,In_423,In_739);
or U394 (N_394,In_917,In_631);
or U395 (N_395,In_80,In_71);
and U396 (N_396,In_531,In_95);
or U397 (N_397,In_543,In_508);
or U398 (N_398,In_770,In_5);
nor U399 (N_399,In_523,In_45);
nor U400 (N_400,In_959,In_642);
or U401 (N_401,In_54,In_673);
nand U402 (N_402,In_661,In_40);
nor U403 (N_403,In_64,In_723);
or U404 (N_404,In_30,In_529);
xnor U405 (N_405,In_837,In_539);
nor U406 (N_406,In_295,In_270);
and U407 (N_407,In_407,In_416);
xnor U408 (N_408,In_429,In_476);
nand U409 (N_409,In_808,In_952);
or U410 (N_410,In_354,In_10);
or U411 (N_411,In_472,In_913);
nand U412 (N_412,In_481,In_871);
nor U413 (N_413,In_35,In_701);
or U414 (N_414,In_102,In_562);
nand U415 (N_415,In_695,In_811);
nor U416 (N_416,In_699,In_315);
nand U417 (N_417,In_101,In_347);
nand U418 (N_418,In_432,In_383);
or U419 (N_419,In_317,In_390);
or U420 (N_420,In_874,In_991);
or U421 (N_421,In_870,In_812);
nor U422 (N_422,In_176,In_222);
or U423 (N_423,In_309,In_381);
nor U424 (N_424,In_594,In_70);
nand U425 (N_425,In_13,In_563);
nor U426 (N_426,In_206,In_14);
nand U427 (N_427,In_791,In_541);
nand U428 (N_428,In_103,In_361);
nor U429 (N_429,In_990,In_170);
nand U430 (N_430,In_706,In_186);
and U431 (N_431,In_574,In_709);
nand U432 (N_432,In_417,In_147);
and U433 (N_433,In_250,In_214);
and U434 (N_434,In_868,In_588);
nor U435 (N_435,In_690,In_134);
nor U436 (N_436,In_685,In_475);
or U437 (N_437,In_546,In_835);
nor U438 (N_438,In_787,In_215);
xnor U439 (N_439,In_493,In_56);
or U440 (N_440,In_985,In_867);
nand U441 (N_441,In_931,In_335);
or U442 (N_442,In_23,In_179);
and U443 (N_443,In_614,In_525);
nand U444 (N_444,In_861,In_406);
and U445 (N_445,In_41,In_957);
or U446 (N_446,In_217,In_144);
or U447 (N_447,In_388,In_617);
or U448 (N_448,In_708,In_267);
and U449 (N_449,In_338,In_199);
nor U450 (N_450,In_612,In_148);
and U451 (N_451,In_651,In_894);
nor U452 (N_452,In_542,In_937);
nand U453 (N_453,In_73,In_942);
or U454 (N_454,In_281,In_968);
nand U455 (N_455,In_455,In_440);
nor U456 (N_456,In_755,In_234);
or U457 (N_457,In_247,In_412);
or U458 (N_458,In_469,In_368);
or U459 (N_459,In_877,In_292);
and U460 (N_460,In_544,In_616);
and U461 (N_461,In_478,In_833);
nor U462 (N_462,In_473,In_141);
nand U463 (N_463,In_760,In_619);
and U464 (N_464,In_993,In_898);
or U465 (N_465,In_265,In_477);
and U466 (N_466,In_684,In_935);
and U467 (N_467,In_246,In_487);
and U468 (N_468,In_55,In_831);
and U469 (N_469,In_150,In_768);
or U470 (N_470,In_318,In_286);
nand U471 (N_471,In_722,In_521);
and U472 (N_472,In_156,In_380);
or U473 (N_473,In_114,In_218);
nand U474 (N_474,In_799,In_786);
or U475 (N_475,In_140,In_111);
and U476 (N_476,In_321,In_557);
nand U477 (N_477,In_515,In_864);
or U478 (N_478,In_893,In_221);
and U479 (N_479,In_174,In_375);
and U480 (N_480,In_693,In_578);
and U481 (N_481,In_216,In_7);
nand U482 (N_482,In_659,In_223);
or U483 (N_483,In_601,In_671);
nand U484 (N_484,In_535,In_284);
nor U485 (N_485,In_820,In_910);
nor U486 (N_486,In_967,In_349);
nand U487 (N_487,In_187,In_988);
nand U488 (N_488,In_997,In_277);
nor U489 (N_489,In_168,In_538);
nor U490 (N_490,In_16,In_886);
or U491 (N_491,In_688,In_445);
or U492 (N_492,In_620,In_97);
nand U493 (N_493,In_818,In_202);
or U494 (N_494,In_136,In_710);
nand U495 (N_495,In_583,In_615);
xor U496 (N_496,In_348,In_668);
nand U497 (N_497,In_322,In_87);
nand U498 (N_498,In_305,In_909);
and U499 (N_499,In_323,In_374);
nor U500 (N_500,In_924,In_983);
and U501 (N_501,In_93,In_205);
and U502 (N_502,In_700,In_606);
nand U503 (N_503,In_90,In_746);
and U504 (N_504,In_929,In_926);
and U505 (N_505,In_351,In_558);
nand U506 (N_506,In_434,In_786);
or U507 (N_507,In_294,In_170);
or U508 (N_508,In_124,In_122);
or U509 (N_509,In_167,In_519);
nor U510 (N_510,In_898,In_960);
nor U511 (N_511,In_771,In_818);
nor U512 (N_512,In_494,In_377);
or U513 (N_513,In_764,In_368);
nand U514 (N_514,In_320,In_194);
nor U515 (N_515,In_770,In_243);
nor U516 (N_516,In_691,In_125);
and U517 (N_517,In_655,In_254);
or U518 (N_518,In_390,In_671);
nor U519 (N_519,In_307,In_425);
and U520 (N_520,In_463,In_117);
nand U521 (N_521,In_827,In_31);
nand U522 (N_522,In_813,In_699);
nor U523 (N_523,In_463,In_177);
nor U524 (N_524,In_641,In_677);
nor U525 (N_525,In_141,In_667);
or U526 (N_526,In_330,In_141);
and U527 (N_527,In_166,In_312);
and U528 (N_528,In_44,In_53);
nor U529 (N_529,In_52,In_64);
and U530 (N_530,In_361,In_172);
and U531 (N_531,In_406,In_171);
or U532 (N_532,In_852,In_829);
and U533 (N_533,In_379,In_655);
or U534 (N_534,In_808,In_146);
nor U535 (N_535,In_264,In_600);
nor U536 (N_536,In_451,In_699);
and U537 (N_537,In_756,In_731);
nor U538 (N_538,In_452,In_843);
or U539 (N_539,In_37,In_842);
nand U540 (N_540,In_791,In_957);
or U541 (N_541,In_661,In_515);
and U542 (N_542,In_419,In_719);
nand U543 (N_543,In_635,In_6);
nor U544 (N_544,In_917,In_34);
or U545 (N_545,In_517,In_494);
nand U546 (N_546,In_184,In_738);
nand U547 (N_547,In_90,In_639);
nor U548 (N_548,In_803,In_271);
and U549 (N_549,In_185,In_871);
and U550 (N_550,In_535,In_381);
or U551 (N_551,In_269,In_408);
and U552 (N_552,In_796,In_783);
and U553 (N_553,In_144,In_580);
nand U554 (N_554,In_708,In_740);
nor U555 (N_555,In_113,In_626);
nor U556 (N_556,In_675,In_181);
and U557 (N_557,In_752,In_750);
nand U558 (N_558,In_632,In_748);
and U559 (N_559,In_378,In_444);
nand U560 (N_560,In_240,In_104);
and U561 (N_561,In_282,In_829);
and U562 (N_562,In_936,In_577);
or U563 (N_563,In_130,In_451);
nor U564 (N_564,In_934,In_594);
nand U565 (N_565,In_546,In_872);
and U566 (N_566,In_895,In_808);
and U567 (N_567,In_530,In_731);
nor U568 (N_568,In_711,In_361);
nor U569 (N_569,In_312,In_476);
and U570 (N_570,In_5,In_61);
nand U571 (N_571,In_884,In_346);
or U572 (N_572,In_309,In_22);
and U573 (N_573,In_521,In_875);
nand U574 (N_574,In_113,In_2);
nand U575 (N_575,In_450,In_740);
and U576 (N_576,In_102,In_467);
and U577 (N_577,In_705,In_816);
nand U578 (N_578,In_261,In_9);
nand U579 (N_579,In_11,In_60);
nand U580 (N_580,In_691,In_321);
or U581 (N_581,In_136,In_572);
or U582 (N_582,In_752,In_797);
and U583 (N_583,In_859,In_551);
or U584 (N_584,In_432,In_563);
and U585 (N_585,In_547,In_76);
nor U586 (N_586,In_765,In_673);
or U587 (N_587,In_211,In_968);
nor U588 (N_588,In_0,In_426);
or U589 (N_589,In_269,In_187);
nand U590 (N_590,In_46,In_511);
nand U591 (N_591,In_653,In_812);
and U592 (N_592,In_134,In_294);
and U593 (N_593,In_617,In_181);
nand U594 (N_594,In_787,In_941);
and U595 (N_595,In_186,In_845);
nor U596 (N_596,In_895,In_839);
or U597 (N_597,In_34,In_509);
nand U598 (N_598,In_613,In_74);
nor U599 (N_599,In_65,In_777);
nand U600 (N_600,In_248,In_283);
and U601 (N_601,In_549,In_361);
nand U602 (N_602,In_118,In_725);
and U603 (N_603,In_377,In_221);
nand U604 (N_604,In_880,In_181);
nand U605 (N_605,In_530,In_94);
nor U606 (N_606,In_853,In_278);
nor U607 (N_607,In_58,In_490);
nand U608 (N_608,In_842,In_389);
nor U609 (N_609,In_475,In_919);
nor U610 (N_610,In_639,In_322);
and U611 (N_611,In_64,In_240);
nor U612 (N_612,In_852,In_88);
or U613 (N_613,In_732,In_141);
nor U614 (N_614,In_648,In_292);
nand U615 (N_615,In_947,In_268);
nor U616 (N_616,In_772,In_717);
or U617 (N_617,In_518,In_242);
nor U618 (N_618,In_105,In_597);
and U619 (N_619,In_269,In_492);
and U620 (N_620,In_192,In_935);
and U621 (N_621,In_748,In_23);
nand U622 (N_622,In_143,In_938);
and U623 (N_623,In_26,In_268);
nor U624 (N_624,In_593,In_992);
and U625 (N_625,In_518,In_659);
nand U626 (N_626,In_832,In_137);
and U627 (N_627,In_936,In_476);
or U628 (N_628,In_158,In_440);
nand U629 (N_629,In_95,In_309);
and U630 (N_630,In_515,In_564);
and U631 (N_631,In_598,In_308);
nor U632 (N_632,In_895,In_615);
and U633 (N_633,In_258,In_915);
and U634 (N_634,In_728,In_269);
or U635 (N_635,In_141,In_829);
or U636 (N_636,In_758,In_264);
nor U637 (N_637,In_209,In_505);
nor U638 (N_638,In_73,In_400);
and U639 (N_639,In_544,In_38);
nor U640 (N_640,In_785,In_568);
nor U641 (N_641,In_498,In_244);
and U642 (N_642,In_88,In_624);
or U643 (N_643,In_940,In_433);
and U644 (N_644,In_188,In_656);
and U645 (N_645,In_748,In_925);
nor U646 (N_646,In_430,In_811);
nand U647 (N_647,In_798,In_66);
and U648 (N_648,In_60,In_680);
xnor U649 (N_649,In_584,In_821);
nand U650 (N_650,In_767,In_588);
nand U651 (N_651,In_168,In_703);
nand U652 (N_652,In_570,In_195);
or U653 (N_653,In_516,In_89);
or U654 (N_654,In_535,In_865);
nand U655 (N_655,In_56,In_435);
and U656 (N_656,In_882,In_160);
xnor U657 (N_657,In_151,In_222);
and U658 (N_658,In_335,In_247);
nor U659 (N_659,In_638,In_880);
and U660 (N_660,In_302,In_408);
and U661 (N_661,In_460,In_617);
or U662 (N_662,In_523,In_338);
nor U663 (N_663,In_682,In_527);
nand U664 (N_664,In_7,In_860);
or U665 (N_665,In_637,In_21);
nor U666 (N_666,In_799,In_912);
or U667 (N_667,In_654,In_557);
nor U668 (N_668,In_282,In_113);
or U669 (N_669,In_393,In_637);
and U670 (N_670,In_46,In_392);
or U671 (N_671,In_215,In_568);
and U672 (N_672,In_938,In_455);
nand U673 (N_673,In_701,In_917);
nor U674 (N_674,In_284,In_863);
nand U675 (N_675,In_926,In_799);
or U676 (N_676,In_842,In_768);
nand U677 (N_677,In_720,In_414);
nor U678 (N_678,In_205,In_731);
or U679 (N_679,In_685,In_370);
or U680 (N_680,In_155,In_824);
and U681 (N_681,In_619,In_735);
and U682 (N_682,In_980,In_343);
and U683 (N_683,In_21,In_989);
nor U684 (N_684,In_362,In_252);
nand U685 (N_685,In_855,In_808);
nand U686 (N_686,In_566,In_272);
or U687 (N_687,In_14,In_87);
nor U688 (N_688,In_447,In_883);
and U689 (N_689,In_315,In_677);
and U690 (N_690,In_766,In_893);
or U691 (N_691,In_241,In_367);
xor U692 (N_692,In_764,In_852);
nor U693 (N_693,In_163,In_281);
or U694 (N_694,In_687,In_456);
or U695 (N_695,In_700,In_15);
or U696 (N_696,In_821,In_778);
and U697 (N_697,In_165,In_380);
nor U698 (N_698,In_7,In_944);
nand U699 (N_699,In_800,In_804);
and U700 (N_700,In_792,In_956);
xor U701 (N_701,In_750,In_901);
or U702 (N_702,In_252,In_436);
and U703 (N_703,In_531,In_90);
nor U704 (N_704,In_223,In_423);
and U705 (N_705,In_331,In_629);
nand U706 (N_706,In_456,In_560);
nor U707 (N_707,In_873,In_915);
nor U708 (N_708,In_950,In_982);
or U709 (N_709,In_378,In_792);
and U710 (N_710,In_767,In_985);
nor U711 (N_711,In_850,In_725);
or U712 (N_712,In_35,In_198);
or U713 (N_713,In_488,In_452);
or U714 (N_714,In_843,In_522);
and U715 (N_715,In_441,In_741);
and U716 (N_716,In_732,In_330);
or U717 (N_717,In_417,In_802);
nor U718 (N_718,In_503,In_958);
nor U719 (N_719,In_543,In_61);
nand U720 (N_720,In_762,In_257);
and U721 (N_721,In_768,In_962);
nand U722 (N_722,In_383,In_309);
nand U723 (N_723,In_303,In_576);
nor U724 (N_724,In_936,In_42);
and U725 (N_725,In_940,In_185);
or U726 (N_726,In_271,In_480);
nand U727 (N_727,In_657,In_599);
nor U728 (N_728,In_782,In_226);
or U729 (N_729,In_186,In_227);
nand U730 (N_730,In_354,In_969);
nor U731 (N_731,In_969,In_534);
and U732 (N_732,In_995,In_594);
nor U733 (N_733,In_365,In_911);
nand U734 (N_734,In_902,In_13);
nand U735 (N_735,In_397,In_949);
nand U736 (N_736,In_714,In_75);
or U737 (N_737,In_628,In_909);
or U738 (N_738,In_382,In_755);
nand U739 (N_739,In_373,In_378);
nor U740 (N_740,In_49,In_96);
and U741 (N_741,In_516,In_804);
nor U742 (N_742,In_747,In_359);
and U743 (N_743,In_87,In_844);
nor U744 (N_744,In_899,In_737);
nor U745 (N_745,In_851,In_911);
and U746 (N_746,In_644,In_807);
nand U747 (N_747,In_30,In_378);
nor U748 (N_748,In_299,In_518);
nor U749 (N_749,In_209,In_868);
or U750 (N_750,In_745,In_918);
and U751 (N_751,In_975,In_886);
nor U752 (N_752,In_158,In_136);
nand U753 (N_753,In_81,In_427);
or U754 (N_754,In_871,In_83);
nand U755 (N_755,In_879,In_381);
nor U756 (N_756,In_331,In_287);
nand U757 (N_757,In_786,In_1);
nand U758 (N_758,In_727,In_905);
and U759 (N_759,In_985,In_390);
nand U760 (N_760,In_159,In_166);
nor U761 (N_761,In_42,In_84);
and U762 (N_762,In_882,In_752);
nor U763 (N_763,In_143,In_334);
and U764 (N_764,In_749,In_637);
nand U765 (N_765,In_238,In_159);
or U766 (N_766,In_121,In_610);
or U767 (N_767,In_829,In_763);
or U768 (N_768,In_547,In_966);
and U769 (N_769,In_960,In_148);
or U770 (N_770,In_887,In_55);
or U771 (N_771,In_980,In_986);
or U772 (N_772,In_920,In_757);
or U773 (N_773,In_902,In_496);
nand U774 (N_774,In_903,In_109);
or U775 (N_775,In_184,In_610);
or U776 (N_776,In_544,In_845);
and U777 (N_777,In_708,In_698);
nor U778 (N_778,In_547,In_39);
nor U779 (N_779,In_628,In_643);
nor U780 (N_780,In_920,In_198);
nand U781 (N_781,In_445,In_237);
and U782 (N_782,In_735,In_315);
nor U783 (N_783,In_673,In_527);
and U784 (N_784,In_245,In_331);
or U785 (N_785,In_873,In_848);
and U786 (N_786,In_206,In_488);
nand U787 (N_787,In_13,In_745);
nand U788 (N_788,In_60,In_366);
nand U789 (N_789,In_634,In_808);
nor U790 (N_790,In_114,In_804);
nand U791 (N_791,In_429,In_519);
nor U792 (N_792,In_96,In_255);
nand U793 (N_793,In_949,In_282);
nand U794 (N_794,In_161,In_793);
and U795 (N_795,In_376,In_595);
nand U796 (N_796,In_138,In_680);
and U797 (N_797,In_741,In_95);
nand U798 (N_798,In_612,In_373);
nor U799 (N_799,In_740,In_738);
and U800 (N_800,In_267,In_280);
and U801 (N_801,In_102,In_758);
nor U802 (N_802,In_41,In_475);
nand U803 (N_803,In_61,In_782);
nand U804 (N_804,In_365,In_962);
nand U805 (N_805,In_21,In_163);
nor U806 (N_806,In_670,In_711);
nor U807 (N_807,In_734,In_663);
and U808 (N_808,In_827,In_977);
nor U809 (N_809,In_918,In_659);
nand U810 (N_810,In_32,In_900);
or U811 (N_811,In_61,In_724);
nor U812 (N_812,In_422,In_882);
nor U813 (N_813,In_347,In_578);
nand U814 (N_814,In_771,In_22);
or U815 (N_815,In_605,In_244);
nand U816 (N_816,In_916,In_497);
or U817 (N_817,In_193,In_257);
and U818 (N_818,In_609,In_683);
nor U819 (N_819,In_29,In_655);
and U820 (N_820,In_899,In_215);
nor U821 (N_821,In_48,In_580);
xnor U822 (N_822,In_602,In_457);
or U823 (N_823,In_2,In_449);
or U824 (N_824,In_577,In_202);
nor U825 (N_825,In_339,In_865);
nand U826 (N_826,In_112,In_225);
or U827 (N_827,In_876,In_163);
or U828 (N_828,In_702,In_126);
and U829 (N_829,In_918,In_594);
and U830 (N_830,In_533,In_975);
nand U831 (N_831,In_985,In_807);
and U832 (N_832,In_292,In_209);
nand U833 (N_833,In_447,In_168);
nor U834 (N_834,In_522,In_756);
nor U835 (N_835,In_228,In_713);
or U836 (N_836,In_144,In_817);
and U837 (N_837,In_621,In_416);
nor U838 (N_838,In_13,In_502);
nor U839 (N_839,In_593,In_18);
or U840 (N_840,In_683,In_309);
or U841 (N_841,In_742,In_993);
and U842 (N_842,In_358,In_999);
xor U843 (N_843,In_323,In_787);
or U844 (N_844,In_485,In_938);
nor U845 (N_845,In_410,In_685);
nor U846 (N_846,In_58,In_718);
and U847 (N_847,In_582,In_549);
nand U848 (N_848,In_948,In_95);
nor U849 (N_849,In_419,In_701);
and U850 (N_850,In_708,In_117);
xor U851 (N_851,In_552,In_308);
or U852 (N_852,In_537,In_365);
or U853 (N_853,In_633,In_509);
nand U854 (N_854,In_233,In_443);
nand U855 (N_855,In_281,In_354);
and U856 (N_856,In_538,In_275);
and U857 (N_857,In_132,In_590);
nor U858 (N_858,In_695,In_817);
nand U859 (N_859,In_930,In_620);
nand U860 (N_860,In_701,In_607);
and U861 (N_861,In_132,In_680);
or U862 (N_862,In_374,In_293);
nand U863 (N_863,In_674,In_779);
and U864 (N_864,In_864,In_891);
nand U865 (N_865,In_605,In_750);
or U866 (N_866,In_931,In_89);
nor U867 (N_867,In_735,In_938);
or U868 (N_868,In_914,In_484);
nor U869 (N_869,In_517,In_793);
nor U870 (N_870,In_200,In_445);
nor U871 (N_871,In_892,In_706);
or U872 (N_872,In_995,In_360);
nand U873 (N_873,In_37,In_149);
or U874 (N_874,In_809,In_454);
or U875 (N_875,In_612,In_92);
nor U876 (N_876,In_845,In_982);
nor U877 (N_877,In_3,In_826);
or U878 (N_878,In_92,In_816);
and U879 (N_879,In_995,In_184);
nor U880 (N_880,In_975,In_98);
and U881 (N_881,In_527,In_983);
nor U882 (N_882,In_156,In_574);
or U883 (N_883,In_873,In_196);
nand U884 (N_884,In_455,In_597);
nand U885 (N_885,In_359,In_114);
and U886 (N_886,In_169,In_260);
nor U887 (N_887,In_995,In_495);
nor U888 (N_888,In_124,In_384);
nand U889 (N_889,In_531,In_427);
nor U890 (N_890,In_907,In_19);
and U891 (N_891,In_925,In_696);
nand U892 (N_892,In_914,In_165);
and U893 (N_893,In_852,In_715);
nor U894 (N_894,In_240,In_437);
nand U895 (N_895,In_632,In_505);
nand U896 (N_896,In_549,In_79);
or U897 (N_897,In_393,In_982);
or U898 (N_898,In_181,In_190);
or U899 (N_899,In_321,In_739);
nor U900 (N_900,In_700,In_533);
or U901 (N_901,In_534,In_551);
nor U902 (N_902,In_18,In_366);
and U903 (N_903,In_147,In_614);
or U904 (N_904,In_844,In_785);
or U905 (N_905,In_580,In_642);
nand U906 (N_906,In_877,In_902);
or U907 (N_907,In_175,In_322);
or U908 (N_908,In_667,In_577);
nor U909 (N_909,In_484,In_234);
nor U910 (N_910,In_710,In_365);
or U911 (N_911,In_433,In_765);
or U912 (N_912,In_275,In_160);
nand U913 (N_913,In_4,In_155);
xor U914 (N_914,In_837,In_504);
and U915 (N_915,In_54,In_907);
nor U916 (N_916,In_772,In_50);
or U917 (N_917,In_298,In_79);
or U918 (N_918,In_621,In_76);
and U919 (N_919,In_600,In_683);
nor U920 (N_920,In_313,In_759);
nor U921 (N_921,In_743,In_702);
and U922 (N_922,In_621,In_760);
nand U923 (N_923,In_410,In_686);
or U924 (N_924,In_281,In_815);
nor U925 (N_925,In_554,In_209);
and U926 (N_926,In_555,In_306);
nand U927 (N_927,In_56,In_755);
or U928 (N_928,In_128,In_109);
and U929 (N_929,In_234,In_337);
or U930 (N_930,In_527,In_537);
nand U931 (N_931,In_513,In_265);
nand U932 (N_932,In_277,In_977);
nor U933 (N_933,In_149,In_160);
or U934 (N_934,In_952,In_827);
xnor U935 (N_935,In_506,In_822);
and U936 (N_936,In_750,In_124);
or U937 (N_937,In_245,In_598);
or U938 (N_938,In_477,In_963);
or U939 (N_939,In_934,In_222);
or U940 (N_940,In_642,In_101);
and U941 (N_941,In_826,In_192);
and U942 (N_942,In_68,In_315);
or U943 (N_943,In_161,In_798);
and U944 (N_944,In_648,In_487);
or U945 (N_945,In_784,In_210);
nor U946 (N_946,In_677,In_837);
nand U947 (N_947,In_45,In_105);
nand U948 (N_948,In_515,In_892);
nor U949 (N_949,In_718,In_601);
nand U950 (N_950,In_120,In_789);
and U951 (N_951,In_474,In_656);
nand U952 (N_952,In_262,In_224);
nor U953 (N_953,In_325,In_898);
nand U954 (N_954,In_559,In_668);
or U955 (N_955,In_837,In_486);
or U956 (N_956,In_351,In_174);
or U957 (N_957,In_775,In_474);
nor U958 (N_958,In_638,In_706);
nor U959 (N_959,In_299,In_278);
or U960 (N_960,In_848,In_172);
nand U961 (N_961,In_437,In_992);
nand U962 (N_962,In_928,In_139);
nand U963 (N_963,In_503,In_141);
or U964 (N_964,In_610,In_648);
and U965 (N_965,In_917,In_188);
or U966 (N_966,In_667,In_127);
nand U967 (N_967,In_494,In_972);
nor U968 (N_968,In_527,In_439);
or U969 (N_969,In_968,In_196);
and U970 (N_970,In_578,In_50);
nor U971 (N_971,In_592,In_915);
or U972 (N_972,In_289,In_221);
or U973 (N_973,In_3,In_851);
nand U974 (N_974,In_174,In_521);
or U975 (N_975,In_823,In_158);
nand U976 (N_976,In_404,In_868);
nor U977 (N_977,In_64,In_927);
nor U978 (N_978,In_329,In_891);
and U979 (N_979,In_424,In_362);
and U980 (N_980,In_68,In_422);
nor U981 (N_981,In_411,In_306);
nor U982 (N_982,In_866,In_83);
nand U983 (N_983,In_832,In_292);
nand U984 (N_984,In_317,In_269);
and U985 (N_985,In_549,In_364);
and U986 (N_986,In_636,In_322);
nor U987 (N_987,In_226,In_596);
nand U988 (N_988,In_356,In_4);
and U989 (N_989,In_997,In_275);
or U990 (N_990,In_97,In_700);
or U991 (N_991,In_11,In_95);
nor U992 (N_992,In_718,In_726);
and U993 (N_993,In_481,In_674);
nand U994 (N_994,In_224,In_755);
nand U995 (N_995,In_517,In_285);
nand U996 (N_996,In_742,In_453);
or U997 (N_997,In_516,In_587);
nor U998 (N_998,In_208,In_288);
nor U999 (N_999,In_474,In_626);
and U1000 (N_1000,In_451,In_995);
or U1001 (N_1001,In_668,In_151);
or U1002 (N_1002,In_984,In_985);
nand U1003 (N_1003,In_126,In_927);
and U1004 (N_1004,In_172,In_338);
nand U1005 (N_1005,In_685,In_798);
or U1006 (N_1006,In_600,In_664);
nand U1007 (N_1007,In_133,In_841);
and U1008 (N_1008,In_114,In_349);
nand U1009 (N_1009,In_507,In_147);
or U1010 (N_1010,In_73,In_527);
nand U1011 (N_1011,In_54,In_28);
nand U1012 (N_1012,In_333,In_843);
nor U1013 (N_1013,In_992,In_655);
and U1014 (N_1014,In_609,In_403);
nand U1015 (N_1015,In_774,In_71);
or U1016 (N_1016,In_770,In_369);
nand U1017 (N_1017,In_697,In_199);
nor U1018 (N_1018,In_352,In_956);
nand U1019 (N_1019,In_540,In_547);
or U1020 (N_1020,In_589,In_222);
nor U1021 (N_1021,In_47,In_111);
or U1022 (N_1022,In_615,In_290);
nand U1023 (N_1023,In_663,In_5);
and U1024 (N_1024,In_35,In_267);
or U1025 (N_1025,In_638,In_432);
nor U1026 (N_1026,In_877,In_913);
nor U1027 (N_1027,In_761,In_236);
nand U1028 (N_1028,In_358,In_730);
or U1029 (N_1029,In_81,In_169);
nand U1030 (N_1030,In_444,In_144);
and U1031 (N_1031,In_420,In_515);
or U1032 (N_1032,In_400,In_231);
nor U1033 (N_1033,In_845,In_981);
xor U1034 (N_1034,In_203,In_382);
nand U1035 (N_1035,In_557,In_747);
and U1036 (N_1036,In_43,In_135);
and U1037 (N_1037,In_968,In_964);
nand U1038 (N_1038,In_276,In_70);
nor U1039 (N_1039,In_761,In_713);
and U1040 (N_1040,In_700,In_601);
and U1041 (N_1041,In_68,In_88);
and U1042 (N_1042,In_814,In_491);
and U1043 (N_1043,In_886,In_393);
and U1044 (N_1044,In_452,In_522);
nand U1045 (N_1045,In_390,In_890);
and U1046 (N_1046,In_688,In_715);
or U1047 (N_1047,In_867,In_438);
and U1048 (N_1048,In_526,In_880);
or U1049 (N_1049,In_528,In_971);
nor U1050 (N_1050,In_512,In_872);
nand U1051 (N_1051,In_483,In_644);
nand U1052 (N_1052,In_663,In_916);
or U1053 (N_1053,In_406,In_619);
nand U1054 (N_1054,In_650,In_199);
and U1055 (N_1055,In_642,In_3);
nor U1056 (N_1056,In_164,In_136);
and U1057 (N_1057,In_203,In_60);
nor U1058 (N_1058,In_859,In_361);
or U1059 (N_1059,In_915,In_382);
and U1060 (N_1060,In_302,In_734);
or U1061 (N_1061,In_80,In_789);
and U1062 (N_1062,In_743,In_396);
nor U1063 (N_1063,In_775,In_645);
nor U1064 (N_1064,In_416,In_365);
and U1065 (N_1065,In_635,In_263);
and U1066 (N_1066,In_550,In_763);
xor U1067 (N_1067,In_307,In_951);
nor U1068 (N_1068,In_239,In_51);
or U1069 (N_1069,In_153,In_131);
nor U1070 (N_1070,In_872,In_342);
nor U1071 (N_1071,In_710,In_653);
or U1072 (N_1072,In_962,In_5);
nand U1073 (N_1073,In_727,In_607);
nor U1074 (N_1074,In_122,In_354);
nor U1075 (N_1075,In_736,In_794);
and U1076 (N_1076,In_325,In_698);
or U1077 (N_1077,In_723,In_762);
nor U1078 (N_1078,In_70,In_896);
and U1079 (N_1079,In_830,In_788);
and U1080 (N_1080,In_798,In_492);
or U1081 (N_1081,In_390,In_769);
nor U1082 (N_1082,In_13,In_525);
nand U1083 (N_1083,In_694,In_873);
and U1084 (N_1084,In_712,In_329);
nor U1085 (N_1085,In_590,In_462);
nand U1086 (N_1086,In_462,In_137);
and U1087 (N_1087,In_715,In_729);
nor U1088 (N_1088,In_848,In_967);
nand U1089 (N_1089,In_506,In_308);
nand U1090 (N_1090,In_640,In_826);
nand U1091 (N_1091,In_568,In_577);
nor U1092 (N_1092,In_880,In_153);
nor U1093 (N_1093,In_796,In_672);
nor U1094 (N_1094,In_675,In_929);
or U1095 (N_1095,In_551,In_274);
nand U1096 (N_1096,In_508,In_339);
nand U1097 (N_1097,In_803,In_757);
or U1098 (N_1098,In_3,In_159);
and U1099 (N_1099,In_498,In_402);
and U1100 (N_1100,In_263,In_880);
or U1101 (N_1101,In_482,In_803);
nand U1102 (N_1102,In_573,In_738);
nand U1103 (N_1103,In_418,In_665);
nand U1104 (N_1104,In_213,In_39);
nand U1105 (N_1105,In_978,In_463);
or U1106 (N_1106,In_724,In_941);
nor U1107 (N_1107,In_903,In_625);
and U1108 (N_1108,In_476,In_864);
nor U1109 (N_1109,In_505,In_803);
or U1110 (N_1110,In_7,In_898);
nor U1111 (N_1111,In_444,In_190);
and U1112 (N_1112,In_206,In_195);
nand U1113 (N_1113,In_51,In_141);
or U1114 (N_1114,In_439,In_799);
or U1115 (N_1115,In_142,In_329);
nand U1116 (N_1116,In_561,In_598);
nor U1117 (N_1117,In_789,In_279);
nor U1118 (N_1118,In_93,In_196);
and U1119 (N_1119,In_685,In_299);
nand U1120 (N_1120,In_119,In_523);
nor U1121 (N_1121,In_692,In_752);
nor U1122 (N_1122,In_269,In_93);
nand U1123 (N_1123,In_146,In_818);
or U1124 (N_1124,In_495,In_540);
and U1125 (N_1125,In_54,In_221);
and U1126 (N_1126,In_237,In_677);
nor U1127 (N_1127,In_1,In_388);
nand U1128 (N_1128,In_890,In_920);
nand U1129 (N_1129,In_983,In_273);
nor U1130 (N_1130,In_142,In_344);
nand U1131 (N_1131,In_596,In_359);
or U1132 (N_1132,In_709,In_861);
nand U1133 (N_1133,In_122,In_127);
nand U1134 (N_1134,In_680,In_869);
nor U1135 (N_1135,In_815,In_394);
and U1136 (N_1136,In_233,In_197);
nor U1137 (N_1137,In_899,In_618);
xor U1138 (N_1138,In_821,In_264);
nor U1139 (N_1139,In_885,In_584);
or U1140 (N_1140,In_346,In_845);
nand U1141 (N_1141,In_24,In_703);
or U1142 (N_1142,In_317,In_177);
and U1143 (N_1143,In_455,In_761);
and U1144 (N_1144,In_327,In_783);
nand U1145 (N_1145,In_446,In_193);
nand U1146 (N_1146,In_418,In_9);
nand U1147 (N_1147,In_511,In_722);
or U1148 (N_1148,In_129,In_469);
or U1149 (N_1149,In_900,In_257);
nand U1150 (N_1150,In_412,In_576);
nand U1151 (N_1151,In_8,In_822);
or U1152 (N_1152,In_626,In_42);
nor U1153 (N_1153,In_262,In_495);
or U1154 (N_1154,In_901,In_853);
nor U1155 (N_1155,In_107,In_422);
nor U1156 (N_1156,In_15,In_2);
and U1157 (N_1157,In_38,In_766);
or U1158 (N_1158,In_970,In_972);
or U1159 (N_1159,In_524,In_612);
nor U1160 (N_1160,In_412,In_306);
or U1161 (N_1161,In_238,In_72);
and U1162 (N_1162,In_418,In_298);
nand U1163 (N_1163,In_622,In_51);
or U1164 (N_1164,In_273,In_973);
nor U1165 (N_1165,In_910,In_575);
nor U1166 (N_1166,In_489,In_979);
or U1167 (N_1167,In_583,In_535);
and U1168 (N_1168,In_674,In_478);
xnor U1169 (N_1169,In_885,In_792);
nor U1170 (N_1170,In_116,In_762);
nor U1171 (N_1171,In_421,In_925);
and U1172 (N_1172,In_523,In_114);
or U1173 (N_1173,In_919,In_729);
nand U1174 (N_1174,In_501,In_80);
nand U1175 (N_1175,In_692,In_481);
nor U1176 (N_1176,In_388,In_921);
nor U1177 (N_1177,In_39,In_572);
or U1178 (N_1178,In_837,In_500);
nand U1179 (N_1179,In_766,In_31);
nand U1180 (N_1180,In_844,In_664);
or U1181 (N_1181,In_304,In_774);
nand U1182 (N_1182,In_205,In_209);
nand U1183 (N_1183,In_312,In_690);
or U1184 (N_1184,In_463,In_504);
nand U1185 (N_1185,In_101,In_994);
nand U1186 (N_1186,In_622,In_193);
or U1187 (N_1187,In_606,In_939);
or U1188 (N_1188,In_9,In_878);
and U1189 (N_1189,In_31,In_721);
and U1190 (N_1190,In_284,In_352);
nor U1191 (N_1191,In_784,In_229);
nand U1192 (N_1192,In_452,In_906);
or U1193 (N_1193,In_40,In_421);
or U1194 (N_1194,In_642,In_183);
and U1195 (N_1195,In_793,In_361);
and U1196 (N_1196,In_268,In_766);
and U1197 (N_1197,In_3,In_719);
or U1198 (N_1198,In_603,In_161);
and U1199 (N_1199,In_31,In_471);
or U1200 (N_1200,In_965,In_162);
or U1201 (N_1201,In_643,In_123);
or U1202 (N_1202,In_591,In_295);
nand U1203 (N_1203,In_718,In_30);
or U1204 (N_1204,In_689,In_283);
nor U1205 (N_1205,In_26,In_50);
nor U1206 (N_1206,In_149,In_967);
and U1207 (N_1207,In_227,In_673);
and U1208 (N_1208,In_280,In_308);
or U1209 (N_1209,In_742,In_830);
nand U1210 (N_1210,In_150,In_29);
or U1211 (N_1211,In_637,In_927);
and U1212 (N_1212,In_781,In_364);
nor U1213 (N_1213,In_799,In_483);
and U1214 (N_1214,In_58,In_689);
and U1215 (N_1215,In_268,In_781);
nand U1216 (N_1216,In_563,In_960);
and U1217 (N_1217,In_295,In_840);
nor U1218 (N_1218,In_917,In_354);
or U1219 (N_1219,In_77,In_993);
and U1220 (N_1220,In_665,In_211);
or U1221 (N_1221,In_580,In_710);
nand U1222 (N_1222,In_701,In_505);
nand U1223 (N_1223,In_522,In_70);
and U1224 (N_1224,In_210,In_863);
or U1225 (N_1225,In_915,In_455);
nand U1226 (N_1226,In_426,In_537);
nor U1227 (N_1227,In_587,In_896);
nand U1228 (N_1228,In_321,In_10);
and U1229 (N_1229,In_934,In_935);
and U1230 (N_1230,In_534,In_312);
nor U1231 (N_1231,In_966,In_942);
nor U1232 (N_1232,In_561,In_775);
nand U1233 (N_1233,In_448,In_107);
nor U1234 (N_1234,In_490,In_314);
nor U1235 (N_1235,In_333,In_834);
nand U1236 (N_1236,In_784,In_8);
nor U1237 (N_1237,In_819,In_926);
xor U1238 (N_1238,In_285,In_844);
or U1239 (N_1239,In_4,In_259);
or U1240 (N_1240,In_133,In_450);
or U1241 (N_1241,In_494,In_705);
nor U1242 (N_1242,In_655,In_864);
nor U1243 (N_1243,In_790,In_73);
and U1244 (N_1244,In_433,In_964);
and U1245 (N_1245,In_88,In_709);
nand U1246 (N_1246,In_528,In_147);
nor U1247 (N_1247,In_400,In_692);
nor U1248 (N_1248,In_978,In_27);
nor U1249 (N_1249,In_874,In_638);
nand U1250 (N_1250,In_283,In_915);
nand U1251 (N_1251,In_676,In_113);
and U1252 (N_1252,In_827,In_162);
nor U1253 (N_1253,In_496,In_6);
nand U1254 (N_1254,In_721,In_796);
nand U1255 (N_1255,In_567,In_303);
nand U1256 (N_1256,In_173,In_311);
and U1257 (N_1257,In_675,In_452);
nor U1258 (N_1258,In_155,In_418);
nor U1259 (N_1259,In_927,In_493);
nand U1260 (N_1260,In_879,In_439);
and U1261 (N_1261,In_830,In_622);
nor U1262 (N_1262,In_470,In_126);
nand U1263 (N_1263,In_679,In_645);
and U1264 (N_1264,In_897,In_548);
nand U1265 (N_1265,In_308,In_282);
nand U1266 (N_1266,In_711,In_608);
nand U1267 (N_1267,In_474,In_5);
nand U1268 (N_1268,In_350,In_98);
nor U1269 (N_1269,In_110,In_206);
nand U1270 (N_1270,In_204,In_419);
nor U1271 (N_1271,In_754,In_156);
and U1272 (N_1272,In_101,In_987);
nor U1273 (N_1273,In_803,In_945);
nor U1274 (N_1274,In_510,In_772);
nand U1275 (N_1275,In_325,In_466);
nor U1276 (N_1276,In_784,In_858);
nand U1277 (N_1277,In_468,In_899);
nand U1278 (N_1278,In_350,In_227);
nor U1279 (N_1279,In_219,In_541);
nand U1280 (N_1280,In_70,In_11);
and U1281 (N_1281,In_910,In_286);
nand U1282 (N_1282,In_483,In_380);
and U1283 (N_1283,In_94,In_616);
or U1284 (N_1284,In_676,In_639);
and U1285 (N_1285,In_665,In_2);
xnor U1286 (N_1286,In_391,In_560);
and U1287 (N_1287,In_39,In_824);
and U1288 (N_1288,In_947,In_181);
or U1289 (N_1289,In_608,In_205);
and U1290 (N_1290,In_155,In_283);
and U1291 (N_1291,In_145,In_810);
and U1292 (N_1292,In_333,In_981);
nor U1293 (N_1293,In_77,In_403);
nor U1294 (N_1294,In_587,In_195);
or U1295 (N_1295,In_145,In_518);
and U1296 (N_1296,In_893,In_461);
nand U1297 (N_1297,In_594,In_839);
nor U1298 (N_1298,In_700,In_460);
or U1299 (N_1299,In_598,In_176);
or U1300 (N_1300,In_39,In_510);
nor U1301 (N_1301,In_541,In_531);
nand U1302 (N_1302,In_46,In_534);
or U1303 (N_1303,In_317,In_160);
nand U1304 (N_1304,In_786,In_245);
nor U1305 (N_1305,In_463,In_943);
nor U1306 (N_1306,In_455,In_72);
nor U1307 (N_1307,In_571,In_316);
or U1308 (N_1308,In_56,In_903);
nand U1309 (N_1309,In_406,In_151);
nor U1310 (N_1310,In_748,In_148);
nand U1311 (N_1311,In_54,In_212);
or U1312 (N_1312,In_71,In_315);
and U1313 (N_1313,In_368,In_172);
and U1314 (N_1314,In_786,In_986);
and U1315 (N_1315,In_716,In_968);
nor U1316 (N_1316,In_468,In_386);
nand U1317 (N_1317,In_983,In_96);
or U1318 (N_1318,In_275,In_75);
nand U1319 (N_1319,In_959,In_407);
or U1320 (N_1320,In_417,In_911);
nor U1321 (N_1321,In_956,In_704);
nor U1322 (N_1322,In_750,In_570);
and U1323 (N_1323,In_833,In_153);
or U1324 (N_1324,In_973,In_963);
nor U1325 (N_1325,In_589,In_398);
and U1326 (N_1326,In_919,In_791);
nand U1327 (N_1327,In_903,In_881);
nor U1328 (N_1328,In_301,In_235);
nor U1329 (N_1329,In_426,In_587);
and U1330 (N_1330,In_944,In_596);
or U1331 (N_1331,In_60,In_158);
nor U1332 (N_1332,In_756,In_466);
or U1333 (N_1333,In_136,In_620);
nor U1334 (N_1334,In_909,In_420);
nand U1335 (N_1335,In_262,In_665);
and U1336 (N_1336,In_623,In_103);
nand U1337 (N_1337,In_991,In_88);
nor U1338 (N_1338,In_370,In_312);
and U1339 (N_1339,In_234,In_903);
or U1340 (N_1340,In_388,In_440);
nor U1341 (N_1341,In_214,In_246);
or U1342 (N_1342,In_27,In_734);
nor U1343 (N_1343,In_274,In_139);
nor U1344 (N_1344,In_688,In_973);
xor U1345 (N_1345,In_262,In_136);
nor U1346 (N_1346,In_331,In_791);
nand U1347 (N_1347,In_644,In_25);
nand U1348 (N_1348,In_754,In_866);
nor U1349 (N_1349,In_29,In_561);
nor U1350 (N_1350,In_945,In_461);
or U1351 (N_1351,In_255,In_955);
and U1352 (N_1352,In_451,In_85);
nor U1353 (N_1353,In_988,In_639);
nor U1354 (N_1354,In_894,In_346);
or U1355 (N_1355,In_766,In_565);
or U1356 (N_1356,In_730,In_63);
nand U1357 (N_1357,In_683,In_105);
and U1358 (N_1358,In_412,In_601);
and U1359 (N_1359,In_398,In_694);
and U1360 (N_1360,In_827,In_171);
nor U1361 (N_1361,In_852,In_785);
nor U1362 (N_1362,In_297,In_516);
nor U1363 (N_1363,In_175,In_545);
and U1364 (N_1364,In_335,In_388);
nor U1365 (N_1365,In_13,In_955);
xnor U1366 (N_1366,In_470,In_895);
and U1367 (N_1367,In_314,In_350);
or U1368 (N_1368,In_271,In_566);
or U1369 (N_1369,In_453,In_410);
nand U1370 (N_1370,In_848,In_559);
or U1371 (N_1371,In_282,In_576);
xnor U1372 (N_1372,In_346,In_278);
nor U1373 (N_1373,In_826,In_550);
xor U1374 (N_1374,In_984,In_175);
and U1375 (N_1375,In_306,In_414);
or U1376 (N_1376,In_356,In_652);
or U1377 (N_1377,In_690,In_983);
and U1378 (N_1378,In_849,In_150);
nor U1379 (N_1379,In_102,In_377);
and U1380 (N_1380,In_449,In_57);
or U1381 (N_1381,In_554,In_565);
or U1382 (N_1382,In_599,In_639);
nor U1383 (N_1383,In_525,In_158);
nor U1384 (N_1384,In_302,In_811);
nand U1385 (N_1385,In_13,In_973);
nand U1386 (N_1386,In_981,In_348);
nand U1387 (N_1387,In_671,In_513);
nor U1388 (N_1388,In_60,In_956);
nor U1389 (N_1389,In_201,In_591);
and U1390 (N_1390,In_369,In_40);
nand U1391 (N_1391,In_175,In_331);
nand U1392 (N_1392,In_209,In_923);
or U1393 (N_1393,In_63,In_182);
and U1394 (N_1394,In_623,In_436);
or U1395 (N_1395,In_429,In_292);
xor U1396 (N_1396,In_454,In_178);
and U1397 (N_1397,In_605,In_598);
or U1398 (N_1398,In_679,In_635);
nand U1399 (N_1399,In_182,In_504);
nand U1400 (N_1400,In_713,In_583);
and U1401 (N_1401,In_419,In_876);
nand U1402 (N_1402,In_305,In_747);
nor U1403 (N_1403,In_146,In_521);
or U1404 (N_1404,In_699,In_867);
nor U1405 (N_1405,In_789,In_21);
and U1406 (N_1406,In_245,In_691);
nor U1407 (N_1407,In_679,In_270);
nor U1408 (N_1408,In_266,In_654);
and U1409 (N_1409,In_213,In_483);
or U1410 (N_1410,In_260,In_822);
or U1411 (N_1411,In_963,In_459);
or U1412 (N_1412,In_844,In_367);
and U1413 (N_1413,In_696,In_490);
nand U1414 (N_1414,In_762,In_761);
or U1415 (N_1415,In_523,In_985);
nor U1416 (N_1416,In_98,In_430);
nand U1417 (N_1417,In_303,In_635);
nand U1418 (N_1418,In_766,In_88);
nor U1419 (N_1419,In_96,In_285);
nor U1420 (N_1420,In_44,In_57);
nand U1421 (N_1421,In_217,In_320);
or U1422 (N_1422,In_765,In_196);
or U1423 (N_1423,In_185,In_61);
and U1424 (N_1424,In_885,In_64);
nand U1425 (N_1425,In_844,In_561);
nand U1426 (N_1426,In_901,In_703);
nor U1427 (N_1427,In_24,In_238);
nand U1428 (N_1428,In_933,In_271);
or U1429 (N_1429,In_58,In_364);
nor U1430 (N_1430,In_551,In_377);
or U1431 (N_1431,In_469,In_130);
nor U1432 (N_1432,In_83,In_154);
or U1433 (N_1433,In_626,In_976);
nor U1434 (N_1434,In_763,In_515);
or U1435 (N_1435,In_905,In_983);
nor U1436 (N_1436,In_151,In_248);
and U1437 (N_1437,In_25,In_361);
and U1438 (N_1438,In_543,In_200);
nand U1439 (N_1439,In_113,In_170);
or U1440 (N_1440,In_705,In_179);
and U1441 (N_1441,In_825,In_953);
or U1442 (N_1442,In_521,In_187);
nand U1443 (N_1443,In_584,In_368);
nor U1444 (N_1444,In_819,In_651);
or U1445 (N_1445,In_44,In_615);
and U1446 (N_1446,In_784,In_837);
nor U1447 (N_1447,In_164,In_218);
nand U1448 (N_1448,In_892,In_699);
xnor U1449 (N_1449,In_187,In_607);
and U1450 (N_1450,In_603,In_375);
nor U1451 (N_1451,In_59,In_28);
nand U1452 (N_1452,In_492,In_966);
and U1453 (N_1453,In_387,In_782);
nand U1454 (N_1454,In_79,In_276);
or U1455 (N_1455,In_463,In_963);
or U1456 (N_1456,In_850,In_446);
and U1457 (N_1457,In_464,In_118);
nor U1458 (N_1458,In_146,In_949);
or U1459 (N_1459,In_504,In_64);
nand U1460 (N_1460,In_130,In_294);
and U1461 (N_1461,In_23,In_417);
and U1462 (N_1462,In_755,In_777);
nand U1463 (N_1463,In_238,In_201);
nor U1464 (N_1464,In_944,In_535);
nor U1465 (N_1465,In_480,In_291);
nor U1466 (N_1466,In_740,In_647);
or U1467 (N_1467,In_140,In_928);
or U1468 (N_1468,In_970,In_554);
nand U1469 (N_1469,In_98,In_950);
and U1470 (N_1470,In_101,In_171);
or U1471 (N_1471,In_579,In_441);
nor U1472 (N_1472,In_909,In_660);
nand U1473 (N_1473,In_35,In_912);
nor U1474 (N_1474,In_533,In_588);
nor U1475 (N_1475,In_784,In_539);
nand U1476 (N_1476,In_249,In_197);
nor U1477 (N_1477,In_133,In_462);
or U1478 (N_1478,In_205,In_698);
or U1479 (N_1479,In_242,In_541);
or U1480 (N_1480,In_674,In_428);
and U1481 (N_1481,In_611,In_817);
nor U1482 (N_1482,In_691,In_47);
and U1483 (N_1483,In_727,In_126);
nand U1484 (N_1484,In_852,In_907);
nor U1485 (N_1485,In_513,In_659);
nand U1486 (N_1486,In_18,In_703);
or U1487 (N_1487,In_640,In_857);
and U1488 (N_1488,In_728,In_891);
or U1489 (N_1489,In_880,In_667);
or U1490 (N_1490,In_244,In_497);
nand U1491 (N_1491,In_511,In_167);
or U1492 (N_1492,In_449,In_499);
nor U1493 (N_1493,In_180,In_445);
nor U1494 (N_1494,In_151,In_325);
nand U1495 (N_1495,In_233,In_987);
or U1496 (N_1496,In_886,In_246);
and U1497 (N_1497,In_807,In_584);
and U1498 (N_1498,In_542,In_268);
nor U1499 (N_1499,In_807,In_542);
and U1500 (N_1500,In_668,In_893);
nor U1501 (N_1501,In_519,In_238);
and U1502 (N_1502,In_113,In_208);
nand U1503 (N_1503,In_235,In_712);
nor U1504 (N_1504,In_883,In_90);
nand U1505 (N_1505,In_738,In_192);
nor U1506 (N_1506,In_833,In_904);
or U1507 (N_1507,In_662,In_425);
nor U1508 (N_1508,In_248,In_664);
nand U1509 (N_1509,In_623,In_122);
and U1510 (N_1510,In_925,In_773);
and U1511 (N_1511,In_327,In_425);
and U1512 (N_1512,In_796,In_469);
or U1513 (N_1513,In_577,In_68);
or U1514 (N_1514,In_815,In_619);
nand U1515 (N_1515,In_667,In_29);
and U1516 (N_1516,In_893,In_859);
nand U1517 (N_1517,In_538,In_894);
and U1518 (N_1518,In_66,In_303);
nor U1519 (N_1519,In_419,In_830);
or U1520 (N_1520,In_710,In_805);
or U1521 (N_1521,In_593,In_519);
and U1522 (N_1522,In_465,In_420);
nand U1523 (N_1523,In_922,In_450);
or U1524 (N_1524,In_637,In_937);
nand U1525 (N_1525,In_312,In_923);
and U1526 (N_1526,In_174,In_516);
nor U1527 (N_1527,In_958,In_103);
nor U1528 (N_1528,In_983,In_288);
and U1529 (N_1529,In_619,In_864);
nor U1530 (N_1530,In_315,In_618);
or U1531 (N_1531,In_738,In_783);
nor U1532 (N_1532,In_728,In_403);
nand U1533 (N_1533,In_790,In_503);
and U1534 (N_1534,In_614,In_890);
or U1535 (N_1535,In_775,In_414);
nand U1536 (N_1536,In_618,In_959);
and U1537 (N_1537,In_527,In_696);
and U1538 (N_1538,In_354,In_265);
nor U1539 (N_1539,In_458,In_37);
nor U1540 (N_1540,In_142,In_909);
nand U1541 (N_1541,In_643,In_808);
and U1542 (N_1542,In_831,In_19);
nand U1543 (N_1543,In_165,In_466);
nor U1544 (N_1544,In_921,In_135);
and U1545 (N_1545,In_509,In_345);
or U1546 (N_1546,In_891,In_723);
and U1547 (N_1547,In_638,In_790);
nand U1548 (N_1548,In_491,In_950);
and U1549 (N_1549,In_770,In_102);
nor U1550 (N_1550,In_775,In_298);
and U1551 (N_1551,In_838,In_158);
nand U1552 (N_1552,In_934,In_332);
and U1553 (N_1553,In_456,In_37);
or U1554 (N_1554,In_39,In_656);
nand U1555 (N_1555,In_408,In_682);
nand U1556 (N_1556,In_970,In_638);
nor U1557 (N_1557,In_706,In_349);
nor U1558 (N_1558,In_479,In_317);
and U1559 (N_1559,In_232,In_890);
and U1560 (N_1560,In_644,In_34);
nand U1561 (N_1561,In_910,In_187);
or U1562 (N_1562,In_256,In_423);
and U1563 (N_1563,In_20,In_121);
nor U1564 (N_1564,In_337,In_360);
or U1565 (N_1565,In_896,In_827);
and U1566 (N_1566,In_137,In_970);
nor U1567 (N_1567,In_854,In_458);
nor U1568 (N_1568,In_492,In_209);
and U1569 (N_1569,In_682,In_790);
nand U1570 (N_1570,In_80,In_49);
or U1571 (N_1571,In_627,In_952);
or U1572 (N_1572,In_127,In_734);
and U1573 (N_1573,In_477,In_231);
and U1574 (N_1574,In_953,In_75);
nor U1575 (N_1575,In_337,In_474);
or U1576 (N_1576,In_810,In_557);
and U1577 (N_1577,In_1,In_202);
and U1578 (N_1578,In_123,In_999);
or U1579 (N_1579,In_765,In_463);
nor U1580 (N_1580,In_273,In_147);
or U1581 (N_1581,In_777,In_645);
or U1582 (N_1582,In_739,In_445);
or U1583 (N_1583,In_655,In_756);
or U1584 (N_1584,In_512,In_831);
nor U1585 (N_1585,In_849,In_315);
nor U1586 (N_1586,In_821,In_25);
nor U1587 (N_1587,In_708,In_922);
and U1588 (N_1588,In_631,In_268);
or U1589 (N_1589,In_114,In_897);
or U1590 (N_1590,In_327,In_125);
or U1591 (N_1591,In_835,In_486);
nand U1592 (N_1592,In_195,In_651);
nor U1593 (N_1593,In_888,In_570);
nor U1594 (N_1594,In_702,In_214);
nor U1595 (N_1595,In_957,In_665);
nor U1596 (N_1596,In_741,In_957);
nand U1597 (N_1597,In_182,In_172);
nor U1598 (N_1598,In_425,In_666);
and U1599 (N_1599,In_196,In_683);
nor U1600 (N_1600,In_894,In_490);
or U1601 (N_1601,In_973,In_714);
xor U1602 (N_1602,In_372,In_4);
nand U1603 (N_1603,In_68,In_314);
nand U1604 (N_1604,In_460,In_892);
or U1605 (N_1605,In_636,In_387);
nand U1606 (N_1606,In_522,In_712);
nor U1607 (N_1607,In_449,In_629);
and U1608 (N_1608,In_8,In_922);
or U1609 (N_1609,In_906,In_699);
nand U1610 (N_1610,In_273,In_315);
and U1611 (N_1611,In_95,In_218);
or U1612 (N_1612,In_378,In_901);
nor U1613 (N_1613,In_454,In_162);
and U1614 (N_1614,In_673,In_296);
and U1615 (N_1615,In_427,In_169);
or U1616 (N_1616,In_654,In_606);
or U1617 (N_1617,In_119,In_499);
or U1618 (N_1618,In_385,In_258);
and U1619 (N_1619,In_679,In_166);
nand U1620 (N_1620,In_53,In_475);
or U1621 (N_1621,In_238,In_863);
and U1622 (N_1622,In_209,In_980);
or U1623 (N_1623,In_523,In_154);
nor U1624 (N_1624,In_675,In_674);
nor U1625 (N_1625,In_537,In_295);
nand U1626 (N_1626,In_428,In_611);
and U1627 (N_1627,In_912,In_632);
and U1628 (N_1628,In_12,In_673);
or U1629 (N_1629,In_154,In_873);
nand U1630 (N_1630,In_86,In_599);
or U1631 (N_1631,In_952,In_413);
and U1632 (N_1632,In_815,In_643);
nor U1633 (N_1633,In_894,In_72);
or U1634 (N_1634,In_986,In_814);
nor U1635 (N_1635,In_345,In_897);
or U1636 (N_1636,In_216,In_541);
nand U1637 (N_1637,In_933,In_275);
nor U1638 (N_1638,In_597,In_727);
and U1639 (N_1639,In_686,In_324);
nand U1640 (N_1640,In_409,In_703);
or U1641 (N_1641,In_947,In_136);
and U1642 (N_1642,In_609,In_514);
nand U1643 (N_1643,In_188,In_672);
nand U1644 (N_1644,In_877,In_765);
nor U1645 (N_1645,In_615,In_311);
nor U1646 (N_1646,In_536,In_89);
nor U1647 (N_1647,In_632,In_771);
and U1648 (N_1648,In_349,In_383);
nor U1649 (N_1649,In_380,In_972);
nand U1650 (N_1650,In_862,In_65);
nor U1651 (N_1651,In_766,In_40);
and U1652 (N_1652,In_93,In_107);
and U1653 (N_1653,In_102,In_912);
xnor U1654 (N_1654,In_212,In_676);
nor U1655 (N_1655,In_958,In_591);
and U1656 (N_1656,In_369,In_411);
nand U1657 (N_1657,In_13,In_56);
nand U1658 (N_1658,In_282,In_926);
or U1659 (N_1659,In_117,In_74);
or U1660 (N_1660,In_359,In_549);
and U1661 (N_1661,In_550,In_848);
or U1662 (N_1662,In_991,In_924);
and U1663 (N_1663,In_678,In_747);
nand U1664 (N_1664,In_326,In_472);
or U1665 (N_1665,In_570,In_691);
nand U1666 (N_1666,In_393,In_959);
nand U1667 (N_1667,In_942,In_266);
and U1668 (N_1668,In_508,In_555);
nand U1669 (N_1669,In_800,In_980);
or U1670 (N_1670,In_196,In_869);
nand U1671 (N_1671,In_994,In_516);
nor U1672 (N_1672,In_736,In_637);
nand U1673 (N_1673,In_884,In_350);
and U1674 (N_1674,In_345,In_387);
nor U1675 (N_1675,In_771,In_813);
and U1676 (N_1676,In_729,In_787);
and U1677 (N_1677,In_693,In_78);
or U1678 (N_1678,In_557,In_901);
or U1679 (N_1679,In_670,In_896);
and U1680 (N_1680,In_465,In_373);
nand U1681 (N_1681,In_565,In_689);
or U1682 (N_1682,In_205,In_817);
or U1683 (N_1683,In_504,In_2);
or U1684 (N_1684,In_318,In_864);
nor U1685 (N_1685,In_141,In_490);
nand U1686 (N_1686,In_473,In_881);
and U1687 (N_1687,In_539,In_295);
nand U1688 (N_1688,In_793,In_235);
nand U1689 (N_1689,In_237,In_37);
or U1690 (N_1690,In_741,In_932);
and U1691 (N_1691,In_376,In_485);
nand U1692 (N_1692,In_499,In_541);
nand U1693 (N_1693,In_910,In_306);
nor U1694 (N_1694,In_433,In_827);
nor U1695 (N_1695,In_359,In_497);
nand U1696 (N_1696,In_308,In_536);
or U1697 (N_1697,In_907,In_236);
and U1698 (N_1698,In_821,In_449);
nor U1699 (N_1699,In_42,In_221);
nand U1700 (N_1700,In_258,In_973);
and U1701 (N_1701,In_352,In_537);
and U1702 (N_1702,In_65,In_758);
nor U1703 (N_1703,In_42,In_672);
and U1704 (N_1704,In_897,In_472);
nand U1705 (N_1705,In_191,In_571);
or U1706 (N_1706,In_142,In_215);
and U1707 (N_1707,In_252,In_485);
nor U1708 (N_1708,In_354,In_98);
nand U1709 (N_1709,In_197,In_604);
or U1710 (N_1710,In_811,In_621);
nor U1711 (N_1711,In_746,In_733);
nand U1712 (N_1712,In_174,In_665);
nand U1713 (N_1713,In_748,In_646);
nand U1714 (N_1714,In_900,In_596);
or U1715 (N_1715,In_588,In_131);
and U1716 (N_1716,In_283,In_837);
and U1717 (N_1717,In_177,In_20);
and U1718 (N_1718,In_717,In_574);
and U1719 (N_1719,In_322,In_521);
nand U1720 (N_1720,In_567,In_410);
nor U1721 (N_1721,In_868,In_795);
nand U1722 (N_1722,In_37,In_880);
nor U1723 (N_1723,In_499,In_865);
nor U1724 (N_1724,In_906,In_708);
or U1725 (N_1725,In_587,In_163);
or U1726 (N_1726,In_829,In_20);
and U1727 (N_1727,In_459,In_878);
or U1728 (N_1728,In_693,In_397);
nand U1729 (N_1729,In_212,In_787);
nor U1730 (N_1730,In_460,In_26);
nor U1731 (N_1731,In_830,In_872);
nor U1732 (N_1732,In_785,In_323);
nand U1733 (N_1733,In_737,In_617);
nor U1734 (N_1734,In_479,In_262);
and U1735 (N_1735,In_989,In_157);
and U1736 (N_1736,In_338,In_830);
or U1737 (N_1737,In_480,In_642);
nand U1738 (N_1738,In_337,In_828);
or U1739 (N_1739,In_853,In_318);
nor U1740 (N_1740,In_470,In_98);
nor U1741 (N_1741,In_531,In_394);
nand U1742 (N_1742,In_942,In_61);
or U1743 (N_1743,In_191,In_684);
and U1744 (N_1744,In_930,In_607);
and U1745 (N_1745,In_587,In_808);
or U1746 (N_1746,In_987,In_604);
and U1747 (N_1747,In_358,In_227);
or U1748 (N_1748,In_228,In_979);
and U1749 (N_1749,In_784,In_486);
or U1750 (N_1750,In_73,In_763);
and U1751 (N_1751,In_398,In_297);
or U1752 (N_1752,In_720,In_309);
nor U1753 (N_1753,In_733,In_879);
and U1754 (N_1754,In_309,In_71);
nand U1755 (N_1755,In_319,In_969);
nor U1756 (N_1756,In_328,In_230);
nand U1757 (N_1757,In_723,In_221);
or U1758 (N_1758,In_790,In_789);
and U1759 (N_1759,In_863,In_970);
or U1760 (N_1760,In_272,In_823);
or U1761 (N_1761,In_759,In_634);
nor U1762 (N_1762,In_370,In_58);
and U1763 (N_1763,In_869,In_319);
and U1764 (N_1764,In_368,In_713);
and U1765 (N_1765,In_682,In_216);
nor U1766 (N_1766,In_293,In_21);
or U1767 (N_1767,In_186,In_194);
nand U1768 (N_1768,In_536,In_309);
nand U1769 (N_1769,In_676,In_882);
xor U1770 (N_1770,In_911,In_67);
nor U1771 (N_1771,In_274,In_695);
nand U1772 (N_1772,In_52,In_843);
nand U1773 (N_1773,In_285,In_641);
nand U1774 (N_1774,In_950,In_940);
nor U1775 (N_1775,In_96,In_744);
and U1776 (N_1776,In_745,In_721);
and U1777 (N_1777,In_403,In_781);
nor U1778 (N_1778,In_696,In_243);
nor U1779 (N_1779,In_34,In_339);
and U1780 (N_1780,In_740,In_892);
nor U1781 (N_1781,In_993,In_7);
nor U1782 (N_1782,In_992,In_274);
and U1783 (N_1783,In_243,In_963);
nand U1784 (N_1784,In_705,In_341);
and U1785 (N_1785,In_113,In_961);
or U1786 (N_1786,In_102,In_551);
or U1787 (N_1787,In_634,In_740);
or U1788 (N_1788,In_889,In_516);
or U1789 (N_1789,In_951,In_892);
nand U1790 (N_1790,In_323,In_562);
nor U1791 (N_1791,In_41,In_598);
or U1792 (N_1792,In_273,In_216);
and U1793 (N_1793,In_325,In_367);
nor U1794 (N_1794,In_632,In_226);
nor U1795 (N_1795,In_417,In_635);
or U1796 (N_1796,In_244,In_590);
nor U1797 (N_1797,In_392,In_671);
nand U1798 (N_1798,In_312,In_105);
or U1799 (N_1799,In_580,In_15);
nor U1800 (N_1800,In_119,In_879);
or U1801 (N_1801,In_132,In_947);
nand U1802 (N_1802,In_65,In_718);
and U1803 (N_1803,In_274,In_917);
nor U1804 (N_1804,In_27,In_664);
nand U1805 (N_1805,In_44,In_196);
and U1806 (N_1806,In_673,In_202);
and U1807 (N_1807,In_837,In_430);
nand U1808 (N_1808,In_408,In_717);
nor U1809 (N_1809,In_124,In_423);
nor U1810 (N_1810,In_173,In_561);
nor U1811 (N_1811,In_285,In_463);
and U1812 (N_1812,In_265,In_739);
nand U1813 (N_1813,In_919,In_641);
nor U1814 (N_1814,In_268,In_135);
and U1815 (N_1815,In_684,In_255);
xnor U1816 (N_1816,In_506,In_32);
nand U1817 (N_1817,In_916,In_687);
and U1818 (N_1818,In_60,In_149);
or U1819 (N_1819,In_736,In_967);
nand U1820 (N_1820,In_676,In_366);
and U1821 (N_1821,In_389,In_26);
nand U1822 (N_1822,In_815,In_629);
and U1823 (N_1823,In_498,In_69);
and U1824 (N_1824,In_245,In_188);
nor U1825 (N_1825,In_425,In_231);
nor U1826 (N_1826,In_373,In_56);
and U1827 (N_1827,In_979,In_632);
and U1828 (N_1828,In_449,In_773);
or U1829 (N_1829,In_998,In_32);
nand U1830 (N_1830,In_693,In_287);
or U1831 (N_1831,In_580,In_787);
nand U1832 (N_1832,In_403,In_267);
nand U1833 (N_1833,In_300,In_913);
or U1834 (N_1834,In_592,In_517);
and U1835 (N_1835,In_149,In_694);
nor U1836 (N_1836,In_367,In_864);
nor U1837 (N_1837,In_550,In_563);
or U1838 (N_1838,In_937,In_695);
and U1839 (N_1839,In_40,In_129);
nor U1840 (N_1840,In_693,In_383);
nand U1841 (N_1841,In_294,In_754);
nor U1842 (N_1842,In_351,In_345);
xor U1843 (N_1843,In_161,In_866);
and U1844 (N_1844,In_267,In_236);
nand U1845 (N_1845,In_164,In_24);
nor U1846 (N_1846,In_113,In_657);
nand U1847 (N_1847,In_964,In_978);
or U1848 (N_1848,In_360,In_331);
or U1849 (N_1849,In_540,In_567);
or U1850 (N_1850,In_505,In_865);
nand U1851 (N_1851,In_334,In_416);
or U1852 (N_1852,In_184,In_112);
nand U1853 (N_1853,In_652,In_920);
or U1854 (N_1854,In_19,In_990);
and U1855 (N_1855,In_889,In_667);
nand U1856 (N_1856,In_244,In_241);
or U1857 (N_1857,In_73,In_302);
nor U1858 (N_1858,In_665,In_930);
and U1859 (N_1859,In_510,In_257);
or U1860 (N_1860,In_267,In_407);
or U1861 (N_1861,In_98,In_771);
nand U1862 (N_1862,In_330,In_295);
or U1863 (N_1863,In_486,In_921);
and U1864 (N_1864,In_956,In_50);
nor U1865 (N_1865,In_830,In_807);
and U1866 (N_1866,In_19,In_721);
nand U1867 (N_1867,In_369,In_423);
nand U1868 (N_1868,In_751,In_291);
nand U1869 (N_1869,In_60,In_847);
nand U1870 (N_1870,In_958,In_677);
and U1871 (N_1871,In_292,In_401);
and U1872 (N_1872,In_81,In_341);
nand U1873 (N_1873,In_483,In_765);
or U1874 (N_1874,In_43,In_213);
nand U1875 (N_1875,In_227,In_871);
or U1876 (N_1876,In_527,In_771);
nor U1877 (N_1877,In_998,In_514);
nor U1878 (N_1878,In_505,In_144);
nor U1879 (N_1879,In_143,In_947);
or U1880 (N_1880,In_362,In_0);
nand U1881 (N_1881,In_408,In_487);
nand U1882 (N_1882,In_125,In_792);
nand U1883 (N_1883,In_568,In_941);
or U1884 (N_1884,In_885,In_683);
nor U1885 (N_1885,In_923,In_839);
nand U1886 (N_1886,In_682,In_995);
and U1887 (N_1887,In_458,In_413);
or U1888 (N_1888,In_999,In_145);
nand U1889 (N_1889,In_983,In_52);
or U1890 (N_1890,In_819,In_622);
or U1891 (N_1891,In_268,In_318);
nand U1892 (N_1892,In_205,In_206);
nor U1893 (N_1893,In_989,In_84);
nand U1894 (N_1894,In_605,In_261);
or U1895 (N_1895,In_668,In_138);
or U1896 (N_1896,In_559,In_342);
and U1897 (N_1897,In_919,In_374);
or U1898 (N_1898,In_182,In_989);
or U1899 (N_1899,In_85,In_311);
nand U1900 (N_1900,In_249,In_339);
nor U1901 (N_1901,In_581,In_728);
nand U1902 (N_1902,In_285,In_720);
or U1903 (N_1903,In_48,In_287);
or U1904 (N_1904,In_606,In_7);
nand U1905 (N_1905,In_830,In_159);
nand U1906 (N_1906,In_830,In_373);
and U1907 (N_1907,In_305,In_934);
and U1908 (N_1908,In_707,In_127);
and U1909 (N_1909,In_316,In_55);
or U1910 (N_1910,In_169,In_493);
and U1911 (N_1911,In_235,In_384);
nor U1912 (N_1912,In_530,In_151);
nand U1913 (N_1913,In_705,In_950);
xor U1914 (N_1914,In_649,In_310);
nand U1915 (N_1915,In_834,In_805);
and U1916 (N_1916,In_833,In_956);
nor U1917 (N_1917,In_649,In_410);
nand U1918 (N_1918,In_828,In_899);
or U1919 (N_1919,In_275,In_190);
nor U1920 (N_1920,In_898,In_822);
nand U1921 (N_1921,In_723,In_546);
xnor U1922 (N_1922,In_238,In_414);
and U1923 (N_1923,In_293,In_216);
or U1924 (N_1924,In_207,In_909);
nand U1925 (N_1925,In_218,In_434);
and U1926 (N_1926,In_246,In_847);
nand U1927 (N_1927,In_417,In_909);
or U1928 (N_1928,In_262,In_731);
and U1929 (N_1929,In_68,In_721);
and U1930 (N_1930,In_679,In_867);
or U1931 (N_1931,In_63,In_815);
nand U1932 (N_1932,In_71,In_877);
nor U1933 (N_1933,In_495,In_280);
or U1934 (N_1934,In_13,In_238);
and U1935 (N_1935,In_202,In_824);
or U1936 (N_1936,In_377,In_977);
nand U1937 (N_1937,In_214,In_403);
or U1938 (N_1938,In_675,In_825);
nor U1939 (N_1939,In_154,In_608);
and U1940 (N_1940,In_851,In_546);
nor U1941 (N_1941,In_387,In_23);
or U1942 (N_1942,In_553,In_547);
nor U1943 (N_1943,In_781,In_674);
nand U1944 (N_1944,In_437,In_955);
xnor U1945 (N_1945,In_540,In_159);
and U1946 (N_1946,In_264,In_191);
or U1947 (N_1947,In_310,In_177);
and U1948 (N_1948,In_704,In_719);
and U1949 (N_1949,In_596,In_989);
nor U1950 (N_1950,In_962,In_761);
nor U1951 (N_1951,In_197,In_224);
nand U1952 (N_1952,In_429,In_975);
or U1953 (N_1953,In_169,In_870);
or U1954 (N_1954,In_649,In_749);
nor U1955 (N_1955,In_433,In_917);
and U1956 (N_1956,In_192,In_142);
nand U1957 (N_1957,In_31,In_159);
nand U1958 (N_1958,In_950,In_485);
nand U1959 (N_1959,In_798,In_355);
and U1960 (N_1960,In_410,In_591);
and U1961 (N_1961,In_939,In_292);
and U1962 (N_1962,In_377,In_524);
nand U1963 (N_1963,In_66,In_763);
or U1964 (N_1964,In_233,In_442);
nand U1965 (N_1965,In_494,In_73);
nor U1966 (N_1966,In_31,In_412);
or U1967 (N_1967,In_683,In_866);
nand U1968 (N_1968,In_214,In_186);
and U1969 (N_1969,In_441,In_168);
nor U1970 (N_1970,In_630,In_45);
nor U1971 (N_1971,In_397,In_371);
nand U1972 (N_1972,In_551,In_592);
nand U1973 (N_1973,In_572,In_90);
nand U1974 (N_1974,In_687,In_979);
and U1975 (N_1975,In_606,In_362);
nand U1976 (N_1976,In_62,In_688);
and U1977 (N_1977,In_767,In_455);
and U1978 (N_1978,In_287,In_440);
nand U1979 (N_1979,In_338,In_226);
nor U1980 (N_1980,In_317,In_537);
nor U1981 (N_1981,In_927,In_901);
nor U1982 (N_1982,In_256,In_477);
and U1983 (N_1983,In_128,In_290);
nand U1984 (N_1984,In_746,In_405);
or U1985 (N_1985,In_229,In_546);
or U1986 (N_1986,In_477,In_54);
nor U1987 (N_1987,In_937,In_833);
or U1988 (N_1988,In_727,In_811);
or U1989 (N_1989,In_222,In_535);
and U1990 (N_1990,In_749,In_835);
and U1991 (N_1991,In_863,In_88);
and U1992 (N_1992,In_811,In_947);
or U1993 (N_1993,In_302,In_939);
nor U1994 (N_1994,In_280,In_338);
nor U1995 (N_1995,In_173,In_213);
and U1996 (N_1996,In_684,In_275);
nand U1997 (N_1997,In_360,In_171);
nand U1998 (N_1998,In_493,In_756);
or U1999 (N_1999,In_470,In_481);
nand U2000 (N_2000,N_25,N_1979);
and U2001 (N_2001,N_309,N_232);
and U2002 (N_2002,N_819,N_766);
or U2003 (N_2003,N_624,N_854);
xnor U2004 (N_2004,N_1635,N_425);
nor U2005 (N_2005,N_932,N_1856);
or U2006 (N_2006,N_851,N_9);
and U2007 (N_2007,N_1265,N_432);
nor U2008 (N_2008,N_1884,N_1093);
nand U2009 (N_2009,N_1398,N_513);
and U2010 (N_2010,N_570,N_1385);
and U2011 (N_2011,N_174,N_1606);
nand U2012 (N_2012,N_848,N_339);
nand U2013 (N_2013,N_588,N_1793);
or U2014 (N_2014,N_180,N_1462);
nor U2015 (N_2015,N_844,N_1255);
nand U2016 (N_2016,N_930,N_1573);
nor U2017 (N_2017,N_1263,N_1951);
and U2018 (N_2018,N_1413,N_1156);
nor U2019 (N_2019,N_716,N_1251);
or U2020 (N_2020,N_1992,N_979);
or U2021 (N_2021,N_95,N_578);
and U2022 (N_2022,N_35,N_1092);
nor U2023 (N_2023,N_1318,N_857);
nand U2024 (N_2024,N_1134,N_293);
and U2025 (N_2025,N_1938,N_1819);
and U2026 (N_2026,N_1923,N_254);
nand U2027 (N_2027,N_1315,N_1408);
and U2028 (N_2028,N_1136,N_236);
or U2029 (N_2029,N_158,N_1441);
nand U2030 (N_2030,N_650,N_303);
or U2031 (N_2031,N_885,N_1839);
and U2032 (N_2032,N_242,N_850);
nand U2033 (N_2033,N_1827,N_1066);
nor U2034 (N_2034,N_1632,N_894);
and U2035 (N_2035,N_1630,N_792);
and U2036 (N_2036,N_1192,N_1191);
or U2037 (N_2037,N_1258,N_1120);
and U2038 (N_2038,N_1763,N_1650);
or U2039 (N_2039,N_1200,N_1718);
and U2040 (N_2040,N_247,N_1533);
nor U2041 (N_2041,N_1905,N_1236);
or U2042 (N_2042,N_780,N_1284);
nor U2043 (N_2043,N_1985,N_1877);
nor U2044 (N_2044,N_1607,N_1813);
or U2045 (N_2045,N_1377,N_1198);
and U2046 (N_2046,N_1727,N_892);
and U2047 (N_2047,N_1154,N_310);
and U2048 (N_2048,N_1729,N_1662);
nand U2049 (N_2049,N_7,N_1799);
or U2050 (N_2050,N_718,N_1971);
nand U2051 (N_2051,N_140,N_1286);
nand U2052 (N_2052,N_586,N_559);
or U2053 (N_2053,N_1340,N_132);
nand U2054 (N_2054,N_1476,N_241);
and U2055 (N_2055,N_1144,N_1464);
nand U2056 (N_2056,N_499,N_1683);
nand U2057 (N_2057,N_1139,N_1062);
nor U2058 (N_2058,N_1453,N_1959);
nor U2059 (N_2059,N_325,N_258);
and U2060 (N_2060,N_1689,N_572);
nor U2061 (N_2061,N_878,N_643);
nand U2062 (N_2062,N_1695,N_552);
nand U2063 (N_2063,N_520,N_873);
and U2064 (N_2064,N_1367,N_667);
nand U2065 (N_2065,N_1007,N_1493);
nor U2066 (N_2066,N_739,N_1457);
nand U2067 (N_2067,N_743,N_164);
and U2068 (N_2068,N_323,N_738);
or U2069 (N_2069,N_429,N_705);
nor U2070 (N_2070,N_218,N_1488);
nor U2071 (N_2071,N_99,N_615);
or U2072 (N_2072,N_1230,N_1085);
nor U2073 (N_2073,N_1392,N_1158);
or U2074 (N_2074,N_267,N_1203);
and U2075 (N_2075,N_67,N_647);
nand U2076 (N_2076,N_16,N_126);
nor U2077 (N_2077,N_243,N_1348);
or U2078 (N_2078,N_379,N_188);
nand U2079 (N_2079,N_1953,N_970);
or U2080 (N_2080,N_1925,N_1922);
or U2081 (N_2081,N_1794,N_1305);
nand U2082 (N_2082,N_637,N_1771);
nor U2083 (N_2083,N_1954,N_675);
nor U2084 (N_2084,N_61,N_1009);
nand U2085 (N_2085,N_929,N_250);
nor U2086 (N_2086,N_210,N_110);
or U2087 (N_2087,N_1436,N_1603);
or U2088 (N_2088,N_708,N_266);
nor U2089 (N_2089,N_934,N_428);
and U2090 (N_2090,N_386,N_220);
nor U2091 (N_2091,N_64,N_1789);
nor U2092 (N_2092,N_1514,N_1547);
or U2093 (N_2093,N_1297,N_1430);
nor U2094 (N_2094,N_665,N_385);
or U2095 (N_2095,N_540,N_1809);
or U2096 (N_2096,N_1157,N_629);
nor U2097 (N_2097,N_1048,N_418);
and U2098 (N_2098,N_1679,N_97);
or U2099 (N_2099,N_451,N_1838);
and U2100 (N_2100,N_1162,N_1122);
or U2101 (N_2101,N_1468,N_1661);
or U2102 (N_2102,N_1282,N_494);
nor U2103 (N_2103,N_461,N_1014);
xnor U2104 (N_2104,N_181,N_1750);
or U2105 (N_2105,N_311,N_173);
and U2106 (N_2106,N_205,N_608);
nor U2107 (N_2107,N_918,N_1023);
nand U2108 (N_2108,N_294,N_1339);
nand U2109 (N_2109,N_1024,N_1015);
xnor U2110 (N_2110,N_92,N_495);
nor U2111 (N_2111,N_512,N_147);
nand U2112 (N_2112,N_1732,N_1072);
or U2113 (N_2113,N_1356,N_13);
and U2114 (N_2114,N_797,N_427);
nand U2115 (N_2115,N_1966,N_1059);
nor U2116 (N_2116,N_1918,N_1902);
nor U2117 (N_2117,N_685,N_1596);
and U2118 (N_2118,N_1345,N_858);
and U2119 (N_2119,N_337,N_1444);
xor U2120 (N_2120,N_605,N_868);
nand U2121 (N_2121,N_237,N_690);
or U2122 (N_2122,N_1990,N_413);
nand U2123 (N_2123,N_1214,N_1842);
nand U2124 (N_2124,N_1113,N_1302);
nand U2125 (N_2125,N_723,N_262);
nor U2126 (N_2126,N_1957,N_621);
or U2127 (N_2127,N_1327,N_1491);
or U2128 (N_2128,N_26,N_627);
and U2129 (N_2129,N_772,N_872);
and U2130 (N_2130,N_1574,N_1290);
or U2131 (N_2131,N_1848,N_435);
and U2132 (N_2132,N_1554,N_1676);
and U2133 (N_2133,N_1527,N_228);
nor U2134 (N_2134,N_1768,N_1640);
nor U2135 (N_2135,N_503,N_693);
and U2136 (N_2136,N_1833,N_1802);
nor U2137 (N_2137,N_815,N_1145);
or U2138 (N_2138,N_617,N_1222);
or U2139 (N_2139,N_369,N_391);
and U2140 (N_2140,N_1897,N_1930);
and U2141 (N_2141,N_353,N_689);
nand U2142 (N_2142,N_573,N_1197);
and U2143 (N_2143,N_1351,N_1455);
nor U2144 (N_2144,N_1396,N_119);
and U2145 (N_2145,N_289,N_421);
and U2146 (N_2146,N_717,N_1347);
or U2147 (N_2147,N_1142,N_457);
and U2148 (N_2148,N_1713,N_742);
or U2149 (N_2149,N_1940,N_1536);
nor U2150 (N_2150,N_424,N_922);
nand U2151 (N_2151,N_721,N_448);
or U2152 (N_2152,N_146,N_1691);
nor U2153 (N_2153,N_749,N_1811);
and U2154 (N_2154,N_980,N_996);
nand U2155 (N_2155,N_1497,N_216);
nor U2156 (N_2156,N_1111,N_155);
and U2157 (N_2157,N_1781,N_1878);
nand U2158 (N_2158,N_745,N_877);
and U2159 (N_2159,N_944,N_998);
or U2160 (N_2160,N_567,N_833);
or U2161 (N_2161,N_1764,N_1804);
and U2162 (N_2162,N_1267,N_1776);
nor U2163 (N_2163,N_1460,N_808);
nor U2164 (N_2164,N_498,N_1636);
and U2165 (N_2165,N_1449,N_886);
nand U2166 (N_2166,N_238,N_985);
nor U2167 (N_2167,N_636,N_1354);
or U2168 (N_2168,N_1107,N_1423);
xor U2169 (N_2169,N_1829,N_838);
and U2170 (N_2170,N_1201,N_1745);
nand U2171 (N_2171,N_449,N_317);
nor U2172 (N_2172,N_1390,N_1323);
and U2173 (N_2173,N_662,N_1098);
nand U2174 (N_2174,N_1866,N_1109);
nor U2175 (N_2175,N_18,N_37);
and U2176 (N_2176,N_56,N_684);
and U2177 (N_2177,N_1049,N_1507);
and U2178 (N_2178,N_1053,N_1761);
xor U2179 (N_2179,N_1765,N_876);
and U2180 (N_2180,N_1993,N_1245);
or U2181 (N_2181,N_1257,N_398);
or U2182 (N_2182,N_1461,N_1767);
or U2183 (N_2183,N_1709,N_328);
and U2184 (N_2184,N_763,N_1946);
nand U2185 (N_2185,N_924,N_1517);
or U2186 (N_2186,N_1097,N_1091);
nand U2187 (N_2187,N_1594,N_1556);
nand U2188 (N_2188,N_1019,N_1983);
nor U2189 (N_2189,N_889,N_547);
nand U2190 (N_2190,N_1341,N_344);
nor U2191 (N_2191,N_1199,N_91);
or U2192 (N_2192,N_41,N_0);
or U2193 (N_2193,N_1981,N_1645);
and U2194 (N_2194,N_1118,N_965);
nor U2195 (N_2195,N_1188,N_1620);
nor U2196 (N_2196,N_1006,N_656);
nand U2197 (N_2197,N_52,N_1279);
or U2198 (N_2198,N_1343,N_810);
nand U2199 (N_2199,N_1090,N_1646);
nand U2200 (N_2200,N_913,N_1688);
nor U2201 (N_2201,N_1686,N_1693);
nor U2202 (N_2202,N_327,N_1889);
or U2203 (N_2203,N_402,N_1361);
nor U2204 (N_2204,N_1314,N_246);
and U2205 (N_2205,N_541,N_156);
and U2206 (N_2206,N_471,N_964);
nand U2207 (N_2207,N_931,N_297);
and U2208 (N_2208,N_1296,N_1880);
nand U2209 (N_2209,N_1963,N_1967);
nand U2210 (N_2210,N_1028,N_816);
nor U2211 (N_2211,N_1939,N_1151);
nand U2212 (N_2212,N_1179,N_1475);
or U2213 (N_2213,N_1784,N_505);
or U2214 (N_2214,N_1836,N_1974);
nand U2215 (N_2215,N_1569,N_312);
or U2216 (N_2216,N_1894,N_224);
nand U2217 (N_2217,N_145,N_1546);
nor U2218 (N_2218,N_1847,N_1772);
nor U2219 (N_2219,N_1416,N_1238);
or U2220 (N_2220,N_23,N_807);
or U2221 (N_2221,N_1037,N_1952);
nand U2222 (N_2222,N_862,N_322);
and U2223 (N_2223,N_804,N_154);
or U2224 (N_2224,N_192,N_691);
and U2225 (N_2225,N_779,N_740);
nand U2226 (N_2226,N_153,N_999);
or U2227 (N_2227,N_888,N_1926);
or U2228 (N_2228,N_925,N_687);
nor U2229 (N_2229,N_343,N_1672);
or U2230 (N_2230,N_698,N_1184);
nor U2231 (N_2231,N_1183,N_1355);
nor U2232 (N_2232,N_1874,N_200);
nor U2233 (N_2233,N_209,N_407);
nor U2234 (N_2234,N_21,N_112);
and U2235 (N_2235,N_275,N_1851);
or U2236 (N_2236,N_383,N_364);
and U2237 (N_2237,N_372,N_426);
nor U2238 (N_2238,N_479,N_839);
nor U2239 (N_2239,N_744,N_829);
nand U2240 (N_2240,N_758,N_522);
and U2241 (N_2241,N_1235,N_329);
and U2242 (N_2242,N_1420,N_1775);
nand U2243 (N_2243,N_20,N_1239);
nand U2244 (N_2244,N_57,N_1885);
and U2245 (N_2245,N_769,N_211);
or U2246 (N_2246,N_890,N_515);
or U2247 (N_2247,N_768,N_1671);
or U2248 (N_2248,N_347,N_342);
nor U2249 (N_2249,N_1432,N_511);
and U2250 (N_2250,N_1247,N_1701);
and U2251 (N_2251,N_579,N_142);
or U2252 (N_2252,N_732,N_855);
nor U2253 (N_2253,N_1575,N_1807);
nand U2254 (N_2254,N_1281,N_406);
nor U2255 (N_2255,N_1526,N_1528);
and U2256 (N_2256,N_361,N_1405);
xor U2257 (N_2257,N_1210,N_350);
nand U2258 (N_2258,N_1855,N_405);
nor U2259 (N_2259,N_1696,N_194);
or U2260 (N_2260,N_923,N_561);
nand U2261 (N_2261,N_1052,N_22);
and U2262 (N_2262,N_1625,N_530);
nand U2263 (N_2263,N_230,N_414);
nand U2264 (N_2264,N_197,N_82);
nor U2265 (N_2265,N_574,N_46);
nor U2266 (N_2266,N_355,N_1599);
nor U2267 (N_2267,N_287,N_86);
nand U2268 (N_2268,N_1309,N_1454);
and U2269 (N_2269,N_371,N_1393);
or U2270 (N_2270,N_504,N_601);
or U2271 (N_2271,N_416,N_442);
nor U2272 (N_2272,N_1753,N_846);
nand U2273 (N_2273,N_1288,N_1754);
nand U2274 (N_2274,N_1038,N_1384);
nand U2275 (N_2275,N_1521,N_1182);
or U2276 (N_2276,N_439,N_731);
and U2277 (N_2277,N_127,N_1433);
nand U2278 (N_2278,N_1699,N_1246);
nand U2279 (N_2279,N_582,N_984);
or U2280 (N_2280,N_938,N_1063);
and U2281 (N_2281,N_956,N_1426);
nor U2282 (N_2282,N_827,N_1806);
or U2283 (N_2283,N_1409,N_787);
and U2284 (N_2284,N_1845,N_377);
xnor U2285 (N_2285,N_186,N_1903);
or U2286 (N_2286,N_1731,N_94);
and U2287 (N_2287,N_234,N_897);
or U2288 (N_2288,N_1116,N_901);
or U2289 (N_2289,N_1796,N_419);
nand U2290 (N_2290,N_196,N_477);
or U2291 (N_2291,N_1602,N_1438);
and U2292 (N_2292,N_120,N_411);
or U2293 (N_2293,N_1896,N_1349);
nand U2294 (N_2294,N_1080,N_367);
and U2295 (N_2295,N_1338,N_1786);
or U2296 (N_2296,N_1823,N_737);
nand U2297 (N_2297,N_460,N_324);
nand U2298 (N_2298,N_1668,N_959);
nand U2299 (N_2299,N_641,N_661);
and U2300 (N_2300,N_1389,N_1648);
and U2301 (N_2301,N_49,N_162);
nand U2302 (N_2302,N_1634,N_1585);
and U2303 (N_2303,N_66,N_883);
or U2304 (N_2304,N_1976,N_939);
nor U2305 (N_2305,N_106,N_51);
nand U2306 (N_2306,N_1562,N_459);
nand U2307 (N_2307,N_300,N_899);
nor U2308 (N_2308,N_1068,N_1774);
nand U2309 (N_2309,N_1899,N_1117);
and U2310 (N_2310,N_456,N_1667);
and U2311 (N_2311,N_397,N_212);
nand U2312 (N_2312,N_1161,N_1410);
and U2313 (N_2313,N_445,N_1872);
or U2314 (N_2314,N_614,N_1081);
and U2315 (N_2315,N_764,N_783);
nor U2316 (N_2316,N_1792,N_936);
and U2317 (N_2317,N_986,N_1178);
nand U2318 (N_2318,N_226,N_651);
xor U2319 (N_2319,N_1466,N_1335);
nand U2320 (N_2320,N_1254,N_229);
nor U2321 (N_2321,N_1443,N_45);
and U2322 (N_2322,N_1143,N_1861);
and U2323 (N_2323,N_593,N_1088);
and U2324 (N_2324,N_169,N_1121);
or U2325 (N_2325,N_1368,N_648);
nand U2326 (N_2326,N_1586,N_1231);
nor U2327 (N_2327,N_235,N_746);
or U2328 (N_2328,N_871,N_1084);
nor U2329 (N_2329,N_910,N_1950);
nand U2330 (N_2330,N_1206,N_671);
or U2331 (N_2331,N_1544,N_949);
nor U2332 (N_2332,N_285,N_1032);
nand U2333 (N_2333,N_463,N_487);
nand U2334 (N_2334,N_1499,N_1463);
nor U2335 (N_2335,N_1707,N_31);
nand U2336 (N_2336,N_1275,N_700);
nor U2337 (N_2337,N_1391,N_1834);
nand U2338 (N_2338,N_748,N_1756);
and U2339 (N_2339,N_1552,N_1291);
nand U2340 (N_2340,N_895,N_507);
nand U2341 (N_2341,N_1034,N_32);
or U2342 (N_2342,N_130,N_542);
or U2343 (N_2343,N_1968,N_1232);
and U2344 (N_2344,N_616,N_893);
or U2345 (N_2345,N_770,N_971);
or U2346 (N_2346,N_1929,N_1702);
nor U2347 (N_2347,N_1808,N_58);
nor U2348 (N_2348,N_1040,N_584);
nor U2349 (N_2349,N_486,N_720);
nor U2350 (N_2350,N_1660,N_905);
nor U2351 (N_2351,N_1945,N_76);
nor U2352 (N_2352,N_248,N_724);
and U2353 (N_2353,N_1193,N_1033);
or U2354 (N_2354,N_96,N_1685);
nand U2355 (N_2355,N_1422,N_1404);
nor U2356 (N_2356,N_453,N_1094);
or U2357 (N_2357,N_767,N_812);
or U2358 (N_2358,N_592,N_587);
or U2359 (N_2359,N_356,N_115);
and U2360 (N_2360,N_1652,N_1989);
nor U2361 (N_2361,N_1705,N_77);
and U2362 (N_2362,N_231,N_1474);
nor U2363 (N_2363,N_1782,N_961);
or U2364 (N_2364,N_444,N_859);
nor U2365 (N_2365,N_1164,N_1079);
nand U2366 (N_2366,N_1213,N_562);
nor U2367 (N_2367,N_1934,N_864);
nor U2368 (N_2368,N_1451,N_784);
or U2369 (N_2369,N_1961,N_368);
or U2370 (N_2370,N_1022,N_1227);
nor U2371 (N_2371,N_251,N_1817);
nor U2372 (N_2372,N_842,N_1259);
and U2373 (N_2373,N_4,N_1492);
nand U2374 (N_2374,N_1417,N_1733);
or U2375 (N_2375,N_707,N_1130);
nor U2376 (N_2376,N_1883,N_103);
or U2377 (N_2377,N_1295,N_1843);
and U2378 (N_2378,N_575,N_945);
nor U2379 (N_2379,N_1743,N_1412);
or U2380 (N_2380,N_1129,N_1627);
nor U2381 (N_2381,N_1657,N_673);
or U2382 (N_2382,N_1555,N_53);
nand U2383 (N_2383,N_902,N_1112);
or U2384 (N_2384,N_943,N_880);
nor U2385 (N_2385,N_1036,N_1977);
and U2386 (N_2386,N_1494,N_1330);
nand U2387 (N_2387,N_652,N_835);
or U2388 (N_2388,N_1402,N_1551);
xnor U2389 (N_2389,N_433,N_1125);
nor U2390 (N_2390,N_1615,N_1788);
nor U2391 (N_2391,N_1260,N_1730);
and U2392 (N_2392,N_1477,N_1736);
nand U2393 (N_2393,N_1955,N_1508);
and U2394 (N_2394,N_431,N_1287);
and U2395 (N_2395,N_60,N_841);
and U2396 (N_2396,N_1637,N_1991);
nand U2397 (N_2397,N_1920,N_726);
nand U2398 (N_2398,N_190,N_1740);
or U2399 (N_2399,N_798,N_580);
and U2400 (N_2400,N_440,N_1293);
and U2401 (N_2401,N_114,N_1876);
nor U2402 (N_2402,N_1956,N_915);
nand U2403 (N_2403,N_304,N_1869);
nand U2404 (N_2404,N_233,N_852);
nor U2405 (N_2405,N_1987,N_947);
nor U2406 (N_2406,N_1893,N_1734);
nand U2407 (N_2407,N_1800,N_1375);
or U2408 (N_2408,N_65,N_536);
and U2409 (N_2409,N_926,N_631);
or U2410 (N_2410,N_482,N_603);
nor U2411 (N_2411,N_1450,N_245);
nor U2412 (N_2412,N_1076,N_1003);
nor U2413 (N_2413,N_1148,N_874);
nor U2414 (N_2414,N_1077,N_741);
and U2415 (N_2415,N_1386,N_1530);
or U2416 (N_2416,N_1021,N_1304);
nor U2417 (N_2417,N_1054,N_1146);
or U2418 (N_2418,N_264,N_1045);
and U2419 (N_2419,N_837,N_1868);
nand U2420 (N_2420,N_1452,N_90);
or U2421 (N_2421,N_1365,N_1172);
nor U2422 (N_2422,N_315,N_83);
or U2423 (N_2423,N_244,N_1739);
nand U2424 (N_2424,N_710,N_1372);
and U2425 (N_2425,N_1030,N_813);
nor U2426 (N_2426,N_138,N_36);
or U2427 (N_2427,N_44,N_610);
nor U2428 (N_2428,N_1888,N_1261);
nor U2429 (N_2429,N_388,N_830);
and U2430 (N_2430,N_141,N_28);
or U2431 (N_2431,N_1057,N_722);
nor U2432 (N_2432,N_1378,N_1500);
and U2433 (N_2433,N_775,N_506);
or U2434 (N_2434,N_1511,N_403);
nor U2435 (N_2435,N_912,N_1886);
nand U2436 (N_2436,N_1320,N_1818);
xor U2437 (N_2437,N_1525,N_755);
nor U2438 (N_2438,N_692,N_800);
and U2439 (N_2439,N_1609,N_734);
or U2440 (N_2440,N_150,N_134);
and U2441 (N_2441,N_1639,N_1659);
nand U2442 (N_2442,N_994,N_178);
or U2443 (N_2443,N_1780,N_600);
nand U2444 (N_2444,N_458,N_320);
nor U2445 (N_2445,N_948,N_472);
nor U2446 (N_2446,N_1519,N_1173);
or U2447 (N_2447,N_360,N_1050);
and U2448 (N_2448,N_79,N_535);
or U2449 (N_2449,N_1058,N_1310);
or U2450 (N_2450,N_989,N_69);
nor U2451 (N_2451,N_272,N_497);
and U2452 (N_2452,N_1857,N_694);
xor U2453 (N_2453,N_882,N_1470);
or U2454 (N_2454,N_394,N_1611);
and U2455 (N_2455,N_1276,N_1269);
nand U2456 (N_2456,N_1933,N_806);
nor U2457 (N_2457,N_1984,N_269);
and U2458 (N_2458,N_1988,N_1316);
and U2459 (N_2459,N_1928,N_63);
or U2460 (N_2460,N_39,N_1181);
and U2461 (N_2461,N_1841,N_551);
or U2462 (N_2462,N_566,N_1783);
nand U2463 (N_2463,N_1505,N_1658);
nor U2464 (N_2464,N_199,N_1518);
or U2465 (N_2465,N_1208,N_1710);
xnor U2466 (N_2466,N_1177,N_306);
and U2467 (N_2467,N_38,N_635);
nor U2468 (N_2468,N_480,N_1099);
nor U2469 (N_2469,N_1051,N_256);
nand U2470 (N_2470,N_831,N_866);
nor U2471 (N_2471,N_171,N_568);
nand U2472 (N_2472,N_219,N_919);
nor U2473 (N_2473,N_1155,N_863);
nor U2474 (N_2474,N_33,N_782);
and U2475 (N_2475,N_1947,N_556);
nand U2476 (N_2476,N_430,N_478);
and U2477 (N_2477,N_319,N_670);
and U2478 (N_2478,N_1949,N_330);
nand U2479 (N_2479,N_1986,N_1755);
nor U2480 (N_2480,N_881,N_1399);
or U2481 (N_2481,N_1835,N_1769);
nand U2482 (N_2482,N_1047,N_607);
xor U2483 (N_2483,N_1478,N_1618);
nor U2484 (N_2484,N_443,N_646);
or U2485 (N_2485,N_351,N_1875);
and U2486 (N_2486,N_184,N_528);
nand U2487 (N_2487,N_124,N_867);
or U2488 (N_2488,N_776,N_563);
or U2489 (N_2489,N_1656,N_1746);
nor U2490 (N_2490,N_1566,N_1434);
and U2491 (N_2491,N_1600,N_1102);
nor U2492 (N_2492,N_861,N_521);
and U2493 (N_2493,N_1026,N_1292);
nor U2494 (N_2494,N_1212,N_564);
nor U2495 (N_2495,N_532,N_252);
nor U2496 (N_2496,N_1858,N_1655);
nor U2497 (N_2497,N_729,N_1728);
or U2498 (N_2498,N_1787,N_1541);
and U2499 (N_2499,N_308,N_382);
or U2500 (N_2500,N_903,N_1317);
xnor U2501 (N_2501,N_1581,N_1010);
or U2502 (N_2502,N_273,N_1278);
nor U2503 (N_2503,N_1941,N_225);
and U2504 (N_2504,N_524,N_778);
nor U2505 (N_2505,N_1397,N_48);
xnor U2506 (N_2506,N_6,N_1906);
nand U2507 (N_2507,N_1678,N_1911);
nor U2508 (N_2508,N_728,N_465);
or U2509 (N_2509,N_1266,N_599);
and U2510 (N_2510,N_1299,N_1004);
or U2511 (N_2511,N_470,N_417);
nand U2512 (N_2512,N_639,N_1801);
nand U2513 (N_2513,N_12,N_1018);
or U2514 (N_2514,N_1582,N_223);
and U2515 (N_2515,N_735,N_1531);
and U2516 (N_2516,N_1969,N_1196);
and U2517 (N_2517,N_696,N_701);
nand U2518 (N_2518,N_338,N_757);
and U2519 (N_2519,N_75,N_129);
nor U2520 (N_2520,N_29,N_589);
and U2521 (N_2521,N_1539,N_1437);
nor U2522 (N_2522,N_1078,N_1943);
and U2523 (N_2523,N_1583,N_1892);
nand U2524 (N_2524,N_1186,N_1913);
and U2525 (N_2525,N_202,N_1604);
or U2526 (N_2526,N_1442,N_774);
and U2527 (N_2527,N_191,N_1229);
nor U2528 (N_2528,N_1970,N_820);
or U2529 (N_2529,N_2,N_1680);
nor U2530 (N_2530,N_1110,N_118);
nand U2531 (N_2531,N_1262,N_1715);
nand U2532 (N_2532,N_712,N_537);
and U2533 (N_2533,N_879,N_577);
and U2534 (N_2534,N_909,N_625);
nor U2535 (N_2535,N_653,N_73);
nor U2536 (N_2536,N_669,N_50);
xor U2537 (N_2537,N_1722,N_270);
nand U2538 (N_2538,N_1523,N_1770);
or U2539 (N_2539,N_1711,N_260);
nand U2540 (N_2540,N_1559,N_968);
nor U2541 (N_2541,N_1115,N_1725);
nand U2542 (N_2542,N_1132,N_1185);
nor U2543 (N_2543,N_1171,N_412);
nor U2544 (N_2544,N_1522,N_571);
and U2545 (N_2545,N_316,N_1482);
and U2546 (N_2546,N_1871,N_1123);
nor U2547 (N_2547,N_113,N_1643);
nand U2548 (N_2548,N_796,N_519);
nor U2549 (N_2549,N_1812,N_1264);
nand U2550 (N_2550,N_525,N_1623);
nor U2551 (N_2551,N_1205,N_1487);
nor U2552 (N_2552,N_920,N_1542);
nand U2553 (N_2553,N_1832,N_1502);
and U2554 (N_2554,N_1055,N_754);
nand U2555 (N_2555,N_1563,N_1737);
and U2556 (N_2556,N_997,N_1325);
or U2557 (N_2557,N_1027,N_549);
nor U2558 (N_2558,N_133,N_1744);
nor U2559 (N_2559,N_274,N_1580);
and U2560 (N_2560,N_1830,N_253);
nand U2561 (N_2561,N_1887,N_674);
nor U2562 (N_2562,N_481,N_387);
nor U2563 (N_2563,N_1854,N_1357);
nor U2564 (N_2564,N_1881,N_341);
and U2565 (N_2565,N_1760,N_489);
nand U2566 (N_2566,N_401,N_509);
xor U2567 (N_2567,N_389,N_1822);
and U2568 (N_2568,N_1243,N_1147);
nand U2569 (N_2569,N_1374,N_1189);
and U2570 (N_2570,N_821,N_1694);
nor U2571 (N_2571,N_917,N_131);
nor U2572 (N_2572,N_953,N_1025);
nand U2573 (N_2573,N_1135,N_1927);
and U2574 (N_2574,N_1104,N_1331);
nand U2575 (N_2575,N_1069,N_363);
and U2576 (N_2576,N_1790,N_1561);
nand U2577 (N_2577,N_825,N_34);
nand U2578 (N_2578,N_175,N_1174);
and U2579 (N_2579,N_1216,N_569);
and U2580 (N_2580,N_299,N_1647);
or U2581 (N_2581,N_1207,N_125);
or U2582 (N_2582,N_326,N_719);
or U2583 (N_2583,N_1864,N_668);
nor U2584 (N_2584,N_618,N_1996);
and U2585 (N_2585,N_814,N_452);
nand U2586 (N_2586,N_976,N_1898);
or U2587 (N_2587,N_1415,N_1075);
nand U2588 (N_2588,N_676,N_172);
and U2589 (N_2589,N_352,N_875);
nor U2590 (N_2590,N_1428,N_1999);
and U2591 (N_2591,N_1752,N_688);
nor U2592 (N_2592,N_1584,N_143);
or U2593 (N_2593,N_1535,N_802);
and U2594 (N_2594,N_682,N_1785);
xnor U2595 (N_2595,N_1717,N_415);
nor U2596 (N_2596,N_1485,N_290);
nand U2597 (N_2597,N_1624,N_822);
nand U2598 (N_2598,N_957,N_27);
and U2599 (N_2599,N_1336,N_314);
nor U2600 (N_2600,N_502,N_1215);
or U2601 (N_2601,N_206,N_1891);
and U2602 (N_2602,N_1306,N_68);
nand U2603 (N_2603,N_1012,N_1844);
nand U2604 (N_2604,N_1598,N_295);
and U2605 (N_2605,N_1828,N_1779);
nand U2606 (N_2606,N_952,N_214);
and U2607 (N_2607,N_1937,N_711);
and U2608 (N_2608,N_399,N_1031);
and U2609 (N_2609,N_239,N_193);
nor U2610 (N_2610,N_1649,N_148);
nor U2611 (N_2611,N_1757,N_11);
or U2612 (N_2612,N_1042,N_207);
nor U2613 (N_2613,N_526,N_657);
and U2614 (N_2614,N_501,N_492);
and U2615 (N_2615,N_1307,N_761);
nor U2616 (N_2616,N_276,N_663);
or U2617 (N_2617,N_1382,N_677);
or U2618 (N_2618,N_151,N_1638);
or U2619 (N_2619,N_1252,N_182);
nor U2620 (N_2620,N_856,N_1101);
and U2621 (N_2621,N_679,N_301);
and U2622 (N_2622,N_1577,N_1641);
and U2623 (N_2623,N_762,N_1587);
nor U2624 (N_2624,N_286,N_1219);
nor U2625 (N_2625,N_1350,N_750);
or U2626 (N_2626,N_1380,N_59);
or U2627 (N_2627,N_978,N_1908);
nand U2628 (N_2628,N_664,N_201);
and U2629 (N_2629,N_714,N_292);
nand U2630 (N_2630,N_853,N_159);
or U2631 (N_2631,N_107,N_1712);
nand U2632 (N_2632,N_799,N_633);
or U2633 (N_2633,N_811,N_422);
nand U2634 (N_2634,N_1414,N_1359);
and U2635 (N_2635,N_271,N_1595);
nor U2636 (N_2636,N_105,N_1225);
nand U2637 (N_2637,N_393,N_654);
and U2638 (N_2638,N_1538,N_89);
nand U2639 (N_2639,N_1268,N_891);
and U2640 (N_2640,N_1588,N_972);
nand U2641 (N_2641,N_1692,N_1860);
nor U2642 (N_2642,N_1366,N_644);
or U2643 (N_2643,N_1593,N_1187);
and U2644 (N_2644,N_1895,N_1273);
and U2645 (N_2645,N_1837,N_703);
or U2646 (N_2646,N_954,N_1997);
or U2647 (N_2647,N_1697,N_362);
or U2648 (N_2648,N_602,N_1272);
nand U2649 (N_2649,N_1418,N_1617);
and U2650 (N_2650,N_706,N_1311);
nor U2651 (N_2651,N_281,N_1612);
nor U2652 (N_2652,N_963,N_927);
or U2653 (N_2653,N_8,N_1619);
nand U2654 (N_2654,N_1778,N_649);
and U2655 (N_2655,N_1202,N_213);
and U2656 (N_2656,N_655,N_1605);
or U2657 (N_2657,N_437,N_791);
or U2658 (N_2658,N_62,N_1863);
nand U2659 (N_2659,N_545,N_436);
nor U2660 (N_2660,N_1509,N_1322);
nor U2661 (N_2661,N_516,N_1654);
or U2662 (N_2662,N_1435,N_1935);
xor U2663 (N_2663,N_904,N_818);
nor U2664 (N_2664,N_1250,N_1901);
and U2665 (N_2665,N_1666,N_1319);
or U2666 (N_2666,N_1553,N_1708);
and U2667 (N_2667,N_638,N_995);
nor U2668 (N_2668,N_1095,N_467);
nand U2669 (N_2669,N_1083,N_346);
and U2670 (N_2670,N_84,N_81);
nand U2671 (N_2671,N_809,N_93);
and U2672 (N_2672,N_642,N_1932);
nand U2673 (N_2673,N_1240,N_1669);
and U2674 (N_2674,N_111,N_139);
nand U2675 (N_2675,N_357,N_611);
or U2676 (N_2676,N_836,N_1008);
nor U2677 (N_2677,N_1545,N_1719);
nand U2678 (N_2678,N_1758,N_55);
and U2679 (N_2679,N_1682,N_1439);
nand U2680 (N_2680,N_546,N_1601);
nand U2681 (N_2681,N_544,N_1687);
or U2682 (N_2682,N_1975,N_14);
nand U2683 (N_2683,N_1994,N_462);
and U2684 (N_2684,N_632,N_1529);
nor U2685 (N_2685,N_860,N_1401);
nand U2686 (N_2686,N_973,N_1741);
and U2687 (N_2687,N_1360,N_381);
and U2688 (N_2688,N_420,N_263);
and U2689 (N_2689,N_1919,N_1370);
nor U2690 (N_2690,N_590,N_527);
nor U2691 (N_2691,N_1484,N_1578);
nor U2692 (N_2692,N_500,N_1879);
nand U2693 (N_2693,N_759,N_937);
or U2694 (N_2694,N_1859,N_1124);
or U2695 (N_2695,N_1334,N_1271);
nand U2696 (N_2696,N_697,N_121);
or U2697 (N_2697,N_983,N_1978);
nor U2698 (N_2698,N_951,N_1333);
xnor U2699 (N_2699,N_1479,N_1572);
or U2700 (N_2700,N_1621,N_1379);
nand U2701 (N_2701,N_1137,N_916);
or U2702 (N_2702,N_1221,N_168);
nand U2703 (N_2703,N_560,N_1289);
and U2704 (N_2704,N_466,N_261);
nand U2705 (N_2705,N_1064,N_681);
or U2706 (N_2706,N_581,N_1628);
or U2707 (N_2707,N_1846,N_1820);
or U2708 (N_2708,N_1924,N_1814);
nor U2709 (N_2709,N_1549,N_1568);
and U2710 (N_2710,N_1082,N_1363);
nand U2711 (N_2711,N_1524,N_1308);
or U2712 (N_2712,N_845,N_1748);
or U2713 (N_2713,N_1960,N_167);
and U2714 (N_2714,N_534,N_977);
and U2715 (N_2715,N_942,N_1);
nor U2716 (N_2716,N_40,N_683);
or U2717 (N_2717,N_410,N_1419);
or U2718 (N_2718,N_380,N_128);
and U2719 (N_2719,N_704,N_709);
or U2720 (N_2720,N_988,N_794);
nand U2721 (N_2721,N_702,N_1169);
nand U2722 (N_2722,N_865,N_100);
nand U2723 (N_2723,N_1564,N_1558);
and U2724 (N_2724,N_1376,N_334);
nor U2725 (N_2725,N_715,N_960);
or U2726 (N_2726,N_1965,N_1766);
nor U2727 (N_2727,N_1294,N_1501);
nand U2728 (N_2728,N_1448,N_1681);
nor U2729 (N_2729,N_1570,N_1067);
nor U2730 (N_2730,N_195,N_543);
and U2731 (N_2731,N_832,N_1504);
nor U2732 (N_2732,N_203,N_166);
nand U2733 (N_2733,N_908,N_278);
nand U2734 (N_2734,N_354,N_1431);
nor U2735 (N_2735,N_1119,N_834);
nand U2736 (N_2736,N_518,N_1421);
and U2737 (N_2737,N_1298,N_773);
nor U2738 (N_2738,N_1283,N_1917);
and U2739 (N_2739,N_928,N_695);
and U2740 (N_2740,N_598,N_1749);
nor U2741 (N_2741,N_484,N_1610);
and U2742 (N_2742,N_1043,N_510);
and U2743 (N_2743,N_1353,N_1029);
nand U2744 (N_2744,N_1096,N_483);
nand U2745 (N_2745,N_455,N_15);
nor U2746 (N_2746,N_375,N_1825);
or U2747 (N_2747,N_1532,N_847);
or U2748 (N_2748,N_1614,N_596);
nand U2749 (N_2749,N_370,N_358);
nor U2750 (N_2750,N_553,N_747);
nor U2751 (N_2751,N_491,N_1810);
nand U2752 (N_2752,N_1915,N_1803);
and U2753 (N_2753,N_1061,N_1622);
nor U2754 (N_2754,N_1700,N_1797);
nand U2755 (N_2755,N_1000,N_1424);
nand U2756 (N_2756,N_619,N_1590);
nand U2757 (N_2757,N_623,N_313);
nand U2758 (N_2758,N_298,N_1329);
nor U2759 (N_2759,N_946,N_736);
nand U2760 (N_2760,N_921,N_1543);
nor U2761 (N_2761,N_1388,N_1300);
nand U2762 (N_2762,N_529,N_1608);
nor U2763 (N_2763,N_378,N_227);
or U2764 (N_2764,N_1597,N_1716);
nor U2765 (N_2765,N_1936,N_1224);
nor U2766 (N_2766,N_1904,N_47);
nor U2767 (N_2767,N_1704,N_781);
nand U2768 (N_2768,N_1473,N_752);
nor U2769 (N_2769,N_1242,N_185);
nor U2770 (N_2770,N_1916,N_137);
and U2771 (N_2771,N_1714,N_88);
nor U2772 (N_2772,N_215,N_1394);
and U2773 (N_2773,N_204,N_1073);
or U2774 (N_2774,N_1510,N_438);
or U2775 (N_2775,N_659,N_1160);
nor U2776 (N_2776,N_1180,N_102);
nor U2777 (N_2777,N_1720,N_1849);
or U2778 (N_2778,N_464,N_887);
or U2779 (N_2779,N_514,N_1087);
or U2780 (N_2780,N_1798,N_950);
and U2781 (N_2781,N_305,N_208);
xnor U2782 (N_2782,N_1973,N_221);
nand U2783 (N_2783,N_493,N_790);
nor U2784 (N_2784,N_1690,N_1862);
or U2785 (N_2785,N_539,N_1332);
nor U2786 (N_2786,N_1742,N_1912);
nor U2787 (N_2787,N_828,N_447);
and U2788 (N_2788,N_1150,N_1791);
nand U2789 (N_2789,N_1469,N_1495);
nor U2790 (N_2790,N_366,N_1313);
nand U2791 (N_2791,N_469,N_1106);
or U2792 (N_2792,N_583,N_1277);
or U2793 (N_2793,N_1204,N_496);
and U2794 (N_2794,N_1850,N_870);
or U2795 (N_2795,N_620,N_548);
and U2796 (N_2796,N_1465,N_1002);
or U2797 (N_2797,N_1406,N_187);
or U2798 (N_2798,N_332,N_604);
or U2799 (N_2799,N_1557,N_1909);
nor U2800 (N_2800,N_454,N_43);
and U2801 (N_2801,N_1995,N_1166);
nor U2802 (N_2802,N_1747,N_1425);
and U2803 (N_2803,N_1910,N_1900);
nor U2804 (N_2804,N_1152,N_1773);
nor U2805 (N_2805,N_558,N_345);
and U2806 (N_2806,N_384,N_1249);
or U2807 (N_2807,N_78,N_793);
or U2808 (N_2808,N_1383,N_1490);
or U2809 (N_2809,N_117,N_554);
nor U2810 (N_2810,N_531,N_1149);
and U2811 (N_2811,N_1190,N_666);
nand U2812 (N_2812,N_585,N_373);
nand U2813 (N_2813,N_803,N_160);
and U2814 (N_2814,N_136,N_400);
nor U2815 (N_2815,N_1211,N_1358);
or U2816 (N_2816,N_476,N_975);
nand U2817 (N_2817,N_1972,N_284);
or U2818 (N_2818,N_1011,N_108);
or U2819 (N_2819,N_1337,N_1105);
or U2820 (N_2820,N_87,N_1613);
or U2821 (N_2821,N_1921,N_179);
nor U2822 (N_2822,N_365,N_789);
nor U2823 (N_2823,N_1560,N_1280);
nor U2824 (N_2824,N_785,N_1127);
nand U2825 (N_2825,N_680,N_1223);
or U2826 (N_2826,N_826,N_217);
nand U2827 (N_2827,N_843,N_1684);
nand U2828 (N_2828,N_279,N_423);
and U2829 (N_2829,N_1579,N_622);
nor U2830 (N_2830,N_1041,N_24);
nor U2831 (N_2831,N_1840,N_686);
and U2832 (N_2832,N_163,N_122);
and U2833 (N_2833,N_713,N_795);
or U2834 (N_2834,N_1020,N_907);
nor U2835 (N_2835,N_640,N_1751);
nor U2836 (N_2836,N_1387,N_1324);
nor U2837 (N_2837,N_1665,N_1724);
nor U2838 (N_2838,N_1017,N_318);
and U2839 (N_2839,N_1429,N_331);
or U2840 (N_2840,N_1456,N_725);
nor U2841 (N_2841,N_1931,N_249);
and U2842 (N_2842,N_1481,N_1567);
nand U2843 (N_2843,N_1070,N_1914);
nor U2844 (N_2844,N_434,N_474);
nand U2845 (N_2845,N_730,N_824);
and U2846 (N_2846,N_282,N_291);
or U2847 (N_2847,N_565,N_1471);
or U2848 (N_2848,N_1060,N_771);
and U2849 (N_2849,N_1346,N_1503);
and U2850 (N_2850,N_1114,N_1506);
or U2851 (N_2851,N_933,N_1865);
or U2852 (N_2852,N_408,N_1565);
or U2853 (N_2853,N_1826,N_1537);
nor U2854 (N_2854,N_1513,N_1515);
or U2855 (N_2855,N_1821,N_80);
or U2856 (N_2856,N_1168,N_1364);
nand U2857 (N_2857,N_634,N_189);
nand U2858 (N_2858,N_176,N_1698);
or U2859 (N_2859,N_1831,N_658);
and U2860 (N_2860,N_1100,N_991);
and U2861 (N_2861,N_359,N_1237);
nand U2862 (N_2862,N_1234,N_336);
or U2863 (N_2863,N_1653,N_222);
and U2864 (N_2864,N_1220,N_1427);
or U2865 (N_2865,N_1138,N_1226);
nand U2866 (N_2866,N_1592,N_958);
or U2867 (N_2867,N_85,N_473);
or U2868 (N_2868,N_1089,N_967);
or U2869 (N_2869,N_1589,N_1440);
and U2870 (N_2870,N_1248,N_1726);
nand U2871 (N_2871,N_1706,N_70);
nand U2872 (N_2872,N_1762,N_1673);
nor U2873 (N_2873,N_533,N_990);
and U2874 (N_2874,N_1131,N_591);
and U2875 (N_2875,N_727,N_348);
nand U2876 (N_2876,N_1167,N_1328);
nor U2877 (N_2877,N_1795,N_1312);
nand U2878 (N_2878,N_177,N_183);
nand U2879 (N_2879,N_823,N_475);
or U2880 (N_2880,N_109,N_157);
nand U2881 (N_2881,N_1815,N_538);
nand U2882 (N_2882,N_1942,N_283);
nor U2883 (N_2883,N_1576,N_302);
nor U2884 (N_2884,N_1472,N_628);
nor U2885 (N_2885,N_1371,N_1039);
or U2886 (N_2886,N_869,N_1633);
nand U2887 (N_2887,N_981,N_152);
or U2888 (N_2888,N_1165,N_1616);
nand U2889 (N_2889,N_1980,N_333);
nor U2890 (N_2890,N_17,N_1870);
nor U2891 (N_2891,N_1344,N_1256);
and U2892 (N_2892,N_450,N_390);
nor U2893 (N_2893,N_1948,N_1458);
nand U2894 (N_2894,N_268,N_1982);
nand U2895 (N_2895,N_307,N_1395);
nor U2896 (N_2896,N_1195,N_1735);
nor U2897 (N_2897,N_1489,N_1944);
nand U2898 (N_2898,N_612,N_557);
nor U2899 (N_2899,N_321,N_1907);
or U2900 (N_2900,N_898,N_1445);
nand U2901 (N_2901,N_396,N_1103);
or U2902 (N_2902,N_1016,N_42);
or U2903 (N_2903,N_374,N_1086);
nand U2904 (N_2904,N_1035,N_760);
nor U2905 (N_2905,N_468,N_1128);
and U2906 (N_2906,N_1321,N_340);
nand U2907 (N_2907,N_786,N_1253);
or U2908 (N_2908,N_1498,N_170);
xor U2909 (N_2909,N_1890,N_1241);
or U2910 (N_2910,N_1642,N_19);
or U2911 (N_2911,N_1108,N_1244);
nand U2912 (N_2912,N_914,N_609);
nor U2913 (N_2913,N_777,N_1548);
nor U2914 (N_2914,N_751,N_1663);
nor U2915 (N_2915,N_1369,N_165);
and U2916 (N_2916,N_1233,N_1550);
and U2917 (N_2917,N_911,N_280);
nand U2918 (N_2918,N_645,N_941);
nor U2919 (N_2919,N_265,N_1209);
nand U2920 (N_2920,N_550,N_1626);
nor U2921 (N_2921,N_1046,N_1274);
or U2922 (N_2922,N_101,N_1400);
nor U2923 (N_2923,N_1303,N_1362);
nand U2924 (N_2924,N_974,N_896);
and U2925 (N_2925,N_404,N_1446);
nor U2926 (N_2926,N_1824,N_523);
or U2927 (N_2927,N_277,N_1675);
or U2928 (N_2928,N_517,N_1194);
nor U2929 (N_2929,N_446,N_630);
or U2930 (N_2930,N_606,N_409);
or U2931 (N_2931,N_1044,N_1816);
and U2932 (N_2932,N_1852,N_817);
nand U2933 (N_2933,N_488,N_788);
nor U2934 (N_2934,N_395,N_1270);
and U2935 (N_2935,N_1591,N_595);
nor U2936 (N_2936,N_257,N_30);
nand U2937 (N_2937,N_1631,N_116);
or U2938 (N_2938,N_1133,N_1170);
nand U2939 (N_2939,N_98,N_240);
or U2940 (N_2940,N_1958,N_1163);
nor U2941 (N_2941,N_259,N_288);
nand U2942 (N_2942,N_733,N_1056);
nand U2943 (N_2943,N_1703,N_1805);
or U2944 (N_2944,N_1218,N_969);
nand U2945 (N_2945,N_849,N_955);
or U2946 (N_2946,N_840,N_594);
nand U2947 (N_2947,N_597,N_765);
and U2948 (N_2948,N_161,N_1867);
nand U2949 (N_2949,N_144,N_884);
and U2950 (N_2950,N_1723,N_1962);
and U2951 (N_2951,N_672,N_123);
nand U2952 (N_2952,N_906,N_555);
nand U2953 (N_2953,N_104,N_441);
and U2954 (N_2954,N_1759,N_349);
nand U2955 (N_2955,N_613,N_1159);
or U2956 (N_2956,N_1651,N_392);
nor U2957 (N_2957,N_1516,N_1459);
and U2958 (N_2958,N_1677,N_805);
or U2959 (N_2959,N_993,N_900);
and U2960 (N_2960,N_1407,N_335);
nand U2961 (N_2961,N_1882,N_376);
nand U2962 (N_2962,N_72,N_1074);
and U2963 (N_2963,N_1964,N_149);
nor U2964 (N_2964,N_940,N_1403);
and U2965 (N_2965,N_1721,N_1483);
nor U2966 (N_2966,N_1140,N_1777);
nor U2967 (N_2967,N_485,N_1381);
nand U2968 (N_2968,N_1005,N_1674);
or U2969 (N_2969,N_1534,N_1141);
and U2970 (N_2970,N_660,N_1065);
and U2971 (N_2971,N_753,N_1467);
nor U2972 (N_2972,N_966,N_1326);
nand U2973 (N_2973,N_1175,N_1664);
nor U2974 (N_2974,N_10,N_1352);
nor U2975 (N_2975,N_1013,N_5);
nand U2976 (N_2976,N_756,N_1480);
nor U2977 (N_2977,N_1217,N_255);
or U2978 (N_2978,N_296,N_1126);
nand U2979 (N_2979,N_1342,N_1285);
nand U2980 (N_2980,N_508,N_198);
or U2981 (N_2981,N_54,N_699);
nor U2982 (N_2982,N_1496,N_1873);
and U2983 (N_2983,N_1411,N_626);
or U2984 (N_2984,N_678,N_1071);
nor U2985 (N_2985,N_1670,N_1373);
nand U2986 (N_2986,N_962,N_74);
or U2987 (N_2987,N_801,N_1629);
nand U2988 (N_2988,N_987,N_135);
nand U2989 (N_2989,N_1738,N_992);
nand U2990 (N_2990,N_1001,N_1486);
nor U2991 (N_2991,N_1520,N_1853);
nand U2992 (N_2992,N_982,N_3);
nor U2993 (N_2993,N_1176,N_1153);
xor U2994 (N_2994,N_1540,N_490);
nor U2995 (N_2995,N_1301,N_1228);
and U2996 (N_2996,N_1644,N_576);
or U2997 (N_2997,N_71,N_1512);
or U2998 (N_2998,N_1571,N_935);
nand U2999 (N_2999,N_1447,N_1998);
or U3000 (N_3000,N_1073,N_361);
nand U3001 (N_3001,N_973,N_1514);
xnor U3002 (N_3002,N_557,N_1747);
or U3003 (N_3003,N_1174,N_944);
nor U3004 (N_3004,N_205,N_569);
and U3005 (N_3005,N_529,N_477);
or U3006 (N_3006,N_884,N_1983);
and U3007 (N_3007,N_508,N_421);
nor U3008 (N_3008,N_1507,N_1255);
and U3009 (N_3009,N_1232,N_724);
xor U3010 (N_3010,N_1108,N_115);
and U3011 (N_3011,N_1069,N_1618);
nor U3012 (N_3012,N_996,N_7);
and U3013 (N_3013,N_1581,N_516);
nor U3014 (N_3014,N_406,N_1000);
or U3015 (N_3015,N_1080,N_1750);
and U3016 (N_3016,N_668,N_295);
nand U3017 (N_3017,N_1939,N_926);
nand U3018 (N_3018,N_533,N_387);
nand U3019 (N_3019,N_1476,N_1931);
and U3020 (N_3020,N_763,N_477);
nor U3021 (N_3021,N_316,N_1732);
and U3022 (N_3022,N_507,N_277);
nand U3023 (N_3023,N_1192,N_217);
or U3024 (N_3024,N_380,N_1446);
or U3025 (N_3025,N_77,N_742);
nand U3026 (N_3026,N_1551,N_271);
nor U3027 (N_3027,N_878,N_1873);
nor U3028 (N_3028,N_26,N_1300);
or U3029 (N_3029,N_903,N_627);
and U3030 (N_3030,N_1496,N_1405);
and U3031 (N_3031,N_512,N_1139);
nor U3032 (N_3032,N_452,N_1626);
or U3033 (N_3033,N_1952,N_104);
nand U3034 (N_3034,N_740,N_312);
and U3035 (N_3035,N_839,N_973);
and U3036 (N_3036,N_702,N_898);
nor U3037 (N_3037,N_525,N_1312);
nor U3038 (N_3038,N_1880,N_576);
nor U3039 (N_3039,N_939,N_866);
and U3040 (N_3040,N_393,N_1529);
nor U3041 (N_3041,N_1156,N_885);
and U3042 (N_3042,N_41,N_1495);
or U3043 (N_3043,N_687,N_568);
and U3044 (N_3044,N_183,N_1341);
nand U3045 (N_3045,N_1939,N_308);
nor U3046 (N_3046,N_692,N_9);
xnor U3047 (N_3047,N_972,N_342);
nor U3048 (N_3048,N_1536,N_532);
nand U3049 (N_3049,N_76,N_121);
and U3050 (N_3050,N_557,N_230);
or U3051 (N_3051,N_697,N_1238);
or U3052 (N_3052,N_1066,N_648);
or U3053 (N_3053,N_1160,N_1613);
nand U3054 (N_3054,N_435,N_371);
or U3055 (N_3055,N_730,N_13);
nand U3056 (N_3056,N_1589,N_466);
nand U3057 (N_3057,N_761,N_385);
nand U3058 (N_3058,N_925,N_39);
nor U3059 (N_3059,N_73,N_1198);
or U3060 (N_3060,N_1300,N_542);
and U3061 (N_3061,N_558,N_726);
nor U3062 (N_3062,N_1723,N_955);
or U3063 (N_3063,N_1640,N_930);
and U3064 (N_3064,N_1368,N_1567);
and U3065 (N_3065,N_1151,N_1407);
nor U3066 (N_3066,N_416,N_1543);
nand U3067 (N_3067,N_1690,N_1117);
and U3068 (N_3068,N_1424,N_1072);
nor U3069 (N_3069,N_1679,N_1817);
nor U3070 (N_3070,N_743,N_1876);
and U3071 (N_3071,N_1348,N_1788);
or U3072 (N_3072,N_1203,N_1484);
nor U3073 (N_3073,N_660,N_1823);
and U3074 (N_3074,N_498,N_1055);
nand U3075 (N_3075,N_1542,N_1610);
and U3076 (N_3076,N_1266,N_1840);
nor U3077 (N_3077,N_610,N_1617);
and U3078 (N_3078,N_1154,N_222);
nand U3079 (N_3079,N_1213,N_977);
and U3080 (N_3080,N_462,N_1530);
or U3081 (N_3081,N_697,N_775);
nor U3082 (N_3082,N_30,N_248);
nand U3083 (N_3083,N_1639,N_1760);
nor U3084 (N_3084,N_1651,N_1974);
nor U3085 (N_3085,N_1609,N_286);
nor U3086 (N_3086,N_1587,N_274);
nand U3087 (N_3087,N_1663,N_1703);
or U3088 (N_3088,N_595,N_786);
nor U3089 (N_3089,N_1709,N_1053);
and U3090 (N_3090,N_1937,N_844);
or U3091 (N_3091,N_222,N_1943);
and U3092 (N_3092,N_1463,N_202);
nor U3093 (N_3093,N_957,N_1716);
nor U3094 (N_3094,N_532,N_1820);
xnor U3095 (N_3095,N_284,N_274);
and U3096 (N_3096,N_404,N_881);
or U3097 (N_3097,N_1005,N_1599);
or U3098 (N_3098,N_162,N_1945);
nand U3099 (N_3099,N_727,N_116);
nor U3100 (N_3100,N_39,N_873);
or U3101 (N_3101,N_1463,N_760);
and U3102 (N_3102,N_820,N_1528);
nor U3103 (N_3103,N_718,N_129);
nor U3104 (N_3104,N_58,N_471);
nor U3105 (N_3105,N_798,N_111);
nor U3106 (N_3106,N_780,N_755);
or U3107 (N_3107,N_88,N_1978);
and U3108 (N_3108,N_1824,N_1041);
and U3109 (N_3109,N_1888,N_1389);
and U3110 (N_3110,N_434,N_1614);
nor U3111 (N_3111,N_1369,N_1475);
nor U3112 (N_3112,N_168,N_1241);
nand U3113 (N_3113,N_1103,N_1174);
nor U3114 (N_3114,N_672,N_743);
xor U3115 (N_3115,N_425,N_912);
or U3116 (N_3116,N_838,N_1254);
or U3117 (N_3117,N_1407,N_878);
and U3118 (N_3118,N_1385,N_505);
nor U3119 (N_3119,N_101,N_785);
nand U3120 (N_3120,N_1164,N_730);
or U3121 (N_3121,N_86,N_845);
nor U3122 (N_3122,N_1532,N_1735);
nand U3123 (N_3123,N_1960,N_1936);
nand U3124 (N_3124,N_1461,N_1739);
nor U3125 (N_3125,N_1979,N_1237);
nand U3126 (N_3126,N_369,N_743);
or U3127 (N_3127,N_584,N_1506);
nand U3128 (N_3128,N_217,N_173);
nor U3129 (N_3129,N_400,N_363);
nor U3130 (N_3130,N_1674,N_1438);
nand U3131 (N_3131,N_1478,N_643);
nor U3132 (N_3132,N_1807,N_685);
nand U3133 (N_3133,N_917,N_1934);
and U3134 (N_3134,N_86,N_1866);
nand U3135 (N_3135,N_1709,N_223);
nand U3136 (N_3136,N_427,N_533);
nand U3137 (N_3137,N_1097,N_859);
or U3138 (N_3138,N_724,N_864);
nor U3139 (N_3139,N_540,N_248);
nand U3140 (N_3140,N_202,N_1032);
and U3141 (N_3141,N_767,N_975);
nor U3142 (N_3142,N_238,N_156);
nor U3143 (N_3143,N_76,N_618);
or U3144 (N_3144,N_827,N_1681);
and U3145 (N_3145,N_201,N_786);
nand U3146 (N_3146,N_1375,N_962);
or U3147 (N_3147,N_257,N_949);
or U3148 (N_3148,N_1033,N_443);
and U3149 (N_3149,N_647,N_1348);
and U3150 (N_3150,N_962,N_1986);
or U3151 (N_3151,N_343,N_1637);
nor U3152 (N_3152,N_1235,N_270);
nor U3153 (N_3153,N_859,N_761);
nand U3154 (N_3154,N_231,N_1082);
nor U3155 (N_3155,N_1937,N_556);
nand U3156 (N_3156,N_896,N_436);
nor U3157 (N_3157,N_682,N_497);
nand U3158 (N_3158,N_316,N_1279);
and U3159 (N_3159,N_1579,N_494);
nand U3160 (N_3160,N_636,N_920);
or U3161 (N_3161,N_1170,N_1222);
nor U3162 (N_3162,N_996,N_576);
or U3163 (N_3163,N_1649,N_1025);
nand U3164 (N_3164,N_1598,N_341);
or U3165 (N_3165,N_581,N_328);
and U3166 (N_3166,N_1983,N_1564);
xnor U3167 (N_3167,N_1014,N_1956);
and U3168 (N_3168,N_1529,N_1450);
nand U3169 (N_3169,N_591,N_1444);
or U3170 (N_3170,N_1301,N_1032);
nor U3171 (N_3171,N_577,N_415);
and U3172 (N_3172,N_1524,N_1445);
nand U3173 (N_3173,N_1646,N_194);
nand U3174 (N_3174,N_1699,N_662);
nand U3175 (N_3175,N_323,N_1446);
and U3176 (N_3176,N_718,N_98);
nor U3177 (N_3177,N_1084,N_1058);
or U3178 (N_3178,N_1920,N_1355);
or U3179 (N_3179,N_984,N_1156);
nor U3180 (N_3180,N_561,N_496);
and U3181 (N_3181,N_141,N_479);
nand U3182 (N_3182,N_669,N_965);
or U3183 (N_3183,N_1489,N_1542);
nor U3184 (N_3184,N_1745,N_439);
nand U3185 (N_3185,N_1432,N_642);
or U3186 (N_3186,N_1394,N_561);
nor U3187 (N_3187,N_497,N_1063);
or U3188 (N_3188,N_70,N_756);
nor U3189 (N_3189,N_1722,N_1388);
and U3190 (N_3190,N_190,N_1237);
and U3191 (N_3191,N_1610,N_1637);
and U3192 (N_3192,N_56,N_1031);
and U3193 (N_3193,N_1095,N_1403);
and U3194 (N_3194,N_1197,N_1461);
and U3195 (N_3195,N_1015,N_1403);
nand U3196 (N_3196,N_1624,N_388);
nand U3197 (N_3197,N_89,N_139);
nor U3198 (N_3198,N_1529,N_574);
nand U3199 (N_3199,N_1140,N_1);
or U3200 (N_3200,N_1660,N_1795);
and U3201 (N_3201,N_1737,N_33);
and U3202 (N_3202,N_236,N_616);
nand U3203 (N_3203,N_1787,N_481);
nand U3204 (N_3204,N_49,N_1125);
nor U3205 (N_3205,N_1550,N_213);
or U3206 (N_3206,N_380,N_1856);
or U3207 (N_3207,N_254,N_673);
nor U3208 (N_3208,N_1720,N_1894);
and U3209 (N_3209,N_911,N_340);
or U3210 (N_3210,N_352,N_290);
xnor U3211 (N_3211,N_1335,N_410);
nor U3212 (N_3212,N_608,N_1186);
nand U3213 (N_3213,N_297,N_689);
nor U3214 (N_3214,N_194,N_335);
nor U3215 (N_3215,N_248,N_1649);
nand U3216 (N_3216,N_884,N_940);
nor U3217 (N_3217,N_1192,N_940);
or U3218 (N_3218,N_240,N_530);
or U3219 (N_3219,N_658,N_140);
and U3220 (N_3220,N_557,N_1935);
or U3221 (N_3221,N_1205,N_439);
or U3222 (N_3222,N_1764,N_555);
or U3223 (N_3223,N_1831,N_1595);
or U3224 (N_3224,N_1495,N_1464);
or U3225 (N_3225,N_1869,N_1111);
nor U3226 (N_3226,N_659,N_1133);
and U3227 (N_3227,N_1696,N_577);
and U3228 (N_3228,N_565,N_519);
nand U3229 (N_3229,N_1622,N_881);
and U3230 (N_3230,N_742,N_1317);
nand U3231 (N_3231,N_1907,N_269);
or U3232 (N_3232,N_1327,N_795);
and U3233 (N_3233,N_1295,N_1744);
nand U3234 (N_3234,N_1392,N_352);
and U3235 (N_3235,N_2,N_307);
and U3236 (N_3236,N_630,N_583);
nor U3237 (N_3237,N_231,N_587);
nor U3238 (N_3238,N_1963,N_1816);
or U3239 (N_3239,N_1454,N_781);
nand U3240 (N_3240,N_214,N_1963);
or U3241 (N_3241,N_1461,N_1215);
and U3242 (N_3242,N_221,N_1873);
or U3243 (N_3243,N_1903,N_370);
and U3244 (N_3244,N_256,N_1892);
or U3245 (N_3245,N_1986,N_1224);
and U3246 (N_3246,N_1629,N_953);
nor U3247 (N_3247,N_124,N_1895);
and U3248 (N_3248,N_1150,N_1282);
nor U3249 (N_3249,N_1864,N_375);
or U3250 (N_3250,N_1401,N_764);
and U3251 (N_3251,N_751,N_1853);
or U3252 (N_3252,N_1020,N_1350);
nor U3253 (N_3253,N_316,N_405);
nand U3254 (N_3254,N_1037,N_1865);
and U3255 (N_3255,N_62,N_440);
and U3256 (N_3256,N_52,N_1835);
nor U3257 (N_3257,N_670,N_1287);
nor U3258 (N_3258,N_913,N_1863);
nand U3259 (N_3259,N_376,N_249);
xnor U3260 (N_3260,N_1631,N_455);
nand U3261 (N_3261,N_1662,N_374);
or U3262 (N_3262,N_453,N_86);
nand U3263 (N_3263,N_1368,N_468);
and U3264 (N_3264,N_478,N_1446);
nand U3265 (N_3265,N_383,N_1293);
xor U3266 (N_3266,N_1369,N_299);
nand U3267 (N_3267,N_834,N_1463);
nor U3268 (N_3268,N_1033,N_1071);
or U3269 (N_3269,N_803,N_331);
or U3270 (N_3270,N_17,N_72);
nor U3271 (N_3271,N_856,N_725);
and U3272 (N_3272,N_1488,N_740);
nor U3273 (N_3273,N_1735,N_1525);
and U3274 (N_3274,N_91,N_230);
nand U3275 (N_3275,N_50,N_943);
and U3276 (N_3276,N_1215,N_971);
nor U3277 (N_3277,N_1642,N_381);
nand U3278 (N_3278,N_243,N_1323);
and U3279 (N_3279,N_475,N_1528);
and U3280 (N_3280,N_1264,N_1433);
or U3281 (N_3281,N_1270,N_465);
nor U3282 (N_3282,N_1243,N_492);
or U3283 (N_3283,N_67,N_641);
nand U3284 (N_3284,N_1976,N_1057);
or U3285 (N_3285,N_1411,N_1546);
nand U3286 (N_3286,N_1511,N_25);
nand U3287 (N_3287,N_925,N_933);
and U3288 (N_3288,N_402,N_1914);
nand U3289 (N_3289,N_1,N_1795);
and U3290 (N_3290,N_1025,N_1174);
nand U3291 (N_3291,N_1939,N_1502);
nor U3292 (N_3292,N_1315,N_1564);
or U3293 (N_3293,N_71,N_1602);
xnor U3294 (N_3294,N_229,N_1515);
or U3295 (N_3295,N_722,N_872);
or U3296 (N_3296,N_329,N_481);
xnor U3297 (N_3297,N_1438,N_1581);
and U3298 (N_3298,N_958,N_1544);
nor U3299 (N_3299,N_1934,N_819);
nand U3300 (N_3300,N_1639,N_1751);
or U3301 (N_3301,N_757,N_724);
and U3302 (N_3302,N_852,N_255);
or U3303 (N_3303,N_412,N_374);
or U3304 (N_3304,N_188,N_1582);
nor U3305 (N_3305,N_11,N_609);
or U3306 (N_3306,N_1832,N_1137);
and U3307 (N_3307,N_1938,N_1673);
nor U3308 (N_3308,N_489,N_1334);
nor U3309 (N_3309,N_915,N_934);
nor U3310 (N_3310,N_747,N_163);
and U3311 (N_3311,N_194,N_92);
and U3312 (N_3312,N_835,N_569);
nand U3313 (N_3313,N_397,N_1584);
nor U3314 (N_3314,N_1769,N_296);
nand U3315 (N_3315,N_1542,N_775);
nor U3316 (N_3316,N_1489,N_1217);
or U3317 (N_3317,N_1984,N_1637);
or U3318 (N_3318,N_1662,N_619);
or U3319 (N_3319,N_1236,N_1445);
or U3320 (N_3320,N_1546,N_668);
and U3321 (N_3321,N_1065,N_590);
or U3322 (N_3322,N_98,N_1387);
nand U3323 (N_3323,N_655,N_1584);
nand U3324 (N_3324,N_9,N_321);
and U3325 (N_3325,N_103,N_286);
and U3326 (N_3326,N_847,N_486);
nor U3327 (N_3327,N_452,N_1592);
nand U3328 (N_3328,N_1814,N_240);
or U3329 (N_3329,N_229,N_1365);
and U3330 (N_3330,N_1942,N_1387);
and U3331 (N_3331,N_718,N_1616);
nand U3332 (N_3332,N_1586,N_280);
nor U3333 (N_3333,N_1192,N_283);
nand U3334 (N_3334,N_1629,N_712);
nand U3335 (N_3335,N_1024,N_1152);
nand U3336 (N_3336,N_114,N_1155);
nand U3337 (N_3337,N_949,N_1161);
xnor U3338 (N_3338,N_1078,N_1075);
and U3339 (N_3339,N_609,N_827);
or U3340 (N_3340,N_456,N_1559);
nand U3341 (N_3341,N_270,N_639);
or U3342 (N_3342,N_1812,N_356);
and U3343 (N_3343,N_658,N_1503);
nand U3344 (N_3344,N_1798,N_1150);
or U3345 (N_3345,N_206,N_666);
nand U3346 (N_3346,N_1645,N_886);
and U3347 (N_3347,N_949,N_526);
nand U3348 (N_3348,N_648,N_85);
nor U3349 (N_3349,N_923,N_819);
nor U3350 (N_3350,N_77,N_974);
nand U3351 (N_3351,N_1773,N_1489);
or U3352 (N_3352,N_1501,N_646);
and U3353 (N_3353,N_970,N_1706);
nor U3354 (N_3354,N_1515,N_50);
nand U3355 (N_3355,N_1749,N_1266);
and U3356 (N_3356,N_270,N_618);
nor U3357 (N_3357,N_1138,N_71);
and U3358 (N_3358,N_1256,N_751);
or U3359 (N_3359,N_1550,N_397);
nor U3360 (N_3360,N_1,N_1996);
or U3361 (N_3361,N_1507,N_1477);
and U3362 (N_3362,N_791,N_1632);
nor U3363 (N_3363,N_18,N_774);
or U3364 (N_3364,N_960,N_1480);
nand U3365 (N_3365,N_396,N_1744);
nor U3366 (N_3366,N_1786,N_1682);
or U3367 (N_3367,N_894,N_1512);
or U3368 (N_3368,N_1485,N_448);
and U3369 (N_3369,N_665,N_765);
nand U3370 (N_3370,N_1944,N_864);
nor U3371 (N_3371,N_1932,N_345);
nand U3372 (N_3372,N_1797,N_1101);
or U3373 (N_3373,N_778,N_827);
nor U3374 (N_3374,N_914,N_1232);
nor U3375 (N_3375,N_365,N_1127);
and U3376 (N_3376,N_1719,N_163);
nor U3377 (N_3377,N_1027,N_719);
nor U3378 (N_3378,N_174,N_509);
nand U3379 (N_3379,N_359,N_1650);
nor U3380 (N_3380,N_1685,N_1802);
or U3381 (N_3381,N_1987,N_1515);
or U3382 (N_3382,N_1325,N_387);
nor U3383 (N_3383,N_1544,N_1499);
nand U3384 (N_3384,N_531,N_1200);
and U3385 (N_3385,N_682,N_258);
and U3386 (N_3386,N_1470,N_1065);
nor U3387 (N_3387,N_384,N_1973);
or U3388 (N_3388,N_1134,N_1881);
or U3389 (N_3389,N_453,N_748);
nand U3390 (N_3390,N_347,N_4);
nor U3391 (N_3391,N_344,N_1601);
nor U3392 (N_3392,N_1083,N_98);
nor U3393 (N_3393,N_603,N_1241);
nand U3394 (N_3394,N_1741,N_890);
nor U3395 (N_3395,N_888,N_1121);
nand U3396 (N_3396,N_979,N_1758);
or U3397 (N_3397,N_1223,N_59);
nor U3398 (N_3398,N_1010,N_855);
and U3399 (N_3399,N_1777,N_659);
nand U3400 (N_3400,N_1526,N_1501);
or U3401 (N_3401,N_467,N_1090);
nand U3402 (N_3402,N_37,N_36);
nor U3403 (N_3403,N_1351,N_1527);
and U3404 (N_3404,N_1841,N_113);
or U3405 (N_3405,N_1386,N_1063);
and U3406 (N_3406,N_1245,N_1069);
or U3407 (N_3407,N_1889,N_1863);
nand U3408 (N_3408,N_1902,N_317);
nor U3409 (N_3409,N_1383,N_1486);
nand U3410 (N_3410,N_567,N_1579);
or U3411 (N_3411,N_40,N_530);
or U3412 (N_3412,N_1592,N_830);
or U3413 (N_3413,N_1076,N_1352);
and U3414 (N_3414,N_1384,N_1673);
or U3415 (N_3415,N_1028,N_83);
nor U3416 (N_3416,N_96,N_1690);
nor U3417 (N_3417,N_1757,N_420);
nor U3418 (N_3418,N_136,N_599);
xor U3419 (N_3419,N_1777,N_1418);
or U3420 (N_3420,N_612,N_210);
and U3421 (N_3421,N_1992,N_476);
nor U3422 (N_3422,N_1146,N_503);
nor U3423 (N_3423,N_1170,N_1105);
or U3424 (N_3424,N_1709,N_327);
nor U3425 (N_3425,N_551,N_1287);
nor U3426 (N_3426,N_417,N_932);
nor U3427 (N_3427,N_1596,N_726);
or U3428 (N_3428,N_1294,N_974);
or U3429 (N_3429,N_955,N_681);
and U3430 (N_3430,N_116,N_1740);
nand U3431 (N_3431,N_1625,N_321);
nand U3432 (N_3432,N_286,N_257);
and U3433 (N_3433,N_377,N_232);
or U3434 (N_3434,N_158,N_578);
and U3435 (N_3435,N_828,N_575);
nand U3436 (N_3436,N_1086,N_1768);
nor U3437 (N_3437,N_1803,N_280);
nor U3438 (N_3438,N_1732,N_1514);
nor U3439 (N_3439,N_785,N_1910);
nor U3440 (N_3440,N_473,N_303);
and U3441 (N_3441,N_1711,N_1598);
or U3442 (N_3442,N_67,N_1261);
nand U3443 (N_3443,N_964,N_846);
nor U3444 (N_3444,N_241,N_195);
or U3445 (N_3445,N_377,N_952);
nor U3446 (N_3446,N_724,N_1283);
and U3447 (N_3447,N_931,N_1187);
nand U3448 (N_3448,N_1457,N_857);
or U3449 (N_3449,N_592,N_1826);
and U3450 (N_3450,N_902,N_1200);
nand U3451 (N_3451,N_1817,N_1846);
or U3452 (N_3452,N_208,N_466);
or U3453 (N_3453,N_1015,N_257);
or U3454 (N_3454,N_1020,N_1618);
and U3455 (N_3455,N_1729,N_1128);
or U3456 (N_3456,N_517,N_473);
and U3457 (N_3457,N_1779,N_1546);
nor U3458 (N_3458,N_377,N_793);
or U3459 (N_3459,N_1574,N_61);
and U3460 (N_3460,N_592,N_1927);
or U3461 (N_3461,N_1327,N_1114);
nand U3462 (N_3462,N_1367,N_1616);
or U3463 (N_3463,N_979,N_1207);
nand U3464 (N_3464,N_506,N_552);
xor U3465 (N_3465,N_851,N_519);
or U3466 (N_3466,N_979,N_896);
and U3467 (N_3467,N_1309,N_1764);
nand U3468 (N_3468,N_193,N_1476);
and U3469 (N_3469,N_444,N_198);
or U3470 (N_3470,N_735,N_371);
or U3471 (N_3471,N_151,N_179);
nor U3472 (N_3472,N_413,N_1734);
and U3473 (N_3473,N_1297,N_1445);
and U3474 (N_3474,N_98,N_653);
and U3475 (N_3475,N_1351,N_723);
and U3476 (N_3476,N_1744,N_466);
nor U3477 (N_3477,N_338,N_68);
nor U3478 (N_3478,N_1434,N_1269);
or U3479 (N_3479,N_1109,N_1990);
or U3480 (N_3480,N_1227,N_1036);
nand U3481 (N_3481,N_795,N_683);
or U3482 (N_3482,N_912,N_792);
xor U3483 (N_3483,N_518,N_529);
nor U3484 (N_3484,N_226,N_892);
nand U3485 (N_3485,N_889,N_962);
or U3486 (N_3486,N_1593,N_1063);
and U3487 (N_3487,N_1537,N_561);
and U3488 (N_3488,N_105,N_1575);
and U3489 (N_3489,N_18,N_315);
or U3490 (N_3490,N_106,N_1545);
or U3491 (N_3491,N_385,N_1297);
or U3492 (N_3492,N_1657,N_1199);
nand U3493 (N_3493,N_1697,N_361);
nand U3494 (N_3494,N_228,N_1799);
nor U3495 (N_3495,N_1859,N_394);
or U3496 (N_3496,N_1640,N_1567);
and U3497 (N_3497,N_1670,N_1682);
nand U3498 (N_3498,N_143,N_1047);
and U3499 (N_3499,N_321,N_1192);
or U3500 (N_3500,N_10,N_1745);
nand U3501 (N_3501,N_694,N_1141);
or U3502 (N_3502,N_1299,N_1873);
nand U3503 (N_3503,N_1840,N_1128);
or U3504 (N_3504,N_531,N_219);
nand U3505 (N_3505,N_1726,N_140);
nor U3506 (N_3506,N_1948,N_815);
or U3507 (N_3507,N_1076,N_112);
and U3508 (N_3508,N_1576,N_1039);
and U3509 (N_3509,N_141,N_796);
or U3510 (N_3510,N_1385,N_1150);
nand U3511 (N_3511,N_1600,N_1453);
or U3512 (N_3512,N_601,N_1867);
nand U3513 (N_3513,N_924,N_191);
nand U3514 (N_3514,N_1731,N_1044);
nand U3515 (N_3515,N_271,N_1187);
or U3516 (N_3516,N_456,N_110);
and U3517 (N_3517,N_975,N_125);
nand U3518 (N_3518,N_1930,N_101);
and U3519 (N_3519,N_936,N_318);
nand U3520 (N_3520,N_644,N_341);
nor U3521 (N_3521,N_1637,N_801);
nand U3522 (N_3522,N_1370,N_450);
nand U3523 (N_3523,N_379,N_1151);
nand U3524 (N_3524,N_1274,N_1920);
nor U3525 (N_3525,N_1029,N_1034);
nand U3526 (N_3526,N_25,N_669);
or U3527 (N_3527,N_583,N_1269);
nor U3528 (N_3528,N_858,N_1818);
nand U3529 (N_3529,N_309,N_87);
nor U3530 (N_3530,N_857,N_1169);
or U3531 (N_3531,N_525,N_1424);
and U3532 (N_3532,N_1261,N_1663);
nor U3533 (N_3533,N_911,N_661);
nor U3534 (N_3534,N_1950,N_956);
or U3535 (N_3535,N_1710,N_1145);
nor U3536 (N_3536,N_385,N_1838);
nor U3537 (N_3537,N_37,N_1464);
and U3538 (N_3538,N_1689,N_257);
and U3539 (N_3539,N_988,N_1841);
xor U3540 (N_3540,N_812,N_1684);
nand U3541 (N_3541,N_1264,N_80);
nand U3542 (N_3542,N_837,N_842);
nor U3543 (N_3543,N_599,N_580);
and U3544 (N_3544,N_1754,N_483);
nor U3545 (N_3545,N_317,N_1665);
nor U3546 (N_3546,N_254,N_274);
xor U3547 (N_3547,N_617,N_1193);
nor U3548 (N_3548,N_604,N_1401);
nand U3549 (N_3549,N_93,N_1407);
or U3550 (N_3550,N_1959,N_1237);
or U3551 (N_3551,N_612,N_1388);
nor U3552 (N_3552,N_1434,N_1059);
nand U3553 (N_3553,N_1200,N_1640);
nor U3554 (N_3554,N_1055,N_1733);
nand U3555 (N_3555,N_268,N_76);
or U3556 (N_3556,N_1929,N_149);
or U3557 (N_3557,N_855,N_1131);
and U3558 (N_3558,N_1361,N_1577);
or U3559 (N_3559,N_1538,N_1095);
nor U3560 (N_3560,N_1908,N_754);
or U3561 (N_3561,N_1609,N_1930);
nand U3562 (N_3562,N_527,N_447);
nor U3563 (N_3563,N_297,N_452);
or U3564 (N_3564,N_1903,N_767);
and U3565 (N_3565,N_1501,N_609);
nor U3566 (N_3566,N_719,N_1708);
or U3567 (N_3567,N_1675,N_1879);
and U3568 (N_3568,N_1865,N_1576);
or U3569 (N_3569,N_211,N_970);
nor U3570 (N_3570,N_1043,N_966);
nor U3571 (N_3571,N_1208,N_460);
nor U3572 (N_3572,N_1246,N_1283);
or U3573 (N_3573,N_1605,N_1095);
or U3574 (N_3574,N_1629,N_1685);
nor U3575 (N_3575,N_893,N_1207);
nand U3576 (N_3576,N_1090,N_801);
nand U3577 (N_3577,N_465,N_1746);
and U3578 (N_3578,N_831,N_1853);
or U3579 (N_3579,N_1022,N_7);
or U3580 (N_3580,N_1766,N_209);
or U3581 (N_3581,N_1360,N_331);
nor U3582 (N_3582,N_1012,N_1380);
and U3583 (N_3583,N_1624,N_964);
or U3584 (N_3584,N_1549,N_739);
nor U3585 (N_3585,N_1768,N_1353);
nand U3586 (N_3586,N_1613,N_794);
nor U3587 (N_3587,N_1631,N_1869);
or U3588 (N_3588,N_1627,N_761);
and U3589 (N_3589,N_4,N_1133);
nand U3590 (N_3590,N_1848,N_822);
or U3591 (N_3591,N_198,N_303);
and U3592 (N_3592,N_901,N_1925);
nor U3593 (N_3593,N_495,N_1532);
or U3594 (N_3594,N_420,N_1014);
nand U3595 (N_3595,N_1784,N_943);
nor U3596 (N_3596,N_1422,N_529);
and U3597 (N_3597,N_1046,N_816);
nor U3598 (N_3598,N_1798,N_1573);
nand U3599 (N_3599,N_612,N_42);
nor U3600 (N_3600,N_122,N_622);
and U3601 (N_3601,N_681,N_390);
and U3602 (N_3602,N_397,N_84);
and U3603 (N_3603,N_344,N_1836);
nand U3604 (N_3604,N_371,N_1490);
or U3605 (N_3605,N_1108,N_754);
xnor U3606 (N_3606,N_46,N_861);
and U3607 (N_3607,N_1936,N_1599);
and U3608 (N_3608,N_797,N_87);
nor U3609 (N_3609,N_899,N_572);
nand U3610 (N_3610,N_837,N_1465);
nand U3611 (N_3611,N_1089,N_721);
nand U3612 (N_3612,N_589,N_422);
nand U3613 (N_3613,N_44,N_1713);
nand U3614 (N_3614,N_1574,N_554);
nor U3615 (N_3615,N_182,N_1235);
and U3616 (N_3616,N_488,N_206);
and U3617 (N_3617,N_1204,N_1223);
or U3618 (N_3618,N_404,N_1589);
nand U3619 (N_3619,N_1254,N_782);
or U3620 (N_3620,N_1100,N_370);
nand U3621 (N_3621,N_1972,N_570);
or U3622 (N_3622,N_563,N_1782);
and U3623 (N_3623,N_425,N_338);
and U3624 (N_3624,N_1026,N_1628);
nor U3625 (N_3625,N_1835,N_1808);
or U3626 (N_3626,N_1212,N_1050);
and U3627 (N_3627,N_1667,N_533);
nand U3628 (N_3628,N_1104,N_1228);
nand U3629 (N_3629,N_1301,N_1629);
and U3630 (N_3630,N_1507,N_168);
or U3631 (N_3631,N_1998,N_1748);
or U3632 (N_3632,N_1702,N_1402);
nor U3633 (N_3633,N_850,N_1495);
nor U3634 (N_3634,N_71,N_1850);
nor U3635 (N_3635,N_1655,N_1541);
nor U3636 (N_3636,N_1405,N_1275);
nor U3637 (N_3637,N_1543,N_1366);
or U3638 (N_3638,N_1126,N_962);
or U3639 (N_3639,N_785,N_1022);
or U3640 (N_3640,N_1405,N_940);
and U3641 (N_3641,N_1577,N_1796);
nor U3642 (N_3642,N_191,N_1697);
and U3643 (N_3643,N_1265,N_1853);
or U3644 (N_3644,N_893,N_1176);
and U3645 (N_3645,N_1044,N_1170);
nor U3646 (N_3646,N_1314,N_548);
nand U3647 (N_3647,N_91,N_1571);
nand U3648 (N_3648,N_175,N_1479);
or U3649 (N_3649,N_1399,N_1870);
nand U3650 (N_3650,N_923,N_1629);
and U3651 (N_3651,N_1829,N_866);
or U3652 (N_3652,N_1365,N_146);
or U3653 (N_3653,N_446,N_416);
and U3654 (N_3654,N_1196,N_1725);
and U3655 (N_3655,N_336,N_1870);
or U3656 (N_3656,N_742,N_813);
or U3657 (N_3657,N_998,N_1726);
nor U3658 (N_3658,N_201,N_167);
and U3659 (N_3659,N_1555,N_870);
nand U3660 (N_3660,N_528,N_134);
nand U3661 (N_3661,N_554,N_486);
nor U3662 (N_3662,N_822,N_623);
and U3663 (N_3663,N_1293,N_1302);
or U3664 (N_3664,N_1574,N_1038);
and U3665 (N_3665,N_1461,N_1299);
nand U3666 (N_3666,N_426,N_1495);
nor U3667 (N_3667,N_1116,N_755);
or U3668 (N_3668,N_1460,N_511);
or U3669 (N_3669,N_319,N_1024);
nand U3670 (N_3670,N_307,N_1305);
nand U3671 (N_3671,N_1722,N_67);
or U3672 (N_3672,N_1329,N_1067);
or U3673 (N_3673,N_1516,N_79);
and U3674 (N_3674,N_1099,N_1342);
nand U3675 (N_3675,N_746,N_1191);
nand U3676 (N_3676,N_1870,N_1019);
and U3677 (N_3677,N_876,N_1526);
nand U3678 (N_3678,N_641,N_1038);
and U3679 (N_3679,N_254,N_43);
and U3680 (N_3680,N_156,N_1189);
nand U3681 (N_3681,N_506,N_191);
nor U3682 (N_3682,N_901,N_697);
nor U3683 (N_3683,N_1353,N_666);
nor U3684 (N_3684,N_1374,N_266);
nand U3685 (N_3685,N_186,N_1052);
nand U3686 (N_3686,N_1082,N_1334);
nand U3687 (N_3687,N_582,N_470);
nand U3688 (N_3688,N_1022,N_159);
or U3689 (N_3689,N_677,N_533);
nand U3690 (N_3690,N_530,N_1994);
nand U3691 (N_3691,N_432,N_943);
and U3692 (N_3692,N_774,N_686);
or U3693 (N_3693,N_1102,N_1831);
nor U3694 (N_3694,N_1136,N_1899);
nand U3695 (N_3695,N_357,N_1716);
nand U3696 (N_3696,N_1430,N_1105);
nand U3697 (N_3697,N_1035,N_840);
and U3698 (N_3698,N_330,N_621);
nand U3699 (N_3699,N_1365,N_1401);
or U3700 (N_3700,N_1648,N_1786);
or U3701 (N_3701,N_654,N_1868);
or U3702 (N_3702,N_1462,N_1873);
and U3703 (N_3703,N_25,N_1068);
and U3704 (N_3704,N_751,N_1881);
and U3705 (N_3705,N_1009,N_131);
nand U3706 (N_3706,N_601,N_781);
and U3707 (N_3707,N_1748,N_208);
nor U3708 (N_3708,N_84,N_1741);
nor U3709 (N_3709,N_561,N_432);
or U3710 (N_3710,N_727,N_765);
and U3711 (N_3711,N_338,N_1061);
and U3712 (N_3712,N_1440,N_106);
nor U3713 (N_3713,N_553,N_822);
nand U3714 (N_3714,N_501,N_25);
nand U3715 (N_3715,N_1049,N_1485);
nand U3716 (N_3716,N_912,N_248);
nand U3717 (N_3717,N_1748,N_479);
nand U3718 (N_3718,N_1418,N_1219);
and U3719 (N_3719,N_1609,N_1004);
xnor U3720 (N_3720,N_972,N_812);
nand U3721 (N_3721,N_1151,N_1372);
nand U3722 (N_3722,N_1253,N_1932);
nor U3723 (N_3723,N_1572,N_890);
nor U3724 (N_3724,N_1295,N_238);
nor U3725 (N_3725,N_76,N_757);
or U3726 (N_3726,N_816,N_1090);
or U3727 (N_3727,N_1455,N_676);
nand U3728 (N_3728,N_7,N_168);
nand U3729 (N_3729,N_82,N_920);
nand U3730 (N_3730,N_1501,N_711);
nand U3731 (N_3731,N_1282,N_1922);
nand U3732 (N_3732,N_666,N_659);
nand U3733 (N_3733,N_778,N_274);
nor U3734 (N_3734,N_249,N_103);
nand U3735 (N_3735,N_716,N_606);
nand U3736 (N_3736,N_419,N_807);
or U3737 (N_3737,N_1352,N_1317);
nor U3738 (N_3738,N_1337,N_1904);
and U3739 (N_3739,N_1305,N_1226);
and U3740 (N_3740,N_1791,N_400);
nand U3741 (N_3741,N_1214,N_583);
and U3742 (N_3742,N_0,N_188);
xor U3743 (N_3743,N_1913,N_1110);
nand U3744 (N_3744,N_1469,N_227);
or U3745 (N_3745,N_603,N_120);
and U3746 (N_3746,N_868,N_1657);
nand U3747 (N_3747,N_642,N_1820);
and U3748 (N_3748,N_809,N_844);
nor U3749 (N_3749,N_195,N_488);
or U3750 (N_3750,N_197,N_446);
nor U3751 (N_3751,N_347,N_566);
and U3752 (N_3752,N_1381,N_1793);
nor U3753 (N_3753,N_1845,N_320);
nand U3754 (N_3754,N_1236,N_57);
and U3755 (N_3755,N_1138,N_1760);
and U3756 (N_3756,N_832,N_1010);
nand U3757 (N_3757,N_1552,N_1337);
or U3758 (N_3758,N_1869,N_880);
or U3759 (N_3759,N_1012,N_1191);
and U3760 (N_3760,N_1702,N_878);
and U3761 (N_3761,N_1597,N_65);
nand U3762 (N_3762,N_1978,N_131);
or U3763 (N_3763,N_817,N_1561);
and U3764 (N_3764,N_522,N_1915);
and U3765 (N_3765,N_114,N_223);
and U3766 (N_3766,N_576,N_1895);
nor U3767 (N_3767,N_1613,N_565);
and U3768 (N_3768,N_1043,N_1117);
and U3769 (N_3769,N_797,N_559);
and U3770 (N_3770,N_1779,N_1763);
and U3771 (N_3771,N_609,N_250);
nand U3772 (N_3772,N_383,N_538);
and U3773 (N_3773,N_1390,N_505);
nor U3774 (N_3774,N_1011,N_1979);
nand U3775 (N_3775,N_266,N_805);
nor U3776 (N_3776,N_1454,N_750);
or U3777 (N_3777,N_1262,N_1935);
and U3778 (N_3778,N_1695,N_318);
nand U3779 (N_3779,N_862,N_1300);
or U3780 (N_3780,N_1274,N_1923);
nand U3781 (N_3781,N_76,N_1540);
and U3782 (N_3782,N_316,N_1804);
and U3783 (N_3783,N_707,N_1794);
nand U3784 (N_3784,N_417,N_134);
and U3785 (N_3785,N_1532,N_829);
nand U3786 (N_3786,N_1523,N_788);
and U3787 (N_3787,N_665,N_583);
and U3788 (N_3788,N_1758,N_598);
and U3789 (N_3789,N_1075,N_161);
or U3790 (N_3790,N_423,N_1977);
nand U3791 (N_3791,N_925,N_1202);
nand U3792 (N_3792,N_1497,N_1220);
nor U3793 (N_3793,N_1401,N_1404);
and U3794 (N_3794,N_124,N_227);
nor U3795 (N_3795,N_73,N_1359);
nor U3796 (N_3796,N_1263,N_1406);
nand U3797 (N_3797,N_860,N_1111);
nand U3798 (N_3798,N_278,N_855);
nand U3799 (N_3799,N_1125,N_1836);
xor U3800 (N_3800,N_753,N_56);
or U3801 (N_3801,N_1974,N_1378);
xnor U3802 (N_3802,N_1902,N_1678);
or U3803 (N_3803,N_1681,N_1006);
or U3804 (N_3804,N_1661,N_197);
or U3805 (N_3805,N_293,N_604);
nand U3806 (N_3806,N_901,N_200);
nor U3807 (N_3807,N_991,N_866);
and U3808 (N_3808,N_1857,N_116);
nand U3809 (N_3809,N_902,N_1140);
nor U3810 (N_3810,N_1205,N_96);
and U3811 (N_3811,N_1084,N_824);
or U3812 (N_3812,N_255,N_1119);
nand U3813 (N_3813,N_208,N_1658);
nor U3814 (N_3814,N_155,N_173);
or U3815 (N_3815,N_1015,N_87);
nand U3816 (N_3816,N_550,N_140);
and U3817 (N_3817,N_1730,N_703);
nand U3818 (N_3818,N_244,N_1503);
and U3819 (N_3819,N_781,N_825);
nor U3820 (N_3820,N_1730,N_142);
and U3821 (N_3821,N_525,N_1665);
nand U3822 (N_3822,N_671,N_266);
nand U3823 (N_3823,N_1887,N_230);
and U3824 (N_3824,N_1119,N_735);
nand U3825 (N_3825,N_956,N_1982);
nand U3826 (N_3826,N_817,N_731);
nor U3827 (N_3827,N_78,N_1156);
nor U3828 (N_3828,N_360,N_1176);
nor U3829 (N_3829,N_107,N_1798);
nor U3830 (N_3830,N_261,N_1269);
and U3831 (N_3831,N_289,N_127);
and U3832 (N_3832,N_1618,N_6);
and U3833 (N_3833,N_1805,N_966);
nand U3834 (N_3834,N_1634,N_1462);
and U3835 (N_3835,N_1730,N_299);
or U3836 (N_3836,N_1642,N_594);
nand U3837 (N_3837,N_599,N_1218);
nand U3838 (N_3838,N_736,N_350);
nor U3839 (N_3839,N_1947,N_1544);
nor U3840 (N_3840,N_1439,N_858);
xnor U3841 (N_3841,N_248,N_924);
nor U3842 (N_3842,N_140,N_5);
nor U3843 (N_3843,N_794,N_1751);
and U3844 (N_3844,N_1524,N_1407);
nand U3845 (N_3845,N_1992,N_205);
and U3846 (N_3846,N_628,N_445);
and U3847 (N_3847,N_1153,N_745);
or U3848 (N_3848,N_867,N_1571);
nand U3849 (N_3849,N_1653,N_1964);
or U3850 (N_3850,N_393,N_1472);
and U3851 (N_3851,N_131,N_1994);
nor U3852 (N_3852,N_1145,N_1457);
and U3853 (N_3853,N_1553,N_1727);
nand U3854 (N_3854,N_390,N_1275);
or U3855 (N_3855,N_1722,N_1147);
or U3856 (N_3856,N_21,N_1394);
nand U3857 (N_3857,N_735,N_1424);
and U3858 (N_3858,N_1364,N_85);
or U3859 (N_3859,N_461,N_757);
or U3860 (N_3860,N_194,N_1172);
and U3861 (N_3861,N_940,N_1623);
nor U3862 (N_3862,N_813,N_128);
nand U3863 (N_3863,N_303,N_928);
nor U3864 (N_3864,N_211,N_1034);
nand U3865 (N_3865,N_1472,N_1245);
and U3866 (N_3866,N_1767,N_408);
or U3867 (N_3867,N_897,N_314);
or U3868 (N_3868,N_1684,N_855);
nor U3869 (N_3869,N_1981,N_1688);
or U3870 (N_3870,N_162,N_1824);
nand U3871 (N_3871,N_1274,N_237);
nor U3872 (N_3872,N_682,N_1464);
nor U3873 (N_3873,N_42,N_1702);
nor U3874 (N_3874,N_222,N_1718);
or U3875 (N_3875,N_1971,N_898);
nor U3876 (N_3876,N_946,N_1193);
and U3877 (N_3877,N_1741,N_1375);
and U3878 (N_3878,N_1595,N_1962);
nor U3879 (N_3879,N_398,N_1028);
nor U3880 (N_3880,N_1958,N_1178);
and U3881 (N_3881,N_1566,N_1759);
and U3882 (N_3882,N_723,N_1845);
or U3883 (N_3883,N_1539,N_985);
and U3884 (N_3884,N_1490,N_209);
nor U3885 (N_3885,N_601,N_1179);
and U3886 (N_3886,N_1303,N_1242);
nand U3887 (N_3887,N_1278,N_211);
and U3888 (N_3888,N_410,N_53);
or U3889 (N_3889,N_227,N_458);
and U3890 (N_3890,N_547,N_1572);
nor U3891 (N_3891,N_206,N_1849);
nor U3892 (N_3892,N_434,N_1117);
or U3893 (N_3893,N_821,N_1852);
and U3894 (N_3894,N_1991,N_1052);
and U3895 (N_3895,N_1448,N_1741);
nor U3896 (N_3896,N_435,N_1863);
or U3897 (N_3897,N_1047,N_457);
nand U3898 (N_3898,N_1561,N_88);
nand U3899 (N_3899,N_1115,N_1769);
nor U3900 (N_3900,N_792,N_1775);
and U3901 (N_3901,N_675,N_274);
nor U3902 (N_3902,N_434,N_681);
or U3903 (N_3903,N_1447,N_1210);
nor U3904 (N_3904,N_1299,N_595);
nand U3905 (N_3905,N_1525,N_1406);
or U3906 (N_3906,N_1056,N_755);
nor U3907 (N_3907,N_704,N_432);
nor U3908 (N_3908,N_1750,N_305);
and U3909 (N_3909,N_777,N_491);
nand U3910 (N_3910,N_55,N_1502);
nand U3911 (N_3911,N_623,N_1522);
nand U3912 (N_3912,N_1281,N_244);
nor U3913 (N_3913,N_1953,N_634);
nor U3914 (N_3914,N_585,N_1160);
nand U3915 (N_3915,N_676,N_1000);
nand U3916 (N_3916,N_985,N_844);
and U3917 (N_3917,N_1524,N_1792);
nor U3918 (N_3918,N_771,N_1210);
nand U3919 (N_3919,N_952,N_1674);
nor U3920 (N_3920,N_1578,N_1088);
nand U3921 (N_3921,N_620,N_1987);
or U3922 (N_3922,N_1213,N_1293);
nor U3923 (N_3923,N_1845,N_337);
nor U3924 (N_3924,N_214,N_201);
nand U3925 (N_3925,N_467,N_1860);
nand U3926 (N_3926,N_1822,N_1220);
nor U3927 (N_3927,N_1342,N_421);
nor U3928 (N_3928,N_126,N_1910);
and U3929 (N_3929,N_1935,N_116);
and U3930 (N_3930,N_157,N_512);
nand U3931 (N_3931,N_1848,N_1678);
and U3932 (N_3932,N_203,N_1779);
nor U3933 (N_3933,N_117,N_1533);
and U3934 (N_3934,N_697,N_1660);
and U3935 (N_3935,N_689,N_1060);
or U3936 (N_3936,N_1812,N_461);
and U3937 (N_3937,N_1856,N_1533);
and U3938 (N_3938,N_838,N_258);
nand U3939 (N_3939,N_931,N_193);
nand U3940 (N_3940,N_1073,N_748);
or U3941 (N_3941,N_1098,N_242);
nor U3942 (N_3942,N_617,N_514);
nor U3943 (N_3943,N_1331,N_1188);
nor U3944 (N_3944,N_1578,N_765);
nor U3945 (N_3945,N_1861,N_1056);
and U3946 (N_3946,N_490,N_1160);
or U3947 (N_3947,N_71,N_968);
nor U3948 (N_3948,N_399,N_454);
or U3949 (N_3949,N_163,N_1834);
or U3950 (N_3950,N_1675,N_325);
nor U3951 (N_3951,N_1764,N_72);
nor U3952 (N_3952,N_340,N_1397);
and U3953 (N_3953,N_707,N_395);
nand U3954 (N_3954,N_401,N_1400);
and U3955 (N_3955,N_617,N_402);
and U3956 (N_3956,N_1955,N_1383);
and U3957 (N_3957,N_83,N_1242);
nor U3958 (N_3958,N_745,N_402);
or U3959 (N_3959,N_1484,N_1579);
and U3960 (N_3960,N_560,N_1570);
or U3961 (N_3961,N_1220,N_246);
and U3962 (N_3962,N_1490,N_286);
or U3963 (N_3963,N_689,N_1821);
nand U3964 (N_3964,N_1728,N_29);
nand U3965 (N_3965,N_219,N_1610);
nand U3966 (N_3966,N_301,N_1222);
or U3967 (N_3967,N_999,N_177);
or U3968 (N_3968,N_1361,N_1738);
and U3969 (N_3969,N_1388,N_974);
nand U3970 (N_3970,N_1612,N_651);
and U3971 (N_3971,N_519,N_357);
nand U3972 (N_3972,N_870,N_1355);
or U3973 (N_3973,N_1309,N_1367);
nor U3974 (N_3974,N_1607,N_651);
nor U3975 (N_3975,N_1959,N_1860);
and U3976 (N_3976,N_1126,N_1953);
nor U3977 (N_3977,N_1855,N_712);
nand U3978 (N_3978,N_852,N_210);
and U3979 (N_3979,N_571,N_1443);
nand U3980 (N_3980,N_1764,N_1459);
nand U3981 (N_3981,N_292,N_875);
and U3982 (N_3982,N_1662,N_561);
nand U3983 (N_3983,N_1478,N_1054);
or U3984 (N_3984,N_1459,N_713);
and U3985 (N_3985,N_753,N_883);
nor U3986 (N_3986,N_298,N_140);
nand U3987 (N_3987,N_1455,N_151);
and U3988 (N_3988,N_1419,N_1874);
or U3989 (N_3989,N_437,N_1253);
and U3990 (N_3990,N_98,N_867);
nor U3991 (N_3991,N_310,N_739);
or U3992 (N_3992,N_1220,N_893);
nand U3993 (N_3993,N_287,N_377);
nor U3994 (N_3994,N_1081,N_1647);
or U3995 (N_3995,N_1747,N_1040);
and U3996 (N_3996,N_96,N_1273);
and U3997 (N_3997,N_1007,N_1027);
nand U3998 (N_3998,N_979,N_1542);
or U3999 (N_3999,N_1123,N_851);
nor U4000 (N_4000,N_2689,N_2589);
and U4001 (N_4001,N_2016,N_2334);
nand U4002 (N_4002,N_3445,N_3397);
or U4003 (N_4003,N_2992,N_2111);
nor U4004 (N_4004,N_2539,N_2506);
or U4005 (N_4005,N_3712,N_2869);
or U4006 (N_4006,N_2791,N_3877);
nand U4007 (N_4007,N_2048,N_2525);
and U4008 (N_4008,N_3178,N_2878);
or U4009 (N_4009,N_2667,N_2756);
nand U4010 (N_4010,N_2021,N_3377);
nand U4011 (N_4011,N_2884,N_3334);
or U4012 (N_4012,N_2768,N_2158);
and U4013 (N_4013,N_3001,N_2957);
nor U4014 (N_4014,N_3073,N_3801);
nand U4015 (N_4015,N_3803,N_2676);
nor U4016 (N_4016,N_3759,N_3161);
and U4017 (N_4017,N_3070,N_3850);
nand U4018 (N_4018,N_2462,N_3513);
or U4019 (N_4019,N_2601,N_2772);
and U4020 (N_4020,N_3711,N_3989);
nor U4021 (N_4021,N_3743,N_2566);
or U4022 (N_4022,N_3926,N_2688);
nor U4023 (N_4023,N_2207,N_3741);
nor U4024 (N_4024,N_2128,N_3565);
nand U4025 (N_4025,N_2340,N_2170);
nand U4026 (N_4026,N_3406,N_2242);
nand U4027 (N_4027,N_2897,N_3627);
nor U4028 (N_4028,N_3853,N_3085);
xor U4029 (N_4029,N_2697,N_3844);
nand U4030 (N_4030,N_2180,N_2874);
or U4031 (N_4031,N_3917,N_3997);
nor U4032 (N_4032,N_3814,N_2445);
and U4033 (N_4033,N_3272,N_3974);
and U4034 (N_4034,N_3179,N_2124);
nor U4035 (N_4035,N_3092,N_3184);
nand U4036 (N_4036,N_2763,N_2121);
nor U4037 (N_4037,N_2999,N_3376);
and U4038 (N_4038,N_2843,N_2101);
or U4039 (N_4039,N_2977,N_3097);
nand U4040 (N_4040,N_3261,N_3133);
or U4041 (N_4041,N_3505,N_3613);
nand U4042 (N_4042,N_3914,N_3698);
and U4043 (N_4043,N_2246,N_2153);
or U4044 (N_4044,N_2820,N_3739);
nor U4045 (N_4045,N_2454,N_3553);
nor U4046 (N_4046,N_2375,N_3177);
nor U4047 (N_4047,N_3436,N_2659);
or U4048 (N_4048,N_2133,N_3316);
or U4049 (N_4049,N_2737,N_2726);
and U4050 (N_4050,N_3125,N_3905);
nor U4051 (N_4051,N_2480,N_2393);
and U4052 (N_4052,N_3274,N_3416);
nand U4053 (N_4053,N_2028,N_2013);
and U4054 (N_4054,N_3715,N_3109);
nand U4055 (N_4055,N_2736,N_2686);
nor U4056 (N_4056,N_2652,N_3754);
xnor U4057 (N_4057,N_2512,N_3495);
nand U4058 (N_4058,N_3786,N_3497);
or U4059 (N_4059,N_2492,N_3636);
nand U4060 (N_4060,N_3017,N_3867);
nand U4061 (N_4061,N_3752,N_2071);
and U4062 (N_4062,N_3313,N_3755);
nand U4063 (N_4063,N_2495,N_2727);
or U4064 (N_4064,N_2455,N_2550);
and U4065 (N_4065,N_2027,N_2298);
nor U4066 (N_4066,N_3170,N_2755);
nand U4067 (N_4067,N_2099,N_2945);
or U4068 (N_4068,N_3821,N_3071);
nand U4069 (N_4069,N_3493,N_2672);
and U4070 (N_4070,N_2493,N_2871);
xnor U4071 (N_4071,N_3387,N_2750);
nor U4072 (N_4072,N_2963,N_2831);
or U4073 (N_4073,N_2534,N_2797);
or U4074 (N_4074,N_2400,N_3560);
xnor U4075 (N_4075,N_2678,N_3175);
nor U4076 (N_4076,N_2287,N_2472);
or U4077 (N_4077,N_2961,N_3536);
or U4078 (N_4078,N_2856,N_3007);
and U4079 (N_4079,N_3064,N_2145);
nor U4080 (N_4080,N_2932,N_2799);
and U4081 (N_4081,N_3310,N_2698);
nand U4082 (N_4082,N_3081,N_3790);
or U4083 (N_4083,N_2279,N_2829);
nor U4084 (N_4084,N_3008,N_2909);
and U4085 (N_4085,N_3537,N_2980);
nor U4086 (N_4086,N_2079,N_2885);
and U4087 (N_4087,N_3768,N_2707);
nand U4088 (N_4088,N_3874,N_3290);
and U4089 (N_4089,N_2709,N_3732);
nand U4090 (N_4090,N_2571,N_2914);
and U4091 (N_4091,N_3471,N_2379);
and U4092 (N_4092,N_2511,N_2155);
and U4093 (N_4093,N_2777,N_3047);
and U4094 (N_4094,N_2708,N_3841);
and U4095 (N_4095,N_2783,N_2494);
nor U4096 (N_4096,N_3222,N_2136);
or U4097 (N_4097,N_2320,N_3681);
and U4098 (N_4098,N_2398,N_2805);
and U4099 (N_4099,N_3697,N_2962);
nor U4100 (N_4100,N_3022,N_2793);
nor U4101 (N_4101,N_2841,N_2625);
nor U4102 (N_4102,N_3656,N_2931);
nand U4103 (N_4103,N_3561,N_2866);
or U4104 (N_4104,N_3442,N_2074);
or U4105 (N_4105,N_3534,N_2024);
and U4106 (N_4106,N_3136,N_2796);
or U4107 (N_4107,N_3117,N_3668);
and U4108 (N_4108,N_2618,N_2801);
and U4109 (N_4109,N_3921,N_2558);
or U4110 (N_4110,N_3903,N_3908);
and U4111 (N_4111,N_2231,N_3729);
nor U4112 (N_4112,N_2030,N_3373);
or U4113 (N_4113,N_3480,N_3542);
nand U4114 (N_4114,N_2792,N_2000);
and U4115 (N_4115,N_3925,N_2463);
and U4116 (N_4116,N_2515,N_2628);
nand U4117 (N_4117,N_2330,N_2461);
nor U4118 (N_4118,N_2129,N_2259);
or U4119 (N_4119,N_2257,N_2836);
xnor U4120 (N_4120,N_2825,N_2468);
nand U4121 (N_4121,N_2517,N_3454);
or U4122 (N_4122,N_2859,N_3153);
or U4123 (N_4123,N_2561,N_3395);
and U4124 (N_4124,N_2953,N_3564);
and U4125 (N_4125,N_3713,N_3127);
nand U4126 (N_4126,N_3937,N_2673);
or U4127 (N_4127,N_2085,N_2491);
nand U4128 (N_4128,N_3082,N_2536);
or U4129 (N_4129,N_2335,N_3095);
or U4130 (N_4130,N_3842,N_3583);
nand U4131 (N_4131,N_3407,N_3393);
nand U4132 (N_4132,N_3916,N_3413);
and U4133 (N_4133,N_3152,N_3275);
or U4134 (N_4134,N_3483,N_3485);
nand U4135 (N_4135,N_2970,N_2409);
and U4136 (N_4136,N_2834,N_3455);
or U4137 (N_4137,N_3329,N_3242);
and U4138 (N_4138,N_2587,N_2091);
or U4139 (N_4139,N_3632,N_2235);
nor U4140 (N_4140,N_2405,N_2657);
nand U4141 (N_4141,N_3060,N_2958);
nor U4142 (N_4142,N_3006,N_3155);
nand U4143 (N_4143,N_2723,N_3492);
nand U4144 (N_4144,N_2993,N_3617);
nand U4145 (N_4145,N_2290,N_3769);
nor U4146 (N_4146,N_2634,N_2413);
nor U4147 (N_4147,N_2386,N_2488);
or U4148 (N_4148,N_2579,N_2478);
nand U4149 (N_4149,N_3321,N_2046);
nand U4150 (N_4150,N_3298,N_2784);
or U4151 (N_4151,N_3730,N_2102);
nand U4152 (N_4152,N_2728,N_3980);
nor U4153 (N_4153,N_2466,N_3646);
or U4154 (N_4154,N_3360,N_2378);
and U4155 (N_4155,N_3602,N_3600);
or U4156 (N_4156,N_3423,N_2865);
nor U4157 (N_4157,N_3389,N_2818);
and U4158 (N_4158,N_3140,N_3106);
and U4159 (N_4159,N_2321,N_3836);
and U4160 (N_4160,N_2949,N_2427);
and U4161 (N_4161,N_3888,N_2292);
nor U4162 (N_4162,N_2918,N_3209);
nor U4163 (N_4163,N_3535,N_2654);
and U4164 (N_4164,N_2045,N_3501);
nand U4165 (N_4165,N_3545,N_2645);
nand U4166 (N_4166,N_2870,N_3009);
or U4167 (N_4167,N_2891,N_3132);
or U4168 (N_4168,N_3327,N_3883);
or U4169 (N_4169,N_3939,N_2985);
and U4170 (N_4170,N_3691,N_3585);
nand U4171 (N_4171,N_2901,N_3453);
nor U4172 (N_4172,N_2842,N_3169);
or U4173 (N_4173,N_3005,N_2191);
nand U4174 (N_4174,N_2329,N_2296);
nor U4175 (N_4175,N_3573,N_2975);
nor U4176 (N_4176,N_3651,N_2019);
nand U4177 (N_4177,N_2274,N_2787);
nand U4178 (N_4178,N_2327,N_2526);
or U4179 (N_4179,N_2267,N_3895);
and U4180 (N_4180,N_2749,N_2058);
and U4181 (N_4181,N_2956,N_2535);
nand U4182 (N_4182,N_2700,N_2118);
nor U4183 (N_4183,N_2623,N_3093);
nor U4184 (N_4184,N_3910,N_2368);
nor U4185 (N_4185,N_2778,N_3748);
nand U4186 (N_4186,N_3578,N_3864);
or U4187 (N_4187,N_3719,N_2720);
or U4188 (N_4188,N_3674,N_3278);
or U4189 (N_4189,N_3918,N_2853);
nor U4190 (N_4190,N_3011,N_3474);
and U4191 (N_4191,N_3685,N_2845);
nand U4192 (N_4192,N_2317,N_3173);
nor U4193 (N_4193,N_3323,N_3577);
and U4194 (N_4194,N_2939,N_3124);
or U4195 (N_4195,N_2036,N_3516);
nor U4196 (N_4196,N_2916,N_2620);
and U4197 (N_4197,N_2766,N_3171);
nand U4198 (N_4198,N_3723,N_3189);
and U4199 (N_4199,N_3662,N_2301);
or U4200 (N_4200,N_2255,N_3760);
and U4201 (N_4201,N_3663,N_3456);
and U4202 (N_4202,N_2471,N_2731);
nor U4203 (N_4203,N_2470,N_3700);
xor U4204 (N_4204,N_3653,N_2621);
or U4205 (N_4205,N_3607,N_2369);
and U4206 (N_4206,N_2713,N_3049);
nand U4207 (N_4207,N_3818,N_2875);
and U4208 (N_4208,N_2883,N_3250);
or U4209 (N_4209,N_2338,N_2230);
nand U4210 (N_4210,N_2675,N_2313);
or U4211 (N_4211,N_3435,N_2912);
nand U4212 (N_4212,N_2575,N_2524);
nor U4213 (N_4213,N_2994,N_3309);
and U4214 (N_4214,N_2234,N_3235);
nor U4215 (N_4215,N_3608,N_3780);
nand U4216 (N_4216,N_2941,N_3640);
and U4217 (N_4217,N_2568,N_2527);
and U4218 (N_4218,N_2115,N_3104);
and U4219 (N_4219,N_3244,N_2984);
xnor U4220 (N_4220,N_3227,N_2161);
nor U4221 (N_4221,N_3985,N_2090);
and U4222 (N_4222,N_2940,N_3750);
and U4223 (N_4223,N_2987,N_2500);
or U4224 (N_4224,N_2607,N_3481);
or U4225 (N_4225,N_3524,N_2100);
nor U4226 (N_4226,N_2339,N_3673);
nand U4227 (N_4227,N_3776,N_3637);
and U4228 (N_4228,N_2811,N_2380);
or U4229 (N_4229,N_2052,N_2276);
or U4230 (N_4230,N_2421,N_3225);
or U4231 (N_4231,N_3402,N_3603);
or U4232 (N_4232,N_3294,N_3188);
nand U4233 (N_4233,N_2294,N_2757);
xor U4234 (N_4234,N_2848,N_3077);
and U4235 (N_4235,N_2410,N_3464);
nor U4236 (N_4236,N_3975,N_3307);
and U4237 (N_4237,N_3671,N_3122);
xnor U4238 (N_4238,N_2862,N_2809);
and U4239 (N_4239,N_3433,N_3913);
nand U4240 (N_4240,N_2574,N_3202);
nor U4241 (N_4241,N_3869,N_3417);
and U4242 (N_4242,N_3625,N_2611);
and U4243 (N_4243,N_2549,N_3447);
nor U4244 (N_4244,N_3199,N_3399);
xor U4245 (N_4245,N_3285,N_2879);
nand U4246 (N_4246,N_2826,N_3030);
nand U4247 (N_4247,N_2489,N_2752);
or U4248 (N_4248,N_2724,N_2564);
or U4249 (N_4249,N_2050,N_2229);
and U4250 (N_4250,N_2997,N_3411);
nor U4251 (N_4251,N_3530,N_3245);
or U4252 (N_4252,N_2254,N_2163);
or U4253 (N_4253,N_2053,N_3830);
nor U4254 (N_4254,N_3142,N_2141);
or U4255 (N_4255,N_2089,N_3486);
nor U4256 (N_4256,N_2840,N_3519);
nand U4257 (N_4257,N_3034,N_3343);
or U4258 (N_4258,N_3894,N_2532);
xor U4259 (N_4259,N_3725,N_3540);
or U4260 (N_4260,N_3158,N_3159);
nor U4261 (N_4261,N_2821,N_2886);
nor U4262 (N_4262,N_2239,N_2671);
nor U4263 (N_4263,N_3183,N_2599);
nand U4264 (N_4264,N_3788,N_3805);
and U4265 (N_4265,N_3851,N_2907);
and U4266 (N_4266,N_3123,N_2670);
and U4267 (N_4267,N_3466,N_3981);
nand U4268 (N_4268,N_2363,N_3504);
nand U4269 (N_4269,N_2224,N_3940);
nand U4270 (N_4270,N_3708,N_2774);
and U4271 (N_4271,N_2241,N_2325);
and U4272 (N_4272,N_3134,N_2804);
or U4273 (N_4273,N_3482,N_3665);
or U4274 (N_4274,N_2819,N_3478);
and U4275 (N_4275,N_2600,N_3872);
or U4276 (N_4276,N_2425,N_2084);
nor U4277 (N_4277,N_3870,N_2808);
nor U4278 (N_4278,N_3388,N_3441);
nor U4279 (N_4279,N_3782,N_2236);
and U4280 (N_4280,N_3410,N_3563);
nor U4281 (N_4281,N_2057,N_2767);
and U4282 (N_4282,N_3088,N_3431);
or U4283 (N_4283,N_2733,N_3051);
or U4284 (N_4284,N_2182,N_2986);
and U4285 (N_4285,N_2633,N_2637);
nand U4286 (N_4286,N_3476,N_2666);
nor U4287 (N_4287,N_2350,N_3138);
or U4288 (N_4288,N_2248,N_3150);
or U4289 (N_4289,N_2098,N_3567);
and U4290 (N_4290,N_2648,N_2245);
or U4291 (N_4291,N_2597,N_3652);
nand U4292 (N_4292,N_3233,N_3231);
nor U4293 (N_4293,N_3210,N_2401);
nand U4294 (N_4294,N_2938,N_3684);
nor U4295 (N_4295,N_2691,N_2031);
and U4296 (N_4296,N_3381,N_2377);
and U4297 (N_4297,N_3054,N_3016);
and U4298 (N_4298,N_2093,N_2020);
nor U4299 (N_4299,N_3689,N_2384);
and U4300 (N_4300,N_2894,N_2919);
and U4301 (N_4301,N_3187,N_2747);
nor U4302 (N_4302,N_2586,N_2603);
or U4303 (N_4303,N_2244,N_3067);
nor U4304 (N_4304,N_2012,N_3165);
or U4305 (N_4305,N_2521,N_3581);
or U4306 (N_4306,N_2982,N_3121);
nor U4307 (N_4307,N_2694,N_2483);
nor U4308 (N_4308,N_3434,N_2920);
or U4309 (N_4309,N_3988,N_2237);
and U4310 (N_4310,N_2927,N_3499);
or U4311 (N_4311,N_3084,N_3021);
and U4312 (N_4312,N_2929,N_3889);
nand U4313 (N_4313,N_3325,N_2559);
or U4314 (N_4314,N_3518,N_2922);
nor U4315 (N_4315,N_3284,N_3770);
or U4316 (N_4316,N_3197,N_3208);
and U4317 (N_4317,N_2433,N_2573);
and U4318 (N_4318,N_2505,N_2520);
nor U4319 (N_4319,N_2469,N_3628);
and U4320 (N_4320,N_3630,N_3962);
nand U4321 (N_4321,N_2125,N_2047);
nand U4322 (N_4322,N_2418,N_3699);
or U4323 (N_4323,N_2215,N_2399);
and U4324 (N_4324,N_2164,N_3773);
nor U4325 (N_4325,N_2703,N_3425);
nor U4326 (N_4326,N_3920,N_3484);
or U4327 (N_4327,N_3606,N_3282);
and U4328 (N_4328,N_2827,N_3463);
and U4329 (N_4329,N_3787,N_2309);
nor U4330 (N_4330,N_2890,N_2198);
nor U4331 (N_4331,N_3449,N_3437);
or U4332 (N_4332,N_2223,N_3828);
nor U4333 (N_4333,N_2417,N_2665);
nor U4334 (N_4334,N_2528,N_3664);
and U4335 (N_4335,N_3429,N_2714);
or U4336 (N_4336,N_2502,N_2277);
nand U4337 (N_4337,N_3907,N_3461);
nand U4338 (N_4338,N_2779,N_3057);
or U4339 (N_4339,N_2943,N_3220);
nand U4340 (N_4340,N_2770,N_3965);
and U4341 (N_4341,N_3252,N_3503);
nor U4342 (N_4342,N_3297,N_3871);
or U4343 (N_4343,N_3766,N_3881);
or U4344 (N_4344,N_3605,N_2314);
and U4345 (N_4345,N_3820,N_2218);
nor U4346 (N_4346,N_3742,N_3228);
or U4347 (N_4347,N_3586,N_2202);
and U4348 (N_4348,N_2188,N_3288);
and U4349 (N_4349,N_2817,N_3837);
nand U4350 (N_4350,N_2194,N_2852);
or U4351 (N_4351,N_3251,N_3614);
nor U4352 (N_4352,N_3459,N_3706);
nand U4353 (N_4353,N_3858,N_3212);
nor U4354 (N_4354,N_2978,N_3108);
nor U4355 (N_4355,N_3315,N_2664);
or U4356 (N_4356,N_3180,N_2426);
or U4357 (N_4357,N_2881,N_3659);
xnor U4358 (N_4358,N_3115,N_3174);
or U4359 (N_4359,N_2570,N_2186);
or U4360 (N_4360,N_3200,N_2569);
or U4361 (N_4361,N_2744,N_3254);
nor U4362 (N_4362,N_2216,N_2991);
or U4363 (N_4363,N_2134,N_2947);
nor U4364 (N_4364,N_2088,N_3896);
or U4365 (N_4365,N_3103,N_2839);
or U4366 (N_4366,N_3749,N_2580);
and U4367 (N_4367,N_2278,N_3075);
or U4368 (N_4368,N_3487,N_3591);
nor U4369 (N_4369,N_3056,N_3357);
xnor U4370 (N_4370,N_2591,N_2269);
nand U4371 (N_4371,N_2452,N_2548);
nor U4372 (N_4372,N_2157,N_2467);
nor U4373 (N_4373,N_2109,N_3544);
or U4374 (N_4374,N_3037,N_3796);
or U4375 (N_4375,N_3500,N_2477);
nor U4376 (N_4376,N_2876,N_2432);
and U4377 (N_4377,N_2106,N_2137);
and U4378 (N_4378,N_3405,N_3181);
or U4379 (N_4379,N_3083,N_2073);
and U4380 (N_4380,N_3308,N_3306);
or U4381 (N_4381,N_2917,N_2765);
and U4382 (N_4382,N_3015,N_3296);
and U4383 (N_4383,N_3264,N_3216);
and U4384 (N_4384,N_3765,N_2360);
nor U4385 (N_4385,N_3554,N_2729);
nor U4386 (N_4386,N_3584,N_3696);
or U4387 (N_4387,N_3206,N_3987);
and U4388 (N_4388,N_3372,N_3059);
nand U4389 (N_4389,N_2078,N_2374);
or U4390 (N_4390,N_2740,N_2120);
nor U4391 (N_4391,N_3777,N_2116);
nor U4392 (N_4392,N_3594,N_3144);
or U4393 (N_4393,N_3816,N_2760);
and U4394 (N_4394,N_2408,N_3784);
nand U4395 (N_4395,N_2882,N_2365);
and U4396 (N_4396,N_2439,N_2872);
nand U4397 (N_4397,N_2913,N_2190);
and U4398 (N_4398,N_3458,N_2172);
nand U4399 (N_4399,N_3078,N_3361);
nand U4400 (N_4400,N_3761,N_2681);
and U4401 (N_4401,N_2509,N_2609);
nor U4402 (N_4402,N_2795,N_2312);
or U4403 (N_4403,N_2928,N_3624);
and U4404 (N_4404,N_2858,N_3824);
nor U4405 (N_4405,N_2451,N_2734);
or U4406 (N_4406,N_2936,N_2403);
nand U4407 (N_4407,N_3215,N_3195);
or U4408 (N_4408,N_2812,N_2132);
nor U4409 (N_4409,N_2072,N_3404);
nor U4410 (N_4410,N_3198,N_2543);
nand U4411 (N_4411,N_2160,N_3817);
or U4412 (N_4412,N_3855,N_3379);
nand U4413 (N_4413,N_3919,N_2954);
or U4414 (N_4414,N_3301,N_2837);
and U4415 (N_4415,N_3969,N_3904);
or U4416 (N_4416,N_3574,N_2391);
nand U4417 (N_4417,N_3621,N_3927);
nand U4418 (N_4418,N_2002,N_3349);
and U4419 (N_4419,N_3514,N_3634);
nand U4420 (N_4420,N_3641,N_2032);
nand U4421 (N_4421,N_3139,N_3300);
and U4422 (N_4422,N_3572,N_3263);
or U4423 (N_4423,N_2303,N_3938);
or U4424 (N_4424,N_2631,N_3695);
or U4425 (N_4425,N_3885,N_2361);
or U4426 (N_4426,N_2226,N_3866);
or U4427 (N_4427,N_2854,N_3356);
nand U4428 (N_4428,N_3477,N_2476);
nor U4429 (N_4429,N_3055,N_3880);
and U4430 (N_4430,N_2266,N_3234);
nand U4431 (N_4431,N_2265,N_3342);
or U4432 (N_4432,N_3924,N_3137);
or U4433 (N_4433,N_3207,N_3146);
nor U4434 (N_4434,N_3094,N_2307);
nand U4435 (N_4435,N_2889,N_3358);
and U4436 (N_4436,N_3116,N_3619);
and U4437 (N_4437,N_2326,N_2473);
and U4438 (N_4438,N_2143,N_3194);
or U4439 (N_4439,N_3676,N_2453);
nor U4440 (N_4440,N_3999,N_2342);
nand U4441 (N_4441,N_2788,N_3400);
or U4442 (N_4442,N_3887,N_3947);
nand U4443 (N_4443,N_3273,N_3570);
or U4444 (N_4444,N_3221,N_3956);
or U4445 (N_4445,N_2632,N_3147);
nand U4446 (N_4446,N_2660,N_2249);
nand U4447 (N_4447,N_3550,N_2646);
nand U4448 (N_4448,N_3330,N_3018);
or U4449 (N_4449,N_3552,N_2144);
nor U4450 (N_4450,N_3906,N_2873);
nand U4451 (N_4451,N_2605,N_3196);
or U4452 (N_4452,N_3604,N_2844);
nand U4453 (N_4453,N_2437,N_2430);
and U4454 (N_4454,N_3185,N_3143);
nand U4455 (N_4455,N_3595,N_2203);
and U4456 (N_4456,N_3912,N_3176);
and U4457 (N_4457,N_3795,N_2014);
and U4458 (N_4458,N_2064,N_2557);
nand U4459 (N_4459,N_2001,N_3677);
and U4460 (N_4460,N_3266,N_2902);
or U4461 (N_4461,N_3967,N_3559);
and U4462 (N_4462,N_2612,N_2286);
or U4463 (N_4463,N_3558,N_2762);
and U4464 (N_4464,N_3509,N_3355);
and U4465 (N_4465,N_2651,N_3638);
nand U4466 (N_4466,N_3807,N_2304);
and U4467 (N_4467,N_2965,N_2122);
or U4468 (N_4468,N_2710,N_3655);
nor U4469 (N_4469,N_3496,N_3710);
nand U4470 (N_4470,N_2759,N_3762);
or U4471 (N_4471,N_3587,N_2197);
nand U4472 (N_4472,N_2175,N_2486);
nand U4473 (N_4473,N_3390,N_3833);
nand U4474 (N_4474,N_2390,N_3168);
nor U4475 (N_4475,N_2967,N_2066);
and U4476 (N_4476,N_3350,N_2411);
or U4477 (N_4477,N_3172,N_3338);
or U4478 (N_4478,N_3230,N_3915);
nand U4479 (N_4479,N_3701,N_3333);
nand U4480 (N_4480,N_3949,N_2771);
nor U4481 (N_4481,N_2263,N_3353);
nand U4482 (N_4482,N_3792,N_2864);
and U4483 (N_4483,N_3238,N_2183);
or U4484 (N_4484,N_3374,N_2114);
and U4485 (N_4485,N_3053,N_2459);
nor U4486 (N_4486,N_3891,N_3690);
nand U4487 (N_4487,N_3031,N_3738);
and U4488 (N_4488,N_3279,N_2112);
nand U4489 (N_4489,N_2850,N_3365);
nor U4490 (N_4490,N_2687,N_3898);
nor U4491 (N_4491,N_3825,N_3110);
or U4492 (N_4492,N_2416,N_3692);
or U4493 (N_4493,N_3922,N_2113);
and U4494 (N_4494,N_3305,N_2923);
or U4495 (N_4495,N_2608,N_2906);
nor U4496 (N_4496,N_2018,N_2285);
nor U4497 (N_4497,N_3951,N_2966);
nor U4498 (N_4498,N_2227,N_3994);
or U4499 (N_4499,N_3396,N_2711);
and U4500 (N_4500,N_2807,N_3348);
nand U4501 (N_4501,N_3317,N_3237);
or U4502 (N_4502,N_2026,N_3512);
nand U4503 (N_4503,N_2552,N_2833);
or U4504 (N_4504,N_2542,N_2316);
and U4505 (N_4505,N_3694,N_3521);
or U4506 (N_4506,N_2178,N_3860);
nand U4507 (N_4507,N_2565,N_2010);
nor U4508 (N_4508,N_3191,N_2715);
nand U4509 (N_4509,N_2076,N_2998);
nor U4510 (N_4510,N_3667,N_2626);
nand U4511 (N_4511,N_2219,N_3953);
and U4512 (N_4512,N_2513,N_3946);
and U4513 (N_4513,N_2960,N_2696);
nor U4514 (N_4514,N_2444,N_3068);
and U4515 (N_4515,N_2773,N_2062);
nand U4516 (N_4516,N_2522,N_3979);
or U4517 (N_4517,N_2800,N_2187);
xnor U4518 (N_4518,N_3468,N_3354);
nand U4519 (N_4519,N_2006,N_2087);
and U4520 (N_4520,N_2077,N_3223);
nand U4521 (N_4521,N_2638,N_3076);
nand U4522 (N_4522,N_2382,N_3048);
and U4523 (N_4523,N_3538,N_3203);
nand U4524 (N_4524,N_3089,N_3046);
nor U4525 (N_4525,N_2617,N_2156);
xnor U4526 (N_4526,N_2541,N_3775);
and U4527 (N_4527,N_3731,N_2606);
nor U4528 (N_4528,N_2684,N_2680);
nand U4529 (N_4529,N_3204,N_2233);
and U4530 (N_4530,N_2171,N_3815);
and U4531 (N_4531,N_3998,N_3601);
and U4532 (N_4532,N_2220,N_3472);
nor U4533 (N_4533,N_2496,N_2450);
or U4534 (N_4534,N_2567,N_3623);
nor U4535 (N_4535,N_3201,N_2937);
nand U4536 (N_4536,N_3639,N_2004);
or U4537 (N_4537,N_2594,N_3582);
nor U4538 (N_4538,N_2465,N_3930);
or U4539 (N_4539,N_2577,N_3794);
and U4540 (N_4540,N_3112,N_2614);
nor U4541 (N_4541,N_2082,N_2518);
or U4542 (N_4542,N_2926,N_3857);
xor U4543 (N_4543,N_3295,N_3414);
and U4544 (N_4544,N_2123,N_3778);
or U4545 (N_4545,N_2682,N_3113);
nor U4546 (N_4546,N_3100,N_2357);
and U4547 (N_4547,N_2781,N_3658);
and U4548 (N_4548,N_3465,N_3438);
nand U4549 (N_4549,N_3383,N_3352);
and U4550 (N_4550,N_3255,N_2025);
and U4551 (N_4551,N_3211,N_2412);
nor U4552 (N_4552,N_2544,N_2785);
or U4553 (N_4553,N_3096,N_3314);
or U4554 (N_4554,N_2860,N_3933);
or U4555 (N_4555,N_2510,N_3703);
nand U4556 (N_4556,N_2256,N_3253);
and U4557 (N_4557,N_3258,N_2653);
or U4558 (N_4558,N_2428,N_2271);
and U4559 (N_4559,N_3522,N_3276);
and U4560 (N_4560,N_3280,N_3840);
and U4561 (N_4561,N_3767,N_3289);
and U4562 (N_4562,N_2322,N_3098);
or U4563 (N_4563,N_3050,N_2039);
nand U4564 (N_4564,N_2165,N_2832);
nor U4565 (N_4565,N_3024,N_3498);
and U4566 (N_4566,N_3102,N_2447);
or U4567 (N_4567,N_2683,N_2639);
and U4568 (N_4568,N_3430,N_3590);
and U4569 (N_4569,N_3822,N_3571);
and U4570 (N_4570,N_2008,N_2964);
or U4571 (N_4571,N_3875,N_2119);
nand U4572 (N_4572,N_3489,N_2899);
nor U4573 (N_4573,N_3576,N_2397);
and U4574 (N_4574,N_3948,N_2622);
and U4575 (N_4575,N_3367,N_3543);
and U4576 (N_4576,N_3517,N_2201);
nor U4577 (N_4577,N_3727,N_3450);
and U4578 (N_4578,N_2748,N_3268);
or U4579 (N_4579,N_3566,N_2551);
and U4580 (N_4580,N_3226,N_2485);
nand U4581 (N_4581,N_2148,N_3328);
or U4582 (N_4582,N_2022,N_2585);
and U4583 (N_4583,N_2150,N_2924);
nand U4584 (N_4584,N_3062,N_3968);
or U4585 (N_4585,N_3592,N_2446);
and U4586 (N_4586,N_3045,N_2861);
and U4587 (N_4587,N_2649,N_2677);
nand U4588 (N_4588,N_3978,N_3157);
nor U4589 (N_4589,N_3687,N_3923);
and U4590 (N_4590,N_2896,N_2166);
nand U4591 (N_4591,N_3763,N_2699);
and U4592 (N_4592,N_2816,N_2996);
nor U4593 (N_4593,N_3611,N_2741);
nor U4594 (N_4594,N_3791,N_2107);
nor U4595 (N_4595,N_2598,N_2097);
or U4596 (N_4596,N_2806,N_2381);
or U4597 (N_4597,N_3529,N_2297);
and U4598 (N_4598,N_3966,N_2578);
nand U4599 (N_4599,N_2212,N_3944);
and U4600 (N_4600,N_3303,N_3368);
and U4601 (N_4601,N_2376,N_2674);
xor U4602 (N_4602,N_2990,N_2971);
nor U4603 (N_4603,N_3675,N_3588);
nand U4604 (N_4604,N_2537,N_3322);
nor U4605 (N_4605,N_2044,N_3479);
nand U4606 (N_4606,N_3863,N_3058);
nand U4607 (N_4607,N_2149,N_3107);
or U4608 (N_4608,N_3422,N_3546);
nor U4609 (N_4609,N_3154,N_3217);
nand U4610 (N_4610,N_2311,N_3774);
or U4611 (N_4611,N_3364,N_2959);
nand U4612 (N_4612,N_2973,N_2595);
and U4613 (N_4613,N_3013,N_2584);
nand U4614 (N_4614,N_3964,N_3494);
and U4615 (N_4615,N_2498,N_2644);
or U4616 (N_4616,N_3375,N_3335);
nor U4617 (N_4617,N_3849,N_3932);
nand U4618 (N_4618,N_3756,N_2988);
and U4619 (N_4619,N_2604,N_2636);
or U4620 (N_4620,N_3243,N_3337);
or U4621 (N_4621,N_3688,N_3452);
nand U4622 (N_4622,N_2042,N_2900);
nand U4623 (N_4623,N_3019,N_2661);
xor U4624 (N_4624,N_2348,N_3539);
nand U4625 (N_4625,N_3631,N_2138);
and U4626 (N_4626,N_2185,N_3911);
or U4627 (N_4627,N_2822,N_3419);
or U4628 (N_4628,N_3044,N_2615);
and U4629 (N_4629,N_3935,N_3846);
nor U4630 (N_4630,N_2331,N_3241);
nor U4631 (N_4631,N_3718,N_3033);
or U4632 (N_4632,N_3959,N_3678);
and U4633 (N_4633,N_3945,N_3789);
nor U4634 (N_4634,N_2258,N_3304);
or U4635 (N_4635,N_2487,N_3745);
and U4636 (N_4636,N_2474,N_2328);
nand U4637 (N_4637,N_3460,N_2293);
nand U4638 (N_4638,N_2624,N_3679);
or U4639 (N_4639,N_2650,N_2009);
or U4640 (N_4640,N_3260,N_2892);
and U4641 (N_4641,N_2023,N_2989);
and U4642 (N_4642,N_2011,N_2067);
or U4643 (N_4643,N_2855,N_2337);
or U4644 (N_4644,N_2262,N_3802);
and U4645 (N_4645,N_2388,N_2921);
nor U4646 (N_4646,N_3683,N_2824);
and U4647 (N_4647,N_3069,N_3737);
nor U4648 (N_4648,N_2782,N_2555);
and U4649 (N_4649,N_3670,N_3873);
nor U4650 (N_4650,N_3385,N_3467);
nand U4651 (N_4651,N_3548,N_2415);
or U4652 (N_4652,N_2596,N_3733);
nand U4653 (N_4653,N_2305,N_2590);
nand U4654 (N_4654,N_3439,N_3366);
and U4655 (N_4655,N_2746,N_3928);
nor U4656 (N_4656,N_3829,N_3508);
and U4657 (N_4657,N_3020,N_2341);
or U4658 (N_4658,N_3808,N_3672);
or U4659 (N_4659,N_2930,N_2456);
or U4660 (N_4660,N_2359,N_3380);
and U4661 (N_4661,N_3819,N_3528);
nand U4662 (N_4662,N_2951,N_3490);
and U4663 (N_4663,N_2556,N_2823);
nand U4664 (N_4664,N_3726,N_3736);
and U4665 (N_4665,N_3654,N_2068);
nor U4666 (N_4666,N_2802,N_2789);
or U4667 (N_4667,N_3074,N_2619);
and U4668 (N_4668,N_2289,N_2503);
nor U4669 (N_4669,N_2193,N_3000);
or U4670 (N_4670,N_3753,N_3473);
and U4671 (N_4671,N_2602,N_3779);
nor U4672 (N_4672,N_3556,N_2888);
xor U4673 (N_4673,N_3163,N_2081);
and U4674 (N_4674,N_2323,N_2969);
nand U4675 (N_4675,N_2830,N_2497);
nand U4676 (N_4676,N_3444,N_2803);
nor U4677 (N_4677,N_2950,N_3014);
or U4678 (N_4678,N_2662,N_2049);
nand U4679 (N_4679,N_2344,N_2238);
nor U4680 (N_4680,N_3823,N_3345);
or U4681 (N_4681,N_2658,N_2208);
nand U4682 (N_4682,N_3488,N_3101);
and U4683 (N_4683,N_2847,N_2704);
and U4684 (N_4684,N_2846,N_2507);
nor U4685 (N_4685,N_3934,N_3457);
nand U4686 (N_4686,N_3281,N_2007);
or U4687 (N_4687,N_3616,N_3426);
nor U4688 (N_4688,N_2968,N_3720);
nand U4689 (N_4689,N_2299,N_3942);
and U4690 (N_4690,N_2828,N_3785);
or U4691 (N_4691,N_2610,N_3635);
nand U4692 (N_4692,N_3292,N_2719);
nand U4693 (N_4693,N_2225,N_3246);
xnor U4694 (N_4694,N_3398,N_3166);
nand U4695 (N_4695,N_2333,N_2404);
and U4696 (N_4696,N_3440,N_2635);
nor U4697 (N_4697,N_3669,N_2204);
nor U4698 (N_4698,N_3448,N_3598);
and U4699 (N_4699,N_3798,N_3239);
and U4700 (N_4700,N_3401,N_2754);
and U4701 (N_4701,N_3371,N_3392);
nand U4702 (N_4702,N_3941,N_2282);
and U4703 (N_4703,N_3156,N_2355);
nand U4704 (N_4704,N_2108,N_2096);
nand U4705 (N_4705,N_2387,N_3995);
and U4706 (N_4706,N_2154,N_2504);
and U4707 (N_4707,N_3557,N_3809);
nor U4708 (N_4708,N_2695,N_3709);
nand U4709 (N_4709,N_3615,N_2441);
nor U4710 (N_4710,N_2366,N_3693);
or U4711 (N_4711,N_3943,N_3757);
or U4712 (N_4712,N_2063,N_3312);
nand U4713 (N_4713,N_2395,N_3262);
or U4714 (N_4714,N_2214,N_2583);
or U4715 (N_4715,N_2656,N_2135);
nor U4716 (N_4716,N_3025,N_3973);
nand U4717 (N_4717,N_2270,N_2692);
and U4718 (N_4718,N_3126,N_2523);
or U4719 (N_4719,N_2668,N_3680);
nand U4720 (N_4720,N_2051,N_3834);
and U4721 (N_4721,N_3451,N_3066);
nor U4722 (N_4722,N_3311,N_2739);
nor U4723 (N_4723,N_3040,N_2540);
and U4724 (N_4724,N_3954,N_2131);
nand U4725 (N_4725,N_3977,N_3645);
or U4726 (N_4726,N_2745,N_3270);
nand U4727 (N_4727,N_2702,N_2995);
and U4728 (N_4728,N_3271,N_2139);
nor U4729 (N_4729,N_3160,N_3469);
or U4730 (N_4730,N_2448,N_2092);
nand U4731 (N_4731,N_2915,N_2300);
and U4732 (N_4732,N_2332,N_3856);
and U4733 (N_4733,N_2253,N_3287);
nor U4734 (N_4734,N_2554,N_2769);
nand U4735 (N_4735,N_3214,N_3847);
or U4736 (N_4736,N_3079,N_3648);
and U4737 (N_4737,N_2038,N_2857);
nand U4738 (N_4738,N_2738,N_2640);
or U4739 (N_4739,N_2056,N_3192);
nand U4740 (N_4740,N_2370,N_2069);
nor U4741 (N_4741,N_3950,N_2147);
and U4742 (N_4742,N_3052,N_3080);
or U4743 (N_4743,N_3131,N_3893);
nor U4744 (N_4744,N_2880,N_3394);
or U4745 (N_4745,N_2798,N_2545);
nor U4746 (N_4746,N_2761,N_2406);
and U4747 (N_4747,N_2434,N_2442);
or U4748 (N_4748,N_2944,N_2275);
nor U4749 (N_4749,N_2252,N_3596);
nor U4750 (N_4750,N_3562,N_2751);
nand U4751 (N_4751,N_2538,N_3409);
nand U4752 (N_4752,N_3130,N_3332);
nor U4753 (N_4753,N_3265,N_2213);
or U4754 (N_4754,N_2060,N_3929);
nand U4755 (N_4755,N_2029,N_2354);
nand U4756 (N_4756,N_2385,N_2440);
and U4757 (N_4757,N_3897,N_2490);
or U4758 (N_4758,N_2431,N_3609);
nor U4759 (N_4759,N_2353,N_3403);
or U4760 (N_4760,N_3714,N_3797);
and U4761 (N_4761,N_3882,N_2281);
and U4762 (N_4762,N_3269,N_3547);
or U4763 (N_4763,N_3072,N_2582);
nor U4764 (N_4764,N_3029,N_3746);
or U4765 (N_4765,N_3415,N_3990);
nand U4766 (N_4766,N_2908,N_3878);
or U4767 (N_4767,N_3004,N_3012);
nor U4768 (N_4768,N_2103,N_2195);
nor U4769 (N_4769,N_2162,N_2372);
nand U4770 (N_4770,N_3506,N_3120);
nor U4771 (N_4771,N_2054,N_2449);
or U4772 (N_4772,N_2813,N_2206);
nor U4773 (N_4773,N_3589,N_2211);
and U4774 (N_4774,N_2429,N_3620);
nand U4775 (N_4775,N_2260,N_2033);
or U4776 (N_4776,N_2501,N_3569);
nor U4777 (N_4777,N_2955,N_3511);
nor U4778 (N_4778,N_2373,N_2389);
or U4779 (N_4779,N_2464,N_3963);
or U4780 (N_4780,N_2291,N_2142);
or U4781 (N_4781,N_3462,N_2629);
or U4782 (N_4782,N_2851,N_3041);
nand U4783 (N_4783,N_3319,N_3164);
nor U4784 (N_4784,N_2576,N_2192);
nand U4785 (N_4785,N_3642,N_3992);
and U4786 (N_4786,N_3764,N_2533);
or U4787 (N_4787,N_2553,N_3347);
and U4788 (N_4788,N_3610,N_3418);
nand U4789 (N_4789,N_3993,N_3002);
nor U4790 (N_4790,N_3541,N_3032);
nor U4791 (N_4791,N_3961,N_2742);
nand U4792 (N_4792,N_2514,N_2250);
nor U4793 (N_4793,N_3035,N_3370);
nor U4794 (N_4794,N_3205,N_2546);
or U4795 (N_4795,N_3470,N_3259);
nor U4796 (N_4796,N_2352,N_2017);
and U4797 (N_4797,N_3859,N_2529);
and U4798 (N_4798,N_3382,N_2716);
nand U4799 (N_4799,N_3734,N_2169);
and U4800 (N_4800,N_2041,N_3428);
and U4801 (N_4801,N_2159,N_2179);
and U4802 (N_4802,N_2283,N_2130);
nor U4803 (N_4803,N_3091,N_3976);
nor U4804 (N_4804,N_2217,N_3900);
nand U4805 (N_4805,N_2942,N_2383);
nand U4806 (N_4806,N_2887,N_2863);
or U4807 (N_4807,N_3722,N_2643);
xor U4808 (N_4808,N_3135,N_2642);
nor U4809 (N_4809,N_3061,N_2306);
nor U4810 (N_4810,N_3386,N_3579);
nor U4811 (N_4811,N_2972,N_2065);
and U4812 (N_4812,N_3800,N_2457);
nand U4813 (N_4813,N_3391,N_2346);
or U4814 (N_4814,N_3065,N_3026);
and U4815 (N_4815,N_3618,N_3751);
and U4816 (N_4816,N_2055,N_2228);
nor U4817 (N_4817,N_2835,N_2780);
and U4818 (N_4818,N_2838,N_3363);
nand U4819 (N_4819,N_2435,N_2877);
nand U4820 (N_4820,N_2952,N_3224);
nor U4821 (N_4821,N_2367,N_2904);
and U4822 (N_4822,N_2392,N_3232);
nand U4823 (N_4823,N_2898,N_2251);
or U4824 (N_4824,N_2460,N_3901);
nor U4825 (N_4825,N_3502,N_3384);
nand U4826 (N_4826,N_3909,N_2310);
nor U4827 (N_4827,N_2616,N_3862);
nor U4828 (N_4828,N_3520,N_2562);
and U4829 (N_4829,N_2423,N_3090);
or U4830 (N_4830,N_2407,N_3848);
and U4831 (N_4831,N_2117,N_2232);
nor U4832 (N_4832,N_3167,N_2394);
or U4833 (N_4833,N_3219,N_3876);
and U4834 (N_4834,N_3593,N_3772);
nor U4835 (N_4835,N_3507,N_2302);
or U4836 (N_4836,N_3813,N_2685);
or U4837 (N_4837,N_2508,N_3023);
nand U4838 (N_4838,N_2560,N_3213);
nand U4839 (N_4839,N_2519,N_2083);
xor U4840 (N_4840,N_2581,N_3575);
or U4841 (N_4841,N_2104,N_2364);
nor U4842 (N_4842,N_2903,N_3649);
and U4843 (N_4843,N_3931,N_2717);
nand U4844 (N_4844,N_3996,N_2221);
nor U4845 (N_4845,N_3555,N_2037);
or U4846 (N_4846,N_2095,N_3186);
nand U4847 (N_4847,N_3747,N_3339);
nand U4848 (N_4848,N_2324,N_2531);
nor U4849 (N_4849,N_3960,N_2240);
or U4850 (N_4850,N_2196,N_3346);
nand U4851 (N_4851,N_2268,N_3705);
nand U4852 (N_4852,N_3510,N_3420);
nand U4853 (N_4853,N_3647,N_2308);
nand U4854 (N_4854,N_2371,N_2070);
or U4855 (N_4855,N_2974,N_3256);
nor U4856 (N_4856,N_3369,N_3533);
nor U4857 (N_4857,N_2725,N_3351);
nand U4858 (N_4858,N_3686,N_3099);
nand U4859 (N_4859,N_2641,N_3835);
nor U4860 (N_4860,N_3955,N_3612);
nand U4861 (N_4861,N_3340,N_3424);
and U4862 (N_4862,N_2110,N_2419);
and U4863 (N_4863,N_2199,N_3657);
and U4864 (N_4864,N_2983,N_3149);
nand U4865 (N_4865,N_3580,N_3119);
or U4866 (N_4866,N_2925,N_3852);
or U4867 (N_4867,N_2284,N_3650);
nor U4868 (N_4868,N_2358,N_2613);
nand U4869 (N_4869,N_2484,N_3982);
nand U4870 (N_4870,N_2592,N_3838);
or U4871 (N_4871,N_2040,N_3523);
nand U4872 (N_4872,N_3843,N_3845);
or U4873 (N_4873,N_2061,N_3936);
and U4874 (N_4874,N_3868,N_3721);
nor U4875 (N_4875,N_2979,N_3597);
or U4876 (N_4876,N_3899,N_2647);
nor U4877 (N_4877,N_2679,N_2593);
nor U4878 (N_4878,N_2396,N_2351);
nand U4879 (N_4879,N_3193,N_3799);
and U4880 (N_4880,N_3970,N_3879);
and U4881 (N_4881,N_2790,N_3038);
or U4882 (N_4882,N_2630,N_2168);
and U4883 (N_4883,N_3884,N_3336);
nand U4884 (N_4884,N_2479,N_3531);
nand U4885 (N_4885,N_2295,N_2043);
or U4886 (N_4886,N_3771,N_3249);
nand U4887 (N_4887,N_2200,N_3740);
nor U4888 (N_4888,N_3291,N_3986);
or U4889 (N_4889,N_2005,N_3568);
nor U4890 (N_4890,N_2261,N_3086);
nor U4891 (N_4891,N_3148,N_3421);
nand U4892 (N_4892,N_2345,N_3983);
nor U4893 (N_4893,N_3331,N_3515);
nor U4894 (N_4894,N_3717,N_2572);
nand U4895 (N_4895,N_2730,N_3551);
or U4896 (N_4896,N_2705,N_2981);
nor U4897 (N_4897,N_3257,N_2499);
nor U4898 (N_4898,N_2758,N_3804);
nand U4899 (N_4899,N_2151,N_3892);
and U4900 (N_4900,N_3028,N_2815);
or U4901 (N_4901,N_2167,N_3633);
or U4902 (N_4902,N_2176,N_2814);
and U4903 (N_4903,N_2086,N_2948);
or U4904 (N_4904,N_3027,N_2356);
and U4905 (N_4905,N_3972,N_3622);
and U4906 (N_4906,N_2722,N_2946);
or U4907 (N_4907,N_2034,N_3865);
and U4908 (N_4908,N_2935,N_3162);
nor U4909 (N_4909,N_3277,N_2243);
nor U4910 (N_4910,N_2209,N_2776);
nand U4911 (N_4911,N_3293,N_2481);
or U4912 (N_4912,N_3118,N_2003);
or U4913 (N_4913,N_3362,N_2152);
and U4914 (N_4914,N_3991,N_2349);
or U4915 (N_4915,N_3491,N_3704);
or U4916 (N_4916,N_2272,N_3043);
or U4917 (N_4917,N_3984,N_2458);
or U4918 (N_4918,N_2712,N_3443);
nand U4919 (N_4919,N_2516,N_3182);
nor U4920 (N_4920,N_3806,N_3003);
or U4921 (N_4921,N_3042,N_3783);
nor U4922 (N_4922,N_2690,N_2205);
nor U4923 (N_4923,N_3236,N_3087);
nand U4924 (N_4924,N_3629,N_2895);
nor U4925 (N_4925,N_2015,N_2706);
or U4926 (N_4926,N_3446,N_2347);
or U4927 (N_4927,N_2424,N_2911);
nor U4928 (N_4928,N_3644,N_2126);
and U4929 (N_4929,N_2735,N_2810);
nor U4930 (N_4930,N_2849,N_3839);
or U4931 (N_4931,N_3318,N_2315);
and U4932 (N_4932,N_2094,N_3666);
nand U4933 (N_4933,N_3957,N_2910);
nand U4934 (N_4934,N_2743,N_2867);
or U4935 (N_4935,N_3527,N_2059);
and U4936 (N_4936,N_2732,N_2786);
or U4937 (N_4937,N_3302,N_3831);
or U4938 (N_4938,N_2933,N_2721);
or U4939 (N_4939,N_2414,N_3341);
or U4940 (N_4940,N_3626,N_3141);
nand U4941 (N_4941,N_2438,N_3781);
and U4942 (N_4942,N_3128,N_2436);
nand U4943 (N_4943,N_3643,N_2318);
or U4944 (N_4944,N_3744,N_2173);
and U4945 (N_4945,N_2127,N_2627);
nor U4946 (N_4946,N_2693,N_2264);
or U4947 (N_4947,N_3971,N_3810);
and U4948 (N_4948,N_3952,N_2080);
xnor U4949 (N_4949,N_3724,N_3248);
or U4950 (N_4950,N_3702,N_3145);
nand U4951 (N_4951,N_3283,N_2181);
or U4952 (N_4952,N_2402,N_3378);
nand U4953 (N_4953,N_3267,N_3812);
nor U4954 (N_4954,N_3105,N_3599);
or U4955 (N_4955,N_3299,N_3707);
and U4956 (N_4956,N_2905,N_2530);
nand U4957 (N_4957,N_3324,N_2146);
nor U4958 (N_4958,N_3716,N_2177);
or U4959 (N_4959,N_2362,N_3240);
nor U4960 (N_4960,N_2035,N_3854);
nand U4961 (N_4961,N_3660,N_2663);
and U4962 (N_4962,N_3286,N_3247);
nor U4963 (N_4963,N_3758,N_3063);
nand U4964 (N_4964,N_3036,N_3229);
or U4965 (N_4965,N_2336,N_2655);
nand U4966 (N_4966,N_3432,N_3218);
nand U4967 (N_4967,N_2764,N_2775);
nand U4968 (N_4968,N_3190,N_2563);
or U4969 (N_4969,N_3320,N_2319);
nand U4970 (N_4970,N_3735,N_2184);
and U4971 (N_4971,N_2247,N_3039);
nor U4972 (N_4972,N_2273,N_3525);
nor U4973 (N_4973,N_3408,N_2174);
xnor U4974 (N_4974,N_3344,N_3114);
nand U4975 (N_4975,N_2893,N_2475);
nor U4976 (N_4976,N_3682,N_2588);
nand U4977 (N_4977,N_2701,N_3532);
nand U4978 (N_4978,N_2422,N_3151);
nor U4979 (N_4979,N_3826,N_3412);
and U4980 (N_4980,N_3129,N_3958);
nor U4981 (N_4981,N_3832,N_2718);
nand U4982 (N_4982,N_2753,N_3526);
xnor U4983 (N_4983,N_2482,N_2669);
and U4984 (N_4984,N_2280,N_3827);
nor U4985 (N_4985,N_2420,N_3359);
and U4986 (N_4986,N_3326,N_2140);
nor U4987 (N_4987,N_2934,N_3661);
nor U4988 (N_4988,N_3902,N_3886);
nand U4989 (N_4989,N_3111,N_2976);
nor U4990 (N_4990,N_3010,N_3890);
nand U4991 (N_4991,N_2075,N_2868);
nor U4992 (N_4992,N_2105,N_2288);
or U4993 (N_4993,N_3861,N_2343);
nand U4994 (N_4994,N_3793,N_2794);
nand U4995 (N_4995,N_2547,N_3475);
and U4996 (N_4996,N_2210,N_2222);
and U4997 (N_4997,N_3427,N_2189);
nor U4998 (N_4998,N_3549,N_3728);
or U4999 (N_4999,N_2443,N_3811);
and U5000 (N_5000,N_3310,N_3457);
nand U5001 (N_5001,N_3288,N_3093);
and U5002 (N_5002,N_3118,N_2390);
nor U5003 (N_5003,N_3103,N_2982);
nor U5004 (N_5004,N_3416,N_2901);
nor U5005 (N_5005,N_3196,N_3847);
or U5006 (N_5006,N_3542,N_3042);
or U5007 (N_5007,N_2105,N_3327);
nor U5008 (N_5008,N_3641,N_2497);
nor U5009 (N_5009,N_2024,N_3933);
or U5010 (N_5010,N_3861,N_2268);
nand U5011 (N_5011,N_3509,N_3722);
and U5012 (N_5012,N_3613,N_2350);
nor U5013 (N_5013,N_2816,N_2305);
or U5014 (N_5014,N_2645,N_2457);
nor U5015 (N_5015,N_3312,N_2703);
or U5016 (N_5016,N_2685,N_3306);
nor U5017 (N_5017,N_2815,N_2839);
nand U5018 (N_5018,N_2018,N_3349);
and U5019 (N_5019,N_3730,N_3169);
nand U5020 (N_5020,N_3979,N_3998);
or U5021 (N_5021,N_3483,N_2810);
and U5022 (N_5022,N_3782,N_3964);
nor U5023 (N_5023,N_2873,N_3976);
xor U5024 (N_5024,N_2365,N_2809);
nand U5025 (N_5025,N_3537,N_3053);
nand U5026 (N_5026,N_3354,N_3957);
nand U5027 (N_5027,N_2061,N_3797);
and U5028 (N_5028,N_3403,N_2670);
or U5029 (N_5029,N_3755,N_2773);
or U5030 (N_5030,N_3611,N_3995);
nand U5031 (N_5031,N_3233,N_3815);
and U5032 (N_5032,N_2119,N_3307);
or U5033 (N_5033,N_2625,N_3164);
nor U5034 (N_5034,N_3730,N_3645);
and U5035 (N_5035,N_3795,N_2577);
and U5036 (N_5036,N_2396,N_2885);
nand U5037 (N_5037,N_2699,N_2506);
nor U5038 (N_5038,N_2764,N_2118);
nand U5039 (N_5039,N_3599,N_2276);
nor U5040 (N_5040,N_2664,N_3751);
nor U5041 (N_5041,N_3977,N_2431);
and U5042 (N_5042,N_2844,N_2050);
and U5043 (N_5043,N_2066,N_2999);
nor U5044 (N_5044,N_3322,N_2462);
nand U5045 (N_5045,N_3585,N_2354);
or U5046 (N_5046,N_2784,N_2160);
or U5047 (N_5047,N_2724,N_2475);
nand U5048 (N_5048,N_2330,N_2255);
nand U5049 (N_5049,N_3764,N_2837);
and U5050 (N_5050,N_2543,N_3799);
and U5051 (N_5051,N_3917,N_3583);
nand U5052 (N_5052,N_3334,N_2397);
nor U5053 (N_5053,N_2788,N_2962);
or U5054 (N_5054,N_2151,N_3578);
nand U5055 (N_5055,N_2638,N_3032);
nor U5056 (N_5056,N_3383,N_3956);
or U5057 (N_5057,N_3643,N_3853);
or U5058 (N_5058,N_2561,N_2608);
nand U5059 (N_5059,N_2588,N_2804);
or U5060 (N_5060,N_3450,N_2312);
or U5061 (N_5061,N_2928,N_3668);
nor U5062 (N_5062,N_2152,N_3572);
nand U5063 (N_5063,N_3155,N_2855);
and U5064 (N_5064,N_3706,N_2302);
nand U5065 (N_5065,N_3126,N_2874);
nand U5066 (N_5066,N_3780,N_2374);
or U5067 (N_5067,N_2734,N_2513);
nor U5068 (N_5068,N_2369,N_3084);
nor U5069 (N_5069,N_3289,N_2944);
or U5070 (N_5070,N_3067,N_2369);
and U5071 (N_5071,N_2913,N_3498);
or U5072 (N_5072,N_3574,N_2619);
or U5073 (N_5073,N_3219,N_2916);
and U5074 (N_5074,N_3643,N_3359);
nor U5075 (N_5075,N_2689,N_3054);
nand U5076 (N_5076,N_2350,N_3773);
and U5077 (N_5077,N_2429,N_2495);
nor U5078 (N_5078,N_3281,N_3901);
and U5079 (N_5079,N_2723,N_3978);
or U5080 (N_5080,N_3366,N_3657);
and U5081 (N_5081,N_2053,N_3351);
and U5082 (N_5082,N_3984,N_3252);
nand U5083 (N_5083,N_2104,N_2175);
nor U5084 (N_5084,N_2580,N_2722);
and U5085 (N_5085,N_2768,N_3526);
nor U5086 (N_5086,N_2544,N_2401);
nor U5087 (N_5087,N_3359,N_3540);
xor U5088 (N_5088,N_2629,N_3245);
or U5089 (N_5089,N_2293,N_3810);
nor U5090 (N_5090,N_2459,N_3087);
or U5091 (N_5091,N_2999,N_2455);
or U5092 (N_5092,N_2707,N_2906);
nor U5093 (N_5093,N_2379,N_3727);
or U5094 (N_5094,N_3755,N_2670);
and U5095 (N_5095,N_3827,N_3842);
and U5096 (N_5096,N_2357,N_3803);
nand U5097 (N_5097,N_2021,N_3515);
or U5098 (N_5098,N_3196,N_2972);
nand U5099 (N_5099,N_3218,N_2781);
and U5100 (N_5100,N_3816,N_3288);
or U5101 (N_5101,N_3838,N_3580);
or U5102 (N_5102,N_3530,N_3359);
nand U5103 (N_5103,N_2169,N_3701);
nand U5104 (N_5104,N_2608,N_2252);
or U5105 (N_5105,N_3426,N_3290);
nor U5106 (N_5106,N_3928,N_2644);
nand U5107 (N_5107,N_3173,N_2447);
or U5108 (N_5108,N_2618,N_3320);
nand U5109 (N_5109,N_2378,N_3244);
nand U5110 (N_5110,N_3063,N_3303);
or U5111 (N_5111,N_3727,N_3635);
xor U5112 (N_5112,N_2421,N_3213);
or U5113 (N_5113,N_3879,N_2686);
xnor U5114 (N_5114,N_3786,N_3342);
and U5115 (N_5115,N_3239,N_2203);
nor U5116 (N_5116,N_3076,N_3916);
nand U5117 (N_5117,N_3227,N_3595);
and U5118 (N_5118,N_3993,N_2316);
and U5119 (N_5119,N_2765,N_2720);
or U5120 (N_5120,N_3820,N_3921);
or U5121 (N_5121,N_2749,N_2004);
or U5122 (N_5122,N_2521,N_2636);
and U5123 (N_5123,N_2981,N_3787);
and U5124 (N_5124,N_3521,N_2294);
and U5125 (N_5125,N_2586,N_2666);
or U5126 (N_5126,N_2507,N_3198);
nor U5127 (N_5127,N_3612,N_3140);
nand U5128 (N_5128,N_3054,N_2134);
nor U5129 (N_5129,N_2768,N_3608);
nor U5130 (N_5130,N_2216,N_2009);
nand U5131 (N_5131,N_2591,N_3672);
or U5132 (N_5132,N_2021,N_2037);
nor U5133 (N_5133,N_2119,N_3226);
or U5134 (N_5134,N_3333,N_3941);
nand U5135 (N_5135,N_3444,N_3354);
nand U5136 (N_5136,N_3936,N_3552);
and U5137 (N_5137,N_2332,N_3324);
and U5138 (N_5138,N_2656,N_3533);
or U5139 (N_5139,N_2110,N_2249);
or U5140 (N_5140,N_3673,N_2472);
and U5141 (N_5141,N_2562,N_2766);
nand U5142 (N_5142,N_3158,N_2716);
nor U5143 (N_5143,N_3838,N_2412);
nor U5144 (N_5144,N_3355,N_2052);
nor U5145 (N_5145,N_2876,N_3837);
or U5146 (N_5146,N_2069,N_3057);
nor U5147 (N_5147,N_2629,N_2375);
nor U5148 (N_5148,N_2786,N_2351);
or U5149 (N_5149,N_3316,N_3951);
or U5150 (N_5150,N_2163,N_3236);
and U5151 (N_5151,N_3016,N_3209);
or U5152 (N_5152,N_2399,N_2091);
or U5153 (N_5153,N_2545,N_2955);
and U5154 (N_5154,N_3681,N_2815);
nor U5155 (N_5155,N_2372,N_2481);
or U5156 (N_5156,N_2213,N_3244);
nor U5157 (N_5157,N_2650,N_2096);
and U5158 (N_5158,N_3806,N_3159);
nand U5159 (N_5159,N_2020,N_3783);
and U5160 (N_5160,N_3937,N_3696);
and U5161 (N_5161,N_2026,N_3536);
nor U5162 (N_5162,N_2744,N_2256);
nor U5163 (N_5163,N_2934,N_2653);
or U5164 (N_5164,N_2264,N_3712);
or U5165 (N_5165,N_3507,N_2613);
or U5166 (N_5166,N_2033,N_2086);
nand U5167 (N_5167,N_3117,N_3129);
and U5168 (N_5168,N_2610,N_2941);
or U5169 (N_5169,N_3158,N_3878);
nand U5170 (N_5170,N_3699,N_2920);
and U5171 (N_5171,N_3393,N_2378);
nand U5172 (N_5172,N_2439,N_3763);
nand U5173 (N_5173,N_2196,N_2462);
and U5174 (N_5174,N_2419,N_2524);
and U5175 (N_5175,N_2579,N_3396);
or U5176 (N_5176,N_3934,N_3012);
nand U5177 (N_5177,N_3023,N_3432);
or U5178 (N_5178,N_2591,N_2294);
nor U5179 (N_5179,N_2871,N_3429);
and U5180 (N_5180,N_2638,N_3140);
xnor U5181 (N_5181,N_2745,N_2459);
and U5182 (N_5182,N_2051,N_3486);
and U5183 (N_5183,N_3485,N_3823);
nand U5184 (N_5184,N_2120,N_2450);
nand U5185 (N_5185,N_3293,N_3839);
or U5186 (N_5186,N_2671,N_3816);
and U5187 (N_5187,N_3239,N_3892);
or U5188 (N_5188,N_3778,N_2731);
and U5189 (N_5189,N_2411,N_3949);
nand U5190 (N_5190,N_2633,N_3452);
and U5191 (N_5191,N_2425,N_2094);
nor U5192 (N_5192,N_3675,N_2417);
or U5193 (N_5193,N_3367,N_2585);
and U5194 (N_5194,N_3419,N_3617);
and U5195 (N_5195,N_3376,N_3960);
nand U5196 (N_5196,N_3535,N_3048);
nand U5197 (N_5197,N_2900,N_3401);
and U5198 (N_5198,N_3094,N_3138);
or U5199 (N_5199,N_2260,N_2577);
or U5200 (N_5200,N_2228,N_2291);
nand U5201 (N_5201,N_2545,N_3736);
nand U5202 (N_5202,N_3559,N_2844);
and U5203 (N_5203,N_3656,N_2652);
or U5204 (N_5204,N_3510,N_3435);
and U5205 (N_5205,N_2975,N_2849);
nand U5206 (N_5206,N_3841,N_2662);
or U5207 (N_5207,N_3707,N_2961);
or U5208 (N_5208,N_3005,N_3650);
nand U5209 (N_5209,N_3755,N_2446);
nand U5210 (N_5210,N_2617,N_2932);
nor U5211 (N_5211,N_3653,N_3111);
nor U5212 (N_5212,N_2920,N_3408);
and U5213 (N_5213,N_2132,N_3288);
and U5214 (N_5214,N_3086,N_3449);
or U5215 (N_5215,N_3453,N_2348);
and U5216 (N_5216,N_2940,N_2846);
nand U5217 (N_5217,N_2017,N_2054);
nand U5218 (N_5218,N_2059,N_2159);
and U5219 (N_5219,N_2852,N_2183);
or U5220 (N_5220,N_2680,N_2854);
nor U5221 (N_5221,N_2780,N_2276);
nand U5222 (N_5222,N_3663,N_3744);
nor U5223 (N_5223,N_2753,N_2975);
nor U5224 (N_5224,N_3186,N_2354);
nand U5225 (N_5225,N_2520,N_2101);
or U5226 (N_5226,N_2039,N_2612);
and U5227 (N_5227,N_3392,N_3527);
xnor U5228 (N_5228,N_2929,N_2646);
nand U5229 (N_5229,N_2405,N_2466);
and U5230 (N_5230,N_3438,N_3065);
and U5231 (N_5231,N_2492,N_3643);
or U5232 (N_5232,N_3332,N_3292);
nand U5233 (N_5233,N_2953,N_3712);
nor U5234 (N_5234,N_3471,N_3507);
nand U5235 (N_5235,N_2196,N_3065);
and U5236 (N_5236,N_2986,N_3220);
nor U5237 (N_5237,N_2996,N_2041);
and U5238 (N_5238,N_3750,N_3305);
nor U5239 (N_5239,N_3066,N_2351);
and U5240 (N_5240,N_2543,N_2407);
and U5241 (N_5241,N_3420,N_3457);
and U5242 (N_5242,N_3138,N_3146);
xnor U5243 (N_5243,N_3534,N_2877);
nor U5244 (N_5244,N_2217,N_2140);
nand U5245 (N_5245,N_2701,N_3461);
or U5246 (N_5246,N_2867,N_2705);
and U5247 (N_5247,N_3930,N_3684);
nor U5248 (N_5248,N_3004,N_3082);
xnor U5249 (N_5249,N_3846,N_3028);
or U5250 (N_5250,N_3414,N_3528);
nand U5251 (N_5251,N_2389,N_3060);
nand U5252 (N_5252,N_2119,N_3296);
nand U5253 (N_5253,N_2840,N_2072);
xor U5254 (N_5254,N_2805,N_2271);
and U5255 (N_5255,N_2691,N_3269);
or U5256 (N_5256,N_3364,N_2863);
nor U5257 (N_5257,N_3988,N_2547);
and U5258 (N_5258,N_2840,N_3205);
nor U5259 (N_5259,N_3878,N_3143);
nor U5260 (N_5260,N_2125,N_2222);
nor U5261 (N_5261,N_2429,N_3670);
xnor U5262 (N_5262,N_3726,N_3866);
or U5263 (N_5263,N_2770,N_3401);
and U5264 (N_5264,N_3190,N_3585);
nor U5265 (N_5265,N_3077,N_3955);
and U5266 (N_5266,N_2447,N_2580);
xor U5267 (N_5267,N_2143,N_2019);
nand U5268 (N_5268,N_2228,N_2924);
and U5269 (N_5269,N_3872,N_3335);
nand U5270 (N_5270,N_2627,N_2688);
nor U5271 (N_5271,N_3505,N_2305);
and U5272 (N_5272,N_3622,N_3339);
nand U5273 (N_5273,N_2139,N_2324);
or U5274 (N_5274,N_3707,N_2206);
and U5275 (N_5275,N_2507,N_2278);
nor U5276 (N_5276,N_2836,N_2337);
and U5277 (N_5277,N_3709,N_3319);
nor U5278 (N_5278,N_3594,N_3827);
or U5279 (N_5279,N_3942,N_3224);
and U5280 (N_5280,N_2169,N_3429);
nor U5281 (N_5281,N_2285,N_3094);
and U5282 (N_5282,N_2837,N_2899);
and U5283 (N_5283,N_3435,N_3911);
nor U5284 (N_5284,N_2422,N_3457);
and U5285 (N_5285,N_2614,N_3378);
nand U5286 (N_5286,N_3792,N_2888);
or U5287 (N_5287,N_2674,N_2391);
nor U5288 (N_5288,N_3146,N_2017);
nor U5289 (N_5289,N_2917,N_3578);
nor U5290 (N_5290,N_3217,N_2690);
or U5291 (N_5291,N_2584,N_2575);
nand U5292 (N_5292,N_3787,N_3703);
nor U5293 (N_5293,N_2500,N_3154);
and U5294 (N_5294,N_3334,N_2681);
nor U5295 (N_5295,N_2722,N_2704);
nor U5296 (N_5296,N_2798,N_3543);
and U5297 (N_5297,N_3878,N_2323);
nor U5298 (N_5298,N_2461,N_2472);
and U5299 (N_5299,N_2211,N_2226);
nor U5300 (N_5300,N_2382,N_2202);
and U5301 (N_5301,N_2991,N_2866);
or U5302 (N_5302,N_2962,N_3320);
nand U5303 (N_5303,N_2837,N_2442);
and U5304 (N_5304,N_3578,N_2527);
and U5305 (N_5305,N_3963,N_3421);
nor U5306 (N_5306,N_3570,N_2811);
or U5307 (N_5307,N_3015,N_2376);
or U5308 (N_5308,N_3352,N_2673);
or U5309 (N_5309,N_2496,N_3521);
nand U5310 (N_5310,N_3135,N_3960);
and U5311 (N_5311,N_2441,N_3077);
nand U5312 (N_5312,N_2981,N_3188);
nor U5313 (N_5313,N_3188,N_3786);
or U5314 (N_5314,N_3956,N_2963);
nor U5315 (N_5315,N_2676,N_2331);
nand U5316 (N_5316,N_3920,N_3236);
or U5317 (N_5317,N_2259,N_2482);
and U5318 (N_5318,N_3143,N_2861);
or U5319 (N_5319,N_2749,N_3972);
nand U5320 (N_5320,N_2542,N_2942);
nor U5321 (N_5321,N_2917,N_2287);
nor U5322 (N_5322,N_3784,N_3393);
nand U5323 (N_5323,N_2614,N_2891);
nand U5324 (N_5324,N_2569,N_3765);
or U5325 (N_5325,N_3078,N_2043);
and U5326 (N_5326,N_2860,N_2834);
nand U5327 (N_5327,N_3880,N_2577);
nand U5328 (N_5328,N_3798,N_2496);
nor U5329 (N_5329,N_2628,N_3761);
and U5330 (N_5330,N_2883,N_2642);
and U5331 (N_5331,N_2371,N_3850);
or U5332 (N_5332,N_3124,N_2637);
and U5333 (N_5333,N_2029,N_2435);
nand U5334 (N_5334,N_3109,N_3103);
or U5335 (N_5335,N_2495,N_3734);
or U5336 (N_5336,N_3210,N_3867);
nor U5337 (N_5337,N_2121,N_3525);
nor U5338 (N_5338,N_3205,N_3016);
and U5339 (N_5339,N_2116,N_2294);
nor U5340 (N_5340,N_3259,N_3870);
nor U5341 (N_5341,N_3015,N_3151);
or U5342 (N_5342,N_3568,N_2672);
nand U5343 (N_5343,N_2382,N_3485);
nor U5344 (N_5344,N_3402,N_3456);
and U5345 (N_5345,N_3141,N_2102);
and U5346 (N_5346,N_3918,N_2513);
nand U5347 (N_5347,N_2486,N_3629);
nand U5348 (N_5348,N_2078,N_2010);
or U5349 (N_5349,N_2211,N_3278);
nand U5350 (N_5350,N_2145,N_2082);
xor U5351 (N_5351,N_3564,N_2658);
nor U5352 (N_5352,N_3725,N_2442);
and U5353 (N_5353,N_3404,N_2784);
nor U5354 (N_5354,N_2567,N_3638);
or U5355 (N_5355,N_3506,N_2020);
and U5356 (N_5356,N_3256,N_3197);
and U5357 (N_5357,N_3613,N_3446);
nand U5358 (N_5358,N_3272,N_2833);
or U5359 (N_5359,N_3665,N_2902);
nor U5360 (N_5360,N_2494,N_3604);
or U5361 (N_5361,N_2936,N_2484);
nand U5362 (N_5362,N_3977,N_2741);
and U5363 (N_5363,N_3542,N_2295);
nor U5364 (N_5364,N_2742,N_3684);
or U5365 (N_5365,N_3839,N_3490);
or U5366 (N_5366,N_2973,N_2924);
or U5367 (N_5367,N_2659,N_2202);
nor U5368 (N_5368,N_2936,N_3334);
or U5369 (N_5369,N_3524,N_3682);
nand U5370 (N_5370,N_3504,N_3484);
nand U5371 (N_5371,N_3570,N_3039);
nand U5372 (N_5372,N_2970,N_3890);
nor U5373 (N_5373,N_3161,N_2507);
nand U5374 (N_5374,N_2603,N_3600);
or U5375 (N_5375,N_2947,N_3614);
and U5376 (N_5376,N_2680,N_2495);
nand U5377 (N_5377,N_2791,N_2429);
and U5378 (N_5378,N_2001,N_2932);
or U5379 (N_5379,N_2419,N_2107);
and U5380 (N_5380,N_2005,N_2545);
xor U5381 (N_5381,N_2669,N_2170);
or U5382 (N_5382,N_2344,N_2156);
nand U5383 (N_5383,N_3945,N_3857);
or U5384 (N_5384,N_2923,N_3574);
or U5385 (N_5385,N_3727,N_3937);
and U5386 (N_5386,N_3295,N_2484);
and U5387 (N_5387,N_3474,N_3304);
and U5388 (N_5388,N_2864,N_3875);
nand U5389 (N_5389,N_2160,N_3198);
nand U5390 (N_5390,N_3505,N_2327);
or U5391 (N_5391,N_2389,N_2572);
nand U5392 (N_5392,N_3989,N_3031);
or U5393 (N_5393,N_3510,N_2025);
nand U5394 (N_5394,N_2581,N_2006);
or U5395 (N_5395,N_3790,N_3051);
and U5396 (N_5396,N_3286,N_3936);
nor U5397 (N_5397,N_2108,N_3263);
and U5398 (N_5398,N_3924,N_3457);
and U5399 (N_5399,N_3564,N_2421);
nand U5400 (N_5400,N_3016,N_2296);
or U5401 (N_5401,N_3692,N_2202);
and U5402 (N_5402,N_3540,N_3175);
nand U5403 (N_5403,N_3939,N_3541);
and U5404 (N_5404,N_3360,N_3786);
and U5405 (N_5405,N_2746,N_2092);
or U5406 (N_5406,N_3685,N_3545);
nand U5407 (N_5407,N_2696,N_2611);
nand U5408 (N_5408,N_2683,N_2666);
and U5409 (N_5409,N_3462,N_2460);
nor U5410 (N_5410,N_2435,N_2756);
or U5411 (N_5411,N_3600,N_2961);
nor U5412 (N_5412,N_3743,N_3360);
nand U5413 (N_5413,N_3126,N_2611);
or U5414 (N_5414,N_2121,N_3802);
nand U5415 (N_5415,N_3992,N_2353);
and U5416 (N_5416,N_3095,N_2307);
or U5417 (N_5417,N_3360,N_2482);
nand U5418 (N_5418,N_2958,N_3715);
nor U5419 (N_5419,N_3291,N_2150);
or U5420 (N_5420,N_2615,N_2139);
and U5421 (N_5421,N_2620,N_2361);
nand U5422 (N_5422,N_2669,N_2273);
nor U5423 (N_5423,N_3751,N_3286);
and U5424 (N_5424,N_2032,N_3033);
or U5425 (N_5425,N_2128,N_2421);
nor U5426 (N_5426,N_3011,N_2391);
and U5427 (N_5427,N_3008,N_3051);
nand U5428 (N_5428,N_2601,N_3986);
or U5429 (N_5429,N_3817,N_3614);
or U5430 (N_5430,N_3464,N_3871);
and U5431 (N_5431,N_3927,N_2192);
nor U5432 (N_5432,N_2828,N_3503);
nor U5433 (N_5433,N_2413,N_3448);
nor U5434 (N_5434,N_2287,N_2939);
and U5435 (N_5435,N_3347,N_2527);
nor U5436 (N_5436,N_2567,N_3236);
and U5437 (N_5437,N_2179,N_2823);
nor U5438 (N_5438,N_3552,N_3581);
or U5439 (N_5439,N_3834,N_2653);
or U5440 (N_5440,N_3642,N_2192);
nor U5441 (N_5441,N_3548,N_2165);
nand U5442 (N_5442,N_3879,N_2950);
and U5443 (N_5443,N_2853,N_3752);
nand U5444 (N_5444,N_2251,N_3414);
or U5445 (N_5445,N_3459,N_3111);
or U5446 (N_5446,N_2560,N_3132);
nor U5447 (N_5447,N_2104,N_3888);
nand U5448 (N_5448,N_2737,N_2029);
and U5449 (N_5449,N_3441,N_2857);
or U5450 (N_5450,N_3697,N_2148);
nor U5451 (N_5451,N_2757,N_2725);
or U5452 (N_5452,N_2011,N_2825);
nor U5453 (N_5453,N_3369,N_3675);
nor U5454 (N_5454,N_2680,N_3355);
or U5455 (N_5455,N_2823,N_2789);
and U5456 (N_5456,N_2096,N_3181);
nor U5457 (N_5457,N_2628,N_2422);
or U5458 (N_5458,N_2417,N_2296);
nor U5459 (N_5459,N_2150,N_2626);
nand U5460 (N_5460,N_2911,N_3909);
nand U5461 (N_5461,N_3708,N_2180);
or U5462 (N_5462,N_2530,N_2769);
or U5463 (N_5463,N_3717,N_3162);
nor U5464 (N_5464,N_3811,N_3265);
and U5465 (N_5465,N_2947,N_3062);
and U5466 (N_5466,N_3167,N_2630);
and U5467 (N_5467,N_2228,N_3194);
and U5468 (N_5468,N_2241,N_3768);
nor U5469 (N_5469,N_3485,N_2215);
nor U5470 (N_5470,N_2960,N_3661);
nand U5471 (N_5471,N_2166,N_3296);
and U5472 (N_5472,N_3988,N_2284);
or U5473 (N_5473,N_2157,N_2807);
nand U5474 (N_5474,N_3457,N_3274);
nand U5475 (N_5475,N_3391,N_3244);
nor U5476 (N_5476,N_2624,N_3456);
or U5477 (N_5477,N_2331,N_2162);
and U5478 (N_5478,N_3457,N_2618);
and U5479 (N_5479,N_2377,N_2075);
or U5480 (N_5480,N_3627,N_3278);
or U5481 (N_5481,N_2558,N_2699);
nor U5482 (N_5482,N_3310,N_3758);
xor U5483 (N_5483,N_2616,N_3772);
or U5484 (N_5484,N_3581,N_2256);
nor U5485 (N_5485,N_2493,N_2063);
nand U5486 (N_5486,N_2934,N_3714);
nand U5487 (N_5487,N_2110,N_2388);
nor U5488 (N_5488,N_3256,N_3339);
or U5489 (N_5489,N_2715,N_3304);
nand U5490 (N_5490,N_3640,N_3161);
and U5491 (N_5491,N_2882,N_3042);
nand U5492 (N_5492,N_3895,N_2469);
nand U5493 (N_5493,N_3029,N_2841);
nor U5494 (N_5494,N_3000,N_2415);
and U5495 (N_5495,N_3665,N_2433);
or U5496 (N_5496,N_2607,N_3939);
nor U5497 (N_5497,N_2455,N_3816);
nor U5498 (N_5498,N_3988,N_3644);
nand U5499 (N_5499,N_3343,N_3650);
nor U5500 (N_5500,N_3295,N_2480);
and U5501 (N_5501,N_3800,N_3402);
and U5502 (N_5502,N_2411,N_3429);
or U5503 (N_5503,N_2598,N_2032);
nor U5504 (N_5504,N_2796,N_2937);
and U5505 (N_5505,N_2689,N_2539);
nor U5506 (N_5506,N_2237,N_3138);
nand U5507 (N_5507,N_3722,N_2435);
nand U5508 (N_5508,N_2974,N_2619);
and U5509 (N_5509,N_3405,N_3860);
and U5510 (N_5510,N_3207,N_2965);
or U5511 (N_5511,N_3466,N_3999);
nor U5512 (N_5512,N_2770,N_2865);
and U5513 (N_5513,N_3384,N_2987);
or U5514 (N_5514,N_3881,N_3903);
nand U5515 (N_5515,N_2795,N_3712);
and U5516 (N_5516,N_2577,N_3135);
nor U5517 (N_5517,N_3120,N_2184);
nand U5518 (N_5518,N_2273,N_2129);
nand U5519 (N_5519,N_3852,N_2348);
and U5520 (N_5520,N_2107,N_3667);
and U5521 (N_5521,N_3524,N_2427);
nor U5522 (N_5522,N_2352,N_3807);
nor U5523 (N_5523,N_3478,N_3547);
or U5524 (N_5524,N_2027,N_3057);
nor U5525 (N_5525,N_3055,N_3556);
or U5526 (N_5526,N_3071,N_3135);
nor U5527 (N_5527,N_3371,N_2858);
nand U5528 (N_5528,N_2524,N_3960);
nand U5529 (N_5529,N_3095,N_2327);
and U5530 (N_5530,N_3067,N_2785);
nor U5531 (N_5531,N_2841,N_3173);
and U5532 (N_5532,N_2121,N_3029);
or U5533 (N_5533,N_3947,N_2560);
or U5534 (N_5534,N_2225,N_2522);
nor U5535 (N_5535,N_3965,N_2107);
nor U5536 (N_5536,N_2203,N_3449);
and U5537 (N_5537,N_2212,N_3242);
and U5538 (N_5538,N_3195,N_2063);
or U5539 (N_5539,N_2704,N_2477);
or U5540 (N_5540,N_3187,N_3030);
nand U5541 (N_5541,N_2169,N_2954);
nor U5542 (N_5542,N_2488,N_3521);
nand U5543 (N_5543,N_2907,N_2960);
and U5544 (N_5544,N_2780,N_3315);
nand U5545 (N_5545,N_2303,N_2484);
nor U5546 (N_5546,N_2238,N_3917);
nor U5547 (N_5547,N_3522,N_3721);
nand U5548 (N_5548,N_2433,N_3841);
nand U5549 (N_5549,N_2061,N_3748);
or U5550 (N_5550,N_2244,N_2818);
nand U5551 (N_5551,N_3849,N_2137);
nand U5552 (N_5552,N_3787,N_2427);
or U5553 (N_5553,N_2353,N_3019);
nor U5554 (N_5554,N_3606,N_2321);
and U5555 (N_5555,N_2710,N_3853);
nor U5556 (N_5556,N_2456,N_2809);
nand U5557 (N_5557,N_2632,N_3085);
or U5558 (N_5558,N_3010,N_3966);
and U5559 (N_5559,N_2806,N_2943);
or U5560 (N_5560,N_3504,N_3496);
nand U5561 (N_5561,N_3090,N_3899);
nand U5562 (N_5562,N_3636,N_3764);
xnor U5563 (N_5563,N_2397,N_3848);
and U5564 (N_5564,N_2418,N_3580);
and U5565 (N_5565,N_2372,N_3014);
and U5566 (N_5566,N_2932,N_2131);
nor U5567 (N_5567,N_3813,N_3815);
nand U5568 (N_5568,N_2467,N_2681);
and U5569 (N_5569,N_2843,N_2195);
and U5570 (N_5570,N_3430,N_2839);
and U5571 (N_5571,N_2911,N_3695);
nor U5572 (N_5572,N_3484,N_2636);
or U5573 (N_5573,N_2635,N_2670);
and U5574 (N_5574,N_2405,N_2591);
and U5575 (N_5575,N_3797,N_3536);
nand U5576 (N_5576,N_2014,N_2957);
nand U5577 (N_5577,N_2344,N_3949);
and U5578 (N_5578,N_3440,N_3266);
or U5579 (N_5579,N_2341,N_3945);
nor U5580 (N_5580,N_2770,N_2491);
nor U5581 (N_5581,N_2558,N_2936);
nor U5582 (N_5582,N_2958,N_3080);
or U5583 (N_5583,N_2523,N_3679);
or U5584 (N_5584,N_3935,N_3453);
or U5585 (N_5585,N_3812,N_3177);
nor U5586 (N_5586,N_3974,N_2359);
nor U5587 (N_5587,N_2879,N_2109);
nor U5588 (N_5588,N_3386,N_3826);
nand U5589 (N_5589,N_3450,N_3400);
and U5590 (N_5590,N_3331,N_2868);
nand U5591 (N_5591,N_3360,N_3594);
or U5592 (N_5592,N_3369,N_2772);
nor U5593 (N_5593,N_2209,N_2897);
nand U5594 (N_5594,N_3997,N_2606);
or U5595 (N_5595,N_3138,N_3506);
or U5596 (N_5596,N_3257,N_3827);
nand U5597 (N_5597,N_2881,N_2605);
or U5598 (N_5598,N_3834,N_3849);
nor U5599 (N_5599,N_3863,N_2116);
nor U5600 (N_5600,N_3035,N_2494);
nand U5601 (N_5601,N_2859,N_2772);
nor U5602 (N_5602,N_3982,N_3244);
and U5603 (N_5603,N_2324,N_3078);
and U5604 (N_5604,N_3013,N_2515);
and U5605 (N_5605,N_3698,N_3190);
or U5606 (N_5606,N_3960,N_2934);
nand U5607 (N_5607,N_2298,N_3970);
or U5608 (N_5608,N_2520,N_2669);
and U5609 (N_5609,N_3494,N_2614);
nor U5610 (N_5610,N_3983,N_2983);
and U5611 (N_5611,N_2190,N_2557);
nand U5612 (N_5612,N_3036,N_2614);
nand U5613 (N_5613,N_3593,N_2233);
or U5614 (N_5614,N_3564,N_3522);
nor U5615 (N_5615,N_3728,N_3871);
and U5616 (N_5616,N_2472,N_2468);
nand U5617 (N_5617,N_2328,N_2056);
and U5618 (N_5618,N_2378,N_3737);
and U5619 (N_5619,N_3891,N_2942);
nor U5620 (N_5620,N_2342,N_2364);
nor U5621 (N_5621,N_2895,N_3328);
or U5622 (N_5622,N_3728,N_2692);
nor U5623 (N_5623,N_2828,N_2656);
and U5624 (N_5624,N_2337,N_2316);
nand U5625 (N_5625,N_3213,N_3795);
and U5626 (N_5626,N_2221,N_3722);
and U5627 (N_5627,N_2702,N_3061);
and U5628 (N_5628,N_2721,N_3089);
or U5629 (N_5629,N_3672,N_3612);
nor U5630 (N_5630,N_2433,N_3756);
nor U5631 (N_5631,N_2335,N_2835);
and U5632 (N_5632,N_3395,N_2641);
and U5633 (N_5633,N_2378,N_3994);
and U5634 (N_5634,N_3462,N_3752);
or U5635 (N_5635,N_3009,N_3415);
xnor U5636 (N_5636,N_3667,N_2947);
or U5637 (N_5637,N_2996,N_3382);
nor U5638 (N_5638,N_2374,N_3353);
and U5639 (N_5639,N_2998,N_3972);
or U5640 (N_5640,N_3122,N_3692);
nor U5641 (N_5641,N_3358,N_2817);
nand U5642 (N_5642,N_2119,N_3424);
nand U5643 (N_5643,N_3786,N_2121);
and U5644 (N_5644,N_3340,N_3250);
nor U5645 (N_5645,N_3468,N_2890);
nand U5646 (N_5646,N_3006,N_3512);
nand U5647 (N_5647,N_3109,N_3183);
and U5648 (N_5648,N_2399,N_2547);
xnor U5649 (N_5649,N_3704,N_2944);
or U5650 (N_5650,N_3848,N_2773);
and U5651 (N_5651,N_2334,N_3327);
nor U5652 (N_5652,N_3997,N_2296);
and U5653 (N_5653,N_2098,N_2772);
or U5654 (N_5654,N_2383,N_2201);
nand U5655 (N_5655,N_3506,N_2687);
nand U5656 (N_5656,N_2495,N_3620);
and U5657 (N_5657,N_2690,N_3143);
and U5658 (N_5658,N_3645,N_3696);
and U5659 (N_5659,N_3631,N_2879);
or U5660 (N_5660,N_2528,N_2790);
or U5661 (N_5661,N_3584,N_3178);
and U5662 (N_5662,N_2740,N_3879);
or U5663 (N_5663,N_3552,N_2292);
or U5664 (N_5664,N_2587,N_3249);
and U5665 (N_5665,N_3478,N_3026);
nor U5666 (N_5666,N_2229,N_3593);
and U5667 (N_5667,N_2115,N_3826);
or U5668 (N_5668,N_3925,N_3615);
nor U5669 (N_5669,N_2176,N_3338);
and U5670 (N_5670,N_2156,N_2226);
and U5671 (N_5671,N_2002,N_2217);
and U5672 (N_5672,N_2047,N_3950);
nand U5673 (N_5673,N_2479,N_3046);
nor U5674 (N_5674,N_3893,N_2899);
nand U5675 (N_5675,N_2039,N_2184);
nor U5676 (N_5676,N_3166,N_3105);
nand U5677 (N_5677,N_2907,N_3890);
and U5678 (N_5678,N_2555,N_3371);
and U5679 (N_5679,N_3278,N_2260);
and U5680 (N_5680,N_2310,N_3069);
and U5681 (N_5681,N_2508,N_3140);
or U5682 (N_5682,N_2456,N_3335);
and U5683 (N_5683,N_3452,N_2893);
nand U5684 (N_5684,N_3544,N_3147);
nand U5685 (N_5685,N_2059,N_3591);
or U5686 (N_5686,N_3359,N_3177);
and U5687 (N_5687,N_2310,N_2495);
and U5688 (N_5688,N_2474,N_3867);
nand U5689 (N_5689,N_3784,N_3323);
or U5690 (N_5690,N_2563,N_3520);
or U5691 (N_5691,N_3596,N_3398);
and U5692 (N_5692,N_3144,N_2497);
or U5693 (N_5693,N_2022,N_3452);
nor U5694 (N_5694,N_2491,N_2223);
nand U5695 (N_5695,N_2384,N_3717);
xor U5696 (N_5696,N_2513,N_2240);
nor U5697 (N_5697,N_2129,N_3753);
nand U5698 (N_5698,N_2295,N_2882);
nor U5699 (N_5699,N_3915,N_2947);
nor U5700 (N_5700,N_3343,N_3002);
nor U5701 (N_5701,N_3935,N_2874);
or U5702 (N_5702,N_2973,N_2080);
or U5703 (N_5703,N_3864,N_2678);
and U5704 (N_5704,N_3586,N_3926);
nor U5705 (N_5705,N_2363,N_2699);
or U5706 (N_5706,N_3130,N_3141);
nand U5707 (N_5707,N_2938,N_2315);
nand U5708 (N_5708,N_3600,N_2102);
and U5709 (N_5709,N_3376,N_3400);
and U5710 (N_5710,N_2496,N_2815);
or U5711 (N_5711,N_2151,N_3454);
or U5712 (N_5712,N_2650,N_3547);
and U5713 (N_5713,N_3184,N_2313);
and U5714 (N_5714,N_2314,N_3308);
nand U5715 (N_5715,N_3371,N_3510);
nor U5716 (N_5716,N_2304,N_2458);
or U5717 (N_5717,N_3410,N_2727);
nand U5718 (N_5718,N_2569,N_2117);
nor U5719 (N_5719,N_2763,N_2368);
or U5720 (N_5720,N_3753,N_3295);
nor U5721 (N_5721,N_2676,N_3717);
nand U5722 (N_5722,N_2304,N_2272);
or U5723 (N_5723,N_2754,N_3644);
nor U5724 (N_5724,N_3161,N_2611);
nand U5725 (N_5725,N_2401,N_3195);
and U5726 (N_5726,N_2189,N_2402);
nand U5727 (N_5727,N_3947,N_3130);
or U5728 (N_5728,N_3124,N_3357);
or U5729 (N_5729,N_2189,N_3170);
nand U5730 (N_5730,N_3710,N_2075);
nand U5731 (N_5731,N_2970,N_2444);
nor U5732 (N_5732,N_2679,N_2398);
nor U5733 (N_5733,N_2840,N_3801);
and U5734 (N_5734,N_2728,N_2588);
nor U5735 (N_5735,N_2185,N_2708);
xnor U5736 (N_5736,N_3743,N_2457);
nand U5737 (N_5737,N_3572,N_3402);
nand U5738 (N_5738,N_3963,N_2794);
nand U5739 (N_5739,N_3780,N_2421);
and U5740 (N_5740,N_2658,N_3393);
nor U5741 (N_5741,N_2065,N_2098);
or U5742 (N_5742,N_2403,N_2046);
or U5743 (N_5743,N_3767,N_2049);
nand U5744 (N_5744,N_2921,N_2409);
and U5745 (N_5745,N_2585,N_3897);
xnor U5746 (N_5746,N_2383,N_3540);
nand U5747 (N_5747,N_2958,N_3341);
nor U5748 (N_5748,N_3564,N_3761);
and U5749 (N_5749,N_2180,N_3629);
nor U5750 (N_5750,N_2279,N_3203);
and U5751 (N_5751,N_3652,N_3856);
and U5752 (N_5752,N_3704,N_2893);
nor U5753 (N_5753,N_2624,N_2114);
or U5754 (N_5754,N_3514,N_3464);
nor U5755 (N_5755,N_2301,N_2409);
or U5756 (N_5756,N_2893,N_3529);
nor U5757 (N_5757,N_3302,N_2104);
or U5758 (N_5758,N_3026,N_3995);
xor U5759 (N_5759,N_3140,N_3274);
or U5760 (N_5760,N_3742,N_3910);
and U5761 (N_5761,N_2871,N_3419);
and U5762 (N_5762,N_3347,N_3056);
xor U5763 (N_5763,N_2579,N_3388);
nor U5764 (N_5764,N_3727,N_2854);
or U5765 (N_5765,N_3057,N_3576);
and U5766 (N_5766,N_2356,N_2101);
nand U5767 (N_5767,N_3458,N_3652);
and U5768 (N_5768,N_2830,N_2745);
nor U5769 (N_5769,N_3798,N_2698);
nand U5770 (N_5770,N_3483,N_3422);
nor U5771 (N_5771,N_2010,N_2847);
nor U5772 (N_5772,N_3665,N_3805);
nor U5773 (N_5773,N_3557,N_3556);
nand U5774 (N_5774,N_3342,N_3389);
and U5775 (N_5775,N_3303,N_2184);
and U5776 (N_5776,N_3083,N_2423);
nor U5777 (N_5777,N_2830,N_3332);
and U5778 (N_5778,N_3696,N_2363);
or U5779 (N_5779,N_3546,N_2736);
or U5780 (N_5780,N_2614,N_2104);
or U5781 (N_5781,N_2060,N_2965);
or U5782 (N_5782,N_3146,N_3556);
nor U5783 (N_5783,N_2781,N_3378);
or U5784 (N_5784,N_2882,N_2131);
nor U5785 (N_5785,N_2110,N_3509);
nand U5786 (N_5786,N_2412,N_3367);
and U5787 (N_5787,N_2990,N_2942);
and U5788 (N_5788,N_2520,N_3242);
or U5789 (N_5789,N_2483,N_2733);
and U5790 (N_5790,N_2679,N_3914);
and U5791 (N_5791,N_3306,N_2105);
nand U5792 (N_5792,N_3485,N_3060);
and U5793 (N_5793,N_2062,N_3420);
nand U5794 (N_5794,N_2692,N_2379);
and U5795 (N_5795,N_3966,N_2127);
and U5796 (N_5796,N_3008,N_2376);
nand U5797 (N_5797,N_2734,N_2436);
and U5798 (N_5798,N_2674,N_3955);
and U5799 (N_5799,N_3831,N_3884);
and U5800 (N_5800,N_3537,N_3398);
and U5801 (N_5801,N_3167,N_3744);
nand U5802 (N_5802,N_2376,N_2095);
xnor U5803 (N_5803,N_3584,N_3883);
nand U5804 (N_5804,N_3044,N_2620);
xor U5805 (N_5805,N_2926,N_3664);
or U5806 (N_5806,N_2345,N_2304);
and U5807 (N_5807,N_2288,N_3560);
nor U5808 (N_5808,N_3230,N_2317);
nor U5809 (N_5809,N_3321,N_2916);
nor U5810 (N_5810,N_3321,N_3889);
and U5811 (N_5811,N_3462,N_2292);
or U5812 (N_5812,N_2043,N_3194);
or U5813 (N_5813,N_3378,N_3288);
nor U5814 (N_5814,N_3156,N_2207);
nor U5815 (N_5815,N_3697,N_3521);
xor U5816 (N_5816,N_3389,N_2281);
and U5817 (N_5817,N_3383,N_3995);
or U5818 (N_5818,N_3024,N_2560);
nand U5819 (N_5819,N_2943,N_2306);
nand U5820 (N_5820,N_2764,N_3270);
nand U5821 (N_5821,N_3046,N_3871);
xor U5822 (N_5822,N_2942,N_3027);
nor U5823 (N_5823,N_2240,N_3101);
or U5824 (N_5824,N_2392,N_2293);
nand U5825 (N_5825,N_2154,N_2309);
and U5826 (N_5826,N_3312,N_3194);
nor U5827 (N_5827,N_3028,N_2614);
nand U5828 (N_5828,N_2681,N_3156);
nor U5829 (N_5829,N_2462,N_3740);
or U5830 (N_5830,N_3268,N_3832);
nor U5831 (N_5831,N_3641,N_2939);
or U5832 (N_5832,N_3463,N_3299);
nand U5833 (N_5833,N_3572,N_2448);
and U5834 (N_5834,N_3326,N_2892);
nand U5835 (N_5835,N_2610,N_2474);
or U5836 (N_5836,N_3989,N_2008);
nand U5837 (N_5837,N_3759,N_2886);
nand U5838 (N_5838,N_3794,N_2351);
nor U5839 (N_5839,N_3946,N_3581);
or U5840 (N_5840,N_2897,N_2121);
or U5841 (N_5841,N_2043,N_3690);
or U5842 (N_5842,N_3541,N_2428);
and U5843 (N_5843,N_3360,N_3517);
or U5844 (N_5844,N_2085,N_3310);
and U5845 (N_5845,N_3914,N_3048);
nand U5846 (N_5846,N_3674,N_3631);
nand U5847 (N_5847,N_2684,N_3652);
or U5848 (N_5848,N_3127,N_2024);
and U5849 (N_5849,N_2098,N_2232);
or U5850 (N_5850,N_3723,N_2453);
and U5851 (N_5851,N_2700,N_2264);
nand U5852 (N_5852,N_3617,N_3732);
and U5853 (N_5853,N_3126,N_3779);
and U5854 (N_5854,N_3088,N_2263);
and U5855 (N_5855,N_2700,N_3838);
or U5856 (N_5856,N_2122,N_2499);
and U5857 (N_5857,N_2670,N_2193);
nand U5858 (N_5858,N_2819,N_3133);
nor U5859 (N_5859,N_3338,N_2191);
xnor U5860 (N_5860,N_2611,N_2457);
and U5861 (N_5861,N_2999,N_3990);
and U5862 (N_5862,N_2347,N_2696);
nand U5863 (N_5863,N_2292,N_3935);
nand U5864 (N_5864,N_3936,N_2108);
or U5865 (N_5865,N_3274,N_2463);
or U5866 (N_5866,N_2990,N_3863);
nand U5867 (N_5867,N_3253,N_3375);
nor U5868 (N_5868,N_3321,N_2856);
or U5869 (N_5869,N_3730,N_2497);
and U5870 (N_5870,N_2188,N_3193);
and U5871 (N_5871,N_2002,N_3465);
nand U5872 (N_5872,N_2427,N_3980);
nor U5873 (N_5873,N_3828,N_3672);
nand U5874 (N_5874,N_2831,N_3025);
nand U5875 (N_5875,N_3669,N_2755);
and U5876 (N_5876,N_2567,N_3429);
nor U5877 (N_5877,N_2968,N_2185);
or U5878 (N_5878,N_2810,N_3105);
nor U5879 (N_5879,N_2095,N_2026);
nor U5880 (N_5880,N_3618,N_2750);
nor U5881 (N_5881,N_2112,N_2852);
or U5882 (N_5882,N_2216,N_2244);
and U5883 (N_5883,N_2563,N_2885);
nand U5884 (N_5884,N_2637,N_2840);
nor U5885 (N_5885,N_3268,N_3139);
nor U5886 (N_5886,N_3821,N_2399);
nand U5887 (N_5887,N_2494,N_3673);
and U5888 (N_5888,N_2952,N_2361);
and U5889 (N_5889,N_3419,N_3516);
and U5890 (N_5890,N_3571,N_3625);
nor U5891 (N_5891,N_2523,N_3361);
or U5892 (N_5892,N_2476,N_2078);
nor U5893 (N_5893,N_2148,N_2664);
nor U5894 (N_5894,N_3122,N_3624);
nand U5895 (N_5895,N_2177,N_3544);
nor U5896 (N_5896,N_3291,N_3039);
nand U5897 (N_5897,N_3332,N_2922);
nor U5898 (N_5898,N_2050,N_2558);
and U5899 (N_5899,N_3079,N_2823);
nor U5900 (N_5900,N_2886,N_3302);
nor U5901 (N_5901,N_2918,N_3254);
nor U5902 (N_5902,N_2226,N_3393);
or U5903 (N_5903,N_2929,N_2506);
nor U5904 (N_5904,N_2964,N_2364);
and U5905 (N_5905,N_3697,N_2171);
or U5906 (N_5906,N_2435,N_2102);
or U5907 (N_5907,N_2444,N_3697);
and U5908 (N_5908,N_2999,N_2976);
nand U5909 (N_5909,N_2251,N_3616);
nor U5910 (N_5910,N_2515,N_2745);
nand U5911 (N_5911,N_2507,N_2018);
or U5912 (N_5912,N_2181,N_2909);
nor U5913 (N_5913,N_3928,N_2490);
nor U5914 (N_5914,N_3362,N_2971);
nor U5915 (N_5915,N_3315,N_3080);
nand U5916 (N_5916,N_2224,N_3116);
or U5917 (N_5917,N_3005,N_3170);
nor U5918 (N_5918,N_2809,N_3180);
and U5919 (N_5919,N_3147,N_3698);
nand U5920 (N_5920,N_2775,N_3321);
nand U5921 (N_5921,N_3506,N_2106);
and U5922 (N_5922,N_3052,N_3480);
and U5923 (N_5923,N_2907,N_3524);
and U5924 (N_5924,N_2323,N_3183);
or U5925 (N_5925,N_2839,N_2766);
nand U5926 (N_5926,N_2178,N_3294);
nand U5927 (N_5927,N_2175,N_3585);
and U5928 (N_5928,N_2527,N_2183);
or U5929 (N_5929,N_3275,N_3012);
or U5930 (N_5930,N_2068,N_3044);
or U5931 (N_5931,N_2502,N_3529);
nor U5932 (N_5932,N_2045,N_2392);
or U5933 (N_5933,N_3124,N_2428);
or U5934 (N_5934,N_2831,N_3750);
nand U5935 (N_5935,N_3832,N_2811);
nor U5936 (N_5936,N_3789,N_3785);
or U5937 (N_5937,N_3576,N_3501);
and U5938 (N_5938,N_3689,N_2833);
and U5939 (N_5939,N_2185,N_3703);
nand U5940 (N_5940,N_3295,N_2382);
nand U5941 (N_5941,N_2481,N_3445);
nand U5942 (N_5942,N_2263,N_2818);
nor U5943 (N_5943,N_3571,N_2029);
nor U5944 (N_5944,N_3789,N_3364);
nor U5945 (N_5945,N_3225,N_3827);
nand U5946 (N_5946,N_3837,N_2096);
nand U5947 (N_5947,N_3702,N_3321);
nand U5948 (N_5948,N_2674,N_3873);
and U5949 (N_5949,N_3502,N_2909);
or U5950 (N_5950,N_2420,N_3720);
nand U5951 (N_5951,N_2563,N_3478);
nor U5952 (N_5952,N_3005,N_3787);
nor U5953 (N_5953,N_3194,N_3667);
xnor U5954 (N_5954,N_3876,N_3559);
nor U5955 (N_5955,N_3526,N_2651);
nand U5956 (N_5956,N_2193,N_2659);
nand U5957 (N_5957,N_2373,N_3595);
nor U5958 (N_5958,N_3546,N_3359);
nand U5959 (N_5959,N_2100,N_2151);
and U5960 (N_5960,N_3931,N_2667);
nor U5961 (N_5961,N_3084,N_3237);
nor U5962 (N_5962,N_3811,N_2204);
nand U5963 (N_5963,N_2453,N_2475);
nor U5964 (N_5964,N_2990,N_3268);
nand U5965 (N_5965,N_3834,N_3594);
and U5966 (N_5966,N_2503,N_3612);
and U5967 (N_5967,N_2802,N_3524);
nor U5968 (N_5968,N_3088,N_3302);
and U5969 (N_5969,N_3828,N_2982);
nor U5970 (N_5970,N_2435,N_2615);
nand U5971 (N_5971,N_3946,N_3180);
or U5972 (N_5972,N_3293,N_3930);
nand U5973 (N_5973,N_3652,N_2620);
nand U5974 (N_5974,N_3416,N_2705);
and U5975 (N_5975,N_2403,N_3199);
nor U5976 (N_5976,N_2997,N_3703);
nand U5977 (N_5977,N_2878,N_3005);
or U5978 (N_5978,N_2498,N_2435);
nand U5979 (N_5979,N_3086,N_3221);
or U5980 (N_5980,N_2619,N_3337);
and U5981 (N_5981,N_2523,N_3539);
nor U5982 (N_5982,N_2823,N_2831);
or U5983 (N_5983,N_3470,N_3982);
nand U5984 (N_5984,N_2236,N_2549);
nor U5985 (N_5985,N_2272,N_3987);
nor U5986 (N_5986,N_2752,N_2919);
or U5987 (N_5987,N_3609,N_3274);
or U5988 (N_5988,N_3589,N_2539);
and U5989 (N_5989,N_3710,N_2450);
and U5990 (N_5990,N_3875,N_2362);
and U5991 (N_5991,N_2616,N_3015);
nand U5992 (N_5992,N_3919,N_2305);
nor U5993 (N_5993,N_2460,N_2569);
nor U5994 (N_5994,N_3445,N_3560);
nor U5995 (N_5995,N_2139,N_3274);
and U5996 (N_5996,N_2007,N_2010);
and U5997 (N_5997,N_2284,N_2882);
nor U5998 (N_5998,N_2331,N_3924);
nor U5999 (N_5999,N_2678,N_2638);
xnor U6000 (N_6000,N_5085,N_4299);
or U6001 (N_6001,N_5268,N_4525);
or U6002 (N_6002,N_5044,N_4827);
and U6003 (N_6003,N_5611,N_4606);
and U6004 (N_6004,N_5278,N_5795);
nor U6005 (N_6005,N_5636,N_4735);
nor U6006 (N_6006,N_5227,N_4098);
and U6007 (N_6007,N_5970,N_5823);
nand U6008 (N_6008,N_4029,N_4520);
nor U6009 (N_6009,N_4773,N_5147);
nor U6010 (N_6010,N_5959,N_4253);
nand U6011 (N_6011,N_4976,N_4708);
nand U6012 (N_6012,N_4000,N_5911);
nand U6013 (N_6013,N_5119,N_5995);
or U6014 (N_6014,N_4276,N_5742);
or U6015 (N_6015,N_5336,N_4433);
or U6016 (N_6016,N_4903,N_4243);
and U6017 (N_6017,N_5866,N_5190);
or U6018 (N_6018,N_4424,N_4593);
nand U6019 (N_6019,N_4836,N_5221);
and U6020 (N_6020,N_5571,N_4596);
or U6021 (N_6021,N_4216,N_5414);
nor U6022 (N_6022,N_5904,N_5038);
nand U6023 (N_6023,N_4712,N_5578);
or U6024 (N_6024,N_4306,N_5667);
nand U6025 (N_6025,N_4034,N_4930);
or U6026 (N_6026,N_4536,N_5416);
nor U6027 (N_6027,N_4585,N_4053);
nor U6028 (N_6028,N_4823,N_5525);
or U6029 (N_6029,N_4274,N_5912);
or U6030 (N_6030,N_5779,N_5099);
nand U6031 (N_6031,N_5367,N_5839);
and U6032 (N_6032,N_4635,N_4790);
and U6033 (N_6033,N_5285,N_5161);
and U6034 (N_6034,N_4666,N_5132);
and U6035 (N_6035,N_5187,N_5537);
and U6036 (N_6036,N_4136,N_5469);
or U6037 (N_6037,N_4899,N_5671);
nand U6038 (N_6038,N_5835,N_5974);
or U6039 (N_6039,N_4463,N_4928);
nor U6040 (N_6040,N_4504,N_4173);
nor U6041 (N_6041,N_5109,N_5164);
nor U6042 (N_6042,N_4428,N_5483);
or U6043 (N_6043,N_4963,N_4788);
nand U6044 (N_6044,N_4115,N_5564);
nor U6045 (N_6045,N_4441,N_5669);
and U6046 (N_6046,N_5720,N_5960);
nand U6047 (N_6047,N_4308,N_5019);
or U6048 (N_6048,N_4415,N_5990);
or U6049 (N_6049,N_4031,N_4335);
or U6050 (N_6050,N_5729,N_4208);
nor U6051 (N_6051,N_5185,N_5282);
or U6052 (N_6052,N_4713,N_5641);
and U6053 (N_6053,N_4512,N_4647);
and U6054 (N_6054,N_5006,N_5819);
nand U6055 (N_6055,N_4990,N_4796);
or U6056 (N_6056,N_5337,N_5951);
and U6057 (N_6057,N_4514,N_5289);
or U6058 (N_6058,N_5873,N_4907);
or U6059 (N_6059,N_5438,N_4317);
and U6060 (N_6060,N_5971,N_4537);
and U6061 (N_6061,N_5957,N_5045);
nor U6062 (N_6062,N_5575,N_5654);
and U6063 (N_6063,N_5486,N_4964);
and U6064 (N_6064,N_4069,N_4180);
nor U6065 (N_6065,N_5073,N_5412);
nand U6066 (N_6066,N_5191,N_4224);
nor U6067 (N_6067,N_4330,N_4456);
or U6068 (N_6068,N_4557,N_5324);
nor U6069 (N_6069,N_4238,N_4252);
and U6070 (N_6070,N_5580,N_5434);
nand U6071 (N_6071,N_5879,N_5939);
or U6072 (N_6072,N_4854,N_4400);
and U6073 (N_6073,N_5308,N_5644);
or U6074 (N_6074,N_4474,N_5950);
nand U6075 (N_6075,N_5521,N_4949);
and U6076 (N_6076,N_5030,N_5747);
and U6077 (N_6077,N_4261,N_4548);
nand U6078 (N_6078,N_5888,N_5850);
and U6079 (N_6079,N_4254,N_5194);
nor U6080 (N_6080,N_5105,N_5152);
and U6081 (N_6081,N_4573,N_5293);
nor U6082 (N_6082,N_4054,N_4088);
and U6083 (N_6083,N_4207,N_5725);
or U6084 (N_6084,N_5909,N_5512);
or U6085 (N_6085,N_4838,N_5601);
and U6086 (N_6086,N_5622,N_4714);
and U6087 (N_6087,N_5093,N_4926);
nor U6088 (N_6088,N_4813,N_5544);
and U6089 (N_6089,N_5963,N_4003);
and U6090 (N_6090,N_4161,N_5347);
nand U6091 (N_6091,N_4383,N_5306);
nand U6092 (N_6092,N_5877,N_4986);
or U6093 (N_6093,N_4526,N_5095);
nor U6094 (N_6094,N_5771,N_4787);
or U6095 (N_6095,N_4966,N_5884);
nor U6096 (N_6096,N_5609,N_5468);
nor U6097 (N_6097,N_5057,N_5067);
nand U6098 (N_6098,N_5917,N_4336);
nor U6099 (N_6099,N_4820,N_5793);
nand U6100 (N_6100,N_4325,N_4211);
nor U6101 (N_6101,N_4333,N_4781);
and U6102 (N_6102,N_5899,N_4910);
nor U6103 (N_6103,N_4695,N_4381);
or U6104 (N_6104,N_4356,N_4795);
or U6105 (N_6105,N_5811,N_5430);
nand U6106 (N_6106,N_5481,N_5903);
or U6107 (N_6107,N_5538,N_4460);
and U6108 (N_6108,N_5373,N_4542);
or U6109 (N_6109,N_5825,N_5479);
and U6110 (N_6110,N_5441,N_4302);
nor U6111 (N_6111,N_4329,N_5966);
nand U6112 (N_6112,N_5344,N_5913);
and U6113 (N_6113,N_5062,N_4832);
nand U6114 (N_6114,N_5024,N_4889);
nand U6115 (N_6115,N_5813,N_4133);
nor U6116 (N_6116,N_5854,N_5660);
or U6117 (N_6117,N_4829,N_5969);
and U6118 (N_6118,N_5606,N_4806);
or U6119 (N_6119,N_4917,N_5954);
or U6120 (N_6120,N_4364,N_4682);
and U6121 (N_6121,N_5645,N_4396);
nor U6122 (N_6122,N_4799,N_4156);
or U6123 (N_6123,N_5902,N_4817);
and U6124 (N_6124,N_5100,N_4532);
or U6125 (N_6125,N_4011,N_4687);
nor U6126 (N_6126,N_4960,N_4097);
or U6127 (N_6127,N_4675,N_5245);
nand U6128 (N_6128,N_4282,N_4915);
or U6129 (N_6129,N_4150,N_5508);
nor U6130 (N_6130,N_4105,N_4545);
nor U6131 (N_6131,N_5698,N_5421);
or U6132 (N_6132,N_4758,N_5688);
nand U6133 (N_6133,N_4495,N_5548);
nand U6134 (N_6134,N_4581,N_5153);
and U6135 (N_6135,N_4511,N_5762);
nand U6136 (N_6136,N_5587,N_4667);
nand U6137 (N_6137,N_4856,N_5397);
and U6138 (N_6138,N_5334,N_4265);
or U6139 (N_6139,N_4849,N_5151);
nand U6140 (N_6140,N_5092,N_5527);
and U6141 (N_6141,N_4108,N_5043);
nor U6142 (N_6142,N_5734,N_4981);
and U6143 (N_6143,N_4255,N_4692);
nand U6144 (N_6144,N_4655,N_4195);
nand U6145 (N_6145,N_4158,N_5160);
or U6146 (N_6146,N_5200,N_5919);
nand U6147 (N_6147,N_5703,N_5203);
nand U6148 (N_6148,N_4703,N_4037);
nor U6149 (N_6149,N_4015,N_4693);
and U6150 (N_6150,N_4867,N_5649);
nor U6151 (N_6151,N_5039,N_5304);
nand U6152 (N_6152,N_4840,N_4443);
nor U6153 (N_6153,N_4215,N_4517);
or U6154 (N_6154,N_5140,N_5033);
nand U6155 (N_6155,N_4578,N_4595);
and U6156 (N_6156,N_5088,N_5847);
and U6157 (N_6157,N_5766,N_5704);
and U6158 (N_6158,N_4489,N_5701);
nand U6159 (N_6159,N_5297,N_5935);
and U6160 (N_6160,N_4058,N_5137);
nand U6161 (N_6161,N_4978,N_5689);
nor U6162 (N_6162,N_4411,N_4194);
or U6163 (N_6163,N_5255,N_5767);
and U6164 (N_6164,N_4529,N_5927);
nor U6165 (N_6165,N_4312,N_4318);
or U6166 (N_6166,N_4860,N_5849);
nor U6167 (N_6167,N_4843,N_5653);
nor U6168 (N_6168,N_4283,N_4995);
nor U6169 (N_6169,N_5712,N_5702);
nand U6170 (N_6170,N_5547,N_4056);
xor U6171 (N_6171,N_5910,N_5215);
nand U6172 (N_6172,N_5391,N_4563);
and U6173 (N_6173,N_5922,N_4081);
and U6174 (N_6174,N_4737,N_5748);
or U6175 (N_6175,N_5615,N_4804);
nor U6176 (N_6176,N_4386,N_5715);
or U6177 (N_6177,N_5112,N_4177);
nor U6178 (N_6178,N_5253,N_4881);
nor U6179 (N_6179,N_4162,N_4125);
nand U6180 (N_6180,N_4858,N_5396);
and U6181 (N_6181,N_5106,N_4240);
nor U6182 (N_6182,N_4142,N_5022);
or U6183 (N_6183,N_5674,N_4920);
or U6184 (N_6184,N_5518,N_5210);
and U6185 (N_6185,N_5064,N_5980);
or U6186 (N_6186,N_5646,N_5376);
nand U6187 (N_6187,N_4237,N_5631);
and U6188 (N_6188,N_5530,N_4146);
or U6189 (N_6189,N_5802,N_5311);
nand U6190 (N_6190,N_5102,N_5249);
and U6191 (N_6191,N_5320,N_5650);
and U6192 (N_6192,N_5830,N_4974);
or U6193 (N_6193,N_5060,N_5485);
nor U6194 (N_6194,N_4614,N_4239);
nor U6195 (N_6195,N_4604,N_5536);
nand U6196 (N_6196,N_4534,N_4061);
or U6197 (N_6197,N_4733,N_5487);
and U6198 (N_6198,N_5368,N_4196);
nand U6199 (N_6199,N_5924,N_5473);
nand U6200 (N_6200,N_5238,N_4670);
nand U6201 (N_6201,N_4445,N_4991);
nand U6202 (N_6202,N_4734,N_4630);
and U6203 (N_6203,N_4609,N_5676);
nor U6204 (N_6204,N_5696,N_5665);
or U6205 (N_6205,N_4159,N_4970);
nand U6206 (N_6206,N_4527,N_5523);
nor U6207 (N_6207,N_4686,N_5244);
nor U6208 (N_6208,N_5007,N_4124);
or U6209 (N_6209,N_5362,N_5419);
or U6210 (N_6210,N_5301,N_5932);
or U6211 (N_6211,N_5893,N_5328);
nand U6212 (N_6212,N_5431,N_4476);
and U6213 (N_6213,N_4837,N_5212);
nor U6214 (N_6214,N_4139,N_5713);
and U6215 (N_6215,N_5018,N_4810);
or U6216 (N_6216,N_5439,N_5625);
nor U6217 (N_6217,N_5568,N_4861);
and U6218 (N_6218,N_4950,N_4886);
nor U6219 (N_6219,N_4199,N_5915);
and U6220 (N_6220,N_5626,N_5063);
nand U6221 (N_6221,N_5372,N_4036);
nand U6222 (N_6222,N_5040,N_4848);
and U6223 (N_6223,N_5517,N_5861);
nor U6224 (N_6224,N_4414,N_4109);
nor U6225 (N_6225,N_5949,N_5407);
and U6226 (N_6226,N_5292,N_5188);
and U6227 (N_6227,N_4524,N_4144);
nand U6228 (N_6228,N_5319,N_4114);
and U6229 (N_6229,N_4185,N_5726);
nor U6230 (N_6230,N_4749,N_5454);
nor U6231 (N_6231,N_5230,N_5484);
and U6232 (N_6232,N_4834,N_4610);
and U6233 (N_6233,N_5716,N_5066);
nor U6234 (N_6234,N_4619,N_5353);
or U6235 (N_6235,N_5058,N_5918);
nand U6236 (N_6236,N_4030,N_5217);
and U6237 (N_6237,N_4281,N_5603);
and U6238 (N_6238,N_4166,N_5448);
xor U6239 (N_6239,N_4882,N_4618);
nand U6240 (N_6240,N_4084,N_5478);
nor U6241 (N_6241,N_4471,N_5429);
and U6242 (N_6242,N_4701,N_5799);
and U6243 (N_6243,N_4353,N_5723);
and U6244 (N_6244,N_5193,N_4519);
nor U6245 (N_6245,N_4946,N_4651);
nor U6246 (N_6246,N_4090,N_4996);
or U6247 (N_6247,N_5504,N_5299);
nand U6248 (N_6248,N_5392,N_5069);
xnor U6249 (N_6249,N_5540,N_5993);
and U6250 (N_6250,N_4902,N_4863);
xnor U6251 (N_6251,N_5179,N_4932);
nand U6252 (N_6252,N_4835,N_5387);
or U6253 (N_6253,N_5305,N_5051);
or U6254 (N_6254,N_4672,N_5141);
and U6255 (N_6255,N_5731,N_5011);
nor U6256 (N_6256,N_5390,N_4155);
nor U6257 (N_6257,N_4769,N_5869);
nand U6258 (N_6258,N_5380,N_5420);
or U6259 (N_6259,N_4797,N_5574);
and U6260 (N_6260,N_5405,N_4762);
and U6261 (N_6261,N_5252,N_5082);
nand U6262 (N_6262,N_5300,N_5488);
and U6263 (N_6263,N_5350,N_4373);
or U6264 (N_6264,N_4597,N_4020);
and U6265 (N_6265,N_4874,N_4959);
and U6266 (N_6266,N_5898,N_4075);
nor U6267 (N_6267,N_4957,N_5156);
and U6268 (N_6268,N_5169,N_5868);
or U6269 (N_6269,N_5424,N_5111);
nor U6270 (N_6270,N_5089,N_4296);
and U6271 (N_6271,N_4560,N_4355);
nor U6272 (N_6272,N_5739,N_5216);
and U6273 (N_6273,N_4492,N_5505);
or U6274 (N_6274,N_5897,N_4116);
nor U6275 (N_6275,N_4498,N_4638);
and U6276 (N_6276,N_4190,N_5510);
or U6277 (N_6277,N_4307,N_4439);
and U6278 (N_6278,N_4467,N_5937);
or U6279 (N_6279,N_4064,N_4540);
nor U6280 (N_6280,N_5843,N_5551);
nor U6281 (N_6281,N_4556,N_4257);
and U6282 (N_6282,N_4006,N_4009);
or U6283 (N_6283,N_4197,N_4392);
or U6284 (N_6284,N_4751,N_4494);
nor U6285 (N_6285,N_5965,N_4262);
and U6286 (N_6286,N_5078,N_4360);
or U6287 (N_6287,N_4931,N_4175);
or U6288 (N_6288,N_4331,N_4592);
nand U6289 (N_6289,N_5047,N_5471);
and U6290 (N_6290,N_4844,N_4664);
nand U6291 (N_6291,N_4576,N_5280);
nand U6292 (N_6292,N_5686,N_4757);
nand U6293 (N_6293,N_4927,N_4406);
nand U6294 (N_6294,N_4879,N_4087);
or U6295 (N_6295,N_5198,N_5853);
and U6296 (N_6296,N_4948,N_4453);
or U6297 (N_6297,N_5800,N_5933);
or U6298 (N_6298,N_5882,N_4673);
nand U6299 (N_6299,N_4232,N_5612);
nor U6300 (N_6300,N_4658,N_5394);
and U6301 (N_6301,N_5340,N_4507);
nand U6302 (N_6302,N_5901,N_4334);
and U6303 (N_6303,N_4706,N_4148);
and U6304 (N_6304,N_5228,N_4273);
nand U6305 (N_6305,N_5466,N_5542);
nor U6306 (N_6306,N_4412,N_5947);
or U6307 (N_6307,N_4072,N_4294);
nand U6308 (N_6308,N_4420,N_5261);
nand U6309 (N_6309,N_4143,N_4582);
nor U6310 (N_6310,N_5201,N_5664);
nor U6311 (N_6311,N_4070,N_4093);
and U6312 (N_6312,N_4755,N_5639);
or U6313 (N_6313,N_4117,N_4226);
or U6314 (N_6314,N_4985,N_4502);
or U6315 (N_6315,N_4342,N_4366);
nor U6316 (N_6316,N_5594,N_5408);
nand U6317 (N_6317,N_4438,N_5700);
nand U6318 (N_6318,N_4914,N_4278);
nor U6319 (N_6319,N_4873,N_5209);
and U6320 (N_6320,N_4685,N_5075);
nor U6321 (N_6321,N_4639,N_4584);
nand U6322 (N_6322,N_4431,N_5605);
nor U6323 (N_6323,N_4750,N_5846);
and U6324 (N_6324,N_4076,N_5316);
nand U6325 (N_6325,N_5894,N_4659);
nor U6326 (N_6326,N_4285,N_4515);
and U6327 (N_6327,N_5535,N_5235);
nand U6328 (N_6328,N_4468,N_4689);
and U6329 (N_6329,N_4455,N_5327);
nor U6330 (N_6330,N_5931,N_5600);
and U6331 (N_6331,N_5275,N_4705);
nand U6332 (N_6332,N_5433,N_5673);
nor U6333 (N_6333,N_5202,N_5361);
or U6334 (N_6334,N_4059,N_5363);
or U6335 (N_6335,N_4892,N_5690);
or U6336 (N_6336,N_4739,N_5355);
nor U6337 (N_6337,N_4661,N_5501);
or U6338 (N_6338,N_5878,N_4370);
and U6339 (N_6339,N_5943,N_5273);
nor U6340 (N_6340,N_5557,N_4071);
and U6341 (N_6341,N_5683,N_5449);
and U6342 (N_6342,N_4033,N_4698);
nand U6343 (N_6343,N_4454,N_5399);
nor U6344 (N_6344,N_4636,N_5080);
nand U6345 (N_6345,N_4483,N_5948);
or U6346 (N_6346,N_4997,N_5074);
nand U6347 (N_6347,N_4246,N_5081);
and U6348 (N_6348,N_4590,N_4677);
and U6349 (N_6349,N_5533,N_4961);
nand U6350 (N_6350,N_4477,N_4895);
and U6351 (N_6351,N_5907,N_4972);
nor U6352 (N_6352,N_4397,N_5335);
xor U6353 (N_6353,N_4671,N_4993);
or U6354 (N_6354,N_4324,N_4496);
nor U6355 (N_6355,N_5150,N_5895);
nor U6356 (N_6356,N_5049,N_4035);
and U6357 (N_6357,N_4186,N_4745);
and U6358 (N_6358,N_5103,N_4247);
nand U6359 (N_6359,N_5678,N_5905);
and U6360 (N_6360,N_5891,N_5956);
nor U6361 (N_6361,N_4611,N_4480);
and U6362 (N_6362,N_4663,N_5826);
and U6363 (N_6363,N_5597,N_5656);
or U6364 (N_6364,N_4711,N_4051);
or U6365 (N_6365,N_5426,N_5632);
nor U6366 (N_6366,N_5384,N_4665);
and U6367 (N_6367,N_4112,N_4181);
xor U6368 (N_6368,N_4074,N_5120);
nand U6369 (N_6369,N_4442,N_4362);
nor U6370 (N_6370,N_5681,N_4890);
and U6371 (N_6371,N_5589,N_5684);
nor U6372 (N_6372,N_4934,N_5012);
and U6373 (N_6373,N_4244,N_4864);
nor U6374 (N_6374,N_4645,N_4316);
nand U6375 (N_6375,N_4736,N_5157);
and U6376 (N_6376,N_4096,N_5008);
or U6377 (N_6377,N_5165,N_4825);
or U6378 (N_6378,N_5329,N_5247);
and U6379 (N_6379,N_5174,N_5068);
nand U6380 (N_6380,N_4038,N_5628);
or U6381 (N_6381,N_4357,N_4937);
nor U6382 (N_6382,N_4089,N_4709);
or U6383 (N_6383,N_4871,N_5647);
or U6384 (N_6384,N_4794,N_5675);
and U6385 (N_6385,N_5999,N_4430);
and U6386 (N_6386,N_4940,N_4883);
nor U6387 (N_6387,N_5822,N_5532);
and U6388 (N_6388,N_5880,N_4933);
and U6389 (N_6389,N_5162,N_4625);
and U6390 (N_6390,N_5699,N_4615);
nand U6391 (N_6391,N_5113,N_5114);
nand U6392 (N_6392,N_4583,N_4696);
nand U6393 (N_6393,N_4140,N_5862);
nand U6394 (N_6394,N_5149,N_5616);
nand U6395 (N_6395,N_5772,N_4017);
nor U6396 (N_6396,N_4862,N_5640);
nor U6397 (N_6397,N_5386,N_4204);
or U6398 (N_6398,N_4405,N_4060);
or U6399 (N_6399,N_5946,N_5596);
and U6400 (N_6400,N_5462,N_5724);
and U6401 (N_6401,N_4968,N_5010);
nor U6402 (N_6402,N_4388,N_5602);
nand U6403 (N_6403,N_5593,N_4616);
or U6404 (N_6404,N_4305,N_4152);
nand U6405 (N_6405,N_5524,N_5315);
nand U6406 (N_6406,N_5930,N_5032);
or U6407 (N_6407,N_4857,N_4925);
or U6408 (N_6408,N_4183,N_4154);
nand U6409 (N_6409,N_4808,N_5941);
and U6410 (N_6410,N_5036,N_4025);
nor U6411 (N_6411,N_4530,N_4007);
nor U6412 (N_6412,N_5001,N_4906);
and U6413 (N_6413,N_5497,N_4451);
nand U6414 (N_6414,N_5923,N_4510);
or U6415 (N_6415,N_4807,N_5129);
and U6416 (N_6416,N_4380,N_5997);
xnor U6417 (N_6417,N_4233,N_4361);
and U6418 (N_6418,N_4831,N_4008);
or U6419 (N_6419,N_5005,N_5511);
nand U6420 (N_6420,N_4942,N_5422);
or U6421 (N_6421,N_4229,N_5296);
nand U6422 (N_6422,N_4176,N_4359);
or U6423 (N_6423,N_4644,N_5056);
nor U6424 (N_6424,N_5541,N_4729);
nor U6425 (N_6425,N_4493,N_5489);
nand U6426 (N_6426,N_5205,N_5783);
nand U6427 (N_6427,N_5741,N_4297);
or U6428 (N_6428,N_4293,N_5549);
nand U6429 (N_6429,N_4044,N_4290);
or U6430 (N_6430,N_4522,N_4027);
or U6431 (N_6431,N_5070,N_4260);
or U6432 (N_6432,N_4800,N_4258);
nand U6433 (N_6433,N_4979,N_4561);
or U6434 (N_6434,N_4632,N_5458);
or U6435 (N_6435,N_5318,N_5756);
nor U6436 (N_6436,N_4032,N_4971);
nand U6437 (N_6437,N_5651,N_4167);
and U6438 (N_6438,N_5094,N_4202);
nand U6439 (N_6439,N_4912,N_5791);
nand U6440 (N_6440,N_4343,N_5727);
or U6441 (N_6441,N_4740,N_4083);
nand U6442 (N_6442,N_4222,N_4878);
nand U6443 (N_6443,N_5638,N_5402);
and U6444 (N_6444,N_5798,N_4572);
nand U6445 (N_6445,N_5427,N_5131);
and U6446 (N_6446,N_4127,N_5709);
nand U6447 (N_6447,N_4752,N_4918);
nor U6448 (N_6448,N_4754,N_4092);
nand U6449 (N_6449,N_4434,N_5495);
and U6450 (N_6450,N_4163,N_4668);
nand U6451 (N_6451,N_5371,N_4945);
nand U6452 (N_6452,N_4805,N_5968);
or U6453 (N_6453,N_4868,N_4019);
or U6454 (N_6454,N_5858,N_5450);
or U6455 (N_6455,N_5262,N_5635);
or U6456 (N_6456,N_4126,N_5021);
nand U6457 (N_6457,N_5617,N_5764);
nand U6458 (N_6458,N_4398,N_5284);
or U6459 (N_6459,N_4102,N_4924);
or U6460 (N_6460,N_4956,N_4780);
or U6461 (N_6461,N_5851,N_4337);
nor U6462 (N_6462,N_4622,N_4602);
nor U6463 (N_6463,N_5534,N_4731);
and U6464 (N_6464,N_4171,N_5176);
nor U6465 (N_6465,N_4549,N_5546);
nand U6466 (N_6466,N_5796,N_5687);
nand U6467 (N_6467,N_5125,N_4779);
nor U6468 (N_6468,N_4016,N_4256);
nand U6469 (N_6469,N_4987,N_4046);
or U6470 (N_6470,N_4271,N_5928);
nand U6471 (N_6471,N_5233,N_5083);
or U6472 (N_6472,N_5052,N_4702);
and U6473 (N_6473,N_5042,N_5254);
or U6474 (N_6474,N_4338,N_4002);
and U6475 (N_6475,N_5998,N_4509);
and U6476 (N_6476,N_5754,N_5477);
and U6477 (N_6477,N_4479,N_5661);
nand U6478 (N_6478,N_4748,N_5740);
nor U6479 (N_6479,N_4322,N_4775);
nor U6480 (N_6480,N_4486,N_5146);
or U6481 (N_6481,N_4219,N_4577);
nand U6482 (N_6482,N_4218,N_4082);
nor U6483 (N_6483,N_4605,N_5531);
nor U6484 (N_6484,N_4168,N_4462);
or U6485 (N_6485,N_4943,N_4694);
nor U6486 (N_6486,N_4328,N_4291);
nor U6487 (N_6487,N_5470,N_4911);
and U6488 (N_6488,N_5586,N_5250);
nand U6489 (N_6489,N_4371,N_5183);
nand U6490 (N_6490,N_4660,N_5592);
xor U6491 (N_6491,N_5451,N_4198);
nor U6492 (N_6492,N_4962,N_5962);
and U6493 (N_6493,N_5810,N_5180);
nand U6494 (N_6494,N_4877,N_5759);
nor U6495 (N_6495,N_5573,N_5845);
nand U6496 (N_6496,N_5652,N_5817);
nor U6497 (N_6497,N_4821,N_5732);
xnor U6498 (N_6498,N_5908,N_4135);
or U6499 (N_6499,N_4209,N_4320);
or U6500 (N_6500,N_5552,N_5621);
nand U6501 (N_6501,N_5809,N_4157);
and U6502 (N_6502,N_4631,N_4588);
and U6503 (N_6503,N_5737,N_5629);
and U6504 (N_6504,N_4321,N_5312);
or U6505 (N_6505,N_5774,N_5122);
and U6506 (N_6506,N_5352,N_5456);
xor U6507 (N_6507,N_4598,N_5581);
nor U6508 (N_6508,N_4352,N_4587);
or U6509 (N_6509,N_5500,N_4500);
and U6510 (N_6510,N_4077,N_4459);
nor U6511 (N_6511,N_4458,N_5782);
and U6512 (N_6512,N_5751,N_5107);
and U6513 (N_6513,N_4063,N_4394);
nand U6514 (N_6514,N_5610,N_5818);
nand U6515 (N_6515,N_4951,N_4580);
nand U6516 (N_6516,N_4384,N_5159);
or U6517 (N_6517,N_5670,N_5290);
nand U6518 (N_6518,N_4189,N_4094);
or U6519 (N_6519,N_4449,N_5442);
nor U6520 (N_6520,N_4633,N_5743);
or U6521 (N_6521,N_4643,N_5513);
nor U6522 (N_6522,N_5964,N_5515);
or U6523 (N_6523,N_5455,N_5657);
and U6524 (N_6524,N_5860,N_5374);
nand U6525 (N_6525,N_5896,N_5692);
or U6526 (N_6526,N_4049,N_5630);
and U6527 (N_6527,N_4248,N_5780);
and U6528 (N_6528,N_4589,N_4768);
nor U6529 (N_6529,N_5116,N_5672);
nand U6530 (N_6530,N_5375,N_5627);
nor U6531 (N_6531,N_5736,N_5303);
nor U6532 (N_6532,N_4547,N_4954);
or U6533 (N_6533,N_5976,N_5643);
or U6534 (N_6534,N_4684,N_4558);
nand U6535 (N_6535,N_4680,N_5357);
nand U6536 (N_6536,N_5170,N_4566);
and U6537 (N_6537,N_5463,N_4936);
or U6538 (N_6538,N_4422,N_5309);
or U6539 (N_6539,N_5220,N_5570);
nand U6540 (N_6540,N_5876,N_5295);
nand U6541 (N_6541,N_5364,N_4579);
or U6542 (N_6542,N_5257,N_5886);
and U6543 (N_6543,N_4921,N_5333);
and U6544 (N_6544,N_4245,N_5265);
nand U6545 (N_6545,N_5404,N_4591);
and U6546 (N_6546,N_4251,N_4111);
or U6547 (N_6547,N_4815,N_4487);
and U6548 (N_6548,N_5857,N_5126);
and U6549 (N_6549,N_5892,N_5117);
or U6550 (N_6550,N_4236,N_4416);
or U6551 (N_6551,N_5718,N_4289);
or U6552 (N_6552,N_4440,N_4681);
or U6553 (N_6553,N_5562,N_5223);
nor U6554 (N_6554,N_5499,N_5750);
nor U6555 (N_6555,N_4028,N_5722);
or U6556 (N_6556,N_4904,N_5475);
nor U6557 (N_6557,N_4410,N_4941);
nor U6558 (N_6558,N_4802,N_4131);
or U6559 (N_6559,N_5134,N_5613);
and U6560 (N_6560,N_4608,N_5031);
and U6561 (N_6561,N_4332,N_4464);
nand U6562 (N_6562,N_5883,N_4523);
nor U6563 (N_6563,N_4726,N_5994);
nand U6564 (N_6564,N_4700,N_4123);
nand U6565 (N_6565,N_5618,N_4662);
nand U6566 (N_6566,N_4756,N_4485);
nor U6567 (N_6567,N_5662,N_4220);
and U6568 (N_6568,N_5246,N_5519);
and U6569 (N_6569,N_4298,N_4269);
nand U6570 (N_6570,N_5815,N_4347);
or U6571 (N_6571,N_5934,N_5714);
or U6572 (N_6572,N_5808,N_4048);
or U6573 (N_6573,N_5269,N_4178);
and U6574 (N_6574,N_5520,N_5940);
nor U6575 (N_6575,N_4106,N_5401);
nand U6576 (N_6576,N_5812,N_4833);
and U6577 (N_6577,N_4551,N_5234);
or U6578 (N_6578,N_4301,N_5385);
and U6579 (N_6579,N_4286,N_5801);
nor U6580 (N_6580,N_5091,N_5506);
or U6581 (N_6581,N_4900,N_5219);
nor U6582 (N_6582,N_5480,N_5775);
and U6583 (N_6583,N_4200,N_5206);
nand U6584 (N_6584,N_5251,N_4704);
xnor U6585 (N_6585,N_4568,N_4674);
or U6586 (N_6586,N_5900,N_5341);
and U6587 (N_6587,N_5398,N_4776);
nor U6588 (N_6588,N_5121,N_4501);
or U6589 (N_6589,N_5967,N_4210);
or U6590 (N_6590,N_4851,N_5359);
and U6591 (N_6591,N_4613,N_4607);
nor U6592 (N_6592,N_5814,N_5369);
or U6593 (N_6593,N_5972,N_4901);
or U6594 (N_6594,N_4351,N_5569);
xor U6595 (N_6595,N_5642,N_4543);
and U6596 (N_6596,N_5821,N_4079);
xor U6597 (N_6597,N_4738,N_5118);
or U6598 (N_6598,N_5016,N_5865);
or U6599 (N_6599,N_4846,N_4022);
or U6600 (N_6600,N_4801,N_5258);
and U6601 (N_6601,N_5072,N_4348);
or U6602 (N_6602,N_4188,N_5204);
nand U6603 (N_6603,N_4992,N_5528);
nand U6604 (N_6604,N_4013,N_4691);
nor U6605 (N_6605,N_4642,N_5757);
nand U6606 (N_6606,N_5824,N_5788);
nor U6607 (N_6607,N_4182,N_4550);
and U6608 (N_6608,N_4021,N_4184);
and U6609 (N_6609,N_5760,N_5749);
nand U6610 (N_6610,N_5379,N_4716);
and U6611 (N_6611,N_4179,N_5027);
nand U6612 (N_6612,N_5332,N_5996);
nor U6613 (N_6613,N_5452,N_5502);
or U6614 (N_6614,N_5071,N_4223);
and U6615 (N_6615,N_4026,N_4852);
or U6616 (N_6616,N_4407,N_5887);
nand U6617 (N_6617,N_4174,N_5467);
nor U6618 (N_6618,N_5286,N_4390);
and U6619 (N_6619,N_4404,N_4759);
nor U6620 (N_6620,N_5437,N_4521);
and U6621 (N_6621,N_5389,N_4137);
nand U6622 (N_6622,N_4771,N_5208);
and U6623 (N_6623,N_5761,N_5985);
and U6624 (N_6624,N_4469,N_4922);
nand U6625 (N_6625,N_4385,N_4923);
nor U6626 (N_6626,N_5582,N_5648);
nor U6627 (N_6627,N_4311,N_4640);
or U6628 (N_6628,N_5167,N_5889);
nand U6629 (N_6629,N_5192,N_5790);
and U6630 (N_6630,N_4811,N_4724);
nor U6631 (N_6631,N_5186,N_5975);
or U6632 (N_6632,N_5348,N_5339);
nand U6633 (N_6633,N_4919,N_4379);
nor U6634 (N_6634,N_5961,N_5841);
or U6635 (N_6635,N_4266,N_4893);
nor U6636 (N_6636,N_5945,N_4929);
or U6637 (N_6637,N_5555,N_4977);
and U6638 (N_6638,N_4612,N_4586);
nand U6639 (N_6639,N_4601,N_4403);
and U6640 (N_6640,N_5553,N_4191);
and U6641 (N_6641,N_5507,N_4938);
or U6642 (N_6642,N_5938,N_4444);
xor U6643 (N_6643,N_4570,N_5566);
or U6644 (N_6644,N_5619,N_5428);
nand U6645 (N_6645,N_4402,N_4192);
or U6646 (N_6646,N_5921,N_5381);
or U6647 (N_6647,N_4818,N_4637);
nor U6648 (N_6648,N_4785,N_5443);
and U6649 (N_6649,N_5242,N_4393);
nand U6650 (N_6650,N_4683,N_5248);
nor U6651 (N_6651,N_4855,N_4850);
or U6652 (N_6652,N_5087,N_5711);
nor U6653 (N_6653,N_4432,N_4953);
nand U6654 (N_6654,N_5526,N_4565);
nand U6655 (N_6655,N_4099,N_5366);
or U6656 (N_6656,N_5464,N_4650);
or U6657 (N_6657,N_4657,N_4418);
nor U6658 (N_6658,N_5411,N_5490);
nand U6659 (N_6659,N_4272,N_5659);
or U6660 (N_6660,N_5086,N_4531);
and U6661 (N_6661,N_5046,N_5181);
nor U6662 (N_6662,N_4341,N_5595);
nand U6663 (N_6663,N_5343,N_5721);
or U6664 (N_6664,N_4544,N_4562);
or U6665 (N_6665,N_5322,N_5222);
and U6666 (N_6666,N_4062,N_5663);
nand U6667 (N_6667,N_4104,N_4354);
nor U6668 (N_6668,N_4472,N_4965);
and U6669 (N_6669,N_4567,N_4481);
or U6670 (N_6670,N_5706,N_5323);
nand U6671 (N_6671,N_5276,N_4626);
and U6672 (N_6672,N_5383,N_5195);
nor U6673 (N_6673,N_4720,N_5079);
and U6674 (N_6674,N_5844,N_4853);
and U6675 (N_6675,N_5837,N_4213);
nand U6676 (N_6676,N_5177,N_4409);
and U6677 (N_6677,N_4784,N_4786);
nor U6678 (N_6678,N_4828,N_4413);
nor U6679 (N_6679,N_5666,N_5133);
and U6680 (N_6680,N_5050,N_5354);
nor U6681 (N_6681,N_5135,N_5567);
nor U6682 (N_6682,N_4730,N_5697);
and U6683 (N_6683,N_4599,N_4967);
and U6684 (N_6684,N_5076,N_5735);
nand U6685 (N_6685,N_5229,N_5979);
or U6686 (N_6686,N_4982,N_4345);
or U6687 (N_6687,N_4710,N_4470);
and U6688 (N_6688,N_4267,N_5313);
or U6689 (N_6689,N_5266,N_4554);
nor U6690 (N_6690,N_5738,N_5881);
and U6691 (N_6691,N_5272,N_5855);
nand U6692 (N_6692,N_5023,N_4149);
nor U6693 (N_6693,N_5307,N_4777);
nor U6694 (N_6694,N_4499,N_5351);
nand U6695 (N_6695,N_4876,N_5952);
nand U6696 (N_6696,N_5777,N_4050);
or U6697 (N_6697,N_5914,N_4043);
nor U6698 (N_6698,N_5459,N_4791);
nor U6699 (N_6699,N_5545,N_5378);
nor U6700 (N_6700,N_5410,N_4078);
and U6701 (N_6701,N_4789,N_5784);
or U6702 (N_6702,N_4201,N_5988);
and U6703 (N_6703,N_4782,N_5172);
nand U6704 (N_6704,N_4344,N_5360);
or U6705 (N_6705,N_4217,N_5096);
nand U6706 (N_6706,N_4376,N_5130);
nand U6707 (N_6707,N_4423,N_4742);
and U6708 (N_6708,N_4284,N_4989);
and U6709 (N_6709,N_4055,N_4457);
nand U6710 (N_6710,N_4482,N_5325);
and U6711 (N_6711,N_5108,N_5987);
nand U6712 (N_6712,N_5166,N_5104);
or U6713 (N_6713,N_4688,N_5287);
nor U6714 (N_6714,N_5758,N_5346);
nor U6715 (N_6715,N_4203,N_5168);
nor U6716 (N_6716,N_4552,N_5781);
nand U6717 (N_6717,N_5763,N_4648);
nor U6718 (N_6718,N_5277,N_4728);
nor U6719 (N_6719,N_5055,N_4944);
nor U6720 (N_6720,N_5281,N_4891);
and U6721 (N_6721,N_4896,N_4103);
nand U6722 (N_6722,N_4365,N_4935);
nand U6723 (N_6723,N_5773,N_4225);
nor U6724 (N_6724,N_5539,N_4100);
or U6725 (N_6725,N_4363,N_4170);
or U6726 (N_6726,N_4327,N_4679);
nor U6727 (N_6727,N_5691,N_5020);
nor U6728 (N_6728,N_5977,N_4513);
nor U6729 (N_6729,N_4617,N_4389);
and U6730 (N_6730,N_4169,N_5693);
nand U6731 (N_6731,N_4490,N_5816);
nor U6732 (N_6732,N_4939,N_4230);
or U6733 (N_6733,N_5563,N_5936);
nor U6734 (N_6734,N_4315,N_5797);
or U6735 (N_6735,N_5746,N_5143);
nand U6736 (N_6736,N_4774,N_4865);
nor U6737 (N_6737,N_5982,N_5393);
nand U6738 (N_6738,N_5171,N_4275);
or U6739 (N_6739,N_4172,N_5719);
nor U6740 (N_6740,N_4042,N_5048);
nor U6741 (N_6741,N_4816,N_4885);
nor U6742 (N_6742,N_4280,N_5867);
or U6743 (N_6743,N_4313,N_5577);
or U6744 (N_6744,N_4913,N_5288);
nor U6745 (N_6745,N_5794,N_5053);
nand U6746 (N_6746,N_4646,N_5842);
or U6747 (N_6747,N_5163,N_4947);
nor U6748 (N_6748,N_4147,N_5457);
or U6749 (N_6749,N_5598,N_4505);
nand U6750 (N_6750,N_5498,N_5634);
and U6751 (N_6751,N_5806,N_5330);
or U6752 (N_6752,N_4629,N_4718);
nand U6753 (N_6753,N_5807,N_4310);
and U6754 (N_6754,N_5831,N_4690);
nor U6755 (N_6755,N_5025,N_4004);
nand U6756 (N_6756,N_4401,N_5981);
or U6757 (N_6757,N_4129,N_4368);
and U6758 (N_6758,N_5241,N_4747);
or U6759 (N_6759,N_5196,N_4969);
nor U6760 (N_6760,N_5279,N_5418);
nor U6761 (N_6761,N_4446,N_4023);
nand U6762 (N_6762,N_5415,N_4847);
or U6763 (N_6763,N_5406,N_4375);
or U6764 (N_6764,N_5682,N_5885);
and U6765 (N_6765,N_5942,N_5365);
and U6766 (N_6766,N_4541,N_4778);
nor U6767 (N_6767,N_4421,N_5243);
nand U6768 (N_6768,N_5509,N_5294);
and U6769 (N_6769,N_4242,N_4653);
and U6770 (N_6770,N_4973,N_5637);
nor U6771 (N_6771,N_5576,N_4277);
nor U6772 (N_6772,N_4452,N_4628);
nand U6773 (N_6773,N_4980,N_5623);
and U6774 (N_6774,N_5789,N_5356);
nand U6775 (N_6775,N_4812,N_5423);
and U6776 (N_6776,N_4326,N_4466);
or U6777 (N_6777,N_4429,N_4719);
or U6778 (N_6778,N_5139,N_5009);
nor U6779 (N_6779,N_5554,N_5302);
nand U6780 (N_6780,N_5776,N_5496);
and U6781 (N_6781,N_4045,N_4518);
nor U6782 (N_6782,N_4721,N_5358);
nor U6783 (N_6783,N_5377,N_5679);
nor U6784 (N_6784,N_5124,N_4160);
or U6785 (N_6785,N_4866,N_4955);
nand U6786 (N_6786,N_5403,N_5925);
nand U6787 (N_6787,N_4374,N_4766);
or U6788 (N_6788,N_5730,N_4066);
nor U6789 (N_6789,N_4086,N_4309);
or U6790 (N_6790,N_4047,N_5446);
and U6791 (N_6791,N_5271,N_5958);
nand U6792 (N_6792,N_5529,N_4484);
and U6793 (N_6793,N_4506,N_4772);
or U6794 (N_6794,N_4450,N_4101);
nand U6795 (N_6795,N_4118,N_5232);
nand U6796 (N_6796,N_4497,N_5607);
nand U6797 (N_6797,N_5349,N_5482);
or U6798 (N_6798,N_5992,N_4304);
or U6799 (N_6799,N_5765,N_5015);
nor U6800 (N_6800,N_5445,N_5769);
and U6801 (N_6801,N_5409,N_5041);
nand U6802 (N_6802,N_4727,N_4998);
and U6803 (N_6803,N_5633,N_5225);
nand U6804 (N_6804,N_5178,N_4952);
nand U6805 (N_6805,N_4753,N_5142);
or U6806 (N_6806,N_5561,N_4888);
and U6807 (N_6807,N_5550,N_5834);
nor U6808 (N_6808,N_4897,N_4249);
and U6809 (N_6809,N_4270,N_4287);
nand U6810 (N_6810,N_4488,N_5155);
or U6811 (N_6811,N_4898,N_5034);
nand U6812 (N_6812,N_4859,N_4654);
and U6813 (N_6813,N_5560,N_5717);
or U6814 (N_6814,N_5207,N_5256);
and U6815 (N_6815,N_4793,N_4107);
nand U6816 (N_6816,N_4761,N_4528);
nand U6817 (N_6817,N_4870,N_5476);
nor U6818 (N_6818,N_5310,N_4187);
nor U6819 (N_6819,N_5984,N_4018);
and U6820 (N_6820,N_5263,N_5828);
or U6821 (N_6821,N_5413,N_5274);
nand U6822 (N_6822,N_5983,N_4732);
nand U6823 (N_6823,N_5224,N_4234);
or U6824 (N_6824,N_4164,N_4760);
or U6825 (N_6825,N_4372,N_5460);
nor U6826 (N_6826,N_5338,N_4594);
nor U6827 (N_6827,N_5110,N_4538);
and U6828 (N_6828,N_5493,N_5065);
and U6829 (N_6829,N_4803,N_4426);
nor U6830 (N_6830,N_4845,N_5744);
and U6831 (N_6831,N_4119,N_4699);
nor U6832 (N_6832,N_4767,N_4508);
and U6833 (N_6833,N_4303,N_4447);
or U6834 (N_6834,N_5778,N_5583);
nor U6835 (N_6835,N_4212,N_5054);
or U6836 (N_6836,N_5077,N_5447);
nand U6837 (N_6837,N_5326,N_5136);
nand U6838 (N_6838,N_5098,N_5331);
and U6839 (N_6839,N_4052,N_4905);
nand U6840 (N_6840,N_5148,N_5599);
nor U6841 (N_6841,N_5875,N_4725);
or U6842 (N_6842,N_4068,N_5514);
nand U6843 (N_6843,N_4193,N_4319);
or U6844 (N_6844,N_4095,N_5084);
and U6845 (N_6845,N_5986,N_4085);
nor U6846 (N_6846,N_4564,N_5792);
and U6847 (N_6847,N_5444,N_4656);
and U6848 (N_6848,N_4999,N_4676);
nand U6849 (N_6849,N_5920,N_4473);
and U6850 (N_6850,N_5097,N_5752);
nand U6851 (N_6851,N_4770,N_4869);
or U6852 (N_6852,N_5184,N_5491);
and U6853 (N_6853,N_4880,N_4288);
and U6854 (N_6854,N_5829,N_5827);
nor U6855 (N_6855,N_4391,N_4437);
nor U6856 (N_6856,N_4707,N_5805);
or U6857 (N_6857,N_4652,N_4887);
and U6858 (N_6858,N_5658,N_4122);
nand U6859 (N_6859,N_5317,N_4340);
nand U6860 (N_6860,N_4145,N_4715);
or U6861 (N_6861,N_4884,N_5342);
nor U6862 (N_6862,N_4349,N_4717);
and U6863 (N_6863,N_4627,N_4448);
nor U6864 (N_6864,N_5214,N_4783);
or U6865 (N_6865,N_5004,N_5856);
nor U6866 (N_6866,N_5035,N_5572);
or U6867 (N_6867,N_4041,N_5991);
nand U6868 (N_6868,N_5259,N_5453);
and U6869 (N_6869,N_4130,N_4574);
nand U6870 (N_6870,N_4040,N_5059);
and U6871 (N_6871,N_4264,N_4292);
xor U6872 (N_6872,N_4516,N_4057);
and U6873 (N_6873,N_4641,N_5264);
and U6874 (N_6874,N_5115,N_5461);
nor U6875 (N_6875,N_5267,N_5000);
nor U6876 (N_6876,N_5028,N_4798);
and U6877 (N_6877,N_4387,N_5465);
nand U6878 (N_6878,N_4012,N_5707);
nor U6879 (N_6879,N_5859,N_4300);
and U6880 (N_6880,N_4744,N_5565);
nor U6881 (N_6881,N_5283,N_5382);
and U6882 (N_6882,N_5090,N_4722);
nor U6883 (N_6883,N_5197,N_4358);
and U6884 (N_6884,N_5840,N_4461);
nor U6885 (N_6885,N_4503,N_5002);
nor U6886 (N_6886,N_4620,N_5753);
and U6887 (N_6887,N_5556,N_5848);
and U6888 (N_6888,N_4872,N_5154);
or U6889 (N_6889,N_4841,N_4830);
or U6890 (N_6890,N_5770,N_4994);
or U6891 (N_6891,N_4165,N_5916);
nand U6892 (N_6892,N_5863,N_5516);
xnor U6893 (N_6893,N_4138,N_4478);
nand U6894 (N_6894,N_4399,N_4417);
nand U6895 (N_6895,N_4231,N_5944);
nor U6896 (N_6896,N_5211,N_5864);
nor U6897 (N_6897,N_4741,N_4826);
and U6898 (N_6898,N_4669,N_4975);
nand U6899 (N_6899,N_5584,N_5708);
nor U6900 (N_6900,N_5145,N_5655);
nor U6901 (N_6901,N_5872,N_4491);
nand U6902 (N_6902,N_4824,N_5953);
nor U6903 (N_6903,N_4228,N_4001);
nor U6904 (N_6904,N_5400,N_4743);
or U6905 (N_6905,N_5144,N_4227);
nor U6906 (N_6906,N_4983,N_5838);
nand U6907 (N_6907,N_5522,N_4792);
and U6908 (N_6908,N_4984,N_4134);
nor U6909 (N_6909,N_5728,N_5436);
nand U6910 (N_6910,N_5929,N_4206);
or U6911 (N_6911,N_5820,N_4141);
xnor U6912 (N_6912,N_5173,N_5345);
or U6913 (N_6913,N_5585,N_5695);
nor U6914 (N_6914,N_4425,N_5624);
and U6915 (N_6915,N_4822,N_4697);
and U6916 (N_6916,N_4575,N_4958);
or U6917 (N_6917,N_5874,N_5890);
nand U6918 (N_6918,N_4539,N_4988);
nand U6919 (N_6919,N_4039,N_5973);
nand U6920 (N_6920,N_5061,N_5240);
nand U6921 (N_6921,N_5182,N_4350);
or U6922 (N_6922,N_4621,N_4151);
or U6923 (N_6923,N_4010,N_4649);
or U6924 (N_6924,N_5768,N_4819);
or U6925 (N_6925,N_4624,N_5440);
or U6926 (N_6926,N_4214,N_4678);
nor U6927 (N_6927,N_5590,N_4065);
nand U6928 (N_6928,N_5472,N_4559);
or U6929 (N_6929,N_5128,N_5494);
nor U6930 (N_6930,N_4295,N_4571);
or U6931 (N_6931,N_4603,N_4005);
nor U6932 (N_6932,N_5604,N_5237);
xnor U6933 (N_6933,N_5614,N_4419);
nor U6934 (N_6934,N_5013,N_4367);
nand U6935 (N_6935,N_5755,N_4623);
nand U6936 (N_6936,N_4024,N_5685);
nand U6937 (N_6937,N_5558,N_5017);
nor U6938 (N_6938,N_4435,N_4809);
nor U6939 (N_6939,N_4073,N_5213);
nand U6940 (N_6940,N_4268,N_4378);
and U6941 (N_6941,N_4875,N_5435);
or U6942 (N_6942,N_5298,N_5158);
nand U6943 (N_6943,N_4314,N_4535);
nand U6944 (N_6944,N_4014,N_5321);
nor U6945 (N_6945,N_4839,N_4128);
nor U6946 (N_6946,N_5314,N_4600);
and U6947 (N_6947,N_5803,N_5029);
nor U6948 (N_6948,N_5836,N_5014);
or U6949 (N_6949,N_5003,N_4408);
and U6950 (N_6950,N_5231,N_4916);
nand U6951 (N_6951,N_5733,N_5492);
and U6952 (N_6952,N_4909,N_5474);
nand U6953 (N_6953,N_5694,N_4723);
or U6954 (N_6954,N_4569,N_4091);
or U6955 (N_6955,N_4153,N_5370);
nand U6956 (N_6956,N_5425,N_4908);
or U6957 (N_6957,N_4814,N_4894);
and U6958 (N_6958,N_5101,N_5906);
and U6959 (N_6959,N_5417,N_5291);
nor U6960 (N_6960,N_4323,N_5787);
and U6961 (N_6961,N_4132,N_5745);
and U6962 (N_6962,N_4221,N_4346);
or U6963 (N_6963,N_5588,N_4763);
nor U6964 (N_6964,N_4369,N_5236);
and U6965 (N_6965,N_5677,N_5832);
and U6966 (N_6966,N_4067,N_4110);
nand U6967 (N_6967,N_5559,N_5175);
nand U6968 (N_6968,N_4427,N_5026);
and U6969 (N_6969,N_5239,N_5989);
nor U6970 (N_6970,N_4764,N_4553);
nor U6971 (N_6971,N_5705,N_5833);
or U6972 (N_6972,N_5926,N_4250);
nor U6973 (N_6973,N_5123,N_4235);
and U6974 (N_6974,N_5270,N_5579);
and U6975 (N_6975,N_5037,N_4121);
or U6976 (N_6976,N_4746,N_5388);
nand U6977 (N_6977,N_5218,N_5127);
and U6978 (N_6978,N_4634,N_4546);
nand U6979 (N_6979,N_4205,N_4120);
and U6980 (N_6980,N_5870,N_4533);
and U6981 (N_6981,N_5395,N_5608);
nand U6982 (N_6982,N_4382,N_5138);
nand U6983 (N_6983,N_5503,N_5710);
nand U6984 (N_6984,N_5852,N_4377);
nand U6985 (N_6985,N_4436,N_4113);
nor U6986 (N_6986,N_4395,N_5543);
or U6987 (N_6987,N_5668,N_5955);
nor U6988 (N_6988,N_4279,N_4555);
and U6989 (N_6989,N_5226,N_5620);
nor U6990 (N_6990,N_5785,N_4339);
and U6991 (N_6991,N_5591,N_5260);
nor U6992 (N_6992,N_4465,N_4842);
nor U6993 (N_6993,N_5189,N_4475);
or U6994 (N_6994,N_4765,N_5871);
and U6995 (N_6995,N_5199,N_4080);
and U6996 (N_6996,N_5978,N_4263);
nor U6997 (N_6997,N_5786,N_5432);
nor U6998 (N_6998,N_5804,N_5680);
nand U6999 (N_6999,N_4241,N_4259);
and U7000 (N_7000,N_5652,N_4152);
or U7001 (N_7001,N_5448,N_5817);
or U7002 (N_7002,N_4542,N_4253);
nand U7003 (N_7003,N_5606,N_5930);
nand U7004 (N_7004,N_5492,N_5417);
nor U7005 (N_7005,N_4031,N_5309);
and U7006 (N_7006,N_5364,N_4802);
and U7007 (N_7007,N_4807,N_5349);
and U7008 (N_7008,N_4018,N_4555);
nand U7009 (N_7009,N_4344,N_5810);
and U7010 (N_7010,N_5995,N_4094);
nor U7011 (N_7011,N_5729,N_5262);
nand U7012 (N_7012,N_5292,N_5963);
nand U7013 (N_7013,N_5230,N_4629);
nor U7014 (N_7014,N_5110,N_5547);
nand U7015 (N_7015,N_4164,N_5456);
and U7016 (N_7016,N_5413,N_4602);
and U7017 (N_7017,N_4533,N_5013);
nor U7018 (N_7018,N_5719,N_5956);
and U7019 (N_7019,N_5324,N_5526);
and U7020 (N_7020,N_4926,N_5666);
nor U7021 (N_7021,N_4765,N_5063);
nor U7022 (N_7022,N_4694,N_4947);
and U7023 (N_7023,N_5459,N_5681);
nor U7024 (N_7024,N_4376,N_4353);
nand U7025 (N_7025,N_4461,N_5383);
nor U7026 (N_7026,N_5868,N_5032);
nor U7027 (N_7027,N_4415,N_4868);
nand U7028 (N_7028,N_5114,N_4299);
nor U7029 (N_7029,N_5560,N_4864);
nor U7030 (N_7030,N_5205,N_5387);
and U7031 (N_7031,N_5023,N_5973);
or U7032 (N_7032,N_5354,N_4322);
nor U7033 (N_7033,N_5954,N_5853);
and U7034 (N_7034,N_5558,N_4845);
and U7035 (N_7035,N_5011,N_5042);
or U7036 (N_7036,N_5314,N_4293);
nand U7037 (N_7037,N_5595,N_4084);
nor U7038 (N_7038,N_4318,N_4917);
nor U7039 (N_7039,N_5401,N_4944);
and U7040 (N_7040,N_5584,N_5167);
or U7041 (N_7041,N_4613,N_5347);
nand U7042 (N_7042,N_5972,N_4472);
and U7043 (N_7043,N_4010,N_4599);
or U7044 (N_7044,N_5520,N_5004);
or U7045 (N_7045,N_5936,N_4018);
nand U7046 (N_7046,N_4684,N_4157);
nand U7047 (N_7047,N_5802,N_5707);
xnor U7048 (N_7048,N_4811,N_4992);
and U7049 (N_7049,N_5741,N_4646);
nand U7050 (N_7050,N_4835,N_5648);
and U7051 (N_7051,N_5335,N_4289);
and U7052 (N_7052,N_4588,N_4542);
and U7053 (N_7053,N_4376,N_5383);
and U7054 (N_7054,N_4876,N_5701);
nor U7055 (N_7055,N_5943,N_4054);
and U7056 (N_7056,N_5715,N_5573);
and U7057 (N_7057,N_5362,N_4758);
or U7058 (N_7058,N_5639,N_4304);
and U7059 (N_7059,N_5091,N_4427);
nor U7060 (N_7060,N_5428,N_4813);
nor U7061 (N_7061,N_5850,N_4559);
or U7062 (N_7062,N_5477,N_4931);
nor U7063 (N_7063,N_4623,N_5996);
and U7064 (N_7064,N_4360,N_4908);
and U7065 (N_7065,N_5571,N_5430);
or U7066 (N_7066,N_4639,N_4227);
nor U7067 (N_7067,N_5506,N_4240);
nor U7068 (N_7068,N_4782,N_5847);
nor U7069 (N_7069,N_4726,N_4631);
nand U7070 (N_7070,N_4894,N_4761);
nand U7071 (N_7071,N_4884,N_4439);
nor U7072 (N_7072,N_5291,N_5232);
nor U7073 (N_7073,N_4618,N_4488);
and U7074 (N_7074,N_4264,N_5780);
nand U7075 (N_7075,N_5553,N_4483);
or U7076 (N_7076,N_5964,N_4931);
nand U7077 (N_7077,N_4246,N_4913);
and U7078 (N_7078,N_5899,N_5386);
nand U7079 (N_7079,N_5289,N_5696);
nand U7080 (N_7080,N_4141,N_5407);
xnor U7081 (N_7081,N_4605,N_4427);
nand U7082 (N_7082,N_4373,N_4340);
or U7083 (N_7083,N_5511,N_5188);
or U7084 (N_7084,N_5615,N_4048);
nand U7085 (N_7085,N_5145,N_4833);
nor U7086 (N_7086,N_4723,N_4196);
nand U7087 (N_7087,N_5383,N_4926);
nor U7088 (N_7088,N_5089,N_5729);
nor U7089 (N_7089,N_5002,N_4799);
and U7090 (N_7090,N_5524,N_4893);
nand U7091 (N_7091,N_4920,N_5617);
nor U7092 (N_7092,N_5984,N_5480);
and U7093 (N_7093,N_5290,N_4687);
or U7094 (N_7094,N_5168,N_4371);
and U7095 (N_7095,N_5941,N_4374);
nand U7096 (N_7096,N_4516,N_4906);
and U7097 (N_7097,N_4102,N_5404);
or U7098 (N_7098,N_5236,N_4901);
or U7099 (N_7099,N_5703,N_5046);
and U7100 (N_7100,N_5608,N_5108);
nand U7101 (N_7101,N_4829,N_5459);
nor U7102 (N_7102,N_5543,N_4609);
nor U7103 (N_7103,N_5706,N_5066);
nor U7104 (N_7104,N_5853,N_4046);
or U7105 (N_7105,N_5742,N_5234);
and U7106 (N_7106,N_5787,N_4089);
and U7107 (N_7107,N_5967,N_4800);
or U7108 (N_7108,N_5095,N_5385);
or U7109 (N_7109,N_4822,N_5964);
nand U7110 (N_7110,N_5583,N_4533);
and U7111 (N_7111,N_5018,N_4171);
and U7112 (N_7112,N_4755,N_4106);
and U7113 (N_7113,N_5157,N_5639);
and U7114 (N_7114,N_4509,N_5934);
nand U7115 (N_7115,N_5471,N_5041);
and U7116 (N_7116,N_5537,N_5025);
nand U7117 (N_7117,N_4487,N_5310);
or U7118 (N_7118,N_5006,N_4133);
or U7119 (N_7119,N_5627,N_5516);
nand U7120 (N_7120,N_5744,N_4949);
xor U7121 (N_7121,N_4999,N_5769);
nor U7122 (N_7122,N_5213,N_5085);
and U7123 (N_7123,N_5468,N_4181);
xor U7124 (N_7124,N_5427,N_5377);
nand U7125 (N_7125,N_5948,N_4339);
nor U7126 (N_7126,N_5963,N_4246);
or U7127 (N_7127,N_4405,N_5798);
nand U7128 (N_7128,N_5921,N_4961);
nand U7129 (N_7129,N_4789,N_5870);
and U7130 (N_7130,N_4252,N_5248);
nand U7131 (N_7131,N_4677,N_5994);
and U7132 (N_7132,N_4269,N_4189);
and U7133 (N_7133,N_4121,N_5796);
nand U7134 (N_7134,N_5094,N_5462);
nand U7135 (N_7135,N_4357,N_4592);
nand U7136 (N_7136,N_4158,N_4073);
or U7137 (N_7137,N_4904,N_5170);
nand U7138 (N_7138,N_5980,N_5073);
nand U7139 (N_7139,N_4669,N_4691);
nor U7140 (N_7140,N_4921,N_5009);
and U7141 (N_7141,N_4909,N_5738);
and U7142 (N_7142,N_4517,N_5380);
nor U7143 (N_7143,N_5643,N_4140);
nor U7144 (N_7144,N_4333,N_5840);
or U7145 (N_7145,N_5109,N_5693);
nand U7146 (N_7146,N_5412,N_5575);
nor U7147 (N_7147,N_4495,N_5442);
and U7148 (N_7148,N_5019,N_4292);
or U7149 (N_7149,N_5422,N_5363);
or U7150 (N_7150,N_5898,N_4394);
or U7151 (N_7151,N_4312,N_4356);
nand U7152 (N_7152,N_5554,N_4379);
or U7153 (N_7153,N_4821,N_5629);
or U7154 (N_7154,N_4605,N_4409);
nand U7155 (N_7155,N_4357,N_5667);
or U7156 (N_7156,N_4944,N_5192);
or U7157 (N_7157,N_5721,N_4743);
or U7158 (N_7158,N_4942,N_5193);
nor U7159 (N_7159,N_4185,N_4460);
and U7160 (N_7160,N_5614,N_5711);
or U7161 (N_7161,N_4106,N_5720);
or U7162 (N_7162,N_5798,N_4551);
and U7163 (N_7163,N_5110,N_5785);
nor U7164 (N_7164,N_4822,N_5488);
and U7165 (N_7165,N_4749,N_5003);
or U7166 (N_7166,N_5072,N_5867);
or U7167 (N_7167,N_5958,N_5077);
and U7168 (N_7168,N_4754,N_5325);
nand U7169 (N_7169,N_5596,N_5240);
nand U7170 (N_7170,N_5587,N_4198);
or U7171 (N_7171,N_4014,N_5135);
nor U7172 (N_7172,N_5977,N_5349);
and U7173 (N_7173,N_4744,N_5747);
and U7174 (N_7174,N_4299,N_5948);
nand U7175 (N_7175,N_4639,N_5630);
nor U7176 (N_7176,N_4742,N_4998);
and U7177 (N_7177,N_5805,N_5138);
and U7178 (N_7178,N_5553,N_5402);
nor U7179 (N_7179,N_4739,N_5450);
nand U7180 (N_7180,N_5677,N_5358);
or U7181 (N_7181,N_4791,N_5363);
nand U7182 (N_7182,N_5956,N_5314);
and U7183 (N_7183,N_4225,N_5643);
nand U7184 (N_7184,N_5847,N_4954);
nor U7185 (N_7185,N_5183,N_4576);
nor U7186 (N_7186,N_4284,N_5922);
xnor U7187 (N_7187,N_4543,N_4048);
nand U7188 (N_7188,N_5938,N_4132);
nor U7189 (N_7189,N_5189,N_4786);
nand U7190 (N_7190,N_4377,N_5665);
and U7191 (N_7191,N_5989,N_4397);
nand U7192 (N_7192,N_5205,N_5862);
nand U7193 (N_7193,N_4941,N_4138);
nand U7194 (N_7194,N_4243,N_5328);
xnor U7195 (N_7195,N_4903,N_5308);
nor U7196 (N_7196,N_5080,N_4266);
or U7197 (N_7197,N_5070,N_5100);
or U7198 (N_7198,N_4154,N_4587);
or U7199 (N_7199,N_4781,N_4389);
xor U7200 (N_7200,N_5886,N_4541);
or U7201 (N_7201,N_5111,N_5739);
nand U7202 (N_7202,N_4777,N_5775);
and U7203 (N_7203,N_5783,N_4816);
nand U7204 (N_7204,N_4055,N_4417);
nand U7205 (N_7205,N_4318,N_4014);
nand U7206 (N_7206,N_4422,N_4770);
or U7207 (N_7207,N_4251,N_5959);
xnor U7208 (N_7208,N_4653,N_4136);
and U7209 (N_7209,N_4228,N_4004);
nand U7210 (N_7210,N_4877,N_4504);
nand U7211 (N_7211,N_5815,N_4579);
or U7212 (N_7212,N_5935,N_4816);
nor U7213 (N_7213,N_5996,N_5352);
or U7214 (N_7214,N_5286,N_5053);
and U7215 (N_7215,N_4959,N_5611);
nor U7216 (N_7216,N_4535,N_5037);
nor U7217 (N_7217,N_5843,N_4932);
or U7218 (N_7218,N_5592,N_4560);
and U7219 (N_7219,N_5961,N_5790);
nand U7220 (N_7220,N_5548,N_5033);
nand U7221 (N_7221,N_4149,N_4130);
or U7222 (N_7222,N_4181,N_5815);
or U7223 (N_7223,N_4968,N_5116);
nor U7224 (N_7224,N_4749,N_5074);
or U7225 (N_7225,N_5282,N_5355);
and U7226 (N_7226,N_4366,N_4441);
nand U7227 (N_7227,N_4819,N_4123);
nand U7228 (N_7228,N_4188,N_5923);
nand U7229 (N_7229,N_5330,N_4510);
and U7230 (N_7230,N_4290,N_4101);
nor U7231 (N_7231,N_4051,N_5410);
nand U7232 (N_7232,N_4463,N_4129);
or U7233 (N_7233,N_5808,N_4436);
or U7234 (N_7234,N_4115,N_4440);
or U7235 (N_7235,N_4510,N_4457);
and U7236 (N_7236,N_4196,N_5676);
nor U7237 (N_7237,N_4765,N_4627);
or U7238 (N_7238,N_4145,N_4299);
or U7239 (N_7239,N_4736,N_5595);
nor U7240 (N_7240,N_4454,N_4958);
or U7241 (N_7241,N_4990,N_5396);
nor U7242 (N_7242,N_4398,N_4149);
nor U7243 (N_7243,N_4228,N_4309);
and U7244 (N_7244,N_4332,N_5551);
nand U7245 (N_7245,N_4906,N_4833);
and U7246 (N_7246,N_5571,N_5735);
nor U7247 (N_7247,N_5996,N_5954);
or U7248 (N_7248,N_5735,N_4568);
nand U7249 (N_7249,N_4512,N_4185);
nor U7250 (N_7250,N_4604,N_4831);
or U7251 (N_7251,N_5680,N_4434);
and U7252 (N_7252,N_4432,N_5842);
and U7253 (N_7253,N_4526,N_4688);
nor U7254 (N_7254,N_4256,N_4561);
nand U7255 (N_7255,N_4498,N_5211);
nand U7256 (N_7256,N_5180,N_5989);
nand U7257 (N_7257,N_5528,N_4879);
nor U7258 (N_7258,N_4800,N_5073);
and U7259 (N_7259,N_4402,N_5106);
or U7260 (N_7260,N_4473,N_5225);
xor U7261 (N_7261,N_5828,N_5295);
or U7262 (N_7262,N_5155,N_4522);
or U7263 (N_7263,N_5663,N_5978);
nor U7264 (N_7264,N_4039,N_4701);
or U7265 (N_7265,N_4217,N_5081);
nand U7266 (N_7266,N_5316,N_4495);
nand U7267 (N_7267,N_5909,N_4704);
and U7268 (N_7268,N_4750,N_4888);
or U7269 (N_7269,N_4535,N_4454);
and U7270 (N_7270,N_4609,N_4344);
nand U7271 (N_7271,N_4212,N_4401);
nand U7272 (N_7272,N_4483,N_5892);
nand U7273 (N_7273,N_5969,N_5086);
nand U7274 (N_7274,N_5465,N_5516);
nand U7275 (N_7275,N_5239,N_4113);
nand U7276 (N_7276,N_5336,N_5239);
or U7277 (N_7277,N_4554,N_5340);
nand U7278 (N_7278,N_4966,N_5510);
or U7279 (N_7279,N_5470,N_4614);
nand U7280 (N_7280,N_5919,N_4547);
nand U7281 (N_7281,N_5213,N_5810);
nand U7282 (N_7282,N_4770,N_5031);
nand U7283 (N_7283,N_5786,N_5737);
and U7284 (N_7284,N_4739,N_4501);
nand U7285 (N_7285,N_5081,N_5426);
nor U7286 (N_7286,N_5060,N_5913);
or U7287 (N_7287,N_4235,N_4713);
or U7288 (N_7288,N_5404,N_5941);
nand U7289 (N_7289,N_4907,N_4967);
and U7290 (N_7290,N_5109,N_5397);
and U7291 (N_7291,N_4274,N_4601);
and U7292 (N_7292,N_4665,N_5522);
nor U7293 (N_7293,N_4930,N_4176);
or U7294 (N_7294,N_4636,N_5419);
or U7295 (N_7295,N_4007,N_4349);
nand U7296 (N_7296,N_4270,N_5814);
and U7297 (N_7297,N_5644,N_5389);
nand U7298 (N_7298,N_5060,N_4474);
or U7299 (N_7299,N_4440,N_5554);
nor U7300 (N_7300,N_4957,N_4471);
and U7301 (N_7301,N_4138,N_4528);
nand U7302 (N_7302,N_5987,N_4186);
nor U7303 (N_7303,N_5710,N_5389);
nand U7304 (N_7304,N_4872,N_5964);
or U7305 (N_7305,N_5623,N_4731);
nand U7306 (N_7306,N_5897,N_5338);
and U7307 (N_7307,N_4661,N_5723);
and U7308 (N_7308,N_5177,N_5530);
and U7309 (N_7309,N_4407,N_5614);
or U7310 (N_7310,N_4108,N_4625);
and U7311 (N_7311,N_5745,N_5571);
xor U7312 (N_7312,N_4423,N_4472);
or U7313 (N_7313,N_4537,N_4459);
and U7314 (N_7314,N_5423,N_5771);
nor U7315 (N_7315,N_4151,N_4840);
and U7316 (N_7316,N_4339,N_4457);
nor U7317 (N_7317,N_5539,N_5524);
or U7318 (N_7318,N_5275,N_5752);
and U7319 (N_7319,N_5089,N_4367);
and U7320 (N_7320,N_5764,N_5780);
nor U7321 (N_7321,N_5150,N_4426);
and U7322 (N_7322,N_4369,N_4958);
and U7323 (N_7323,N_5895,N_5280);
or U7324 (N_7324,N_5954,N_5779);
nand U7325 (N_7325,N_4894,N_4589);
or U7326 (N_7326,N_4656,N_5270);
and U7327 (N_7327,N_5299,N_4249);
nand U7328 (N_7328,N_4808,N_5729);
and U7329 (N_7329,N_4431,N_5681);
nand U7330 (N_7330,N_4639,N_4708);
nand U7331 (N_7331,N_5610,N_5169);
nor U7332 (N_7332,N_4810,N_4575);
nand U7333 (N_7333,N_4467,N_5258);
nand U7334 (N_7334,N_5637,N_5399);
nand U7335 (N_7335,N_5637,N_5623);
nand U7336 (N_7336,N_5187,N_5561);
nand U7337 (N_7337,N_4963,N_5030);
or U7338 (N_7338,N_4828,N_5997);
or U7339 (N_7339,N_5669,N_5426);
and U7340 (N_7340,N_4350,N_5474);
and U7341 (N_7341,N_5616,N_5743);
or U7342 (N_7342,N_5461,N_5116);
nand U7343 (N_7343,N_4797,N_4160);
nand U7344 (N_7344,N_5273,N_5928);
nor U7345 (N_7345,N_5527,N_5882);
or U7346 (N_7346,N_4393,N_5800);
xor U7347 (N_7347,N_5976,N_5088);
nor U7348 (N_7348,N_5965,N_4012);
or U7349 (N_7349,N_5766,N_4051);
nand U7350 (N_7350,N_4429,N_5956);
and U7351 (N_7351,N_4737,N_5424);
nand U7352 (N_7352,N_5712,N_5233);
or U7353 (N_7353,N_4585,N_5625);
or U7354 (N_7354,N_5348,N_4788);
nor U7355 (N_7355,N_5900,N_5361);
nand U7356 (N_7356,N_4448,N_4482);
nor U7357 (N_7357,N_4056,N_5763);
or U7358 (N_7358,N_4565,N_4208);
and U7359 (N_7359,N_5880,N_5159);
nand U7360 (N_7360,N_5529,N_5171);
and U7361 (N_7361,N_5738,N_5232);
nand U7362 (N_7362,N_4538,N_4346);
nand U7363 (N_7363,N_4104,N_5001);
nand U7364 (N_7364,N_4704,N_5066);
or U7365 (N_7365,N_4469,N_5473);
or U7366 (N_7366,N_4997,N_4637);
nand U7367 (N_7367,N_5743,N_5745);
nor U7368 (N_7368,N_5461,N_5989);
xor U7369 (N_7369,N_5880,N_5279);
and U7370 (N_7370,N_5167,N_5242);
and U7371 (N_7371,N_5363,N_4276);
nand U7372 (N_7372,N_4920,N_4407);
nand U7373 (N_7373,N_4687,N_5701);
or U7374 (N_7374,N_4579,N_5001);
nor U7375 (N_7375,N_5716,N_5762);
or U7376 (N_7376,N_5613,N_4090);
nand U7377 (N_7377,N_5139,N_5851);
nor U7378 (N_7378,N_4889,N_4480);
or U7379 (N_7379,N_4552,N_5495);
nor U7380 (N_7380,N_5423,N_4228);
or U7381 (N_7381,N_5414,N_5741);
nor U7382 (N_7382,N_4308,N_4469);
or U7383 (N_7383,N_4426,N_4039);
nand U7384 (N_7384,N_4498,N_4327);
and U7385 (N_7385,N_4020,N_5369);
nand U7386 (N_7386,N_4590,N_4729);
nand U7387 (N_7387,N_4015,N_5787);
nand U7388 (N_7388,N_5476,N_5922);
nor U7389 (N_7389,N_4135,N_5683);
nand U7390 (N_7390,N_4484,N_4112);
and U7391 (N_7391,N_4783,N_5866);
nand U7392 (N_7392,N_4700,N_5910);
and U7393 (N_7393,N_4467,N_4704);
nor U7394 (N_7394,N_5424,N_4379);
nand U7395 (N_7395,N_4647,N_4956);
and U7396 (N_7396,N_4393,N_4870);
or U7397 (N_7397,N_5157,N_5958);
and U7398 (N_7398,N_5157,N_5015);
nand U7399 (N_7399,N_5497,N_4856);
and U7400 (N_7400,N_4259,N_4329);
and U7401 (N_7401,N_4293,N_5436);
nand U7402 (N_7402,N_4492,N_4315);
nor U7403 (N_7403,N_5517,N_4824);
or U7404 (N_7404,N_4326,N_4894);
nand U7405 (N_7405,N_4968,N_4035);
or U7406 (N_7406,N_5682,N_4090);
nor U7407 (N_7407,N_4765,N_5610);
nand U7408 (N_7408,N_5073,N_4894);
nand U7409 (N_7409,N_5212,N_4681);
nand U7410 (N_7410,N_4823,N_5337);
nand U7411 (N_7411,N_4824,N_4097);
nor U7412 (N_7412,N_4322,N_4652);
nor U7413 (N_7413,N_4016,N_4664);
or U7414 (N_7414,N_5488,N_4278);
nor U7415 (N_7415,N_5010,N_4679);
nor U7416 (N_7416,N_5917,N_5328);
xnor U7417 (N_7417,N_5529,N_5133);
and U7418 (N_7418,N_5808,N_4618);
nor U7419 (N_7419,N_5041,N_4518);
nor U7420 (N_7420,N_5547,N_5945);
or U7421 (N_7421,N_5441,N_5299);
nor U7422 (N_7422,N_4353,N_5620);
nor U7423 (N_7423,N_5857,N_5353);
nor U7424 (N_7424,N_4279,N_4722);
and U7425 (N_7425,N_5370,N_4113);
nor U7426 (N_7426,N_4776,N_4256);
or U7427 (N_7427,N_5786,N_4889);
nor U7428 (N_7428,N_5117,N_4312);
nor U7429 (N_7429,N_4750,N_4292);
nor U7430 (N_7430,N_5459,N_5042);
nor U7431 (N_7431,N_5278,N_4295);
and U7432 (N_7432,N_4972,N_5519);
or U7433 (N_7433,N_4023,N_4865);
or U7434 (N_7434,N_5087,N_4334);
nand U7435 (N_7435,N_5181,N_5014);
nor U7436 (N_7436,N_5374,N_4708);
nand U7437 (N_7437,N_5893,N_5455);
nand U7438 (N_7438,N_5850,N_4413);
or U7439 (N_7439,N_4260,N_4513);
and U7440 (N_7440,N_4134,N_5159);
and U7441 (N_7441,N_4561,N_5617);
nand U7442 (N_7442,N_4845,N_4648);
or U7443 (N_7443,N_4428,N_4039);
or U7444 (N_7444,N_4226,N_4516);
and U7445 (N_7445,N_4064,N_4126);
nor U7446 (N_7446,N_5052,N_4019);
nand U7447 (N_7447,N_5421,N_5381);
nand U7448 (N_7448,N_4313,N_5238);
nand U7449 (N_7449,N_4726,N_5626);
and U7450 (N_7450,N_4859,N_5366);
or U7451 (N_7451,N_5157,N_4123);
and U7452 (N_7452,N_4521,N_5565);
nor U7453 (N_7453,N_5406,N_4310);
nor U7454 (N_7454,N_5368,N_5928);
or U7455 (N_7455,N_4753,N_5275);
and U7456 (N_7456,N_5868,N_5585);
or U7457 (N_7457,N_4257,N_4289);
and U7458 (N_7458,N_5478,N_5734);
nand U7459 (N_7459,N_4850,N_5462);
nor U7460 (N_7460,N_5498,N_4988);
nand U7461 (N_7461,N_5163,N_5985);
or U7462 (N_7462,N_4639,N_4257);
nor U7463 (N_7463,N_5169,N_4211);
and U7464 (N_7464,N_4580,N_5172);
nand U7465 (N_7465,N_5744,N_5503);
and U7466 (N_7466,N_5184,N_5277);
or U7467 (N_7467,N_4102,N_4014);
and U7468 (N_7468,N_4670,N_4049);
and U7469 (N_7469,N_4230,N_4058);
nor U7470 (N_7470,N_4517,N_4406);
nor U7471 (N_7471,N_5221,N_5359);
nand U7472 (N_7472,N_5423,N_4081);
and U7473 (N_7473,N_5929,N_5835);
or U7474 (N_7474,N_4407,N_4717);
nand U7475 (N_7475,N_5765,N_5672);
nand U7476 (N_7476,N_4474,N_5561);
or U7477 (N_7477,N_5627,N_4748);
nor U7478 (N_7478,N_5332,N_4889);
or U7479 (N_7479,N_5155,N_5805);
nor U7480 (N_7480,N_4628,N_5052);
nor U7481 (N_7481,N_5059,N_5736);
nand U7482 (N_7482,N_5325,N_4907);
or U7483 (N_7483,N_4868,N_5009);
and U7484 (N_7484,N_4267,N_5852);
or U7485 (N_7485,N_5881,N_4161);
or U7486 (N_7486,N_4404,N_5707);
nand U7487 (N_7487,N_5595,N_4052);
and U7488 (N_7488,N_4228,N_4784);
nor U7489 (N_7489,N_4181,N_4546);
nor U7490 (N_7490,N_4215,N_4401);
nand U7491 (N_7491,N_4987,N_4425);
and U7492 (N_7492,N_5658,N_5671);
or U7493 (N_7493,N_5944,N_5219);
nor U7494 (N_7494,N_5273,N_5775);
and U7495 (N_7495,N_5092,N_4328);
or U7496 (N_7496,N_5353,N_5596);
nand U7497 (N_7497,N_4005,N_4846);
nand U7498 (N_7498,N_4293,N_4219);
nor U7499 (N_7499,N_4590,N_5359);
nand U7500 (N_7500,N_5737,N_4406);
nor U7501 (N_7501,N_4933,N_5128);
nor U7502 (N_7502,N_5733,N_5717);
or U7503 (N_7503,N_4026,N_4546);
or U7504 (N_7504,N_4877,N_5614);
nor U7505 (N_7505,N_4711,N_4900);
nand U7506 (N_7506,N_5088,N_5545);
or U7507 (N_7507,N_4579,N_4815);
and U7508 (N_7508,N_4939,N_4428);
or U7509 (N_7509,N_4024,N_5054);
and U7510 (N_7510,N_4697,N_4947);
nor U7511 (N_7511,N_5297,N_5242);
or U7512 (N_7512,N_4302,N_4806);
nand U7513 (N_7513,N_5448,N_5857);
nand U7514 (N_7514,N_5177,N_4890);
nand U7515 (N_7515,N_4371,N_4063);
nand U7516 (N_7516,N_4854,N_5780);
and U7517 (N_7517,N_5553,N_5526);
nor U7518 (N_7518,N_5680,N_4670);
and U7519 (N_7519,N_5265,N_4132);
nand U7520 (N_7520,N_4775,N_5085);
nor U7521 (N_7521,N_4911,N_5327);
nor U7522 (N_7522,N_4960,N_4683);
and U7523 (N_7523,N_5764,N_4150);
nand U7524 (N_7524,N_4051,N_4016);
and U7525 (N_7525,N_5057,N_4687);
or U7526 (N_7526,N_4599,N_5543);
or U7527 (N_7527,N_5117,N_4539);
and U7528 (N_7528,N_4929,N_5570);
or U7529 (N_7529,N_4053,N_5780);
and U7530 (N_7530,N_5857,N_5026);
nand U7531 (N_7531,N_5012,N_4907);
nand U7532 (N_7532,N_5150,N_5902);
or U7533 (N_7533,N_4460,N_5034);
nand U7534 (N_7534,N_4202,N_4756);
nor U7535 (N_7535,N_4400,N_4132);
nand U7536 (N_7536,N_4839,N_5526);
nand U7537 (N_7537,N_4456,N_4409);
nand U7538 (N_7538,N_4281,N_5077);
and U7539 (N_7539,N_4227,N_4570);
nand U7540 (N_7540,N_4305,N_5446);
xnor U7541 (N_7541,N_4078,N_5406);
nand U7542 (N_7542,N_4284,N_4283);
nor U7543 (N_7543,N_5990,N_4225);
nand U7544 (N_7544,N_4567,N_4296);
or U7545 (N_7545,N_4390,N_5009);
nor U7546 (N_7546,N_4354,N_4584);
and U7547 (N_7547,N_5332,N_5288);
and U7548 (N_7548,N_4886,N_4628);
nand U7549 (N_7549,N_5610,N_5033);
nor U7550 (N_7550,N_5145,N_4323);
xor U7551 (N_7551,N_5593,N_5827);
and U7552 (N_7552,N_5343,N_4994);
nor U7553 (N_7553,N_5925,N_5780);
nand U7554 (N_7554,N_5022,N_5468);
nor U7555 (N_7555,N_4535,N_5212);
nor U7556 (N_7556,N_4253,N_5476);
or U7557 (N_7557,N_5366,N_5077);
nand U7558 (N_7558,N_5191,N_5251);
nand U7559 (N_7559,N_5228,N_4734);
or U7560 (N_7560,N_4513,N_4662);
nor U7561 (N_7561,N_5198,N_5177);
or U7562 (N_7562,N_5697,N_5338);
or U7563 (N_7563,N_4414,N_5360);
nand U7564 (N_7564,N_4082,N_5485);
nand U7565 (N_7565,N_4124,N_5699);
nor U7566 (N_7566,N_4907,N_5277);
and U7567 (N_7567,N_5021,N_4833);
nand U7568 (N_7568,N_5014,N_4184);
or U7569 (N_7569,N_5373,N_4272);
or U7570 (N_7570,N_5221,N_5961);
and U7571 (N_7571,N_4126,N_4253);
xnor U7572 (N_7572,N_5981,N_4173);
nand U7573 (N_7573,N_5374,N_5029);
nand U7574 (N_7574,N_4155,N_5237);
and U7575 (N_7575,N_4716,N_5108);
or U7576 (N_7576,N_4840,N_5467);
nand U7577 (N_7577,N_5853,N_4966);
or U7578 (N_7578,N_4242,N_5213);
nor U7579 (N_7579,N_4823,N_4129);
nand U7580 (N_7580,N_4110,N_5219);
nand U7581 (N_7581,N_5582,N_4814);
or U7582 (N_7582,N_4657,N_4956);
nand U7583 (N_7583,N_5928,N_5853);
and U7584 (N_7584,N_4359,N_5019);
or U7585 (N_7585,N_4803,N_4885);
nand U7586 (N_7586,N_4778,N_5635);
nand U7587 (N_7587,N_5825,N_5795);
and U7588 (N_7588,N_5502,N_4430);
or U7589 (N_7589,N_5921,N_4180);
nand U7590 (N_7590,N_4656,N_5720);
or U7591 (N_7591,N_5321,N_5433);
and U7592 (N_7592,N_4902,N_5143);
nor U7593 (N_7593,N_4354,N_5101);
and U7594 (N_7594,N_5694,N_4664);
and U7595 (N_7595,N_5297,N_4036);
or U7596 (N_7596,N_5149,N_4172);
and U7597 (N_7597,N_5418,N_5918);
nor U7598 (N_7598,N_4684,N_4514);
nand U7599 (N_7599,N_4121,N_5099);
nand U7600 (N_7600,N_4540,N_5914);
or U7601 (N_7601,N_4187,N_5627);
nand U7602 (N_7602,N_5080,N_5658);
or U7603 (N_7603,N_4468,N_5603);
and U7604 (N_7604,N_5021,N_4606);
nor U7605 (N_7605,N_4865,N_4244);
or U7606 (N_7606,N_5762,N_4588);
or U7607 (N_7607,N_5203,N_4987);
nor U7608 (N_7608,N_4657,N_5406);
nor U7609 (N_7609,N_5984,N_4700);
nor U7610 (N_7610,N_4078,N_4498);
and U7611 (N_7611,N_5983,N_4936);
nor U7612 (N_7612,N_5827,N_5318);
or U7613 (N_7613,N_4316,N_5136);
and U7614 (N_7614,N_4185,N_4462);
and U7615 (N_7615,N_5212,N_5530);
nor U7616 (N_7616,N_4449,N_4391);
nand U7617 (N_7617,N_4466,N_5293);
nand U7618 (N_7618,N_5519,N_4799);
or U7619 (N_7619,N_4235,N_5021);
or U7620 (N_7620,N_4215,N_4300);
or U7621 (N_7621,N_4912,N_4796);
and U7622 (N_7622,N_5931,N_4530);
or U7623 (N_7623,N_5903,N_4644);
nor U7624 (N_7624,N_5014,N_5003);
or U7625 (N_7625,N_5768,N_4644);
nor U7626 (N_7626,N_5306,N_4996);
nor U7627 (N_7627,N_5324,N_4978);
nand U7628 (N_7628,N_4980,N_4376);
and U7629 (N_7629,N_4413,N_5866);
and U7630 (N_7630,N_5155,N_4773);
nand U7631 (N_7631,N_4932,N_5443);
and U7632 (N_7632,N_5054,N_5396);
nand U7633 (N_7633,N_5204,N_5810);
and U7634 (N_7634,N_5677,N_5712);
nand U7635 (N_7635,N_4075,N_5811);
and U7636 (N_7636,N_4401,N_5146);
and U7637 (N_7637,N_5198,N_5502);
and U7638 (N_7638,N_5534,N_5228);
or U7639 (N_7639,N_4071,N_4472);
and U7640 (N_7640,N_5903,N_4421);
nand U7641 (N_7641,N_5680,N_5828);
and U7642 (N_7642,N_5371,N_4508);
nor U7643 (N_7643,N_5522,N_5683);
nand U7644 (N_7644,N_5964,N_4146);
or U7645 (N_7645,N_4232,N_4815);
nor U7646 (N_7646,N_4835,N_5518);
nor U7647 (N_7647,N_4615,N_5441);
and U7648 (N_7648,N_4960,N_4500);
nor U7649 (N_7649,N_5562,N_5361);
or U7650 (N_7650,N_5093,N_4356);
and U7651 (N_7651,N_5625,N_5544);
nor U7652 (N_7652,N_4993,N_4058);
nor U7653 (N_7653,N_4231,N_5792);
or U7654 (N_7654,N_4758,N_4186);
or U7655 (N_7655,N_5890,N_4999);
nand U7656 (N_7656,N_5394,N_5659);
and U7657 (N_7657,N_5164,N_5710);
and U7658 (N_7658,N_4507,N_5711);
or U7659 (N_7659,N_5346,N_5780);
and U7660 (N_7660,N_5898,N_5015);
nand U7661 (N_7661,N_4570,N_5627);
or U7662 (N_7662,N_5307,N_4204);
and U7663 (N_7663,N_5618,N_4393);
or U7664 (N_7664,N_5283,N_4995);
nor U7665 (N_7665,N_4913,N_5870);
or U7666 (N_7666,N_5665,N_4086);
nand U7667 (N_7667,N_5959,N_4611);
nand U7668 (N_7668,N_5645,N_5015);
nor U7669 (N_7669,N_4558,N_4658);
nand U7670 (N_7670,N_5111,N_4997);
nand U7671 (N_7671,N_4483,N_4816);
and U7672 (N_7672,N_4014,N_5760);
or U7673 (N_7673,N_4076,N_4665);
or U7674 (N_7674,N_5013,N_4184);
nand U7675 (N_7675,N_5537,N_5439);
or U7676 (N_7676,N_4958,N_4303);
nor U7677 (N_7677,N_5510,N_5052);
nand U7678 (N_7678,N_4284,N_4723);
nor U7679 (N_7679,N_4536,N_5512);
or U7680 (N_7680,N_4532,N_5520);
nor U7681 (N_7681,N_5241,N_4661);
and U7682 (N_7682,N_5509,N_4189);
nand U7683 (N_7683,N_4728,N_5371);
and U7684 (N_7684,N_5689,N_4614);
xnor U7685 (N_7685,N_5440,N_4504);
or U7686 (N_7686,N_5705,N_4654);
and U7687 (N_7687,N_5358,N_5008);
or U7688 (N_7688,N_5867,N_4627);
and U7689 (N_7689,N_4778,N_4719);
and U7690 (N_7690,N_5312,N_5989);
nor U7691 (N_7691,N_5372,N_5751);
or U7692 (N_7692,N_4097,N_4667);
nand U7693 (N_7693,N_4301,N_4585);
or U7694 (N_7694,N_4186,N_5269);
nand U7695 (N_7695,N_5902,N_4312);
and U7696 (N_7696,N_4040,N_4737);
or U7697 (N_7697,N_4288,N_4754);
or U7698 (N_7698,N_4813,N_5302);
nand U7699 (N_7699,N_5067,N_4295);
nand U7700 (N_7700,N_4200,N_4932);
or U7701 (N_7701,N_5693,N_4856);
nor U7702 (N_7702,N_4760,N_5736);
or U7703 (N_7703,N_4509,N_4920);
and U7704 (N_7704,N_4406,N_4313);
and U7705 (N_7705,N_4963,N_5040);
or U7706 (N_7706,N_4125,N_4714);
nor U7707 (N_7707,N_4249,N_5896);
nand U7708 (N_7708,N_5037,N_4051);
nor U7709 (N_7709,N_4164,N_5941);
nor U7710 (N_7710,N_5043,N_4385);
and U7711 (N_7711,N_5126,N_5587);
nand U7712 (N_7712,N_5897,N_4466);
nor U7713 (N_7713,N_5233,N_5099);
nand U7714 (N_7714,N_4973,N_4142);
nor U7715 (N_7715,N_4013,N_5921);
nor U7716 (N_7716,N_5429,N_5412);
nor U7717 (N_7717,N_5593,N_4130);
or U7718 (N_7718,N_4819,N_4968);
or U7719 (N_7719,N_4001,N_5217);
nand U7720 (N_7720,N_5805,N_4536);
and U7721 (N_7721,N_4308,N_5157);
nor U7722 (N_7722,N_5532,N_4862);
and U7723 (N_7723,N_4921,N_4046);
or U7724 (N_7724,N_4224,N_5687);
nand U7725 (N_7725,N_5058,N_4171);
nand U7726 (N_7726,N_5617,N_4816);
xor U7727 (N_7727,N_4254,N_4400);
or U7728 (N_7728,N_4264,N_4113);
or U7729 (N_7729,N_4803,N_4785);
nand U7730 (N_7730,N_5407,N_5570);
nand U7731 (N_7731,N_5158,N_4008);
nand U7732 (N_7732,N_5457,N_4853);
and U7733 (N_7733,N_5699,N_4079);
nand U7734 (N_7734,N_4777,N_4251);
and U7735 (N_7735,N_4884,N_4424);
and U7736 (N_7736,N_5526,N_5285);
nand U7737 (N_7737,N_5991,N_4168);
nand U7738 (N_7738,N_4356,N_4781);
nand U7739 (N_7739,N_4993,N_4507);
nand U7740 (N_7740,N_4155,N_5253);
and U7741 (N_7741,N_5554,N_4472);
nor U7742 (N_7742,N_5254,N_4565);
or U7743 (N_7743,N_4891,N_5686);
or U7744 (N_7744,N_5014,N_4077);
and U7745 (N_7745,N_4542,N_4590);
nor U7746 (N_7746,N_5994,N_5627);
nor U7747 (N_7747,N_5248,N_4160);
nand U7748 (N_7748,N_4684,N_4241);
nand U7749 (N_7749,N_4068,N_4878);
nand U7750 (N_7750,N_4239,N_4933);
and U7751 (N_7751,N_4942,N_4049);
nor U7752 (N_7752,N_5468,N_5513);
or U7753 (N_7753,N_5929,N_4846);
or U7754 (N_7754,N_4175,N_4923);
nand U7755 (N_7755,N_4392,N_5499);
nand U7756 (N_7756,N_4312,N_5743);
or U7757 (N_7757,N_5505,N_5058);
and U7758 (N_7758,N_5154,N_4256);
and U7759 (N_7759,N_5376,N_4630);
nand U7760 (N_7760,N_5801,N_4218);
nand U7761 (N_7761,N_4040,N_4610);
nand U7762 (N_7762,N_4310,N_4890);
nor U7763 (N_7763,N_4642,N_5538);
and U7764 (N_7764,N_4961,N_5027);
and U7765 (N_7765,N_4635,N_5219);
and U7766 (N_7766,N_4905,N_4131);
nor U7767 (N_7767,N_5469,N_4530);
and U7768 (N_7768,N_4131,N_5311);
or U7769 (N_7769,N_4479,N_5449);
and U7770 (N_7770,N_5590,N_4120);
nand U7771 (N_7771,N_5098,N_5113);
nor U7772 (N_7772,N_5571,N_4530);
and U7773 (N_7773,N_4535,N_4146);
nor U7774 (N_7774,N_5438,N_5060);
nand U7775 (N_7775,N_5317,N_4322);
nand U7776 (N_7776,N_4030,N_4376);
or U7777 (N_7777,N_4228,N_5794);
nor U7778 (N_7778,N_5924,N_4639);
or U7779 (N_7779,N_5709,N_4215);
nand U7780 (N_7780,N_5276,N_5703);
or U7781 (N_7781,N_5848,N_4032);
and U7782 (N_7782,N_4940,N_4616);
nand U7783 (N_7783,N_5568,N_4339);
and U7784 (N_7784,N_4776,N_4450);
or U7785 (N_7785,N_4830,N_4452);
and U7786 (N_7786,N_4769,N_4286);
nand U7787 (N_7787,N_5835,N_4741);
or U7788 (N_7788,N_4334,N_5632);
or U7789 (N_7789,N_4233,N_5998);
and U7790 (N_7790,N_5551,N_5899);
or U7791 (N_7791,N_5440,N_5536);
nand U7792 (N_7792,N_4485,N_5957);
and U7793 (N_7793,N_5757,N_5834);
xnor U7794 (N_7794,N_5909,N_4204);
and U7795 (N_7795,N_4593,N_5645);
or U7796 (N_7796,N_4339,N_4985);
and U7797 (N_7797,N_4744,N_5475);
nor U7798 (N_7798,N_5494,N_4281);
nand U7799 (N_7799,N_5881,N_5418);
or U7800 (N_7800,N_4128,N_4543);
and U7801 (N_7801,N_4608,N_5795);
or U7802 (N_7802,N_5597,N_4997);
nand U7803 (N_7803,N_5693,N_5553);
nor U7804 (N_7804,N_4818,N_5772);
nor U7805 (N_7805,N_5456,N_5745);
or U7806 (N_7806,N_5949,N_4324);
and U7807 (N_7807,N_5188,N_4982);
nand U7808 (N_7808,N_4152,N_4544);
nand U7809 (N_7809,N_5078,N_5409);
nand U7810 (N_7810,N_4298,N_4570);
nand U7811 (N_7811,N_4028,N_4410);
and U7812 (N_7812,N_4322,N_4381);
or U7813 (N_7813,N_4260,N_5169);
or U7814 (N_7814,N_5683,N_5337);
or U7815 (N_7815,N_4689,N_5443);
or U7816 (N_7816,N_4515,N_5586);
or U7817 (N_7817,N_5295,N_5831);
and U7818 (N_7818,N_4687,N_5646);
and U7819 (N_7819,N_5338,N_5724);
nand U7820 (N_7820,N_4900,N_4080);
or U7821 (N_7821,N_5214,N_5774);
or U7822 (N_7822,N_4543,N_5402);
or U7823 (N_7823,N_4791,N_5943);
nor U7824 (N_7824,N_4661,N_4105);
and U7825 (N_7825,N_4821,N_4632);
nand U7826 (N_7826,N_5807,N_5428);
and U7827 (N_7827,N_4105,N_5142);
nand U7828 (N_7828,N_5405,N_4209);
and U7829 (N_7829,N_4232,N_5462);
nor U7830 (N_7830,N_5237,N_4752);
nand U7831 (N_7831,N_4993,N_4453);
nor U7832 (N_7832,N_4400,N_4281);
nand U7833 (N_7833,N_5499,N_5577);
and U7834 (N_7834,N_4428,N_4958);
nor U7835 (N_7835,N_4042,N_4937);
or U7836 (N_7836,N_4329,N_4134);
or U7837 (N_7837,N_4980,N_5887);
or U7838 (N_7838,N_4888,N_4004);
nand U7839 (N_7839,N_4287,N_4852);
nor U7840 (N_7840,N_4462,N_4868);
or U7841 (N_7841,N_4985,N_4371);
nor U7842 (N_7842,N_4548,N_4704);
and U7843 (N_7843,N_4334,N_4052);
and U7844 (N_7844,N_4890,N_4785);
nor U7845 (N_7845,N_4350,N_4753);
nand U7846 (N_7846,N_4431,N_5732);
nor U7847 (N_7847,N_5615,N_4123);
and U7848 (N_7848,N_5277,N_4483);
nand U7849 (N_7849,N_5887,N_5178);
and U7850 (N_7850,N_4835,N_4833);
nor U7851 (N_7851,N_5741,N_5343);
nor U7852 (N_7852,N_5954,N_4650);
or U7853 (N_7853,N_4992,N_5034);
or U7854 (N_7854,N_4128,N_4326);
and U7855 (N_7855,N_5340,N_5147);
or U7856 (N_7856,N_4720,N_5520);
nor U7857 (N_7857,N_4776,N_4037);
and U7858 (N_7858,N_5692,N_5025);
and U7859 (N_7859,N_5401,N_4780);
nor U7860 (N_7860,N_5296,N_4684);
or U7861 (N_7861,N_5479,N_4647);
nand U7862 (N_7862,N_4347,N_5917);
or U7863 (N_7863,N_5534,N_5886);
nand U7864 (N_7864,N_5956,N_5389);
nor U7865 (N_7865,N_5105,N_5834);
and U7866 (N_7866,N_5640,N_4673);
and U7867 (N_7867,N_5438,N_5283);
nand U7868 (N_7868,N_4369,N_5285);
and U7869 (N_7869,N_4431,N_5401);
nand U7870 (N_7870,N_4841,N_4463);
nor U7871 (N_7871,N_5322,N_5822);
nand U7872 (N_7872,N_4717,N_5070);
nor U7873 (N_7873,N_5407,N_4307);
or U7874 (N_7874,N_5998,N_5586);
and U7875 (N_7875,N_5161,N_5443);
nor U7876 (N_7876,N_5931,N_4765);
nand U7877 (N_7877,N_5144,N_5085);
nand U7878 (N_7878,N_5307,N_4961);
or U7879 (N_7879,N_5659,N_4588);
and U7880 (N_7880,N_5864,N_5035);
nand U7881 (N_7881,N_4054,N_5385);
and U7882 (N_7882,N_5734,N_4522);
and U7883 (N_7883,N_4296,N_4582);
and U7884 (N_7884,N_5997,N_5157);
nand U7885 (N_7885,N_5948,N_4187);
nand U7886 (N_7886,N_5662,N_5581);
nor U7887 (N_7887,N_5654,N_5970);
nand U7888 (N_7888,N_4404,N_5038);
or U7889 (N_7889,N_5601,N_4836);
and U7890 (N_7890,N_4672,N_4932);
nor U7891 (N_7891,N_4013,N_5745);
nand U7892 (N_7892,N_4253,N_5835);
xnor U7893 (N_7893,N_4882,N_5456);
nor U7894 (N_7894,N_4343,N_5111);
or U7895 (N_7895,N_5805,N_4515);
nand U7896 (N_7896,N_5641,N_5174);
and U7897 (N_7897,N_5126,N_5726);
or U7898 (N_7898,N_4366,N_5650);
nor U7899 (N_7899,N_5395,N_4159);
and U7900 (N_7900,N_4034,N_5542);
and U7901 (N_7901,N_5048,N_5851);
and U7902 (N_7902,N_4509,N_5926);
and U7903 (N_7903,N_4895,N_4673);
and U7904 (N_7904,N_5064,N_4732);
or U7905 (N_7905,N_4969,N_4583);
nand U7906 (N_7906,N_4233,N_4178);
nand U7907 (N_7907,N_5411,N_5838);
and U7908 (N_7908,N_5437,N_4847);
and U7909 (N_7909,N_4992,N_5594);
nor U7910 (N_7910,N_5534,N_4709);
nor U7911 (N_7911,N_5484,N_4998);
and U7912 (N_7912,N_5989,N_5388);
or U7913 (N_7913,N_4000,N_4589);
nand U7914 (N_7914,N_4137,N_4252);
or U7915 (N_7915,N_5119,N_5721);
or U7916 (N_7916,N_4313,N_5479);
and U7917 (N_7917,N_5182,N_4435);
and U7918 (N_7918,N_4355,N_5210);
nand U7919 (N_7919,N_4677,N_5565);
nor U7920 (N_7920,N_5163,N_5002);
nand U7921 (N_7921,N_5003,N_5286);
or U7922 (N_7922,N_4162,N_5785);
and U7923 (N_7923,N_5450,N_5548);
and U7924 (N_7924,N_4120,N_4565);
nor U7925 (N_7925,N_5987,N_4549);
nor U7926 (N_7926,N_4690,N_5074);
nand U7927 (N_7927,N_4158,N_4981);
nand U7928 (N_7928,N_5933,N_4182);
and U7929 (N_7929,N_5121,N_5512);
nor U7930 (N_7930,N_4367,N_5786);
nand U7931 (N_7931,N_5726,N_5548);
nand U7932 (N_7932,N_5976,N_4746);
or U7933 (N_7933,N_5032,N_4435);
nor U7934 (N_7934,N_4466,N_5860);
and U7935 (N_7935,N_5134,N_5481);
nand U7936 (N_7936,N_4361,N_5320);
nor U7937 (N_7937,N_5583,N_4449);
and U7938 (N_7938,N_4429,N_5454);
and U7939 (N_7939,N_4247,N_4526);
and U7940 (N_7940,N_5134,N_5951);
nand U7941 (N_7941,N_5886,N_5920);
or U7942 (N_7942,N_5313,N_5350);
or U7943 (N_7943,N_5752,N_5306);
nor U7944 (N_7944,N_5141,N_5040);
nor U7945 (N_7945,N_5636,N_5559);
or U7946 (N_7946,N_5524,N_5771);
and U7947 (N_7947,N_5521,N_5671);
or U7948 (N_7948,N_5229,N_5364);
nand U7949 (N_7949,N_5616,N_4250);
and U7950 (N_7950,N_4394,N_5502);
nand U7951 (N_7951,N_4625,N_4278);
or U7952 (N_7952,N_5565,N_4999);
and U7953 (N_7953,N_5801,N_5974);
or U7954 (N_7954,N_5259,N_5052);
nand U7955 (N_7955,N_5694,N_4484);
xor U7956 (N_7956,N_4345,N_5791);
and U7957 (N_7957,N_4856,N_4401);
nor U7958 (N_7958,N_4086,N_4030);
nor U7959 (N_7959,N_5605,N_5621);
and U7960 (N_7960,N_4449,N_5033);
nand U7961 (N_7961,N_5165,N_5405);
nor U7962 (N_7962,N_5737,N_4992);
nand U7963 (N_7963,N_5684,N_5961);
nor U7964 (N_7964,N_4853,N_5829);
nand U7965 (N_7965,N_5579,N_4726);
nand U7966 (N_7966,N_4039,N_4737);
nand U7967 (N_7967,N_4251,N_5784);
nor U7968 (N_7968,N_5511,N_4412);
nand U7969 (N_7969,N_4805,N_4447);
and U7970 (N_7970,N_5440,N_5874);
nor U7971 (N_7971,N_5149,N_5567);
and U7972 (N_7972,N_5493,N_4269);
and U7973 (N_7973,N_4148,N_4371);
nand U7974 (N_7974,N_5333,N_5614);
or U7975 (N_7975,N_4804,N_5394);
nand U7976 (N_7976,N_5230,N_5206);
or U7977 (N_7977,N_5461,N_4207);
or U7978 (N_7978,N_4985,N_5424);
nand U7979 (N_7979,N_5361,N_5866);
nand U7980 (N_7980,N_5571,N_4152);
nand U7981 (N_7981,N_4904,N_4582);
nor U7982 (N_7982,N_5259,N_4826);
and U7983 (N_7983,N_5445,N_5348);
and U7984 (N_7984,N_4484,N_5466);
and U7985 (N_7985,N_5517,N_4077);
or U7986 (N_7986,N_5994,N_4446);
nor U7987 (N_7987,N_4719,N_4648);
or U7988 (N_7988,N_5676,N_4962);
nor U7989 (N_7989,N_4742,N_5793);
nor U7990 (N_7990,N_5487,N_4259);
and U7991 (N_7991,N_4027,N_5459);
nor U7992 (N_7992,N_4727,N_5130);
nor U7993 (N_7993,N_5089,N_5046);
or U7994 (N_7994,N_5639,N_5712);
xor U7995 (N_7995,N_5129,N_5862);
and U7996 (N_7996,N_5024,N_5758);
nand U7997 (N_7997,N_4341,N_4563);
nand U7998 (N_7998,N_5617,N_5982);
or U7999 (N_7999,N_5025,N_4980);
or U8000 (N_8000,N_7444,N_7276);
or U8001 (N_8001,N_6306,N_6135);
nor U8002 (N_8002,N_7707,N_7975);
nand U8003 (N_8003,N_7840,N_6323);
nor U8004 (N_8004,N_7824,N_7381);
nand U8005 (N_8005,N_6100,N_7647);
nor U8006 (N_8006,N_6949,N_6997);
or U8007 (N_8007,N_6687,N_7581);
or U8008 (N_8008,N_6378,N_6620);
and U8009 (N_8009,N_6325,N_7194);
nand U8010 (N_8010,N_7821,N_6231);
or U8011 (N_8011,N_7281,N_6817);
nor U8012 (N_8012,N_7916,N_6393);
nand U8013 (N_8013,N_7905,N_6748);
nand U8014 (N_8014,N_6136,N_6326);
or U8015 (N_8015,N_7611,N_7861);
nand U8016 (N_8016,N_7051,N_6489);
nor U8017 (N_8017,N_7668,N_6626);
and U8018 (N_8018,N_6822,N_7961);
or U8019 (N_8019,N_7208,N_6712);
and U8020 (N_8020,N_6920,N_6149);
nor U8021 (N_8021,N_6153,N_7950);
nor U8022 (N_8022,N_7206,N_6941);
nand U8023 (N_8023,N_7620,N_7676);
and U8024 (N_8024,N_6007,N_7778);
nor U8025 (N_8025,N_7241,N_6563);
nand U8026 (N_8026,N_6459,N_7776);
and U8027 (N_8027,N_7130,N_6856);
or U8028 (N_8028,N_6988,N_6892);
and U8029 (N_8029,N_7742,N_7610);
and U8030 (N_8030,N_7990,N_6940);
nand U8031 (N_8031,N_6963,N_7511);
nand U8032 (N_8032,N_6357,N_6075);
nand U8033 (N_8033,N_6667,N_7459);
and U8034 (N_8034,N_6810,N_7586);
or U8035 (N_8035,N_7013,N_6658);
nor U8036 (N_8036,N_6505,N_7080);
or U8037 (N_8037,N_7212,N_6590);
or U8038 (N_8038,N_6257,N_6099);
and U8039 (N_8039,N_7407,N_6072);
nor U8040 (N_8040,N_6118,N_7797);
nor U8041 (N_8041,N_6982,N_7273);
and U8042 (N_8042,N_6453,N_6446);
nand U8043 (N_8043,N_6368,N_7551);
nor U8044 (N_8044,N_7657,N_6581);
nor U8045 (N_8045,N_7790,N_7526);
or U8046 (N_8046,N_6643,N_7417);
nor U8047 (N_8047,N_6280,N_6918);
and U8048 (N_8048,N_7992,N_6558);
nor U8049 (N_8049,N_6797,N_7057);
or U8050 (N_8050,N_6370,N_6957);
and U8051 (N_8051,N_6783,N_6681);
nand U8052 (N_8052,N_7901,N_6033);
nand U8053 (N_8053,N_6874,N_7897);
nand U8054 (N_8054,N_6058,N_6556);
nand U8055 (N_8055,N_6343,N_6604);
or U8056 (N_8056,N_6862,N_6485);
and U8057 (N_8057,N_6221,N_6288);
or U8058 (N_8058,N_6532,N_6763);
nand U8059 (N_8059,N_7794,N_6480);
nand U8060 (N_8060,N_7884,N_6371);
nand U8061 (N_8061,N_7005,N_6899);
and U8062 (N_8062,N_7072,N_6971);
nand U8063 (N_8063,N_7556,N_7464);
and U8064 (N_8064,N_7059,N_6601);
and U8065 (N_8065,N_6450,N_6452);
or U8066 (N_8066,N_7758,N_6800);
nor U8067 (N_8067,N_6644,N_6247);
and U8068 (N_8068,N_7148,N_7078);
and U8069 (N_8069,N_6352,N_6400);
nand U8070 (N_8070,N_6967,N_7492);
or U8071 (N_8071,N_6169,N_6269);
nor U8072 (N_8072,N_6397,N_7593);
nand U8073 (N_8073,N_6197,N_7224);
and U8074 (N_8074,N_7687,N_7822);
nor U8075 (N_8075,N_7675,N_6860);
or U8076 (N_8076,N_6811,N_7356);
or U8077 (N_8077,N_6973,N_6905);
and U8078 (N_8078,N_7086,N_7041);
or U8079 (N_8079,N_6493,N_7736);
nor U8080 (N_8080,N_7465,N_7389);
and U8081 (N_8081,N_7164,N_7106);
or U8082 (N_8082,N_7738,N_6394);
nor U8083 (N_8083,N_7554,N_6939);
or U8084 (N_8084,N_7857,N_6781);
nand U8085 (N_8085,N_6396,N_6185);
and U8086 (N_8086,N_6143,N_6752);
or U8087 (N_8087,N_6463,N_6747);
and U8088 (N_8088,N_7355,N_7344);
or U8089 (N_8089,N_6888,N_6403);
nor U8090 (N_8090,N_7984,N_7823);
or U8091 (N_8091,N_7484,N_6422);
nor U8092 (N_8092,N_6542,N_7649);
nand U8093 (N_8093,N_6282,N_6116);
or U8094 (N_8094,N_7560,N_7777);
and U8095 (N_8095,N_6663,N_6836);
nand U8096 (N_8096,N_7798,N_7878);
or U8097 (N_8097,N_6142,N_7795);
and U8098 (N_8098,N_6666,N_6354);
or U8099 (N_8099,N_7203,N_6914);
or U8100 (N_8100,N_6826,N_6027);
nor U8101 (N_8101,N_7483,N_6517);
and U8102 (N_8102,N_6160,N_7504);
nand U8103 (N_8103,N_7945,N_6235);
nor U8104 (N_8104,N_7490,N_6555);
or U8105 (N_8105,N_7955,N_7998);
or U8106 (N_8106,N_7153,N_6835);
and U8107 (N_8107,N_7262,N_7412);
nand U8108 (N_8108,N_6108,N_7686);
nand U8109 (N_8109,N_6533,N_6829);
nor U8110 (N_8110,N_7832,N_7266);
nand U8111 (N_8111,N_7301,N_6546);
nor U8112 (N_8112,N_6779,N_7100);
nand U8113 (N_8113,N_6004,N_6219);
nor U8114 (N_8114,N_6233,N_7022);
nand U8115 (N_8115,N_7708,N_7793);
or U8116 (N_8116,N_7226,N_7493);
nand U8117 (N_8117,N_6936,N_6304);
and U8118 (N_8118,N_7382,N_7835);
nor U8119 (N_8119,N_7644,N_7801);
nor U8120 (N_8120,N_6106,N_7545);
nor U8121 (N_8121,N_7002,N_6676);
and U8122 (N_8122,N_7980,N_6910);
nand U8123 (N_8123,N_7722,N_6208);
or U8124 (N_8124,N_6430,N_6972);
or U8125 (N_8125,N_6353,N_7540);
and U8126 (N_8126,N_7792,N_7746);
or U8127 (N_8127,N_6691,N_7678);
and U8128 (N_8128,N_6695,N_6682);
nor U8129 (N_8129,N_6039,N_7847);
and U8130 (N_8130,N_6999,N_6125);
nor U8131 (N_8131,N_6868,N_7639);
nor U8132 (N_8132,N_7062,N_6750);
or U8133 (N_8133,N_7590,N_6605);
nand U8134 (N_8134,N_7527,N_7911);
nand U8135 (N_8135,N_7594,N_7159);
and U8136 (N_8136,N_7350,N_7168);
or U8137 (N_8137,N_7683,N_6757);
nor U8138 (N_8138,N_7142,N_6591);
nand U8139 (N_8139,N_7514,N_6021);
and U8140 (N_8140,N_7084,N_6220);
nand U8141 (N_8141,N_7513,N_7079);
and U8142 (N_8142,N_6170,N_7378);
nor U8143 (N_8143,N_6129,N_6907);
nand U8144 (N_8144,N_6365,N_7519);
or U8145 (N_8145,N_6637,N_6030);
nand U8146 (N_8146,N_7383,N_7103);
and U8147 (N_8147,N_7028,N_7116);
nor U8148 (N_8148,N_7634,N_7946);
nand U8149 (N_8149,N_6863,N_6504);
or U8150 (N_8150,N_7928,N_7374);
or U8151 (N_8151,N_6240,N_6557);
nor U8152 (N_8152,N_7141,N_6031);
or U8153 (N_8153,N_7803,N_7120);
nand U8154 (N_8154,N_6207,N_7769);
nand U8155 (N_8155,N_6420,N_7403);
nor U8156 (N_8156,N_7914,N_6413);
nor U8157 (N_8157,N_7447,N_7697);
and U8158 (N_8158,N_7095,N_6080);
nand U8159 (N_8159,N_6568,N_7176);
and U8160 (N_8160,N_6174,N_6273);
nand U8161 (N_8161,N_7138,N_7297);
nand U8162 (N_8162,N_6122,N_7235);
or U8163 (N_8163,N_6548,N_7489);
and U8164 (N_8164,N_7991,N_7468);
nor U8165 (N_8165,N_6646,N_6794);
nand U8166 (N_8166,N_6579,N_6733);
or U8167 (N_8167,N_7993,N_7966);
nor U8168 (N_8168,N_7827,N_6424);
and U8169 (N_8169,N_6383,N_6270);
nand U8170 (N_8170,N_7023,N_6491);
nor U8171 (N_8171,N_6986,N_6989);
nand U8172 (N_8172,N_7162,N_7307);
nand U8173 (N_8173,N_6315,N_7645);
and U8174 (N_8174,N_6974,N_6886);
nor U8175 (N_8175,N_6613,N_6902);
nand U8176 (N_8176,N_6102,N_7733);
nand U8177 (N_8177,N_6770,N_6839);
nor U8178 (N_8178,N_6188,N_6764);
and U8179 (N_8179,N_7898,N_6977);
nor U8180 (N_8180,N_7342,N_7020);
nand U8181 (N_8181,N_7037,N_7693);
and U8182 (N_8182,N_6859,N_6571);
and U8183 (N_8183,N_7316,N_7569);
nor U8184 (N_8184,N_6402,N_6380);
nor U8185 (N_8185,N_6520,N_6968);
or U8186 (N_8186,N_6212,N_6052);
and U8187 (N_8187,N_6434,N_7729);
and U8188 (N_8188,N_7404,N_6717);
nor U8189 (N_8189,N_7152,N_7236);
nand U8190 (N_8190,N_7418,N_6332);
or U8191 (N_8191,N_7770,N_7300);
xnor U8192 (N_8192,N_7548,N_7365);
and U8193 (N_8193,N_6922,N_7615);
nand U8194 (N_8194,N_7575,N_6206);
or U8195 (N_8195,N_7060,N_7274);
xor U8196 (N_8196,N_7727,N_6363);
and U8197 (N_8197,N_7045,N_7666);
and U8198 (N_8198,N_7191,N_6291);
nand U8199 (N_8199,N_6024,N_6087);
nor U8200 (N_8200,N_7091,N_6164);
or U8201 (N_8201,N_6871,N_6069);
or U8202 (N_8202,N_7573,N_7582);
nor U8203 (N_8203,N_7825,N_6001);
or U8204 (N_8204,N_7361,N_7082);
xnor U8205 (N_8205,N_7136,N_7114);
and U8206 (N_8206,N_6372,N_7664);
nor U8207 (N_8207,N_7395,N_7263);
and U8208 (N_8208,N_7195,N_6896);
and U8209 (N_8209,N_6182,N_6580);
or U8210 (N_8210,N_6617,N_6970);
or U8211 (N_8211,N_6791,N_6569);
nand U8212 (N_8212,N_6248,N_6301);
or U8213 (N_8213,N_6909,N_7949);
nor U8214 (N_8214,N_7846,N_6084);
and U8215 (N_8215,N_6753,N_6882);
nand U8216 (N_8216,N_7609,N_7684);
nor U8217 (N_8217,N_7599,N_6689);
or U8218 (N_8218,N_7458,N_6724);
nand U8219 (N_8219,N_7939,N_6311);
or U8220 (N_8220,N_7848,N_7362);
and U8221 (N_8221,N_7938,N_7563);
and U8222 (N_8222,N_7123,N_7854);
and U8223 (N_8223,N_6384,N_6692);
and U8224 (N_8224,N_7872,N_6037);
or U8225 (N_8225,N_7624,N_7583);
nand U8226 (N_8226,N_7133,N_7819);
nor U8227 (N_8227,N_7189,N_6376);
or U8228 (N_8228,N_7070,N_7920);
or U8229 (N_8229,N_6851,N_6036);
and U8230 (N_8230,N_7786,N_6611);
nand U8231 (N_8231,N_6561,N_7783);
nor U8232 (N_8232,N_6466,N_7303);
nor U8233 (N_8233,N_7039,N_6211);
or U8234 (N_8234,N_6958,N_6017);
nand U8235 (N_8235,N_6848,N_6776);
nand U8236 (N_8236,N_6883,N_7927);
nor U8237 (N_8237,N_6870,N_6509);
nand U8238 (N_8238,N_6677,N_7474);
and U8239 (N_8239,N_7498,N_7376);
nor U8240 (N_8240,N_7791,N_6404);
or U8241 (N_8241,N_6565,N_6576);
or U8242 (N_8242,N_7944,N_7882);
nand U8243 (N_8243,N_7043,N_7113);
nand U8244 (N_8244,N_7674,N_7743);
and U8245 (N_8245,N_6911,N_6297);
and U8246 (N_8246,N_7280,N_7895);
and U8247 (N_8247,N_6103,N_7319);
and U8248 (N_8248,N_7537,N_6865);
and U8249 (N_8249,N_6503,N_7217);
or U8250 (N_8250,N_7277,N_7717);
and U8251 (N_8251,N_7867,N_6831);
and U8252 (N_8252,N_7341,N_7174);
nor U8253 (N_8253,N_7284,N_7055);
nand U8254 (N_8254,N_7698,N_6980);
nand U8255 (N_8255,N_7036,N_7211);
nand U8256 (N_8256,N_7748,N_6664);
nand U8257 (N_8257,N_6885,N_7773);
nor U8258 (N_8258,N_7117,N_7957);
nor U8259 (N_8259,N_7310,N_7544);
or U8260 (N_8260,N_7098,N_6684);
nor U8261 (N_8261,N_6648,N_7083);
and U8262 (N_8262,N_6840,N_6731);
nand U8263 (N_8263,N_6082,N_6098);
and U8264 (N_8264,N_6716,N_6602);
nor U8265 (N_8265,N_6405,N_6540);
and U8266 (N_8266,N_6732,N_6864);
xnor U8267 (N_8267,N_6095,N_6670);
nand U8268 (N_8268,N_7906,N_7885);
nand U8269 (N_8269,N_7663,N_6554);
or U8270 (N_8270,N_7128,N_7877);
nand U8271 (N_8271,N_7097,N_7440);
nor U8272 (N_8272,N_6093,N_6227);
nor U8273 (N_8273,N_6994,N_6702);
xor U8274 (N_8274,N_7816,N_6127);
nor U8275 (N_8275,N_6015,N_6067);
and U8276 (N_8276,N_7628,N_7962);
nor U8277 (N_8277,N_6529,N_6693);
or U8278 (N_8278,N_7452,N_6199);
nor U8279 (N_8279,N_7171,N_6573);
nand U8280 (N_8280,N_7173,N_7363);
and U8281 (N_8281,N_6209,N_6333);
nand U8282 (N_8282,N_6823,N_7588);
nor U8283 (N_8283,N_6657,N_6388);
and U8284 (N_8284,N_6408,N_6736);
or U8285 (N_8285,N_7478,N_7431);
or U8286 (N_8286,N_7050,N_7602);
or U8287 (N_8287,N_6144,N_7077);
nand U8288 (N_8288,N_7390,N_6538);
or U8289 (N_8289,N_6975,N_7163);
nor U8290 (N_8290,N_6893,N_6739);
or U8291 (N_8291,N_6046,N_7058);
nor U8292 (N_8292,N_7186,N_7405);
and U8293 (N_8293,N_6313,N_6518);
nand U8294 (N_8294,N_6916,N_6312);
or U8295 (N_8295,N_6410,N_6651);
and U8296 (N_8296,N_7069,N_7971);
nor U8297 (N_8297,N_7669,N_7345);
and U8298 (N_8298,N_6417,N_7087);
and U8299 (N_8299,N_6409,N_6214);
and U8300 (N_8300,N_7011,N_6536);
and U8301 (N_8301,N_7196,N_7889);
or U8302 (N_8302,N_6537,N_7338);
nand U8303 (N_8303,N_6832,N_6578);
and U8304 (N_8304,N_6005,N_6166);
nand U8305 (N_8305,N_6161,N_7505);
or U8306 (N_8306,N_7838,N_7237);
nor U8307 (N_8307,N_6419,N_7909);
or U8308 (N_8308,N_6189,N_6908);
and U8309 (N_8309,N_6850,N_7425);
nor U8310 (N_8310,N_6193,N_6824);
and U8311 (N_8311,N_7988,N_7497);
nor U8312 (N_8312,N_6965,N_6079);
and U8313 (N_8313,N_7398,N_7258);
nor U8314 (N_8314,N_7388,N_6869);
nand U8315 (N_8315,N_7324,N_6109);
or U8316 (N_8316,N_6924,N_7725);
or U8317 (N_8317,N_6196,N_6168);
nor U8318 (N_8318,N_6350,N_6351);
xnor U8319 (N_8319,N_6066,N_7391);
and U8320 (N_8320,N_7225,N_7879);
or U8321 (N_8321,N_6841,N_6232);
nand U8322 (N_8322,N_7205,N_6321);
or U8323 (N_8323,N_6609,N_7700);
nand U8324 (N_8324,N_6259,N_7750);
or U8325 (N_8325,N_7844,N_7601);
nor U8326 (N_8326,N_6076,N_7373);
nor U8327 (N_8327,N_7000,N_6034);
and U8328 (N_8328,N_6307,N_7930);
nand U8329 (N_8329,N_7432,N_6872);
and U8330 (N_8330,N_7446,N_7562);
nor U8331 (N_8331,N_6745,N_7886);
and U8332 (N_8332,N_7534,N_7044);
and U8333 (N_8333,N_6205,N_7288);
nand U8334 (N_8334,N_6152,N_7377);
and U8335 (N_8335,N_6141,N_6302);
and U8336 (N_8336,N_7541,N_7073);
xor U8337 (N_8337,N_7127,N_7807);
nand U8338 (N_8338,N_6993,N_7616);
nor U8339 (N_8339,N_7646,N_6049);
and U8340 (N_8340,N_7640,N_7605);
or U8341 (N_8341,N_7001,N_7681);
and U8342 (N_8342,N_6179,N_7054);
xnor U8343 (N_8343,N_6726,N_7530);
or U8344 (N_8344,N_7275,N_7680);
nor U8345 (N_8345,N_7475,N_7311);
nor U8346 (N_8346,N_6022,N_6488);
and U8347 (N_8347,N_7299,N_7227);
and U8348 (N_8348,N_6043,N_7401);
nand U8349 (N_8349,N_7970,N_6768);
nand U8350 (N_8350,N_6110,N_7243);
and U8351 (N_8351,N_6254,N_7109);
and U8352 (N_8352,N_6636,N_6395);
nand U8353 (N_8353,N_6283,N_6614);
or U8354 (N_8354,N_6891,N_6204);
or U8355 (N_8355,N_7953,N_6761);
nor U8356 (N_8356,N_7564,N_6582);
nor U8357 (N_8357,N_7175,N_7528);
nand U8358 (N_8358,N_6877,N_7485);
nand U8359 (N_8359,N_6669,N_6592);
nand U8360 (N_8360,N_7248,N_6173);
nor U8361 (N_8361,N_6482,N_6654);
nand U8362 (N_8362,N_7337,N_6583);
and U8363 (N_8363,N_6597,N_6317);
nand U8364 (N_8364,N_6392,N_6696);
nor U8365 (N_8365,N_6157,N_7892);
nand U8366 (N_8366,N_6156,N_7435);
and U8367 (N_8367,N_7691,N_6600);
nor U8368 (N_8368,N_7917,N_7856);
nand U8369 (N_8369,N_6431,N_6526);
or U8370 (N_8370,N_7826,N_7653);
or U8371 (N_8371,N_7524,N_7529);
or U8372 (N_8372,N_7500,N_7146);
or U8373 (N_8373,N_6339,N_6132);
or U8374 (N_8374,N_7312,N_7744);
nor U8375 (N_8375,N_7298,N_6790);
nor U8376 (N_8376,N_7421,N_6203);
or U8377 (N_8377,N_7333,N_6701);
nand U8378 (N_8378,N_6155,N_7557);
nor U8379 (N_8379,N_7591,N_7009);
nand U8380 (N_8380,N_6038,N_6112);
xnor U8381 (N_8381,N_7397,N_6713);
nand U8382 (N_8382,N_6063,N_6956);
or U8383 (N_8383,N_6861,N_6566);
and U8384 (N_8384,N_6213,N_6338);
nand U8385 (N_8385,N_7234,N_7088);
nor U8386 (N_8386,N_6081,N_7935);
or U8387 (N_8387,N_7019,N_7240);
nand U8388 (N_8388,N_6460,N_6310);
and U8389 (N_8389,N_6479,N_7034);
nand U8390 (N_8390,N_6194,N_6292);
nor U8391 (N_8391,N_7201,N_7149);
nand U8392 (N_8392,N_6992,N_6470);
nor U8393 (N_8393,N_7071,N_7913);
nand U8394 (N_8394,N_6806,N_6570);
nor U8395 (N_8395,N_7660,N_6433);
and U8396 (N_8396,N_6456,N_7025);
nor U8397 (N_8397,N_7812,N_6454);
nand U8398 (N_8398,N_6073,N_6202);
and U8399 (N_8399,N_7782,N_6531);
xor U8400 (N_8400,N_7936,N_6749);
nand U8401 (N_8401,N_6314,N_6927);
or U8402 (N_8402,N_6318,N_6020);
or U8403 (N_8403,N_6145,N_6966);
and U8404 (N_8404,N_7637,N_7295);
or U8405 (N_8405,N_7134,N_6077);
or U8406 (N_8406,N_6525,N_7566);
nor U8407 (N_8407,N_6198,N_6290);
nand U8408 (N_8408,N_7147,N_6437);
nor U8409 (N_8409,N_7018,N_7730);
and U8410 (N_8410,N_6813,N_6337);
nand U8411 (N_8411,N_7033,N_7291);
or U8412 (N_8412,N_6074,N_7251);
nand U8413 (N_8413,N_7181,N_6278);
and U8414 (N_8414,N_6718,N_6490);
nand U8415 (N_8415,N_6465,N_7860);
and U8416 (N_8416,N_7294,N_7029);
nor U8417 (N_8417,N_7124,N_6336);
nor U8418 (N_8418,N_7780,N_7340);
nor U8419 (N_8419,N_7679,N_7249);
nand U8420 (N_8420,N_6512,N_6678);
nand U8421 (N_8421,N_7253,N_7942);
or U8422 (N_8422,N_7233,N_7215);
and U8423 (N_8423,N_6596,N_6846);
and U8424 (N_8424,N_6552,N_7552);
or U8425 (N_8425,N_7155,N_7967);
nand U8426 (N_8426,N_6711,N_6543);
nor U8427 (N_8427,N_7445,N_7597);
or U8428 (N_8428,N_6071,N_7614);
nand U8429 (N_8429,N_7542,N_7104);
nor U8430 (N_8430,N_7065,N_7042);
nor U8431 (N_8431,N_6625,N_7399);
and U8432 (N_8432,N_7659,N_7327);
or U8433 (N_8433,N_7625,N_7932);
and U8434 (N_8434,N_6180,N_6527);
or U8435 (N_8435,N_6086,N_7496);
or U8436 (N_8436,N_6070,N_6461);
nand U8437 (N_8437,N_7688,N_6471);
or U8438 (N_8438,N_7053,N_7958);
or U8439 (N_8439,N_6171,N_6652);
nor U8440 (N_8440,N_6000,N_6029);
and U8441 (N_8441,N_7549,N_6700);
xor U8442 (N_8442,N_7813,N_6873);
nor U8443 (N_8443,N_7330,N_6847);
and U8444 (N_8444,N_6755,N_7238);
and U8445 (N_8445,N_6035,N_6659);
nor U8446 (N_8446,N_6961,N_6187);
or U8447 (N_8447,N_7749,N_6476);
or U8448 (N_8448,N_7713,N_7461);
nor U8449 (N_8449,N_7703,N_6842);
and U8450 (N_8450,N_6705,N_7919);
or U8451 (N_8451,N_7242,N_6499);
or U8452 (N_8452,N_6500,N_6191);
nor U8453 (N_8453,N_7427,N_6633);
or U8454 (N_8454,N_7460,N_6260);
xor U8455 (N_8455,N_7306,N_6722);
or U8456 (N_8456,N_7842,N_6765);
nor U8457 (N_8457,N_6373,N_7256);
nand U8458 (N_8458,N_6513,N_7204);
nand U8459 (N_8459,N_6316,N_6258);
nand U8460 (N_8460,N_6134,N_6358);
and U8461 (N_8461,N_7546,N_7449);
or U8462 (N_8462,N_7305,N_6725);
or U8463 (N_8463,N_7859,N_6042);
and U8464 (N_8464,N_6932,N_7260);
nor U8465 (N_8465,N_6820,N_7855);
or U8466 (N_8466,N_7494,N_7996);
or U8467 (N_8467,N_6229,N_6983);
and U8468 (N_8468,N_6867,N_7580);
nand U8469 (N_8469,N_7038,N_6821);
nand U8470 (N_8470,N_7170,N_6688);
and U8471 (N_8471,N_6898,N_7165);
or U8472 (N_8472,N_6016,N_6721);
nor U8473 (N_8473,N_6128,N_6680);
nand U8474 (N_8474,N_7969,N_7705);
or U8475 (N_8475,N_7244,N_6787);
or U8476 (N_8476,N_7899,N_6827);
xnor U8477 (N_8477,N_7015,N_7166);
nand U8478 (N_8478,N_7190,N_7193);
or U8479 (N_8479,N_6364,N_6423);
and U8480 (N_8480,N_7735,N_6065);
nand U8481 (N_8481,N_7851,N_6401);
or U8482 (N_8482,N_7032,N_6981);
nor U8483 (N_8483,N_7523,N_6594);
nand U8484 (N_8484,N_7482,N_7745);
nor U8485 (N_8485,N_7600,N_6026);
or U8486 (N_8486,N_6060,N_7987);
nand U8487 (N_8487,N_7151,N_6250);
and U8488 (N_8488,N_7555,N_6342);
and U8489 (N_8489,N_7751,N_6694);
or U8490 (N_8490,N_7207,N_7161);
or U8491 (N_8491,N_7918,N_7760);
nand U8492 (N_8492,N_6044,N_6629);
nor U8493 (N_8493,N_6309,N_6758);
nand U8494 (N_8494,N_6151,N_7623);
nor U8495 (N_8495,N_6876,N_7766);
or U8496 (N_8496,N_6427,N_6040);
nand U8497 (N_8497,N_7759,N_6945);
or U8498 (N_8498,N_6855,N_6389);
or U8499 (N_8499,N_7156,N_7671);
or U8500 (N_8500,N_6635,N_7763);
nor U8501 (N_8501,N_6190,N_7102);
and U8502 (N_8502,N_6496,N_6964);
and U8503 (N_8503,N_7140,N_6878);
nor U8504 (N_8504,N_6119,N_7384);
nor U8505 (N_8505,N_7869,N_6524);
nand U8506 (N_8506,N_6107,N_6263);
or U8507 (N_8507,N_6150,N_7008);
and U8508 (N_8508,N_6774,N_7279);
nand U8509 (N_8509,N_7290,N_6715);
and U8510 (N_8510,N_6929,N_7308);
nor U8511 (N_8511,N_7952,N_6706);
nand U8512 (N_8512,N_7820,N_7880);
nor U8513 (N_8513,N_6275,N_7111);
and U8514 (N_8514,N_7030,N_6559);
or U8515 (N_8515,N_6090,N_7802);
nand U8516 (N_8516,N_6277,N_7108);
or U8517 (N_8517,N_7239,N_6464);
or U8518 (N_8518,N_6475,N_7613);
nand U8519 (N_8519,N_6528,N_7642);
or U8520 (N_8520,N_6737,N_7396);
nor U8521 (N_8521,N_7137,N_7866);
nand U8522 (N_8522,N_6729,N_6146);
and U8523 (N_8523,N_6172,N_6088);
and U8524 (N_8524,N_7213,N_7463);
and U8525 (N_8525,N_7979,N_6854);
or U8526 (N_8526,N_7883,N_7247);
or U8527 (N_8527,N_7451,N_7006);
and U8528 (N_8528,N_7232,N_6225);
and U8529 (N_8529,N_7121,N_6849);
and U8530 (N_8530,N_7817,N_6650);
nand U8531 (N_8531,N_7910,N_7754);
nand U8532 (N_8532,N_6131,N_7818);
nand U8533 (N_8533,N_6616,N_6830);
and U8534 (N_8534,N_6222,N_6195);
and U8535 (N_8535,N_7925,N_6006);
and U8536 (N_8536,N_6133,N_6544);
nand U8537 (N_8537,N_7716,N_7915);
nand U8538 (N_8538,N_6756,N_6445);
nand U8539 (N_8539,N_7360,N_6900);
nor U8540 (N_8540,N_7003,N_6183);
or U8541 (N_8541,N_6775,N_6786);
nor U8542 (N_8542,N_7423,N_6952);
and U8543 (N_8543,N_7902,N_6279);
nand U8544 (N_8544,N_6449,N_6385);
xnor U8545 (N_8545,N_6418,N_7473);
nor U8546 (N_8546,N_6991,N_7499);
nand U8547 (N_8547,N_7652,N_6938);
and U8548 (N_8548,N_7135,N_7182);
nor U8549 (N_8549,N_7420,N_7891);
or U8550 (N_8550,N_6299,N_7771);
or U8551 (N_8551,N_6857,N_6011);
or U8552 (N_8552,N_7286,N_7265);
nand U8553 (N_8553,N_7040,N_6359);
nand U8554 (N_8554,N_7929,N_6115);
or U8555 (N_8555,N_6838,N_6507);
nand U8556 (N_8556,N_7441,N_7983);
or U8557 (N_8557,N_6064,N_6577);
nor U8558 (N_8558,N_6553,N_6121);
and U8559 (N_8559,N_6508,N_6412);
xnor U8560 (N_8560,N_7347,N_6665);
or U8561 (N_8561,N_7257,N_7696);
nand U8562 (N_8562,N_6539,N_6382);
and U8563 (N_8563,N_6943,N_6615);
or U8564 (N_8564,N_7630,N_7568);
or U8565 (N_8565,N_6502,N_7480);
nor U8566 (N_8566,N_6697,N_7223);
and U8567 (N_8567,N_7710,N_7129);
nand U8568 (N_8568,N_6224,N_6124);
nor U8569 (N_8569,N_7858,N_7626);
and U8570 (N_8570,N_6634,N_6432);
nor U8571 (N_8571,N_7516,N_7804);
and U8572 (N_8572,N_7629,N_7467);
nor U8573 (N_8573,N_6623,N_6362);
or U8574 (N_8574,N_6300,N_6535);
nor U8575 (N_8575,N_7951,N_6439);
nor U8576 (N_8576,N_6606,N_6638);
nand U8577 (N_8577,N_6407,N_6281);
nand U8578 (N_8578,N_7656,N_7508);
nor U8579 (N_8579,N_6541,N_7584);
and U8580 (N_8580,N_6773,N_6295);
or U8581 (N_8581,N_6467,N_6218);
nor U8582 (N_8582,N_7372,N_6675);
and U8583 (N_8583,N_6398,N_6327);
nor U8584 (N_8584,N_6484,N_7809);
or U8585 (N_8585,N_7326,N_6906);
nor U8586 (N_8586,N_6950,N_6054);
and U8587 (N_8587,N_6979,N_6486);
nor U8588 (N_8588,N_6200,N_7115);
and U8589 (N_8589,N_6897,N_6951);
nand U8590 (N_8590,N_7387,N_7638);
nor U8591 (N_8591,N_7027,N_7665);
nor U8592 (N_8592,N_6708,N_6511);
and U8593 (N_8593,N_7789,N_6661);
or U8594 (N_8594,N_6628,N_7662);
nand U8595 (N_8595,N_6996,N_6656);
or U8596 (N_8596,N_7393,N_7565);
or U8597 (N_8597,N_6349,N_7606);
and U8598 (N_8598,N_7908,N_6771);
nand U8599 (N_8599,N_7558,N_7849);
and U8600 (N_8600,N_7456,N_7462);
nor U8601 (N_8601,N_7336,N_7364);
nor U8602 (N_8602,N_7926,N_6276);
nor U8603 (N_8603,N_6728,N_7608);
and U8604 (N_8604,N_6147,N_7035);
and U8605 (N_8605,N_7785,N_6335);
xnor U8606 (N_8606,N_6130,N_7607);
nand U8607 (N_8607,N_7837,N_6723);
nor U8608 (N_8608,N_7617,N_7479);
and U8609 (N_8609,N_6734,N_6047);
or U8610 (N_8610,N_7429,N_7090);
nand U8611 (N_8611,N_7874,N_6101);
and U8612 (N_8612,N_7370,N_7261);
or U8613 (N_8613,N_6639,N_6759);
and U8614 (N_8614,N_6884,N_6933);
nand U8615 (N_8615,N_6686,N_6621);
or U8616 (N_8616,N_7413,N_6969);
nand U8617 (N_8617,N_7655,N_7443);
and U8618 (N_8618,N_7948,N_6707);
and U8619 (N_8619,N_6506,N_7799);
or U8620 (N_8620,N_6477,N_6441);
and U8621 (N_8621,N_7673,N_7457);
nand U8622 (N_8622,N_6990,N_7654);
nand U8623 (N_8623,N_6550,N_7650);
nor U8624 (N_8624,N_7787,N_7353);
or U8625 (N_8625,N_7559,N_7329);
and U8626 (N_8626,N_6780,N_6244);
nand U8627 (N_8627,N_6426,N_6762);
nor U8628 (N_8628,N_7368,N_7410);
nor U8629 (N_8629,N_7711,N_7941);
or U8630 (N_8630,N_7017,N_7419);
nand U8631 (N_8631,N_7198,N_7535);
and U8632 (N_8632,N_7392,N_6930);
and U8633 (N_8633,N_6285,N_7981);
nor U8634 (N_8634,N_6751,N_6251);
or U8635 (N_8635,N_7978,N_6799);
and U8636 (N_8636,N_6735,N_7278);
nand U8637 (N_8637,N_7864,N_7199);
nand U8638 (N_8638,N_6322,N_7469);
nor U8639 (N_8639,N_7553,N_6890);
nor U8640 (N_8640,N_6416,N_6560);
nand U8641 (N_8641,N_7621,N_7092);
and U8642 (N_8642,N_7328,N_7343);
nand U8643 (N_8643,N_7254,N_6925);
and U8644 (N_8644,N_6085,N_6953);
nor U8645 (N_8645,N_6947,N_7982);
and U8646 (N_8646,N_6853,N_6369);
and U8647 (N_8647,N_6167,N_6334);
and U8648 (N_8648,N_6719,N_7651);
nand U8649 (N_8649,N_6094,N_6754);
and U8650 (N_8650,N_6631,N_7839);
or U8651 (N_8651,N_7571,N_7989);
nor U8652 (N_8652,N_6880,N_7567);
nor U8653 (N_8653,N_7539,N_6266);
nor U8654 (N_8654,N_6575,N_7139);
nor U8655 (N_8655,N_6903,N_7543);
nand U8656 (N_8656,N_7061,N_6843);
nand U8657 (N_8657,N_7570,N_6057);
nand U8658 (N_8658,N_6744,N_7436);
nand U8659 (N_8659,N_7335,N_6782);
nor U8660 (N_8660,N_6881,N_6858);
nand U8661 (N_8661,N_6012,N_7648);
nand U8662 (N_8662,N_7550,N_7016);
and U8663 (N_8663,N_7752,N_7442);
and U8664 (N_8664,N_6595,N_7314);
or U8665 (N_8665,N_6495,N_6455);
nor U8666 (N_8666,N_6778,N_6672);
or U8667 (N_8667,N_7753,N_6448);
and U8668 (N_8668,N_7331,N_7995);
nor U8669 (N_8669,N_6624,N_6547);
or U8670 (N_8670,N_7230,N_6545);
nand U8671 (N_8671,N_6018,N_6904);
nand U8672 (N_8672,N_6092,N_6305);
and U8673 (N_8673,N_7547,N_6483);
and U8674 (N_8674,N_7110,N_7250);
xnor U8675 (N_8675,N_6487,N_6662);
nor U8676 (N_8676,N_7695,N_7246);
nand U8677 (N_8677,N_7118,N_7784);
nor U8678 (N_8678,N_6743,N_7576);
nand U8679 (N_8679,N_6261,N_6727);
nand U8680 (N_8680,N_6120,N_7049);
or U8681 (N_8681,N_6608,N_7439);
nor U8682 (N_8682,N_7408,N_6328);
nand U8683 (N_8683,N_7810,N_6055);
and U8684 (N_8684,N_6645,N_7887);
nor U8685 (N_8685,N_7532,N_6837);
and U8686 (N_8686,N_6415,N_7068);
nor U8687 (N_8687,N_7800,N_7976);
or U8688 (N_8688,N_6913,N_6704);
nor U8689 (N_8689,N_6009,N_7046);
nand U8690 (N_8690,N_6809,N_7269);
or U8691 (N_8691,N_7229,N_7216);
or U8692 (N_8692,N_6954,N_6078);
and U8693 (N_8693,N_7903,N_7767);
nor U8694 (N_8694,N_6866,N_7619);
and U8695 (N_8695,N_7672,N_7487);
and U8696 (N_8696,N_7075,N_7723);
nor U8697 (N_8697,N_7172,N_6056);
nor U8698 (N_8698,N_6668,N_6348);
or U8699 (N_8699,N_6679,N_7453);
nor U8700 (N_8700,N_6361,N_6478);
nor U8701 (N_8701,N_7202,N_6298);
nand U8702 (N_8702,N_7788,N_7047);
nand U8703 (N_8703,N_7325,N_7862);
and U8704 (N_8704,N_6562,N_7380);
nor U8705 (N_8705,N_6216,N_6429);
nand U8706 (N_8706,N_7985,N_6215);
or U8707 (N_8707,N_6447,N_7183);
nor U8708 (N_8708,N_7682,N_7781);
nand U8709 (N_8709,N_6324,N_7627);
or U8710 (N_8710,N_7209,N_7385);
nor U8711 (N_8711,N_7093,N_6051);
or U8712 (N_8712,N_6111,N_6767);
and U8713 (N_8713,N_6641,N_6375);
nor U8714 (N_8714,N_6519,N_6028);
nor U8715 (N_8715,N_7536,N_7997);
and U8716 (N_8716,N_6653,N_6807);
nor U8717 (N_8717,N_7426,N_6572);
or U8718 (N_8718,N_6825,N_7709);
nor U8719 (N_8719,N_7252,N_7589);
nor U8720 (N_8720,N_7574,N_6391);
xnor U8721 (N_8721,N_6845,N_7177);
nor U8722 (N_8722,N_7369,N_6923);
nand U8723 (N_8723,N_6032,N_7888);
or U8724 (N_8724,N_6802,N_6462);
nor U8725 (N_8725,N_6795,N_7815);
or U8726 (N_8726,N_7160,N_6564);
and U8727 (N_8727,N_7107,N_7685);
nand U8728 (N_8728,N_7012,N_6272);
or U8729 (N_8729,N_7200,N_7636);
and U8730 (N_8730,N_6948,N_6386);
nand U8731 (N_8731,N_6137,N_7346);
or U8732 (N_8732,N_7210,N_7409);
nand U8733 (N_8733,N_7371,N_7264);
and U8734 (N_8734,N_6162,N_7066);
or U8735 (N_8735,N_7667,N_6804);
nand U8736 (N_8736,N_6710,N_7415);
or U8737 (N_8737,N_7964,N_7512);
nand U8738 (N_8738,N_7491,N_7150);
and U8739 (N_8739,N_7119,N_6955);
xor U8740 (N_8740,N_7105,N_6901);
nor U8741 (N_8741,N_6236,N_6816);
or U8742 (N_8742,N_6045,N_6245);
or U8743 (N_8743,N_6228,N_7348);
or U8744 (N_8744,N_6366,N_7334);
or U8745 (N_8745,N_7868,N_7633);
and U8746 (N_8746,N_6053,N_6289);
or U8747 (N_8747,N_6674,N_7402);
and U8748 (N_8748,N_7282,N_7271);
or U8749 (N_8749,N_6274,N_6003);
and U8750 (N_8750,N_6068,N_7761);
nand U8751 (N_8751,N_6798,N_6444);
xor U8752 (N_8752,N_6912,N_6379);
nor U8753 (N_8753,N_7477,N_6264);
nor U8754 (N_8754,N_7219,N_7578);
and U8755 (N_8755,N_6390,N_7359);
nand U8756 (N_8756,N_7907,N_6089);
and U8757 (N_8757,N_7267,N_7577);
nor U8758 (N_8758,N_6234,N_7702);
or U8759 (N_8759,N_7999,N_6050);
or U8760 (N_8760,N_7450,N_7721);
nand U8761 (N_8761,N_6303,N_7658);
or U8762 (N_8762,N_6421,N_6978);
or U8763 (N_8763,N_6117,N_7924);
nor U8764 (N_8764,N_7214,N_6655);
and U8765 (N_8765,N_7747,N_6443);
nand U8766 (N_8766,N_6630,N_6436);
xor U8767 (N_8767,N_7741,N_7222);
and U8768 (N_8768,N_7870,N_7694);
nand U8769 (N_8769,N_6741,N_7831);
xor U8770 (N_8770,N_6223,N_6457);
and U8771 (N_8771,N_7954,N_6158);
or U8772 (N_8772,N_7283,N_7455);
or U8773 (N_8773,N_7400,N_6574);
nand U8774 (N_8774,N_6640,N_7287);
and U8775 (N_8775,N_6919,N_6915);
nor U8776 (N_8776,N_6243,N_6340);
or U8777 (N_8777,N_7712,N_6320);
nor U8778 (N_8778,N_7180,N_7520);
or U8779 (N_8779,N_6319,N_7768);
and U8780 (N_8780,N_6714,N_7959);
or U8781 (N_8781,N_6230,N_7692);
and U8782 (N_8782,N_7833,N_6492);
and U8783 (N_8783,N_6083,N_7304);
and U8784 (N_8784,N_7533,N_7853);
and U8785 (N_8785,N_7157,N_7231);
nand U8786 (N_8786,N_6796,N_6360);
or U8787 (N_8787,N_6114,N_6331);
nand U8788 (N_8788,N_6186,N_6329);
nand U8789 (N_8789,N_6458,N_6819);
and U8790 (N_8790,N_6126,N_7808);
and U8791 (N_8791,N_6284,N_6887);
nor U8792 (N_8792,N_6494,N_6514);
nand U8793 (N_8793,N_7486,N_7438);
nor U8794 (N_8794,N_7968,N_6041);
and U8795 (N_8795,N_7437,N_6262);
or U8796 (N_8796,N_6159,N_7755);
nor U8797 (N_8797,N_6875,N_6019);
and U8798 (N_8798,N_7732,N_7943);
nor U8799 (N_8799,N_7004,N_6374);
nand U8800 (N_8800,N_7873,N_6917);
and U8801 (N_8801,N_6803,N_6255);
and U8802 (N_8802,N_7131,N_6061);
xnor U8803 (N_8803,N_7900,N_7495);
and U8804 (N_8804,N_6256,N_6510);
or U8805 (N_8805,N_7126,N_6789);
nor U8806 (N_8806,N_6140,N_7318);
xor U8807 (N_8807,N_6181,N_7933);
nand U8808 (N_8808,N_7321,N_7339);
and U8809 (N_8809,N_6889,N_6660);
or U8810 (N_8810,N_7912,N_6497);
or U8811 (N_8811,N_6138,N_6995);
nor U8812 (N_8812,N_7197,N_7572);
and U8813 (N_8813,N_6766,N_7502);
and U8814 (N_8814,N_6772,N_7689);
nor U8815 (N_8815,N_6246,N_7192);
or U8816 (N_8816,N_7416,N_7292);
and U8817 (N_8817,N_6344,N_6599);
xnor U8818 (N_8818,N_6976,N_7448);
nand U8819 (N_8819,N_6879,N_7184);
nand U8820 (N_8820,N_6801,N_6703);
nor U8821 (N_8821,N_7424,N_6627);
and U8822 (N_8822,N_6760,N_7245);
and U8823 (N_8823,N_6746,N_7704);
nor U8824 (N_8824,N_7701,N_6473);
and U8825 (N_8825,N_7167,N_7220);
and U8826 (N_8826,N_7470,N_7865);
nor U8827 (N_8827,N_7185,N_7357);
nand U8828 (N_8828,N_6175,N_7507);
nor U8829 (N_8829,N_6287,N_6742);
and U8830 (N_8830,N_7940,N_6738);
nor U8831 (N_8831,N_7579,N_7690);
and U8832 (N_8832,N_6474,N_7852);
or U8833 (N_8833,N_6730,N_6237);
nand U8834 (N_8834,N_7814,N_6113);
nor U8835 (N_8835,N_7728,N_7454);
nor U8836 (N_8836,N_7010,N_6105);
or U8837 (N_8837,N_6217,N_6619);
nor U8838 (N_8838,N_7890,N_6091);
or U8839 (N_8839,N_6698,N_7904);
nor U8840 (N_8840,N_7965,N_6176);
xnor U8841 (N_8841,N_6451,N_7635);
nor U8842 (N_8842,N_7972,N_7661);
and U8843 (N_8843,N_7433,N_6610);
nor U8844 (N_8844,N_7293,N_7351);
nand U8845 (N_8845,N_7125,N_7764);
or U8846 (N_8846,N_7285,N_7158);
nor U8847 (N_8847,N_6844,N_7255);
and U8848 (N_8848,N_7796,N_6534);
or U8849 (N_8849,N_6242,N_7896);
or U8850 (N_8850,N_7525,N_6249);
or U8851 (N_8851,N_7937,N_6673);
nor U8852 (N_8852,N_7719,N_6647);
nand U8853 (N_8853,N_7850,N_7805);
or U8854 (N_8854,N_7947,N_6808);
nor U8855 (N_8855,N_6699,N_6008);
and U8856 (N_8856,N_7026,N_7302);
nand U8857 (N_8857,N_7612,N_7734);
nand U8858 (N_8858,N_6013,N_7739);
nor U8859 (N_8859,N_7772,N_7221);
and U8860 (N_8860,N_6632,N_7596);
nor U8861 (N_8861,N_7358,N_7332);
nand U8862 (N_8862,N_6347,N_6814);
or U8863 (N_8863,N_6649,N_7268);
nor U8864 (N_8864,N_7922,N_6367);
and U8865 (N_8865,N_7169,N_7871);
nand U8866 (N_8866,N_7367,N_6834);
nand U8867 (N_8867,N_6607,N_7322);
or U8868 (N_8868,N_6946,N_7834);
nor U8869 (N_8869,N_7428,N_6330);
and U8870 (N_8870,N_6253,N_7757);
or U8871 (N_8871,N_7934,N_7259);
nor U8872 (N_8872,N_6165,N_6252);
or U8873 (N_8873,N_6346,N_6481);
nor U8874 (N_8874,N_6792,N_7506);
nor U8875 (N_8875,N_6926,N_7587);
nor U8876 (N_8876,N_6984,N_6201);
or U8877 (N_8877,N_6059,N_6515);
and U8878 (N_8878,N_6784,N_7354);
nand U8879 (N_8879,N_6598,N_7931);
xor U8880 (N_8880,N_7021,N_6406);
and U8881 (N_8881,N_6294,N_6345);
and U8882 (N_8882,N_7320,N_6935);
nand U8883 (N_8883,N_6818,N_7187);
and U8884 (N_8884,N_6267,N_7323);
nor U8885 (N_8885,N_7923,N_7737);
or U8886 (N_8886,N_6585,N_6428);
and U8887 (N_8887,N_6271,N_6785);
or U8888 (N_8888,N_6468,N_7828);
and U8889 (N_8889,N_6210,N_7488);
and U8890 (N_8890,N_6308,N_7406);
nor U8891 (N_8891,N_7740,N_6944);
and U8892 (N_8892,N_6438,N_7089);
and U8893 (N_8893,N_7394,N_6683);
or U8894 (N_8894,N_7618,N_7099);
nor U8895 (N_8895,N_6720,N_7963);
and U8896 (N_8896,N_7956,N_7270);
or U8897 (N_8897,N_7056,N_6293);
nor U8898 (N_8898,N_7604,N_7517);
or U8899 (N_8899,N_6931,N_7228);
or U8900 (N_8900,N_7096,N_7379);
nand U8901 (N_8901,N_7218,N_7411);
and U8902 (N_8902,N_6567,N_7806);
and U8903 (N_8903,N_6411,N_7081);
or U8904 (N_8904,N_7875,N_6593);
and U8905 (N_8905,N_7598,N_7414);
or U8906 (N_8906,N_7366,N_7622);
nor U8907 (N_8907,N_6959,N_6472);
nor U8908 (N_8908,N_6805,N_6010);
or U8909 (N_8909,N_6671,N_6442);
and U8910 (N_8910,N_7977,N_7762);
nor U8911 (N_8911,N_7841,N_6622);
or U8912 (N_8912,N_7811,N_7881);
or U8913 (N_8913,N_6777,N_7585);
nor U8914 (N_8914,N_7466,N_6960);
and U8915 (N_8915,N_6588,N_6425);
nand U8916 (N_8916,N_7836,N_7503);
and U8917 (N_8917,N_6793,N_6241);
nor U8918 (N_8918,N_6239,N_6618);
and U8919 (N_8919,N_6177,N_7699);
and U8920 (N_8920,N_6226,N_6387);
nor U8921 (N_8921,N_6852,N_7756);
and U8922 (N_8922,N_6551,N_6815);
and U8923 (N_8923,N_7349,N_6265);
nand U8924 (N_8924,N_7188,N_7561);
nor U8925 (N_8925,N_7845,N_6709);
and U8926 (N_8926,N_6828,N_7731);
nor U8927 (N_8927,N_7518,N_7112);
nand U8928 (N_8928,N_7522,N_7094);
nand U8929 (N_8929,N_7531,N_7779);
and U8930 (N_8930,N_7509,N_7048);
nor U8931 (N_8931,N_7434,N_7724);
or U8932 (N_8932,N_6498,N_7643);
nor U8933 (N_8933,N_7829,N_6516);
nand U8934 (N_8934,N_6894,N_7677);
or U8935 (N_8935,N_6685,N_6937);
nand U8936 (N_8936,N_7893,N_6414);
nand U8937 (N_8937,N_6381,N_7632);
or U8938 (N_8938,N_6962,N_6549);
or U8939 (N_8939,N_7422,N_7843);
nand U8940 (N_8940,N_6521,N_6139);
nand U8941 (N_8941,N_7132,N_7960);
or U8942 (N_8942,N_6469,N_6987);
or U8943 (N_8943,N_7085,N_6355);
nand U8944 (N_8944,N_6928,N_6501);
or U8945 (N_8945,N_7714,N_6268);
or U8946 (N_8946,N_7076,N_6377);
or U8947 (N_8947,N_7863,N_7476);
nor U8948 (N_8948,N_6178,N_6589);
nor U8949 (N_8949,N_6104,N_6123);
or U8950 (N_8950,N_7670,N_6097);
and U8951 (N_8951,N_7631,N_6440);
or U8952 (N_8952,N_6812,N_7720);
or U8953 (N_8953,N_6286,N_6014);
nor U8954 (N_8954,N_6934,N_7052);
nand U8955 (N_8955,N_7774,N_6587);
nand U8956 (N_8956,N_7375,N_7122);
nand U8957 (N_8957,N_7178,N_6740);
nor U8958 (N_8958,N_6985,N_7603);
or U8959 (N_8959,N_6163,N_6522);
or U8960 (N_8960,N_7775,N_7313);
and U8961 (N_8961,N_7143,N_7309);
or U8962 (N_8962,N_7031,N_6192);
nand U8963 (N_8963,N_6062,N_7101);
nor U8964 (N_8964,N_7074,N_7386);
or U8965 (N_8965,N_7317,N_6895);
nand U8966 (N_8966,N_7024,N_6154);
xnor U8967 (N_8967,N_7592,N_7521);
and U8968 (N_8968,N_7154,N_6048);
or U8969 (N_8969,N_6356,N_6921);
and U8970 (N_8970,N_7994,N_6435);
nor U8971 (N_8971,N_7986,N_6399);
nor U8972 (N_8972,N_7352,N_7715);
nand U8973 (N_8973,N_7501,N_6584);
nor U8974 (N_8974,N_6238,N_6023);
or U8975 (N_8975,N_6942,N_6612);
and U8976 (N_8976,N_6148,N_7144);
nor U8977 (N_8977,N_7145,N_6530);
and U8978 (N_8978,N_6002,N_7315);
xnor U8979 (N_8979,N_7014,N_7179);
nor U8980 (N_8980,N_7515,N_7974);
nand U8981 (N_8981,N_7706,N_6998);
nor U8982 (N_8982,N_6603,N_7472);
nand U8983 (N_8983,N_6296,N_6184);
or U8984 (N_8984,N_7726,N_7272);
and U8985 (N_8985,N_7538,N_7921);
nand U8986 (N_8986,N_7641,N_7510);
nand U8987 (N_8987,N_7064,N_6586);
nor U8988 (N_8988,N_6096,N_7973);
nor U8989 (N_8989,N_7007,N_6341);
nor U8990 (N_8990,N_6833,N_7718);
nor U8991 (N_8991,N_7063,N_6788);
nor U8992 (N_8992,N_7430,N_7296);
nand U8993 (N_8993,N_7595,N_7481);
or U8994 (N_8994,N_7471,N_7830);
nand U8995 (N_8995,N_6769,N_7289);
or U8996 (N_8996,N_7894,N_6642);
nor U8997 (N_8997,N_6523,N_6025);
nor U8998 (N_8998,N_7765,N_6690);
or U8999 (N_8999,N_7067,N_7876);
and U9000 (N_9000,N_7195,N_7899);
and U9001 (N_9001,N_6434,N_7721);
or U9002 (N_9002,N_7089,N_7613);
nand U9003 (N_9003,N_6220,N_7967);
and U9004 (N_9004,N_7944,N_6720);
or U9005 (N_9005,N_7602,N_7126);
nor U9006 (N_9006,N_7151,N_7051);
nor U9007 (N_9007,N_6431,N_6878);
nor U9008 (N_9008,N_6045,N_7518);
and U9009 (N_9009,N_6023,N_7120);
and U9010 (N_9010,N_6904,N_6823);
and U9011 (N_9011,N_6838,N_6622);
nor U9012 (N_9012,N_6460,N_7861);
and U9013 (N_9013,N_7145,N_7935);
and U9014 (N_9014,N_6242,N_6679);
and U9015 (N_9015,N_6035,N_6981);
and U9016 (N_9016,N_6756,N_6935);
and U9017 (N_9017,N_7863,N_6378);
nand U9018 (N_9018,N_6557,N_6142);
and U9019 (N_9019,N_6210,N_6267);
nor U9020 (N_9020,N_6105,N_7486);
nand U9021 (N_9021,N_6606,N_6134);
nand U9022 (N_9022,N_6251,N_7226);
nand U9023 (N_9023,N_6689,N_6625);
nand U9024 (N_9024,N_7302,N_6999);
nand U9025 (N_9025,N_7703,N_7994);
or U9026 (N_9026,N_6052,N_6168);
nor U9027 (N_9027,N_7131,N_7371);
and U9028 (N_9028,N_7088,N_6553);
nor U9029 (N_9029,N_6861,N_7669);
nor U9030 (N_9030,N_7394,N_6573);
xnor U9031 (N_9031,N_6691,N_7193);
or U9032 (N_9032,N_6540,N_6648);
nand U9033 (N_9033,N_6601,N_6342);
and U9034 (N_9034,N_6851,N_7342);
and U9035 (N_9035,N_6389,N_7858);
nor U9036 (N_9036,N_7392,N_7476);
and U9037 (N_9037,N_6433,N_6639);
or U9038 (N_9038,N_6169,N_6774);
nand U9039 (N_9039,N_6030,N_7686);
nor U9040 (N_9040,N_7619,N_7871);
nand U9041 (N_9041,N_6471,N_7463);
nor U9042 (N_9042,N_6833,N_6216);
and U9043 (N_9043,N_6690,N_7016);
or U9044 (N_9044,N_7031,N_6412);
nand U9045 (N_9045,N_6153,N_6821);
and U9046 (N_9046,N_6676,N_6802);
nor U9047 (N_9047,N_6339,N_6836);
nand U9048 (N_9048,N_7695,N_6808);
nor U9049 (N_9049,N_7253,N_6628);
and U9050 (N_9050,N_6972,N_6857);
nand U9051 (N_9051,N_6343,N_6492);
and U9052 (N_9052,N_7694,N_6497);
or U9053 (N_9053,N_7423,N_7654);
nand U9054 (N_9054,N_6120,N_6668);
and U9055 (N_9055,N_6429,N_7319);
nand U9056 (N_9056,N_7322,N_7276);
and U9057 (N_9057,N_6546,N_6859);
nor U9058 (N_9058,N_7738,N_7926);
or U9059 (N_9059,N_6237,N_7577);
or U9060 (N_9060,N_6159,N_6274);
nor U9061 (N_9061,N_7481,N_6403);
nand U9062 (N_9062,N_6980,N_7110);
nand U9063 (N_9063,N_6139,N_6552);
nand U9064 (N_9064,N_7432,N_7444);
and U9065 (N_9065,N_7729,N_7928);
or U9066 (N_9066,N_6751,N_7768);
and U9067 (N_9067,N_7335,N_6774);
or U9068 (N_9068,N_6434,N_6220);
nand U9069 (N_9069,N_6827,N_6341);
nor U9070 (N_9070,N_7983,N_6842);
nand U9071 (N_9071,N_6781,N_7295);
and U9072 (N_9072,N_7520,N_6262);
or U9073 (N_9073,N_7606,N_7101);
nor U9074 (N_9074,N_7957,N_6187);
xnor U9075 (N_9075,N_6044,N_7262);
and U9076 (N_9076,N_6033,N_7524);
nand U9077 (N_9077,N_6238,N_7719);
nor U9078 (N_9078,N_6666,N_6098);
nand U9079 (N_9079,N_6205,N_6762);
nor U9080 (N_9080,N_7706,N_6162);
and U9081 (N_9081,N_6099,N_7025);
nor U9082 (N_9082,N_6323,N_7664);
or U9083 (N_9083,N_7869,N_6003);
nor U9084 (N_9084,N_7129,N_7604);
and U9085 (N_9085,N_7571,N_7906);
and U9086 (N_9086,N_7801,N_6456);
or U9087 (N_9087,N_6247,N_7674);
and U9088 (N_9088,N_7912,N_7538);
xnor U9089 (N_9089,N_6485,N_7527);
nor U9090 (N_9090,N_7821,N_6773);
and U9091 (N_9091,N_6769,N_6954);
nand U9092 (N_9092,N_6704,N_7004);
nor U9093 (N_9093,N_6717,N_7749);
and U9094 (N_9094,N_7236,N_7525);
nand U9095 (N_9095,N_6924,N_6847);
nand U9096 (N_9096,N_6327,N_6197);
nand U9097 (N_9097,N_6080,N_6016);
nand U9098 (N_9098,N_6700,N_6961);
nor U9099 (N_9099,N_6599,N_7392);
nor U9100 (N_9100,N_6317,N_7831);
and U9101 (N_9101,N_6950,N_6192);
or U9102 (N_9102,N_6179,N_6642);
and U9103 (N_9103,N_7492,N_6862);
nand U9104 (N_9104,N_7736,N_7441);
or U9105 (N_9105,N_7452,N_7691);
and U9106 (N_9106,N_7651,N_6561);
nand U9107 (N_9107,N_7952,N_7266);
or U9108 (N_9108,N_6118,N_6815);
nand U9109 (N_9109,N_7624,N_6693);
and U9110 (N_9110,N_6237,N_7673);
nor U9111 (N_9111,N_7881,N_6199);
or U9112 (N_9112,N_6368,N_6998);
and U9113 (N_9113,N_7728,N_6331);
or U9114 (N_9114,N_7482,N_6075);
and U9115 (N_9115,N_6647,N_7808);
nor U9116 (N_9116,N_6213,N_7287);
or U9117 (N_9117,N_7203,N_7737);
nor U9118 (N_9118,N_7156,N_7776);
nand U9119 (N_9119,N_6814,N_7445);
nor U9120 (N_9120,N_6817,N_6112);
xor U9121 (N_9121,N_7185,N_6502);
and U9122 (N_9122,N_7158,N_6287);
or U9123 (N_9123,N_7261,N_7604);
or U9124 (N_9124,N_7877,N_7229);
or U9125 (N_9125,N_6411,N_6675);
or U9126 (N_9126,N_6427,N_6418);
and U9127 (N_9127,N_6957,N_7458);
nor U9128 (N_9128,N_6712,N_6447);
and U9129 (N_9129,N_7308,N_7976);
nor U9130 (N_9130,N_7211,N_6940);
and U9131 (N_9131,N_7638,N_6903);
or U9132 (N_9132,N_6205,N_7090);
nand U9133 (N_9133,N_7758,N_7152);
or U9134 (N_9134,N_7243,N_6345);
or U9135 (N_9135,N_7965,N_6888);
nor U9136 (N_9136,N_7812,N_7681);
nand U9137 (N_9137,N_7545,N_6972);
nor U9138 (N_9138,N_7827,N_7068);
nor U9139 (N_9139,N_7895,N_7624);
or U9140 (N_9140,N_7432,N_6659);
and U9141 (N_9141,N_7036,N_7367);
nor U9142 (N_9142,N_6990,N_6789);
or U9143 (N_9143,N_6228,N_6328);
and U9144 (N_9144,N_7686,N_6279);
and U9145 (N_9145,N_6672,N_7389);
nor U9146 (N_9146,N_6858,N_7609);
or U9147 (N_9147,N_6159,N_6353);
and U9148 (N_9148,N_6485,N_6559);
and U9149 (N_9149,N_6988,N_6672);
nor U9150 (N_9150,N_7242,N_7337);
or U9151 (N_9151,N_6738,N_7647);
nor U9152 (N_9152,N_6217,N_7298);
and U9153 (N_9153,N_6603,N_7509);
and U9154 (N_9154,N_6275,N_6825);
nor U9155 (N_9155,N_7671,N_6548);
or U9156 (N_9156,N_6392,N_6315);
and U9157 (N_9157,N_7955,N_6754);
or U9158 (N_9158,N_6664,N_6973);
or U9159 (N_9159,N_6359,N_6363);
nor U9160 (N_9160,N_6020,N_6472);
or U9161 (N_9161,N_7740,N_7874);
nand U9162 (N_9162,N_7334,N_7170);
and U9163 (N_9163,N_7664,N_6908);
nor U9164 (N_9164,N_6787,N_7291);
and U9165 (N_9165,N_7250,N_6629);
or U9166 (N_9166,N_6866,N_7638);
and U9167 (N_9167,N_6602,N_6708);
nand U9168 (N_9168,N_7870,N_6506);
nor U9169 (N_9169,N_6030,N_7030);
nor U9170 (N_9170,N_6469,N_7827);
nor U9171 (N_9171,N_6041,N_7317);
nand U9172 (N_9172,N_6384,N_6431);
nand U9173 (N_9173,N_7259,N_6112);
or U9174 (N_9174,N_7756,N_7059);
and U9175 (N_9175,N_6359,N_7868);
nor U9176 (N_9176,N_6491,N_7548);
nand U9177 (N_9177,N_7091,N_7353);
and U9178 (N_9178,N_6171,N_7169);
nor U9179 (N_9179,N_7855,N_7130);
or U9180 (N_9180,N_6846,N_7420);
xor U9181 (N_9181,N_6697,N_7683);
and U9182 (N_9182,N_7644,N_6916);
nor U9183 (N_9183,N_7689,N_7793);
nand U9184 (N_9184,N_7789,N_7306);
nor U9185 (N_9185,N_6926,N_6868);
or U9186 (N_9186,N_7599,N_7397);
nand U9187 (N_9187,N_7403,N_7842);
and U9188 (N_9188,N_7708,N_6334);
nand U9189 (N_9189,N_7716,N_7195);
nor U9190 (N_9190,N_7452,N_7507);
nand U9191 (N_9191,N_6157,N_7228);
and U9192 (N_9192,N_6995,N_7850);
nand U9193 (N_9193,N_7573,N_7023);
nor U9194 (N_9194,N_6952,N_6019);
and U9195 (N_9195,N_7546,N_6777);
nor U9196 (N_9196,N_6432,N_6161);
or U9197 (N_9197,N_7974,N_7232);
nor U9198 (N_9198,N_7282,N_7046);
xnor U9199 (N_9199,N_6157,N_6911);
and U9200 (N_9200,N_7313,N_7119);
or U9201 (N_9201,N_6518,N_7579);
nor U9202 (N_9202,N_6838,N_7013);
xnor U9203 (N_9203,N_6612,N_6670);
and U9204 (N_9204,N_7172,N_6566);
or U9205 (N_9205,N_7862,N_7079);
nand U9206 (N_9206,N_6734,N_7989);
nor U9207 (N_9207,N_7635,N_6939);
nand U9208 (N_9208,N_7728,N_7664);
nor U9209 (N_9209,N_7664,N_7241);
nand U9210 (N_9210,N_6717,N_7966);
nand U9211 (N_9211,N_6153,N_7022);
nor U9212 (N_9212,N_6582,N_6665);
and U9213 (N_9213,N_6143,N_6485);
nand U9214 (N_9214,N_7441,N_6270);
and U9215 (N_9215,N_6614,N_6960);
nor U9216 (N_9216,N_6350,N_7412);
nand U9217 (N_9217,N_7886,N_7998);
nor U9218 (N_9218,N_7419,N_7289);
and U9219 (N_9219,N_6914,N_6526);
nand U9220 (N_9220,N_7120,N_6077);
nor U9221 (N_9221,N_6408,N_7440);
and U9222 (N_9222,N_7551,N_6606);
and U9223 (N_9223,N_6227,N_6012);
or U9224 (N_9224,N_6059,N_6793);
nor U9225 (N_9225,N_6053,N_7520);
or U9226 (N_9226,N_6466,N_7447);
nand U9227 (N_9227,N_7195,N_7517);
nor U9228 (N_9228,N_7628,N_6526);
or U9229 (N_9229,N_7093,N_6871);
nand U9230 (N_9230,N_6413,N_6766);
and U9231 (N_9231,N_7612,N_6805);
or U9232 (N_9232,N_7554,N_6845);
or U9233 (N_9233,N_7266,N_6803);
nand U9234 (N_9234,N_7654,N_6864);
nand U9235 (N_9235,N_6965,N_7962);
and U9236 (N_9236,N_7614,N_7564);
nand U9237 (N_9237,N_7551,N_6338);
or U9238 (N_9238,N_6857,N_7948);
or U9239 (N_9239,N_7317,N_7638);
nor U9240 (N_9240,N_7227,N_6625);
nor U9241 (N_9241,N_6021,N_7147);
nor U9242 (N_9242,N_6783,N_6147);
nor U9243 (N_9243,N_7524,N_7984);
nand U9244 (N_9244,N_6631,N_7298);
nor U9245 (N_9245,N_6381,N_7845);
nor U9246 (N_9246,N_7709,N_7757);
or U9247 (N_9247,N_6593,N_7846);
and U9248 (N_9248,N_7037,N_7332);
and U9249 (N_9249,N_6314,N_6327);
and U9250 (N_9250,N_7599,N_6739);
and U9251 (N_9251,N_7297,N_7772);
nand U9252 (N_9252,N_7301,N_6965);
and U9253 (N_9253,N_7614,N_6028);
and U9254 (N_9254,N_7302,N_6393);
and U9255 (N_9255,N_6516,N_7388);
nand U9256 (N_9256,N_6849,N_6248);
xnor U9257 (N_9257,N_7752,N_7117);
and U9258 (N_9258,N_7536,N_6183);
nand U9259 (N_9259,N_6236,N_7701);
and U9260 (N_9260,N_6666,N_6856);
or U9261 (N_9261,N_6205,N_6383);
nand U9262 (N_9262,N_7225,N_7244);
and U9263 (N_9263,N_6869,N_7786);
nor U9264 (N_9264,N_6148,N_7077);
or U9265 (N_9265,N_6629,N_7431);
or U9266 (N_9266,N_7882,N_6965);
nor U9267 (N_9267,N_6540,N_6487);
or U9268 (N_9268,N_6857,N_7566);
nand U9269 (N_9269,N_7991,N_7772);
or U9270 (N_9270,N_7127,N_7100);
or U9271 (N_9271,N_6052,N_6291);
nand U9272 (N_9272,N_7992,N_6757);
or U9273 (N_9273,N_7722,N_6975);
or U9274 (N_9274,N_7525,N_7074);
xnor U9275 (N_9275,N_7720,N_7189);
and U9276 (N_9276,N_7079,N_7228);
nand U9277 (N_9277,N_6114,N_6783);
and U9278 (N_9278,N_7945,N_7730);
nand U9279 (N_9279,N_6354,N_6408);
nand U9280 (N_9280,N_7598,N_6622);
nor U9281 (N_9281,N_7576,N_6794);
or U9282 (N_9282,N_6329,N_7892);
xnor U9283 (N_9283,N_7510,N_7504);
nand U9284 (N_9284,N_6022,N_7100);
and U9285 (N_9285,N_7226,N_7245);
and U9286 (N_9286,N_6374,N_7255);
nand U9287 (N_9287,N_7323,N_6694);
nor U9288 (N_9288,N_6839,N_7194);
nand U9289 (N_9289,N_7347,N_6679);
and U9290 (N_9290,N_7037,N_6033);
or U9291 (N_9291,N_7282,N_6491);
and U9292 (N_9292,N_7201,N_7974);
or U9293 (N_9293,N_6092,N_6482);
nor U9294 (N_9294,N_7523,N_6959);
nand U9295 (N_9295,N_7632,N_7612);
or U9296 (N_9296,N_6544,N_7224);
nand U9297 (N_9297,N_6410,N_7602);
or U9298 (N_9298,N_6531,N_6084);
or U9299 (N_9299,N_7990,N_7200);
and U9300 (N_9300,N_6089,N_6941);
nor U9301 (N_9301,N_6815,N_7172);
and U9302 (N_9302,N_7123,N_7792);
and U9303 (N_9303,N_6689,N_6094);
and U9304 (N_9304,N_7059,N_6057);
nor U9305 (N_9305,N_7037,N_6600);
and U9306 (N_9306,N_7502,N_6426);
nor U9307 (N_9307,N_6439,N_6332);
and U9308 (N_9308,N_7919,N_6786);
nor U9309 (N_9309,N_6181,N_7583);
and U9310 (N_9310,N_7822,N_6700);
or U9311 (N_9311,N_7712,N_6806);
nand U9312 (N_9312,N_7100,N_6467);
and U9313 (N_9313,N_6035,N_7350);
nor U9314 (N_9314,N_6857,N_7685);
or U9315 (N_9315,N_7299,N_7980);
or U9316 (N_9316,N_6713,N_6326);
or U9317 (N_9317,N_7906,N_7752);
or U9318 (N_9318,N_6688,N_7005);
nor U9319 (N_9319,N_6539,N_7705);
or U9320 (N_9320,N_7097,N_6441);
nand U9321 (N_9321,N_6869,N_6957);
nand U9322 (N_9322,N_6731,N_7518);
and U9323 (N_9323,N_6683,N_6436);
or U9324 (N_9324,N_6794,N_7097);
nand U9325 (N_9325,N_7329,N_7927);
nor U9326 (N_9326,N_7707,N_6314);
nand U9327 (N_9327,N_6284,N_6256);
and U9328 (N_9328,N_6649,N_7903);
nor U9329 (N_9329,N_6831,N_6649);
nand U9330 (N_9330,N_7495,N_6801);
nor U9331 (N_9331,N_7791,N_7017);
nor U9332 (N_9332,N_6819,N_7165);
nor U9333 (N_9333,N_6300,N_7047);
and U9334 (N_9334,N_7654,N_6908);
nand U9335 (N_9335,N_7218,N_7314);
nand U9336 (N_9336,N_6323,N_6313);
nor U9337 (N_9337,N_6436,N_6813);
nor U9338 (N_9338,N_7526,N_6981);
nand U9339 (N_9339,N_7924,N_7658);
nor U9340 (N_9340,N_6296,N_6525);
or U9341 (N_9341,N_7359,N_6883);
nor U9342 (N_9342,N_6031,N_7222);
or U9343 (N_9343,N_7273,N_6100);
and U9344 (N_9344,N_7209,N_6432);
nand U9345 (N_9345,N_7305,N_7911);
nand U9346 (N_9346,N_6050,N_7387);
nand U9347 (N_9347,N_6282,N_6532);
and U9348 (N_9348,N_7932,N_7610);
nand U9349 (N_9349,N_6701,N_6369);
or U9350 (N_9350,N_7509,N_7596);
nand U9351 (N_9351,N_6226,N_7998);
or U9352 (N_9352,N_6101,N_7582);
nand U9353 (N_9353,N_7817,N_6561);
and U9354 (N_9354,N_7380,N_6929);
or U9355 (N_9355,N_6164,N_6543);
or U9356 (N_9356,N_6873,N_7199);
and U9357 (N_9357,N_7578,N_6109);
and U9358 (N_9358,N_7808,N_7528);
xnor U9359 (N_9359,N_6414,N_6656);
nor U9360 (N_9360,N_6116,N_7130);
or U9361 (N_9361,N_6336,N_7286);
nor U9362 (N_9362,N_6557,N_7336);
and U9363 (N_9363,N_6072,N_6820);
and U9364 (N_9364,N_6262,N_6517);
or U9365 (N_9365,N_6711,N_6081);
and U9366 (N_9366,N_7733,N_6766);
nand U9367 (N_9367,N_7769,N_7951);
nand U9368 (N_9368,N_7055,N_6628);
nand U9369 (N_9369,N_7242,N_7101);
nor U9370 (N_9370,N_6670,N_6723);
nor U9371 (N_9371,N_7304,N_6311);
nand U9372 (N_9372,N_6798,N_7204);
nand U9373 (N_9373,N_6445,N_6774);
nand U9374 (N_9374,N_7830,N_6838);
nand U9375 (N_9375,N_6450,N_6541);
nor U9376 (N_9376,N_6563,N_7107);
and U9377 (N_9377,N_7660,N_6359);
nand U9378 (N_9378,N_7203,N_6552);
nand U9379 (N_9379,N_7818,N_6127);
nor U9380 (N_9380,N_6813,N_6839);
nand U9381 (N_9381,N_6510,N_7071);
nor U9382 (N_9382,N_7365,N_7528);
nand U9383 (N_9383,N_7046,N_7248);
and U9384 (N_9384,N_6710,N_6112);
or U9385 (N_9385,N_7137,N_7163);
and U9386 (N_9386,N_6444,N_7494);
or U9387 (N_9387,N_6394,N_6016);
nor U9388 (N_9388,N_6705,N_7650);
and U9389 (N_9389,N_7650,N_7976);
nor U9390 (N_9390,N_6250,N_7497);
or U9391 (N_9391,N_6403,N_7492);
and U9392 (N_9392,N_7176,N_6105);
nor U9393 (N_9393,N_7273,N_7838);
nand U9394 (N_9394,N_7585,N_7351);
or U9395 (N_9395,N_6567,N_6696);
and U9396 (N_9396,N_7842,N_6179);
nor U9397 (N_9397,N_7842,N_7333);
or U9398 (N_9398,N_6036,N_6840);
nand U9399 (N_9399,N_7061,N_6882);
and U9400 (N_9400,N_7672,N_6618);
nor U9401 (N_9401,N_6822,N_6018);
and U9402 (N_9402,N_7465,N_6507);
nand U9403 (N_9403,N_6695,N_6877);
nor U9404 (N_9404,N_6084,N_6528);
nor U9405 (N_9405,N_7355,N_7235);
or U9406 (N_9406,N_7736,N_6468);
xnor U9407 (N_9407,N_7568,N_6918);
or U9408 (N_9408,N_6759,N_7761);
or U9409 (N_9409,N_7586,N_7837);
nor U9410 (N_9410,N_7070,N_6636);
or U9411 (N_9411,N_6525,N_7030);
nor U9412 (N_9412,N_7725,N_7481);
or U9413 (N_9413,N_7347,N_6565);
or U9414 (N_9414,N_7241,N_6965);
nor U9415 (N_9415,N_6437,N_7457);
and U9416 (N_9416,N_7498,N_7077);
nand U9417 (N_9417,N_7605,N_7896);
or U9418 (N_9418,N_6838,N_6834);
nor U9419 (N_9419,N_6786,N_7632);
nand U9420 (N_9420,N_6879,N_6419);
and U9421 (N_9421,N_6495,N_7841);
and U9422 (N_9422,N_7902,N_6950);
or U9423 (N_9423,N_7421,N_6152);
or U9424 (N_9424,N_6591,N_7593);
and U9425 (N_9425,N_6472,N_7227);
nor U9426 (N_9426,N_6219,N_7685);
or U9427 (N_9427,N_6339,N_7774);
and U9428 (N_9428,N_7849,N_7299);
or U9429 (N_9429,N_7312,N_6560);
nand U9430 (N_9430,N_7707,N_7617);
nor U9431 (N_9431,N_7606,N_7168);
nand U9432 (N_9432,N_6170,N_7008);
or U9433 (N_9433,N_6224,N_7046);
nor U9434 (N_9434,N_6898,N_6194);
and U9435 (N_9435,N_7744,N_6346);
nand U9436 (N_9436,N_7708,N_6658);
and U9437 (N_9437,N_6402,N_7285);
xor U9438 (N_9438,N_7676,N_7600);
and U9439 (N_9439,N_7251,N_6099);
or U9440 (N_9440,N_6548,N_7864);
nor U9441 (N_9441,N_6947,N_7970);
and U9442 (N_9442,N_7555,N_6743);
nor U9443 (N_9443,N_6092,N_7056);
and U9444 (N_9444,N_6388,N_7107);
nor U9445 (N_9445,N_7081,N_7470);
nand U9446 (N_9446,N_6415,N_7720);
nand U9447 (N_9447,N_7501,N_7699);
nand U9448 (N_9448,N_7209,N_7633);
nor U9449 (N_9449,N_7316,N_6713);
nand U9450 (N_9450,N_6644,N_7922);
nand U9451 (N_9451,N_7081,N_6641);
nand U9452 (N_9452,N_6193,N_6305);
nand U9453 (N_9453,N_6340,N_6956);
nand U9454 (N_9454,N_6273,N_6570);
or U9455 (N_9455,N_7226,N_7745);
nor U9456 (N_9456,N_7429,N_7098);
or U9457 (N_9457,N_6733,N_6565);
or U9458 (N_9458,N_6203,N_7998);
and U9459 (N_9459,N_6764,N_7104);
or U9460 (N_9460,N_6548,N_6143);
nand U9461 (N_9461,N_6564,N_7473);
or U9462 (N_9462,N_6239,N_6431);
nand U9463 (N_9463,N_7678,N_7599);
nor U9464 (N_9464,N_6491,N_6913);
or U9465 (N_9465,N_6339,N_6642);
nand U9466 (N_9466,N_7625,N_6615);
nor U9467 (N_9467,N_6623,N_6810);
nand U9468 (N_9468,N_6563,N_7549);
and U9469 (N_9469,N_6365,N_6311);
and U9470 (N_9470,N_7863,N_6401);
and U9471 (N_9471,N_7490,N_6283);
nand U9472 (N_9472,N_6673,N_7727);
or U9473 (N_9473,N_6589,N_6705);
nand U9474 (N_9474,N_7701,N_6676);
nor U9475 (N_9475,N_6059,N_6866);
nor U9476 (N_9476,N_7682,N_6182);
nor U9477 (N_9477,N_7164,N_6836);
and U9478 (N_9478,N_6973,N_6967);
or U9479 (N_9479,N_6594,N_7686);
nor U9480 (N_9480,N_6908,N_7743);
or U9481 (N_9481,N_7508,N_7118);
or U9482 (N_9482,N_6184,N_7159);
and U9483 (N_9483,N_7399,N_7755);
nand U9484 (N_9484,N_7891,N_6534);
nand U9485 (N_9485,N_6565,N_6739);
nand U9486 (N_9486,N_7933,N_6958);
nand U9487 (N_9487,N_6691,N_7865);
or U9488 (N_9488,N_6294,N_6489);
nor U9489 (N_9489,N_7071,N_7804);
or U9490 (N_9490,N_6328,N_6996);
and U9491 (N_9491,N_6143,N_7772);
or U9492 (N_9492,N_6006,N_6900);
nor U9493 (N_9493,N_6232,N_6253);
or U9494 (N_9494,N_7476,N_6858);
or U9495 (N_9495,N_7606,N_7958);
or U9496 (N_9496,N_7103,N_6867);
and U9497 (N_9497,N_7918,N_6309);
nand U9498 (N_9498,N_7896,N_6955);
and U9499 (N_9499,N_6945,N_6041);
nor U9500 (N_9500,N_6021,N_6058);
nor U9501 (N_9501,N_7244,N_7080);
or U9502 (N_9502,N_7814,N_6953);
nor U9503 (N_9503,N_6603,N_6041);
nand U9504 (N_9504,N_7556,N_7749);
nand U9505 (N_9505,N_7952,N_7892);
or U9506 (N_9506,N_7113,N_7973);
and U9507 (N_9507,N_7353,N_6858);
and U9508 (N_9508,N_6304,N_6579);
or U9509 (N_9509,N_7376,N_7757);
nor U9510 (N_9510,N_6809,N_7895);
nor U9511 (N_9511,N_7515,N_7326);
nand U9512 (N_9512,N_7732,N_6780);
nand U9513 (N_9513,N_7643,N_6334);
and U9514 (N_9514,N_7941,N_6120);
nor U9515 (N_9515,N_6028,N_7455);
or U9516 (N_9516,N_6350,N_6585);
nand U9517 (N_9517,N_6853,N_6648);
or U9518 (N_9518,N_6308,N_6941);
and U9519 (N_9519,N_7283,N_7604);
or U9520 (N_9520,N_6945,N_7945);
nand U9521 (N_9521,N_6266,N_7139);
or U9522 (N_9522,N_7845,N_6402);
and U9523 (N_9523,N_6394,N_6702);
nor U9524 (N_9524,N_6339,N_7816);
nand U9525 (N_9525,N_6576,N_6368);
or U9526 (N_9526,N_7403,N_6617);
nand U9527 (N_9527,N_6422,N_7873);
nand U9528 (N_9528,N_7269,N_7822);
nor U9529 (N_9529,N_6984,N_6465);
or U9530 (N_9530,N_6658,N_7880);
nor U9531 (N_9531,N_7491,N_6891);
and U9532 (N_9532,N_6858,N_7442);
and U9533 (N_9533,N_6797,N_6942);
or U9534 (N_9534,N_6098,N_7502);
or U9535 (N_9535,N_7043,N_7921);
or U9536 (N_9536,N_7465,N_6343);
and U9537 (N_9537,N_6169,N_6124);
or U9538 (N_9538,N_6902,N_6753);
and U9539 (N_9539,N_6077,N_6044);
or U9540 (N_9540,N_7225,N_6319);
nand U9541 (N_9541,N_6639,N_6028);
nor U9542 (N_9542,N_6693,N_6123);
or U9543 (N_9543,N_6300,N_6359);
and U9544 (N_9544,N_6331,N_7112);
and U9545 (N_9545,N_6345,N_7099);
nand U9546 (N_9546,N_6348,N_6328);
or U9547 (N_9547,N_7101,N_7974);
or U9548 (N_9548,N_7254,N_6238);
nor U9549 (N_9549,N_6951,N_7647);
nand U9550 (N_9550,N_6142,N_6901);
nand U9551 (N_9551,N_6731,N_7166);
and U9552 (N_9552,N_6206,N_6806);
or U9553 (N_9553,N_6995,N_6400);
or U9554 (N_9554,N_6848,N_7681);
nor U9555 (N_9555,N_7347,N_7643);
nand U9556 (N_9556,N_7343,N_6305);
nor U9557 (N_9557,N_7228,N_7508);
and U9558 (N_9558,N_6926,N_7886);
nand U9559 (N_9559,N_6273,N_7721);
nand U9560 (N_9560,N_7130,N_6091);
nor U9561 (N_9561,N_7822,N_7424);
nand U9562 (N_9562,N_7862,N_7351);
nor U9563 (N_9563,N_6289,N_7933);
nor U9564 (N_9564,N_6003,N_6806);
nand U9565 (N_9565,N_7950,N_6127);
nand U9566 (N_9566,N_7933,N_7849);
or U9567 (N_9567,N_7545,N_7855);
nand U9568 (N_9568,N_6391,N_7058);
and U9569 (N_9569,N_7937,N_7437);
nand U9570 (N_9570,N_6131,N_7648);
nand U9571 (N_9571,N_7015,N_7130);
nor U9572 (N_9572,N_7314,N_6080);
or U9573 (N_9573,N_7022,N_6860);
nand U9574 (N_9574,N_7802,N_7969);
nand U9575 (N_9575,N_7599,N_7714);
nand U9576 (N_9576,N_7666,N_7158);
nor U9577 (N_9577,N_6810,N_6043);
and U9578 (N_9578,N_7546,N_6492);
nand U9579 (N_9579,N_6417,N_7537);
nor U9580 (N_9580,N_6471,N_7772);
and U9581 (N_9581,N_7258,N_6887);
nand U9582 (N_9582,N_7971,N_7574);
and U9583 (N_9583,N_6740,N_6116);
and U9584 (N_9584,N_6738,N_6955);
nor U9585 (N_9585,N_7316,N_7157);
and U9586 (N_9586,N_6618,N_6146);
or U9587 (N_9587,N_7766,N_7202);
or U9588 (N_9588,N_6173,N_6597);
nand U9589 (N_9589,N_7158,N_6299);
nor U9590 (N_9590,N_7012,N_7690);
or U9591 (N_9591,N_6020,N_6133);
and U9592 (N_9592,N_7804,N_6700);
nor U9593 (N_9593,N_7837,N_7782);
and U9594 (N_9594,N_7323,N_7780);
or U9595 (N_9595,N_7674,N_7497);
or U9596 (N_9596,N_7316,N_6366);
nor U9597 (N_9597,N_6945,N_6356);
and U9598 (N_9598,N_7564,N_7857);
or U9599 (N_9599,N_6181,N_6284);
nor U9600 (N_9600,N_6626,N_7354);
and U9601 (N_9601,N_7597,N_7019);
or U9602 (N_9602,N_7418,N_7521);
or U9603 (N_9603,N_6583,N_7280);
and U9604 (N_9604,N_7706,N_6197);
and U9605 (N_9605,N_7949,N_6967);
nor U9606 (N_9606,N_6755,N_6665);
and U9607 (N_9607,N_7118,N_6443);
or U9608 (N_9608,N_7688,N_7572);
or U9609 (N_9609,N_6132,N_7379);
or U9610 (N_9610,N_6867,N_6651);
and U9611 (N_9611,N_6596,N_7720);
and U9612 (N_9612,N_6727,N_7488);
and U9613 (N_9613,N_6353,N_6276);
nor U9614 (N_9614,N_7699,N_6953);
xor U9615 (N_9615,N_7224,N_6437);
nand U9616 (N_9616,N_7739,N_6203);
and U9617 (N_9617,N_6340,N_6199);
nor U9618 (N_9618,N_7768,N_7597);
nor U9619 (N_9619,N_7295,N_7792);
nand U9620 (N_9620,N_7283,N_7089);
or U9621 (N_9621,N_7999,N_7160);
nand U9622 (N_9622,N_6804,N_6977);
and U9623 (N_9623,N_7430,N_6097);
nand U9624 (N_9624,N_6075,N_7486);
and U9625 (N_9625,N_6901,N_7629);
nor U9626 (N_9626,N_6733,N_6239);
xnor U9627 (N_9627,N_6186,N_7218);
and U9628 (N_9628,N_6280,N_6818);
and U9629 (N_9629,N_6868,N_7011);
nor U9630 (N_9630,N_6366,N_6522);
or U9631 (N_9631,N_6336,N_6895);
or U9632 (N_9632,N_7669,N_7726);
xor U9633 (N_9633,N_6822,N_6380);
and U9634 (N_9634,N_6225,N_6362);
nand U9635 (N_9635,N_6452,N_7881);
nand U9636 (N_9636,N_6902,N_6233);
and U9637 (N_9637,N_7490,N_7021);
or U9638 (N_9638,N_6352,N_7502);
and U9639 (N_9639,N_7442,N_7631);
and U9640 (N_9640,N_7434,N_7095);
and U9641 (N_9641,N_7166,N_6965);
or U9642 (N_9642,N_6721,N_6256);
and U9643 (N_9643,N_7305,N_6458);
nand U9644 (N_9644,N_7958,N_7648);
nand U9645 (N_9645,N_6540,N_6472);
nand U9646 (N_9646,N_7603,N_6461);
and U9647 (N_9647,N_7822,N_6546);
and U9648 (N_9648,N_7564,N_6186);
and U9649 (N_9649,N_7346,N_7478);
and U9650 (N_9650,N_6389,N_7347);
and U9651 (N_9651,N_7163,N_7986);
and U9652 (N_9652,N_6847,N_6876);
or U9653 (N_9653,N_6088,N_6470);
or U9654 (N_9654,N_7326,N_6949);
and U9655 (N_9655,N_7576,N_7324);
nor U9656 (N_9656,N_7518,N_6371);
and U9657 (N_9657,N_7299,N_7107);
nor U9658 (N_9658,N_7428,N_7844);
nor U9659 (N_9659,N_6009,N_6651);
nand U9660 (N_9660,N_7699,N_7116);
xor U9661 (N_9661,N_7846,N_6050);
and U9662 (N_9662,N_7861,N_7907);
or U9663 (N_9663,N_7623,N_7091);
or U9664 (N_9664,N_6844,N_7018);
nor U9665 (N_9665,N_7368,N_7045);
nand U9666 (N_9666,N_6733,N_6497);
nor U9667 (N_9667,N_6722,N_7799);
nand U9668 (N_9668,N_7544,N_6259);
and U9669 (N_9669,N_7248,N_7931);
and U9670 (N_9670,N_6934,N_7675);
or U9671 (N_9671,N_7901,N_7448);
nand U9672 (N_9672,N_7516,N_6770);
or U9673 (N_9673,N_7926,N_7241);
nor U9674 (N_9674,N_6204,N_6399);
nand U9675 (N_9675,N_6544,N_7118);
or U9676 (N_9676,N_6010,N_6946);
nor U9677 (N_9677,N_6031,N_6162);
nand U9678 (N_9678,N_6244,N_7832);
nor U9679 (N_9679,N_6073,N_7328);
or U9680 (N_9680,N_7242,N_7338);
nand U9681 (N_9681,N_6133,N_6444);
and U9682 (N_9682,N_6524,N_7030);
nand U9683 (N_9683,N_7190,N_7260);
and U9684 (N_9684,N_6931,N_7479);
or U9685 (N_9685,N_7978,N_6084);
and U9686 (N_9686,N_6710,N_6164);
nor U9687 (N_9687,N_6000,N_7907);
nand U9688 (N_9688,N_7486,N_7357);
nor U9689 (N_9689,N_6314,N_7548);
and U9690 (N_9690,N_7879,N_7279);
nor U9691 (N_9691,N_6743,N_7560);
nor U9692 (N_9692,N_7902,N_7195);
nand U9693 (N_9693,N_7969,N_7977);
or U9694 (N_9694,N_7489,N_7803);
or U9695 (N_9695,N_7734,N_6792);
and U9696 (N_9696,N_7370,N_6716);
nor U9697 (N_9697,N_7701,N_6583);
nor U9698 (N_9698,N_7875,N_6530);
nand U9699 (N_9699,N_7944,N_6730);
or U9700 (N_9700,N_7218,N_6525);
nand U9701 (N_9701,N_7817,N_6198);
and U9702 (N_9702,N_7972,N_6058);
nand U9703 (N_9703,N_7576,N_6175);
nand U9704 (N_9704,N_6348,N_6909);
nand U9705 (N_9705,N_6280,N_6061);
and U9706 (N_9706,N_6288,N_7480);
nor U9707 (N_9707,N_7966,N_6590);
nand U9708 (N_9708,N_6164,N_6292);
and U9709 (N_9709,N_7066,N_7853);
nor U9710 (N_9710,N_7918,N_6670);
nor U9711 (N_9711,N_6438,N_7607);
or U9712 (N_9712,N_6863,N_6114);
nand U9713 (N_9713,N_6191,N_7855);
and U9714 (N_9714,N_7702,N_6575);
xor U9715 (N_9715,N_7338,N_7468);
nand U9716 (N_9716,N_7835,N_7376);
nand U9717 (N_9717,N_7392,N_6784);
nor U9718 (N_9718,N_7357,N_7308);
and U9719 (N_9719,N_7588,N_6607);
nand U9720 (N_9720,N_7093,N_7842);
nor U9721 (N_9721,N_7029,N_6495);
and U9722 (N_9722,N_6239,N_7084);
nand U9723 (N_9723,N_6846,N_7730);
nand U9724 (N_9724,N_6632,N_7169);
or U9725 (N_9725,N_6817,N_7369);
nand U9726 (N_9726,N_7833,N_6367);
or U9727 (N_9727,N_6194,N_6067);
nand U9728 (N_9728,N_7293,N_7687);
nor U9729 (N_9729,N_6033,N_6947);
or U9730 (N_9730,N_7108,N_6720);
nor U9731 (N_9731,N_7034,N_6729);
nand U9732 (N_9732,N_7067,N_6121);
or U9733 (N_9733,N_6192,N_6590);
and U9734 (N_9734,N_6961,N_7653);
nand U9735 (N_9735,N_6185,N_6181);
nand U9736 (N_9736,N_6819,N_6917);
nor U9737 (N_9737,N_7253,N_7035);
nand U9738 (N_9738,N_7123,N_6863);
nand U9739 (N_9739,N_7345,N_7231);
and U9740 (N_9740,N_7469,N_6234);
and U9741 (N_9741,N_7167,N_7848);
nand U9742 (N_9742,N_6680,N_7495);
nor U9743 (N_9743,N_7666,N_6524);
nand U9744 (N_9744,N_6508,N_6353);
nand U9745 (N_9745,N_7434,N_6103);
nand U9746 (N_9746,N_6702,N_7976);
nor U9747 (N_9747,N_6821,N_7142);
or U9748 (N_9748,N_7726,N_7121);
xor U9749 (N_9749,N_6062,N_7411);
nor U9750 (N_9750,N_7673,N_6811);
or U9751 (N_9751,N_6500,N_7196);
nand U9752 (N_9752,N_6311,N_6297);
nor U9753 (N_9753,N_7893,N_6276);
nor U9754 (N_9754,N_7884,N_7756);
or U9755 (N_9755,N_6638,N_7755);
nor U9756 (N_9756,N_6333,N_6260);
nand U9757 (N_9757,N_6007,N_7469);
nand U9758 (N_9758,N_7360,N_6302);
nor U9759 (N_9759,N_7777,N_6725);
nor U9760 (N_9760,N_6019,N_7860);
and U9761 (N_9761,N_6915,N_6918);
and U9762 (N_9762,N_6679,N_7546);
nor U9763 (N_9763,N_6374,N_6603);
and U9764 (N_9764,N_7908,N_6293);
nand U9765 (N_9765,N_6038,N_7718);
and U9766 (N_9766,N_7106,N_6353);
and U9767 (N_9767,N_6359,N_6829);
or U9768 (N_9768,N_7792,N_7868);
nor U9769 (N_9769,N_7995,N_7460);
nand U9770 (N_9770,N_7850,N_7665);
and U9771 (N_9771,N_6379,N_7977);
nand U9772 (N_9772,N_7118,N_6974);
nand U9773 (N_9773,N_7436,N_7118);
nand U9774 (N_9774,N_7262,N_7880);
or U9775 (N_9775,N_6587,N_6958);
nor U9776 (N_9776,N_7619,N_7630);
and U9777 (N_9777,N_7150,N_6517);
nor U9778 (N_9778,N_6802,N_6259);
and U9779 (N_9779,N_7496,N_7704);
nor U9780 (N_9780,N_6632,N_6631);
nand U9781 (N_9781,N_7297,N_7599);
nor U9782 (N_9782,N_7434,N_7175);
nor U9783 (N_9783,N_7897,N_6674);
nor U9784 (N_9784,N_7061,N_6153);
nor U9785 (N_9785,N_6420,N_7728);
and U9786 (N_9786,N_7308,N_7613);
nor U9787 (N_9787,N_7038,N_6781);
nand U9788 (N_9788,N_7120,N_6715);
nor U9789 (N_9789,N_7348,N_7835);
and U9790 (N_9790,N_6669,N_7226);
nor U9791 (N_9791,N_6449,N_7725);
or U9792 (N_9792,N_6912,N_7168);
and U9793 (N_9793,N_6407,N_6838);
or U9794 (N_9794,N_6374,N_6869);
nand U9795 (N_9795,N_6261,N_6408);
or U9796 (N_9796,N_6299,N_6420);
or U9797 (N_9797,N_6437,N_6323);
nand U9798 (N_9798,N_7600,N_7782);
nand U9799 (N_9799,N_6979,N_6620);
nand U9800 (N_9800,N_6446,N_7313);
nor U9801 (N_9801,N_7390,N_7342);
or U9802 (N_9802,N_7124,N_7725);
nand U9803 (N_9803,N_6436,N_6873);
nand U9804 (N_9804,N_6982,N_6801);
and U9805 (N_9805,N_6730,N_7690);
nand U9806 (N_9806,N_6843,N_6373);
and U9807 (N_9807,N_6697,N_6014);
nor U9808 (N_9808,N_6253,N_6423);
and U9809 (N_9809,N_6015,N_6865);
nor U9810 (N_9810,N_7705,N_6746);
nand U9811 (N_9811,N_6643,N_7090);
and U9812 (N_9812,N_6666,N_6716);
and U9813 (N_9813,N_6155,N_7413);
or U9814 (N_9814,N_7924,N_7153);
and U9815 (N_9815,N_7114,N_6407);
and U9816 (N_9816,N_6975,N_6296);
nor U9817 (N_9817,N_7246,N_7680);
nor U9818 (N_9818,N_6873,N_7745);
and U9819 (N_9819,N_6294,N_7727);
nand U9820 (N_9820,N_7344,N_6704);
nor U9821 (N_9821,N_6261,N_6452);
and U9822 (N_9822,N_7605,N_7804);
or U9823 (N_9823,N_7093,N_7086);
and U9824 (N_9824,N_7097,N_6222);
and U9825 (N_9825,N_7207,N_7856);
and U9826 (N_9826,N_6806,N_6860);
nand U9827 (N_9827,N_6141,N_6246);
and U9828 (N_9828,N_7269,N_6103);
and U9829 (N_9829,N_6199,N_7290);
nand U9830 (N_9830,N_7510,N_7860);
or U9831 (N_9831,N_6543,N_6821);
nor U9832 (N_9832,N_7056,N_7093);
nor U9833 (N_9833,N_6633,N_7783);
or U9834 (N_9834,N_6902,N_7298);
or U9835 (N_9835,N_6268,N_7817);
nor U9836 (N_9836,N_7825,N_7905);
nor U9837 (N_9837,N_6800,N_7273);
or U9838 (N_9838,N_6207,N_7056);
and U9839 (N_9839,N_6325,N_6520);
and U9840 (N_9840,N_7289,N_6584);
nor U9841 (N_9841,N_6206,N_7731);
nand U9842 (N_9842,N_7997,N_6652);
or U9843 (N_9843,N_6089,N_6824);
nor U9844 (N_9844,N_6012,N_7987);
nor U9845 (N_9845,N_7877,N_6010);
or U9846 (N_9846,N_6320,N_7959);
or U9847 (N_9847,N_6502,N_7417);
or U9848 (N_9848,N_6359,N_6930);
or U9849 (N_9849,N_7183,N_6957);
nor U9850 (N_9850,N_6231,N_6431);
nand U9851 (N_9851,N_7543,N_6592);
nand U9852 (N_9852,N_7954,N_7613);
nand U9853 (N_9853,N_6667,N_6108);
and U9854 (N_9854,N_6360,N_6410);
nand U9855 (N_9855,N_7272,N_6747);
and U9856 (N_9856,N_6325,N_6611);
nand U9857 (N_9857,N_6349,N_7936);
nor U9858 (N_9858,N_6591,N_7427);
nor U9859 (N_9859,N_7783,N_6835);
nor U9860 (N_9860,N_7583,N_7611);
nand U9861 (N_9861,N_6648,N_6597);
nand U9862 (N_9862,N_7639,N_7320);
nand U9863 (N_9863,N_7178,N_6739);
or U9864 (N_9864,N_7686,N_6095);
and U9865 (N_9865,N_6837,N_7628);
and U9866 (N_9866,N_6978,N_7624);
xor U9867 (N_9867,N_7072,N_6272);
or U9868 (N_9868,N_6545,N_6362);
nor U9869 (N_9869,N_7053,N_7635);
nor U9870 (N_9870,N_7771,N_6888);
and U9871 (N_9871,N_6140,N_7700);
or U9872 (N_9872,N_6102,N_6150);
nand U9873 (N_9873,N_6790,N_7121);
nand U9874 (N_9874,N_7134,N_7019);
and U9875 (N_9875,N_6050,N_6200);
nor U9876 (N_9876,N_6591,N_7459);
nor U9877 (N_9877,N_7486,N_6154);
and U9878 (N_9878,N_7600,N_7346);
nand U9879 (N_9879,N_6726,N_7057);
or U9880 (N_9880,N_7655,N_6116);
nand U9881 (N_9881,N_7419,N_7220);
and U9882 (N_9882,N_7509,N_7882);
or U9883 (N_9883,N_6530,N_6402);
nor U9884 (N_9884,N_7882,N_7983);
nor U9885 (N_9885,N_7507,N_7001);
nor U9886 (N_9886,N_7297,N_6036);
and U9887 (N_9887,N_6087,N_7067);
or U9888 (N_9888,N_7629,N_6335);
and U9889 (N_9889,N_6547,N_7991);
and U9890 (N_9890,N_6153,N_7780);
and U9891 (N_9891,N_7809,N_6537);
or U9892 (N_9892,N_7859,N_6587);
nor U9893 (N_9893,N_6592,N_6422);
nand U9894 (N_9894,N_7060,N_7320);
nand U9895 (N_9895,N_6008,N_7518);
nor U9896 (N_9896,N_6723,N_6374);
and U9897 (N_9897,N_6381,N_6557);
nand U9898 (N_9898,N_7426,N_7506);
or U9899 (N_9899,N_6614,N_7354);
nand U9900 (N_9900,N_6941,N_7532);
and U9901 (N_9901,N_6816,N_6247);
nand U9902 (N_9902,N_6973,N_7794);
and U9903 (N_9903,N_7800,N_6241);
or U9904 (N_9904,N_6578,N_7253);
or U9905 (N_9905,N_6717,N_7453);
nor U9906 (N_9906,N_7377,N_6197);
and U9907 (N_9907,N_7794,N_6012);
and U9908 (N_9908,N_7011,N_6953);
nor U9909 (N_9909,N_6139,N_7034);
or U9910 (N_9910,N_6806,N_6770);
nand U9911 (N_9911,N_6957,N_6656);
nand U9912 (N_9912,N_6561,N_6478);
nand U9913 (N_9913,N_7934,N_6018);
or U9914 (N_9914,N_7101,N_7994);
nand U9915 (N_9915,N_6359,N_7928);
or U9916 (N_9916,N_6333,N_6418);
and U9917 (N_9917,N_6813,N_7024);
nor U9918 (N_9918,N_7939,N_7625);
and U9919 (N_9919,N_6315,N_7613);
nand U9920 (N_9920,N_6899,N_7801);
or U9921 (N_9921,N_7490,N_7969);
or U9922 (N_9922,N_7446,N_7428);
or U9923 (N_9923,N_7598,N_7344);
nand U9924 (N_9924,N_6510,N_7702);
nor U9925 (N_9925,N_6474,N_7772);
and U9926 (N_9926,N_7715,N_7264);
nand U9927 (N_9927,N_6566,N_6812);
and U9928 (N_9928,N_7830,N_7848);
xor U9929 (N_9929,N_7764,N_7803);
or U9930 (N_9930,N_6911,N_6296);
nor U9931 (N_9931,N_7465,N_6210);
nand U9932 (N_9932,N_6935,N_6548);
nor U9933 (N_9933,N_6860,N_6193);
or U9934 (N_9934,N_6269,N_7655);
nand U9935 (N_9935,N_6367,N_7539);
nand U9936 (N_9936,N_6633,N_6954);
nor U9937 (N_9937,N_6111,N_6479);
nor U9938 (N_9938,N_6640,N_7199);
nand U9939 (N_9939,N_6478,N_6727);
nand U9940 (N_9940,N_6317,N_6024);
nand U9941 (N_9941,N_7849,N_6790);
or U9942 (N_9942,N_6174,N_7997);
and U9943 (N_9943,N_6263,N_7546);
nor U9944 (N_9944,N_7398,N_7620);
nand U9945 (N_9945,N_6032,N_7632);
nand U9946 (N_9946,N_6685,N_7997);
and U9947 (N_9947,N_7220,N_7992);
and U9948 (N_9948,N_6944,N_7644);
nand U9949 (N_9949,N_7188,N_7172);
nor U9950 (N_9950,N_7526,N_6412);
nor U9951 (N_9951,N_6730,N_6100);
nand U9952 (N_9952,N_7582,N_6590);
and U9953 (N_9953,N_6380,N_6409);
nor U9954 (N_9954,N_6709,N_7521);
nor U9955 (N_9955,N_7546,N_7772);
or U9956 (N_9956,N_7485,N_7895);
and U9957 (N_9957,N_6395,N_6857);
nor U9958 (N_9958,N_7660,N_6349);
and U9959 (N_9959,N_6876,N_7912);
or U9960 (N_9960,N_6151,N_6823);
or U9961 (N_9961,N_6943,N_6427);
nand U9962 (N_9962,N_6991,N_6649);
or U9963 (N_9963,N_6479,N_6664);
and U9964 (N_9964,N_7731,N_7824);
or U9965 (N_9965,N_7204,N_7785);
and U9966 (N_9966,N_6957,N_6303);
nor U9967 (N_9967,N_7370,N_6659);
and U9968 (N_9968,N_6625,N_7351);
nor U9969 (N_9969,N_7360,N_6421);
nand U9970 (N_9970,N_6259,N_7510);
or U9971 (N_9971,N_7266,N_7892);
nand U9972 (N_9972,N_7992,N_6803);
and U9973 (N_9973,N_6389,N_6619);
or U9974 (N_9974,N_6880,N_6767);
nand U9975 (N_9975,N_7328,N_7536);
nand U9976 (N_9976,N_7863,N_7702);
or U9977 (N_9977,N_6523,N_7830);
and U9978 (N_9978,N_7363,N_6616);
and U9979 (N_9979,N_6088,N_6199);
and U9980 (N_9980,N_7735,N_6803);
nor U9981 (N_9981,N_7918,N_7495);
nand U9982 (N_9982,N_7460,N_6844);
or U9983 (N_9983,N_7287,N_6839);
nand U9984 (N_9984,N_6041,N_6363);
and U9985 (N_9985,N_6463,N_6723);
nor U9986 (N_9986,N_6252,N_7696);
and U9987 (N_9987,N_6477,N_6081);
nand U9988 (N_9988,N_6660,N_7625);
or U9989 (N_9989,N_7609,N_6927);
or U9990 (N_9990,N_7479,N_7246);
or U9991 (N_9991,N_6727,N_6209);
nand U9992 (N_9992,N_6119,N_6088);
nor U9993 (N_9993,N_6633,N_7808);
nor U9994 (N_9994,N_6400,N_6764);
or U9995 (N_9995,N_6161,N_7619);
and U9996 (N_9996,N_7047,N_7797);
and U9997 (N_9997,N_7742,N_7277);
and U9998 (N_9998,N_6700,N_7611);
nand U9999 (N_9999,N_6485,N_6938);
or UO_0 (O_0,N_8996,N_8581);
nand UO_1 (O_1,N_8349,N_9261);
or UO_2 (O_2,N_9058,N_9866);
xor UO_3 (O_3,N_8547,N_9322);
nor UO_4 (O_4,N_9264,N_8337);
or UO_5 (O_5,N_9103,N_9265);
or UO_6 (O_6,N_9359,N_8392);
nand UO_7 (O_7,N_8338,N_8640);
nand UO_8 (O_8,N_8666,N_9581);
nor UO_9 (O_9,N_9721,N_9541);
and UO_10 (O_10,N_9251,N_8642);
nand UO_11 (O_11,N_9670,N_8423);
or UO_12 (O_12,N_8010,N_9075);
or UO_13 (O_13,N_8638,N_9214);
nand UO_14 (O_14,N_8112,N_8750);
nor UO_15 (O_15,N_9512,N_9782);
and UO_16 (O_16,N_9767,N_9733);
or UO_17 (O_17,N_8936,N_9196);
nand UO_18 (O_18,N_9057,N_9718);
nor UO_19 (O_19,N_8465,N_9814);
nor UO_20 (O_20,N_8830,N_9337);
or UO_21 (O_21,N_9557,N_8751);
nor UO_22 (O_22,N_9854,N_8565);
nand UO_23 (O_23,N_9491,N_9786);
nand UO_24 (O_24,N_8851,N_9945);
and UO_25 (O_25,N_8167,N_8102);
nand UO_26 (O_26,N_9259,N_8314);
nand UO_27 (O_27,N_8671,N_8635);
or UO_28 (O_28,N_9112,N_9817);
nand UO_29 (O_29,N_8089,N_8842);
xnor UO_30 (O_30,N_8364,N_8162);
or UO_31 (O_31,N_8962,N_8829);
nand UO_32 (O_32,N_8561,N_8676);
and UO_33 (O_33,N_9100,N_8446);
nor UO_34 (O_34,N_9440,N_9929);
and UO_35 (O_35,N_9883,N_9566);
nor UO_36 (O_36,N_9136,N_8807);
nand UO_37 (O_37,N_8459,N_9799);
nand UO_38 (O_38,N_9098,N_8692);
nor UO_39 (O_39,N_9620,N_8563);
or UO_40 (O_40,N_9878,N_8186);
nand UO_41 (O_41,N_8616,N_8659);
nand UO_42 (O_42,N_8513,N_9138);
nand UO_43 (O_43,N_9730,N_8536);
and UO_44 (O_44,N_9683,N_9912);
and UO_45 (O_45,N_9589,N_9231);
nand UO_46 (O_46,N_9971,N_9630);
nand UO_47 (O_47,N_9082,N_9919);
or UO_48 (O_48,N_9710,N_9356);
nand UO_49 (O_49,N_8597,N_9188);
and UO_50 (O_50,N_9821,N_8199);
or UO_51 (O_51,N_8460,N_9219);
or UO_52 (O_52,N_9524,N_8366);
nor UO_53 (O_53,N_9225,N_9441);
nor UO_54 (O_54,N_8045,N_9542);
or UO_55 (O_55,N_9385,N_9033);
nand UO_56 (O_56,N_8703,N_9508);
and UO_57 (O_57,N_9378,N_9333);
and UO_58 (O_58,N_8971,N_9619);
and UO_59 (O_59,N_9494,N_8852);
nor UO_60 (O_60,N_8189,N_9975);
or UO_61 (O_61,N_8206,N_9626);
and UO_62 (O_62,N_9108,N_9160);
and UO_63 (O_63,N_8694,N_9607);
nand UO_64 (O_64,N_8663,N_8400);
or UO_65 (O_65,N_9092,N_9806);
and UO_66 (O_66,N_8789,N_9674);
nor UO_67 (O_67,N_8797,N_8422);
or UO_68 (O_68,N_9200,N_8428);
nor UO_69 (O_69,N_8307,N_8450);
nand UO_70 (O_70,N_8557,N_8974);
or UO_71 (O_71,N_8231,N_8661);
nor UO_72 (O_72,N_9977,N_9723);
nand UO_73 (O_73,N_9563,N_9282);
nand UO_74 (O_74,N_8504,N_9064);
nor UO_75 (O_75,N_9744,N_8600);
nor UO_76 (O_76,N_8135,N_8864);
nor UO_77 (O_77,N_8887,N_8488);
nand UO_78 (O_78,N_8124,N_9640);
and UO_79 (O_79,N_8689,N_9102);
nor UO_80 (O_80,N_9737,N_8788);
xnor UO_81 (O_81,N_9292,N_9882);
and UO_82 (O_82,N_8628,N_9164);
nand UO_83 (O_83,N_9686,N_9353);
or UO_84 (O_84,N_9689,N_8246);
nor UO_85 (O_85,N_9756,N_9496);
nand UO_86 (O_86,N_9849,N_8986);
nor UO_87 (O_87,N_8786,N_9157);
or UO_88 (O_88,N_9437,N_9382);
xor UO_89 (O_89,N_8675,N_9435);
or UO_90 (O_90,N_8437,N_8526);
or UO_91 (O_91,N_9871,N_8662);
nor UO_92 (O_92,N_9379,N_8012);
and UO_93 (O_93,N_9747,N_8335);
nor UO_94 (O_94,N_8092,N_8716);
nand UO_95 (O_95,N_9964,N_8497);
nand UO_96 (O_96,N_9933,N_8906);
or UO_97 (O_97,N_8781,N_8458);
and UO_98 (O_98,N_9503,N_8668);
and UO_99 (O_99,N_9816,N_9019);
nand UO_100 (O_100,N_9600,N_9249);
and UO_101 (O_101,N_9865,N_8311);
nor UO_102 (O_102,N_8858,N_8268);
and UO_103 (O_103,N_9227,N_9997);
and UO_104 (O_104,N_8782,N_9071);
nand UO_105 (O_105,N_9008,N_8795);
nand UO_106 (O_106,N_8179,N_9067);
nor UO_107 (O_107,N_9675,N_9995);
and UO_108 (O_108,N_9586,N_9388);
and UO_109 (O_109,N_8910,N_8806);
nand UO_110 (O_110,N_9065,N_9545);
nand UO_111 (O_111,N_9870,N_8129);
nor UO_112 (O_112,N_8274,N_9603);
or UO_113 (O_113,N_9109,N_8696);
or UO_114 (O_114,N_8753,N_8241);
nor UO_115 (O_115,N_8578,N_9362);
or UO_116 (O_116,N_8277,N_9829);
nand UO_117 (O_117,N_8941,N_9484);
nor UO_118 (O_118,N_9089,N_8273);
and UO_119 (O_119,N_9860,N_9266);
and UO_120 (O_120,N_9434,N_9281);
or UO_121 (O_121,N_9988,N_8104);
nand UO_122 (O_122,N_8072,N_8327);
or UO_123 (O_123,N_9198,N_9384);
nand UO_124 (O_124,N_8907,N_8850);
nand UO_125 (O_125,N_9592,N_8454);
nor UO_126 (O_126,N_8982,N_9775);
or UO_127 (O_127,N_9624,N_8903);
or UO_128 (O_128,N_8574,N_8918);
nor UO_129 (O_129,N_8677,N_9344);
nor UO_130 (O_130,N_8679,N_9587);
nand UO_131 (O_131,N_8521,N_9294);
nand UO_132 (O_132,N_8049,N_9915);
nand UO_133 (O_133,N_9241,N_9408);
nor UO_134 (O_134,N_8190,N_9203);
nand UO_135 (O_135,N_8059,N_9880);
nor UO_136 (O_136,N_9147,N_9955);
and UO_137 (O_137,N_8947,N_8391);
nor UO_138 (O_138,N_8594,N_8888);
nand UO_139 (O_139,N_9633,N_8007);
or UO_140 (O_140,N_8163,N_9646);
nand UO_141 (O_141,N_9239,N_8954);
nor UO_142 (O_142,N_8582,N_8406);
and UO_143 (O_143,N_9725,N_9952);
nor UO_144 (O_144,N_8834,N_9923);
or UO_145 (O_145,N_8761,N_9951);
nand UO_146 (O_146,N_8394,N_9698);
nand UO_147 (O_147,N_9778,N_9088);
nor UO_148 (O_148,N_9968,N_8260);
nand UO_149 (O_149,N_8644,N_9820);
nor UO_150 (O_150,N_9431,N_8515);
nor UO_151 (O_151,N_8719,N_9490);
and UO_152 (O_152,N_9208,N_8576);
or UO_153 (O_153,N_9146,N_8375);
or UO_154 (O_154,N_9350,N_8478);
and UO_155 (O_155,N_8434,N_8025);
and UO_156 (O_156,N_9343,N_8047);
and UO_157 (O_157,N_8331,N_8997);
nor UO_158 (O_158,N_9234,N_8549);
nand UO_159 (O_159,N_9326,N_8849);
or UO_160 (O_160,N_8461,N_9787);
or UO_161 (O_161,N_9256,N_9529);
or UO_162 (O_162,N_8258,N_8057);
nor UO_163 (O_163,N_8343,N_9514);
nand UO_164 (O_164,N_9391,N_9580);
and UO_165 (O_165,N_8425,N_9414);
nand UO_166 (O_166,N_8038,N_8382);
and UO_167 (O_167,N_9156,N_9528);
nand UO_168 (O_168,N_9453,N_8747);
nor UO_169 (O_169,N_8736,N_9792);
nand UO_170 (O_170,N_8933,N_9447);
or UO_171 (O_171,N_8944,N_9218);
nor UO_172 (O_172,N_8820,N_9038);
or UO_173 (O_173,N_8207,N_9117);
nand UO_174 (O_174,N_9360,N_9056);
or UO_175 (O_175,N_8840,N_8681);
and UO_176 (O_176,N_8360,N_9332);
and UO_177 (O_177,N_8397,N_9536);
and UO_178 (O_178,N_9780,N_9789);
nand UO_179 (O_179,N_8950,N_8605);
nand UO_180 (O_180,N_9277,N_9895);
and UO_181 (O_181,N_8188,N_8160);
and UO_182 (O_182,N_9896,N_8291);
and UO_183 (O_183,N_9983,N_9304);
nor UO_184 (O_184,N_9315,N_9931);
nand UO_185 (O_185,N_9258,N_9825);
and UO_186 (O_186,N_8253,N_8093);
nor UO_187 (O_187,N_8552,N_8953);
nand UO_188 (O_188,N_9495,N_8281);
and UO_189 (O_189,N_9847,N_9111);
or UO_190 (O_190,N_8749,N_8094);
nand UO_191 (O_191,N_8617,N_9090);
or UO_192 (O_192,N_9819,N_8921);
nor UO_193 (O_193,N_9921,N_8882);
and UO_194 (O_194,N_8440,N_9749);
or UO_195 (O_195,N_9289,N_8499);
nor UO_196 (O_196,N_9396,N_8211);
or UO_197 (O_197,N_8344,N_9776);
or UO_198 (O_198,N_9811,N_9436);
nor UO_199 (O_199,N_9760,N_8546);
and UO_200 (O_200,N_9472,N_8618);
or UO_201 (O_201,N_8278,N_9300);
nor UO_202 (O_202,N_8376,N_9504);
nand UO_203 (O_203,N_8090,N_9096);
or UO_204 (O_204,N_9593,N_8218);
nand UO_205 (O_205,N_9175,N_8005);
and UO_206 (O_206,N_8031,N_9573);
nor UO_207 (O_207,N_8035,N_9734);
and UO_208 (O_208,N_9290,N_9761);
and UO_209 (O_209,N_9009,N_8388);
nor UO_210 (O_210,N_9910,N_9901);
nand UO_211 (O_211,N_8336,N_9695);
nor UO_212 (O_212,N_9942,N_9837);
or UO_213 (O_213,N_9086,N_8509);
or UO_214 (O_214,N_8091,N_9052);
nor UO_215 (O_215,N_8949,N_9370);
nand UO_216 (O_216,N_8200,N_8027);
nand UO_217 (O_217,N_9855,N_9069);
or UO_218 (O_218,N_8774,N_9862);
nand UO_219 (O_219,N_9363,N_8303);
nand UO_220 (O_220,N_9576,N_8627);
xnor UO_221 (O_221,N_8988,N_8995);
or UO_222 (O_222,N_8229,N_9470);
and UO_223 (O_223,N_9331,N_8152);
or UO_224 (O_224,N_9002,N_9874);
and UO_225 (O_225,N_8529,N_9739);
and UO_226 (O_226,N_8474,N_9766);
nand UO_227 (O_227,N_9115,N_9110);
or UO_228 (O_228,N_9349,N_8649);
nand UO_229 (O_229,N_8491,N_8288);
nor UO_230 (O_230,N_8224,N_9890);
xor UO_231 (O_231,N_9308,N_8014);
nor UO_232 (O_232,N_9313,N_8340);
and UO_233 (O_233,N_8151,N_8734);
or UO_234 (O_234,N_8203,N_8646);
or UO_235 (O_235,N_8743,N_8214);
nor UO_236 (O_236,N_8046,N_8026);
nor UO_237 (O_237,N_9003,N_8911);
nor UO_238 (O_238,N_9368,N_8776);
nor UO_239 (O_239,N_8855,N_8523);
or UO_240 (O_240,N_9533,N_9544);
xor UO_241 (O_241,N_8016,N_8081);
nor UO_242 (O_242,N_8353,N_8379);
nor UO_243 (O_243,N_8613,N_8656);
nor UO_244 (O_244,N_9455,N_8481);
nand UO_245 (O_245,N_8191,N_9918);
and UO_246 (O_246,N_8687,N_8300);
and UO_247 (O_247,N_8096,N_9822);
and UO_248 (O_248,N_8518,N_9812);
nor UO_249 (O_249,N_8873,N_8466);
nor UO_250 (O_250,N_9850,N_9482);
or UO_251 (O_251,N_8276,N_9417);
nand UO_252 (O_252,N_8725,N_8126);
and UO_253 (O_253,N_8609,N_8069);
nand UO_254 (O_254,N_9255,N_9220);
or UO_255 (O_255,N_9891,N_9232);
nand UO_256 (O_256,N_8589,N_9583);
and UO_257 (O_257,N_8181,N_9209);
nor UO_258 (O_258,N_9978,N_9719);
and UO_259 (O_259,N_8136,N_8505);
nor UO_260 (O_260,N_8614,N_8028);
nor UO_261 (O_261,N_9848,N_8899);
nor UO_262 (O_262,N_9041,N_9663);
nor UO_263 (O_263,N_9608,N_8972);
nor UO_264 (O_264,N_8295,N_8674);
nor UO_265 (O_265,N_8170,N_9014);
or UO_266 (O_266,N_9622,N_8139);
nor UO_267 (O_267,N_9247,N_9920);
and UO_268 (O_268,N_9894,N_9692);
or UO_269 (O_269,N_8752,N_9170);
nor UO_270 (O_270,N_8402,N_8275);
nand UO_271 (O_271,N_8943,N_8922);
and UO_272 (O_272,N_9042,N_8871);
or UO_273 (O_273,N_8817,N_8886);
nor UO_274 (O_274,N_8150,N_9423);
nor UO_275 (O_275,N_8821,N_8877);
and UO_276 (O_276,N_9355,N_9969);
or UO_277 (O_277,N_8371,N_8990);
nor UO_278 (O_278,N_8109,N_8097);
nor UO_279 (O_279,N_9764,N_8545);
and UO_280 (O_280,N_8583,N_9714);
or UO_281 (O_281,N_8452,N_8427);
or UO_282 (O_282,N_8495,N_9571);
nand UO_283 (O_283,N_8044,N_9158);
or UO_284 (O_284,N_8639,N_8631);
and UO_285 (O_285,N_9937,N_8965);
nand UO_286 (O_286,N_8413,N_8236);
nor UO_287 (O_287,N_9167,N_9818);
nand UO_288 (O_288,N_9401,N_9779);
xnor UO_289 (O_289,N_9452,N_8937);
and UO_290 (O_290,N_9206,N_8836);
or UO_291 (O_291,N_8060,N_8926);
nor UO_292 (O_292,N_9987,N_8118);
nand UO_293 (O_293,N_8946,N_8658);
or UO_294 (O_294,N_8204,N_9048);
and UO_295 (O_295,N_8739,N_8527);
nor UO_296 (O_296,N_8634,N_8122);
nand UO_297 (O_297,N_9742,N_8680);
and UO_298 (O_298,N_9924,N_8449);
nor UO_299 (O_299,N_8368,N_8257);
nor UO_300 (O_300,N_9960,N_8977);
nand UO_301 (O_301,N_9123,N_9476);
nand UO_302 (O_302,N_8810,N_9879);
nand UO_303 (O_303,N_8370,N_9549);
nor UO_304 (O_304,N_8664,N_9715);
or UO_305 (O_305,N_8232,N_9420);
nand UO_306 (O_306,N_8956,N_9438);
nor UO_307 (O_307,N_8475,N_8467);
nor UO_308 (O_308,N_9028,N_8172);
nand UO_309 (O_309,N_8021,N_9336);
or UO_310 (O_310,N_9297,N_8827);
nand UO_311 (O_311,N_9973,N_8429);
nor UO_312 (O_312,N_8164,N_8980);
or UO_313 (O_313,N_9369,N_9141);
nand UO_314 (O_314,N_9301,N_9129);
nor UO_315 (O_315,N_9424,N_9690);
nor UO_316 (O_316,N_8714,N_9507);
and UO_317 (O_317,N_9150,N_9253);
xnor UO_318 (O_318,N_8942,N_8436);
nor UO_319 (O_319,N_9076,N_8711);
or UO_320 (O_320,N_9467,N_8123);
nor UO_321 (O_321,N_9319,N_9627);
nand UO_322 (O_322,N_8512,N_9442);
or UO_323 (O_323,N_9552,N_8348);
nor UO_324 (O_324,N_9163,N_8904);
or UO_325 (O_325,N_8915,N_8473);
nor UO_326 (O_326,N_8399,N_9653);
nor UO_327 (O_327,N_8978,N_8064);
nand UO_328 (O_328,N_8496,N_9900);
nand UO_329 (O_329,N_9276,N_9296);
nand UO_330 (O_330,N_9976,N_8726);
or UO_331 (O_331,N_9183,N_9464);
and UO_332 (O_332,N_9285,N_9897);
nor UO_333 (O_333,N_8893,N_9853);
or UO_334 (O_334,N_8020,N_8269);
nor UO_335 (O_335,N_8217,N_9909);
or UO_336 (O_336,N_8477,N_8367);
and UO_337 (O_337,N_9047,N_9244);
nor UO_338 (O_338,N_9947,N_8322);
nand UO_339 (O_339,N_8468,N_8121);
nor UO_340 (O_340,N_8519,N_9902);
nor UO_341 (O_341,N_9867,N_8721);
or UO_342 (O_342,N_9687,N_8329);
and UO_343 (O_343,N_9892,N_8809);
nand UO_344 (O_344,N_9280,N_9194);
nor UO_345 (O_345,N_9181,N_9757);
and UO_346 (O_346,N_9735,N_8532);
nor UO_347 (O_347,N_8223,N_9207);
xor UO_348 (O_348,N_9016,N_9425);
or UO_349 (O_349,N_8879,N_8048);
nor UO_350 (O_350,N_8177,N_9119);
and UO_351 (O_351,N_9543,N_9572);
or UO_352 (O_352,N_8347,N_8174);
nand UO_353 (O_353,N_9212,N_9613);
nand UO_354 (O_354,N_9531,N_9796);
nand UO_355 (O_355,N_8602,N_9238);
nor UO_356 (O_356,N_9905,N_8285);
nand UO_357 (O_357,N_9753,N_9461);
nor UO_358 (O_358,N_8908,N_9925);
and UO_359 (O_359,N_9358,N_8571);
or UO_360 (O_360,N_8053,N_9843);
and UO_361 (O_361,N_9649,N_9638);
nor UO_362 (O_362,N_8356,N_9506);
nand UO_363 (O_363,N_9813,N_9996);
or UO_364 (O_364,N_8629,N_9966);
or UO_365 (O_365,N_9400,N_9906);
and UO_366 (O_366,N_9211,N_9998);
nor UO_367 (O_367,N_8178,N_8516);
or UO_368 (O_368,N_8352,N_9985);
nor UO_369 (O_369,N_9582,N_9036);
and UO_370 (O_370,N_8451,N_8158);
nor UO_371 (O_371,N_8418,N_8125);
and UO_372 (O_372,N_8845,N_9224);
nor UO_373 (O_373,N_8407,N_9527);
or UO_374 (O_374,N_9795,N_9990);
or UO_375 (O_375,N_9515,N_8645);
nand UO_376 (O_376,N_8404,N_9099);
nor UO_377 (O_377,N_9804,N_8487);
or UO_378 (O_378,N_8783,N_9323);
or UO_379 (O_379,N_9834,N_9155);
or UO_380 (O_380,N_9974,N_9768);
and UO_381 (O_381,N_9981,N_9132);
nand UO_382 (O_382,N_9781,N_8248);
nand UO_383 (O_383,N_8585,N_9520);
or UO_384 (O_384,N_8401,N_9445);
and UO_385 (O_385,N_9287,N_8592);
and UO_386 (O_386,N_8612,N_8417);
nand UO_387 (O_387,N_9027,N_9696);
and UO_388 (O_388,N_8002,N_8993);
and UO_389 (O_389,N_8134,N_9204);
or UO_390 (O_390,N_9650,N_9137);
nor UO_391 (O_391,N_8040,N_9116);
nand UO_392 (O_392,N_9798,N_9387);
nor UO_393 (O_393,N_9943,N_9283);
nand UO_394 (O_394,N_8746,N_8119);
nand UO_395 (O_395,N_9429,N_9433);
nand UO_396 (O_396,N_9868,N_9351);
nand UO_397 (O_397,N_8175,N_9273);
nor UO_398 (O_398,N_9660,N_9934);
nand UO_399 (O_399,N_9532,N_8324);
or UO_400 (O_400,N_9307,N_8626);
nor UO_401 (O_401,N_8857,N_9748);
and UO_402 (O_402,N_8885,N_8447);
and UO_403 (O_403,N_8839,N_8983);
and UO_404 (O_404,N_9221,N_9623);
nand UO_405 (O_405,N_9801,N_8462);
nand UO_406 (O_406,N_9035,N_8952);
and UO_407 (O_407,N_8917,N_9645);
or UO_408 (O_408,N_9432,N_8313);
nor UO_409 (O_409,N_9410,N_8430);
nand UO_410 (O_410,N_9252,N_9073);
or UO_411 (O_411,N_8854,N_8165);
nor UO_412 (O_412,N_9015,N_9199);
nand UO_413 (O_413,N_8441,N_8559);
nor UO_414 (O_414,N_8610,N_8989);
nand UO_415 (O_415,N_8283,N_8372);
nand UO_416 (O_416,N_8867,N_9957);
nor UO_417 (O_417,N_9320,N_9959);
or UO_418 (O_418,N_9202,N_9371);
nor UO_419 (O_419,N_8769,N_8138);
and UO_420 (O_420,N_8586,N_8087);
and UO_421 (O_421,N_9126,N_9270);
nor UO_422 (O_422,N_8745,N_9752);
and UO_423 (O_423,N_9539,N_9584);
and UO_424 (O_424,N_9736,N_8884);
nand UO_425 (O_425,N_8963,N_9195);
and UO_426 (O_426,N_8182,N_8794);
and UO_427 (O_427,N_9325,N_9389);
and UO_428 (O_428,N_8067,N_9805);
nor UO_429 (O_429,N_8587,N_8648);
and UO_430 (O_430,N_8575,N_9070);
nor UO_431 (O_431,N_8267,N_8479);
nor UO_432 (O_432,N_9707,N_8100);
nand UO_433 (O_433,N_8606,N_9676);
nor UO_434 (O_434,N_9815,N_9222);
nand UO_435 (O_435,N_9335,N_9050);
and UO_436 (O_436,N_8762,N_8813);
nand UO_437 (O_437,N_8970,N_9629);
and UO_438 (O_438,N_8308,N_8744);
nor UO_439 (O_439,N_9373,N_8350);
nor UO_440 (O_440,N_9835,N_8448);
and UO_441 (O_441,N_8991,N_9877);
nor UO_442 (O_442,N_9392,N_9914);
and UO_443 (O_443,N_8408,N_9553);
nand UO_444 (O_444,N_8271,N_9046);
or UO_445 (O_445,N_8772,N_8976);
nand UO_446 (O_446,N_8715,N_9021);
nor UO_447 (O_447,N_8924,N_8506);
nor UO_448 (O_448,N_9006,N_9093);
xnor UO_449 (O_449,N_9450,N_8927);
or UO_450 (O_450,N_9554,N_9873);
or UO_451 (O_451,N_9500,N_9302);
nor UO_452 (O_452,N_8334,N_8374);
or UO_453 (O_453,N_8078,N_8708);
nand UO_454 (O_454,N_8984,N_9628);
nor UO_455 (O_455,N_8101,N_8779);
or UO_456 (O_456,N_8560,N_8050);
or UO_457 (O_457,N_8691,N_8568);
or UO_458 (O_458,N_9190,N_8202);
nand UO_459 (O_459,N_9139,N_8856);
nor UO_460 (O_460,N_9886,N_9658);
nor UO_461 (O_461,N_9081,N_8255);
or UO_462 (O_462,N_9361,N_9858);
nand UO_463 (O_463,N_8534,N_9967);
or UO_464 (O_464,N_8395,N_8082);
nand UO_465 (O_465,N_9210,N_9130);
nand UO_466 (O_466,N_9519,N_8685);
or UO_467 (O_467,N_8737,N_9448);
nand UO_468 (O_468,N_9596,N_9732);
and UO_469 (O_469,N_9128,N_9979);
nand UO_470 (O_470,N_9956,N_9497);
nor UO_471 (O_471,N_9758,N_8455);
nand UO_472 (O_472,N_8525,N_8106);
or UO_473 (O_473,N_8732,N_9338);
and UO_474 (O_474,N_8380,N_8480);
nand UO_475 (O_475,N_8219,N_9097);
and UO_476 (O_476,N_8405,N_9426);
nor UO_477 (O_477,N_9932,N_8416);
and UO_478 (O_478,N_8443,N_9637);
or UO_479 (O_479,N_9648,N_8168);
and UO_480 (O_480,N_9994,N_8790);
or UO_481 (O_481,N_9380,N_8695);
nand UO_482 (O_482,N_8660,N_9314);
or UO_483 (O_483,N_8419,N_8598);
nand UO_484 (O_484,N_9980,N_9309);
and UO_485 (O_485,N_8905,N_9665);
or UO_486 (O_486,N_8470,N_9295);
and UO_487 (O_487,N_9765,N_8265);
and UO_488 (O_488,N_9888,N_9334);
or UO_489 (O_489,N_8256,N_9406);
nor UO_490 (O_490,N_8961,N_9644);
nand UO_491 (O_491,N_9286,N_9347);
and UO_492 (O_492,N_9101,N_8572);
and UO_493 (O_493,N_9963,N_8483);
nand UO_494 (O_494,N_9079,N_8816);
nand UO_495 (O_495,N_9965,N_8538);
nand UO_496 (O_496,N_9235,N_8290);
and UO_497 (O_497,N_9794,N_9446);
nor UO_498 (O_498,N_9298,N_8320);
or UO_499 (O_499,N_8043,N_8292);
nand UO_500 (O_500,N_9060,N_9634);
and UO_501 (O_501,N_9226,N_8233);
or UO_502 (O_502,N_8147,N_8008);
and UO_503 (O_503,N_8312,N_8865);
nor UO_504 (O_504,N_8748,N_9953);
and UO_505 (O_505,N_9029,N_9738);
nand UO_506 (O_506,N_8740,N_9559);
nand UO_507 (O_507,N_8321,N_8891);
nand UO_508 (O_508,N_8039,N_8951);
or UO_509 (O_509,N_9625,N_8573);
or UO_510 (O_510,N_8832,N_8862);
and UO_511 (O_511,N_8342,N_9066);
or UO_512 (O_512,N_8244,N_9824);
and UO_513 (O_513,N_9340,N_8615);
xor UO_514 (O_514,N_9122,N_9237);
nand UO_515 (O_515,N_9762,N_9104);
nand UO_516 (O_516,N_9186,N_9394);
and UO_517 (O_517,N_9927,N_9262);
nor UO_518 (O_518,N_8381,N_8247);
nand UO_519 (O_519,N_9405,N_8383);
nor UO_520 (O_520,N_8641,N_8522);
or UO_521 (O_521,N_9165,N_8564);
nor UO_522 (O_522,N_9944,N_8712);
nor UO_523 (O_523,N_9242,N_8317);
nand UO_524 (O_524,N_9004,N_8758);
nor UO_525 (O_525,N_9059,N_9427);
nor UO_526 (O_526,N_8835,N_8968);
nor UO_527 (O_527,N_8800,N_8928);
or UO_528 (O_528,N_8599,N_9562);
nor UO_529 (O_529,N_9946,N_8154);
nand UO_530 (O_530,N_8524,N_8608);
xnor UO_531 (O_531,N_8542,N_8923);
nor UO_532 (O_532,N_9745,N_9493);
or UO_533 (O_533,N_9777,N_8755);
and UO_534 (O_534,N_9422,N_9560);
or UO_535 (O_535,N_9399,N_8230);
nand UO_536 (O_536,N_8895,N_8486);
nand UO_537 (O_537,N_9936,N_8171);
nor UO_538 (O_538,N_8270,N_9474);
nor UO_539 (O_539,N_9677,N_8143);
nand UO_540 (O_540,N_8011,N_8869);
nand UO_541 (O_541,N_9993,N_9662);
nor UO_542 (O_542,N_8262,N_9121);
nand UO_543 (O_543,N_9898,N_9513);
nand UO_544 (O_544,N_8601,N_9032);
or UO_545 (O_545,N_8117,N_8630);
and UO_546 (O_546,N_9664,N_9107);
nand UO_547 (O_547,N_8259,N_9024);
nand UO_548 (O_548,N_8294,N_9085);
nand UO_549 (O_549,N_9381,N_8055);
nand UO_550 (O_550,N_8034,N_8874);
or UO_551 (O_551,N_8914,N_9726);
or UO_552 (O_552,N_9612,N_9468);
nand UO_553 (O_553,N_8570,N_9178);
nand UO_554 (O_554,N_8588,N_9706);
or UO_555 (O_555,N_9030,N_8250);
nand UO_556 (O_556,N_8555,N_8464);
nand UO_557 (O_557,N_8205,N_9475);
and UO_558 (O_558,N_9045,N_8411);
nor UO_559 (O_559,N_8814,N_9383);
nor UO_560 (O_560,N_9248,N_8520);
or UO_561 (O_561,N_8272,N_9588);
or UO_562 (O_562,N_8912,N_9773);
and UO_563 (O_563,N_9546,N_8878);
nor UO_564 (O_564,N_9454,N_9372);
and UO_565 (O_565,N_9316,N_9498);
nand UO_566 (O_566,N_9217,N_8185);
or UO_567 (O_567,N_9246,N_9278);
and UO_568 (O_568,N_8720,N_9666);
nand UO_569 (O_569,N_9142,N_8332);
or UO_570 (O_570,N_8785,N_9859);
and UO_571 (O_571,N_8226,N_8741);
nor UO_572 (O_572,N_9279,N_9610);
nor UO_573 (O_573,N_8004,N_9023);
xnor UO_574 (O_574,N_9169,N_8051);
nand UO_575 (O_575,N_8445,N_9823);
and UO_576 (O_576,N_9376,N_8757);
nor UO_577 (O_577,N_9166,N_9949);
nor UO_578 (O_578,N_9161,N_8697);
nor UO_579 (O_579,N_8667,N_8805);
and UO_580 (O_580,N_9750,N_8647);
or UO_581 (O_581,N_9785,N_9530);
or UO_582 (O_582,N_8279,N_9601);
nand UO_583 (O_583,N_9377,N_9680);
or UO_584 (O_584,N_9039,N_8760);
and UO_585 (O_585,N_8355,N_8540);
nand UO_586 (O_586,N_9598,N_8073);
and UO_587 (O_587,N_8088,N_8153);
nor UO_588 (O_588,N_8442,N_9148);
nand UO_589 (O_589,N_9463,N_8209);
or UO_590 (O_590,N_9852,N_8201);
or UO_591 (O_591,N_8316,N_9026);
or UO_592 (O_592,N_9257,N_8302);
or UO_593 (O_593,N_9451,N_8728);
nor UO_594 (O_594,N_9489,N_9274);
nand UO_595 (O_595,N_9005,N_8710);
and UO_596 (O_596,N_8144,N_8239);
and UO_597 (O_597,N_9134,N_9803);
nor UO_598 (O_598,N_9499,N_9611);
and UO_599 (O_599,N_8566,N_9061);
nor UO_600 (O_600,N_8433,N_9348);
nand UO_601 (O_601,N_9904,N_9517);
and UO_602 (O_602,N_9018,N_9861);
or UO_603 (O_603,N_8133,N_9774);
nor UO_604 (O_604,N_9917,N_9615);
or UO_605 (O_605,N_9044,N_8930);
nand UO_606 (O_606,N_9413,N_9275);
nand UO_607 (O_607,N_8363,N_9538);
and UO_608 (O_608,N_9842,N_9153);
and UO_609 (O_609,N_8113,N_9930);
and UO_610 (O_610,N_9411,N_9679);
xnor UO_611 (O_611,N_8841,N_8297);
nand UO_612 (O_612,N_9105,N_8503);
or UO_613 (O_613,N_9828,N_8222);
nand UO_614 (O_614,N_8120,N_9703);
or UO_615 (O_615,N_8717,N_9174);
nor UO_616 (O_616,N_9250,N_9564);
or UO_617 (O_617,N_8764,N_8359);
and UO_618 (O_618,N_9189,N_8890);
nand UO_619 (O_619,N_9617,N_8860);
or UO_620 (O_620,N_9473,N_8919);
and UO_621 (O_621,N_9230,N_8421);
and UO_622 (O_622,N_8420,N_8080);
or UO_623 (O_623,N_8880,N_9223);
or UO_624 (O_624,N_9051,N_9022);
nand UO_625 (O_625,N_8386,N_9522);
nor UO_626 (O_626,N_9317,N_8981);
nor UO_627 (O_627,N_8149,N_9305);
or UO_628 (O_628,N_8593,N_8768);
nor UO_629 (O_629,N_8137,N_9565);
nor UO_630 (O_630,N_8554,N_9568);
nand UO_631 (O_631,N_8196,N_8193);
nor UO_632 (O_632,N_8861,N_8304);
xnor UO_633 (O_633,N_9864,N_8531);
nand UO_634 (O_634,N_8077,N_9135);
and UO_635 (O_635,N_8310,N_8994);
nand UO_636 (O_636,N_8530,N_8920);
nand UO_637 (O_637,N_8114,N_9312);
nand UO_638 (O_638,N_9404,N_8221);
or UO_639 (O_639,N_9618,N_8898);
nand UO_640 (O_640,N_9839,N_9151);
or UO_641 (O_641,N_8632,N_8457);
nand UO_642 (O_642,N_8622,N_9352);
or UO_643 (O_643,N_9632,N_8843);
xnor UO_644 (O_644,N_9578,N_8492);
nor UO_645 (O_645,N_9673,N_9641);
and UO_646 (O_646,N_9713,N_9365);
nor UO_647 (O_647,N_8289,N_8654);
nor UO_648 (O_648,N_9691,N_8183);
nand UO_649 (O_649,N_9688,N_9685);
nor UO_650 (O_650,N_8365,N_9062);
and UO_651 (O_651,N_9197,N_8998);
and UO_652 (O_652,N_8973,N_9084);
and UO_653 (O_653,N_8876,N_9783);
nor UO_654 (O_654,N_9970,N_8590);
nor UO_655 (O_655,N_8580,N_8403);
and UO_656 (O_656,N_8558,N_8713);
or UO_657 (O_657,N_9481,N_8894);
or UO_658 (O_658,N_9439,N_8770);
or UO_659 (O_659,N_8058,N_8799);
or UO_660 (O_660,N_9324,N_8979);
and UO_661 (O_661,N_8225,N_8935);
or UO_662 (O_662,N_9131,N_9831);
nand UO_663 (O_663,N_8655,N_8426);
and UO_664 (O_664,N_9409,N_8727);
and UO_665 (O_665,N_9486,N_9851);
and UO_666 (O_666,N_8176,N_9555);
nor UO_667 (O_667,N_8700,N_8625);
or UO_668 (O_668,N_8085,N_8280);
nor UO_669 (O_669,N_8902,N_9727);
nand UO_670 (O_670,N_8195,N_8543);
nand UO_671 (O_671,N_9791,N_8637);
nor UO_672 (O_672,N_9213,N_9595);
or UO_673 (O_673,N_8409,N_8837);
and UO_674 (O_674,N_8387,N_9263);
nand UO_675 (O_675,N_9844,N_9020);
or UO_676 (O_676,N_8784,N_8187);
and UO_677 (O_677,N_8929,N_8931);
nor UO_678 (O_678,N_8415,N_9072);
or UO_679 (O_679,N_9621,N_9709);
nand UO_680 (O_680,N_8471,N_9254);
and UO_681 (O_681,N_8730,N_8036);
nand UO_682 (O_682,N_8684,N_9537);
or UO_683 (O_683,N_8619,N_9216);
nand UO_684 (O_684,N_9299,N_9885);
and UO_685 (O_685,N_8484,N_8900);
nand UO_686 (O_686,N_8550,N_9342);
nor UO_687 (O_687,N_8916,N_8326);
and UO_688 (O_688,N_9605,N_9567);
and UO_689 (O_689,N_9982,N_9011);
nor UO_690 (O_690,N_9339,N_8987);
nand UO_691 (O_691,N_8323,N_8643);
or UO_692 (O_692,N_8000,N_9836);
and UO_693 (O_693,N_9899,N_9182);
and UO_694 (O_694,N_9184,N_9228);
nand UO_695 (O_695,N_9561,N_9682);
nand UO_696 (O_696,N_8037,N_8301);
nand UO_697 (O_697,N_8017,N_9291);
nor UO_698 (O_698,N_8286,N_8015);
nand UO_699 (O_699,N_8607,N_8603);
and UO_700 (O_700,N_8315,N_9989);
nor UO_701 (O_701,N_9655,N_8535);
nand UO_702 (O_702,N_8508,N_8897);
nand UO_703 (O_703,N_8116,N_9288);
and UO_704 (O_704,N_8939,N_8141);
nor UO_705 (O_705,N_8579,N_9125);
nor UO_706 (O_706,N_8263,N_9466);
or UO_707 (O_707,N_9616,N_8705);
or UO_708 (O_708,N_9661,N_9728);
nand UO_709 (O_709,N_8148,N_8108);
nor UO_710 (O_710,N_8682,N_9485);
and UO_711 (O_711,N_8238,N_9577);
or UO_712 (O_712,N_9540,N_8688);
nor UO_713 (O_713,N_8665,N_9916);
or UO_714 (O_714,N_9741,N_9152);
and UO_715 (O_715,N_9911,N_8013);
nand UO_716 (O_716,N_8494,N_9928);
or UO_717 (O_717,N_8553,N_9374);
or UO_718 (O_718,N_8960,N_9856);
or UO_719 (O_719,N_8424,N_9055);
nor UO_720 (O_720,N_9771,N_8815);
or UO_721 (O_721,N_9731,N_9972);
nand UO_722 (O_722,N_9143,N_8132);
and UO_723 (O_723,N_8673,N_8870);
nor UO_724 (O_724,N_9551,N_9479);
nor UO_725 (O_725,N_8393,N_9604);
or UO_726 (O_726,N_9269,N_8701);
or UO_727 (O_727,N_9826,N_9913);
nor UO_728 (O_728,N_8729,N_8544);
and UO_729 (O_729,N_8511,N_9443);
or UO_730 (O_730,N_9159,N_8686);
or UO_731 (O_731,N_8940,N_8333);
or UO_732 (O_732,N_9701,N_8373);
nand UO_733 (O_733,N_9800,N_8731);
nand UO_734 (O_734,N_9293,N_9310);
and UO_735 (O_735,N_8775,N_9366);
and UO_736 (O_736,N_9594,N_9412);
and UO_737 (O_737,N_9631,N_9133);
or UO_738 (O_738,N_8934,N_9702);
or UO_739 (O_739,N_9074,N_8489);
nor UO_740 (O_740,N_8161,N_9705);
and UO_741 (O_741,N_8215,N_8969);
nand UO_742 (O_742,N_8330,N_9367);
nand UO_743 (O_743,N_8029,N_9176);
and UO_744 (O_744,N_9810,N_8825);
and UO_745 (O_745,N_8115,N_9000);
nand UO_746 (O_746,N_8653,N_9841);
and UO_747 (O_747,N_8432,N_8107);
or UO_748 (O_748,N_9318,N_9458);
or UO_749 (O_749,N_9832,N_8192);
nand UO_750 (O_750,N_8620,N_9284);
nand UO_751 (O_751,N_9144,N_9881);
nor UO_752 (O_752,N_9205,N_8932);
or UO_753 (O_753,N_8318,N_8052);
and UO_754 (O_754,N_8061,N_8444);
nand UO_755 (O_755,N_9478,N_9171);
or UO_756 (O_756,N_9053,N_8157);
and UO_757 (O_757,N_9729,N_8812);
nor UO_758 (O_758,N_9063,N_9037);
nor UO_759 (O_759,N_9267,N_8251);
nor UO_760 (O_760,N_9191,N_9863);
nor UO_761 (O_761,N_8099,N_9659);
nand UO_762 (O_762,N_8838,N_8453);
or UO_763 (O_763,N_8958,N_9652);
and UO_764 (O_764,N_8070,N_9321);
nand UO_765 (O_765,N_8704,N_8844);
and UO_766 (O_766,N_9693,N_9243);
nand UO_767 (O_767,N_8155,N_8098);
and UO_768 (O_768,N_9579,N_9303);
nor UO_769 (O_769,N_9642,N_9386);
or UO_770 (O_770,N_9869,N_8651);
and UO_771 (O_771,N_8056,N_8140);
xor UO_772 (O_772,N_8463,N_8808);
nand UO_773 (O_773,N_8683,N_9407);
nor UO_774 (O_774,N_8822,N_8242);
or UO_775 (O_775,N_8778,N_8282);
or UO_776 (O_776,N_9654,N_9077);
nand UO_777 (O_777,N_9547,N_9459);
xor UO_778 (O_778,N_8009,N_9460);
nand UO_779 (O_779,N_8826,N_8227);
or UO_780 (O_780,N_8672,N_9162);
nor UO_781 (O_781,N_9657,N_9550);
nand UO_782 (O_782,N_9720,N_9872);
nor UO_783 (O_783,N_9948,N_9875);
nand UO_784 (O_784,N_8621,N_9054);
and UO_785 (O_785,N_8068,N_8724);
or UO_786 (O_786,N_9570,N_8957);
nand UO_787 (O_787,N_8999,N_9233);
and UO_788 (O_788,N_9068,N_8325);
nand UO_789 (O_789,N_9395,N_9516);
nand UO_790 (O_790,N_9712,N_9492);
or UO_791 (O_791,N_8735,N_9525);
nand UO_792 (O_792,N_8022,N_8252);
and UO_793 (O_793,N_9311,N_9669);
nand UO_794 (O_794,N_8967,N_9511);
and UO_795 (O_795,N_9330,N_9480);
nand UO_796 (O_796,N_9185,N_9755);
or UO_797 (O_797,N_8824,N_8003);
or UO_798 (O_798,N_8213,N_9488);
or UO_799 (O_799,N_8868,N_9083);
nand UO_800 (O_800,N_9449,N_8261);
or UO_801 (O_801,N_9802,N_9954);
nor UO_802 (O_802,N_9236,N_8084);
nor UO_803 (O_803,N_9180,N_8079);
and UO_804 (O_804,N_8818,N_8398);
and UO_805 (O_805,N_8299,N_9941);
nor UO_806 (O_806,N_8210,N_8142);
nor UO_807 (O_807,N_9769,N_8319);
nor UO_808 (O_808,N_8018,N_8959);
and UO_809 (O_809,N_9087,N_8131);
and UO_810 (O_810,N_9651,N_8074);
nor UO_811 (O_811,N_9699,N_9502);
nor UO_812 (O_812,N_9636,N_8243);
and UO_813 (O_813,N_8693,N_8309);
nand UO_814 (O_814,N_9421,N_8485);
nor UO_815 (O_815,N_9694,N_9724);
and UO_816 (O_816,N_8128,N_8237);
or UO_817 (O_817,N_9574,N_9830);
nand UO_818 (O_818,N_9501,N_8065);
nor UO_819 (O_819,N_9704,N_9746);
nor UO_820 (O_820,N_9784,N_9215);
nand UO_821 (O_821,N_8633,N_8853);
nand UO_822 (O_822,N_9154,N_8848);
or UO_823 (O_823,N_9419,N_9845);
and UO_824 (O_824,N_9124,N_9606);
nand UO_825 (O_825,N_9935,N_8771);
or UO_826 (O_826,N_9609,N_8948);
nand UO_827 (O_827,N_8362,N_9416);
nor UO_828 (O_828,N_8657,N_8803);
or UO_829 (O_829,N_8498,N_8591);
nand UO_830 (O_830,N_9120,N_8145);
and UO_831 (O_831,N_9656,N_8831);
and UO_832 (O_832,N_9788,N_8083);
nand UO_833 (O_833,N_8528,N_8298);
and UO_834 (O_834,N_9684,N_9526);
nand UO_835 (O_835,N_8234,N_9884);
and UO_836 (O_836,N_8293,N_9523);
nand UO_837 (O_837,N_9145,N_8006);
nand UO_838 (O_838,N_8110,N_8156);
and UO_839 (O_839,N_8611,N_9759);
nand UO_840 (O_840,N_8792,N_9172);
nand UO_841 (O_841,N_8507,N_9922);
or UO_842 (O_842,N_9418,N_9556);
nand UO_843 (O_843,N_9149,N_9754);
nand UO_844 (O_844,N_9770,N_8537);
or UO_845 (O_845,N_9668,N_9229);
nor UO_846 (O_846,N_9271,N_9846);
or UO_847 (O_847,N_9095,N_8819);
or UO_848 (O_848,N_8001,N_9509);
nor UO_849 (O_849,N_9672,N_9114);
or UO_850 (O_850,N_8881,N_9403);
or UO_851 (O_851,N_9639,N_9958);
nand UO_852 (O_852,N_8604,N_9245);
or UO_853 (O_853,N_8105,N_9456);
or UO_854 (O_854,N_9007,N_8500);
nor UO_855 (O_855,N_9986,N_9678);
or UO_856 (O_856,N_8569,N_8377);
and UO_857 (O_857,N_9797,N_8476);
nand UO_858 (O_858,N_9708,N_9260);
nor UO_859 (O_859,N_9667,N_8863);
nor UO_860 (O_860,N_9364,N_8847);
nor UO_861 (O_861,N_9827,N_8896);
nor UO_862 (O_862,N_9569,N_9575);
or UO_863 (O_863,N_8410,N_9393);
or UO_864 (O_864,N_8964,N_9034);
or UO_865 (O_865,N_9192,N_8041);
or UO_866 (O_866,N_8228,N_9711);
and UO_867 (O_867,N_8369,N_8596);
nand UO_868 (O_868,N_8062,N_8889);
or UO_869 (O_869,N_8354,N_9457);
or UO_870 (O_870,N_9597,N_9716);
nand UO_871 (O_871,N_8777,N_8184);
or UO_872 (O_872,N_8556,N_8111);
or UO_873 (O_873,N_8567,N_8548);
or UO_874 (O_874,N_8913,N_9012);
and UO_875 (O_875,N_9118,N_8698);
and UO_876 (O_876,N_9268,N_8063);
nand UO_877 (O_877,N_8828,N_9397);
or UO_878 (O_878,N_9740,N_9043);
and UO_879 (O_879,N_9505,N_9521);
or UO_880 (O_880,N_8690,N_8669);
or UO_881 (O_881,N_8780,N_8264);
nor UO_882 (O_882,N_8254,N_8702);
or UO_883 (O_883,N_8742,N_8767);
and UO_884 (O_884,N_8456,N_8945);
and UO_885 (O_885,N_8216,N_8636);
nor UO_886 (O_886,N_8955,N_9049);
and UO_887 (O_887,N_8765,N_9984);
and UO_888 (O_888,N_8541,N_8284);
nand UO_889 (O_889,N_9614,N_9469);
and UO_890 (O_890,N_8197,N_8357);
or UO_891 (O_891,N_8412,N_9017);
nand UO_892 (O_892,N_8146,N_9398);
or UO_893 (O_893,N_9833,N_9201);
or UO_894 (O_894,N_9173,N_9177);
or UO_895 (O_895,N_9722,N_9889);
or UO_896 (O_896,N_8414,N_8482);
nor UO_897 (O_897,N_9428,N_8389);
nand UO_898 (O_898,N_9510,N_8802);
and UO_899 (O_899,N_8220,N_8076);
or UO_900 (O_900,N_9809,N_9487);
nand UO_901 (O_901,N_9430,N_8539);
and UO_902 (O_902,N_9179,N_8823);
and UO_903 (O_903,N_8562,N_8901);
nor UO_904 (O_904,N_8517,N_8624);
and UO_905 (O_905,N_8296,N_8019);
and UO_906 (O_906,N_9345,N_8551);
nor UO_907 (O_907,N_8966,N_8670);
nand UO_908 (O_908,N_8328,N_9793);
or UO_909 (O_909,N_8756,N_9840);
nand UO_910 (O_910,N_9857,N_8801);
nand UO_911 (O_911,N_8909,N_8925);
and UO_912 (O_912,N_8127,N_9940);
nor UO_913 (O_913,N_9390,N_8169);
or UO_914 (O_914,N_8212,N_9306);
nor UO_915 (O_915,N_8345,N_8235);
nand UO_916 (O_916,N_9462,N_8510);
nand UO_917 (O_917,N_8846,N_8791);
and UO_918 (O_918,N_9193,N_9962);
and UO_919 (O_919,N_8472,N_9354);
nand UO_920 (O_920,N_9743,N_9991);
xnor UO_921 (O_921,N_9328,N_9031);
and UO_922 (O_922,N_9635,N_8208);
nor UO_923 (O_923,N_9807,N_8787);
nor UO_924 (O_924,N_9908,N_8159);
or UO_925 (O_925,N_8763,N_8872);
or UO_926 (O_926,N_8071,N_8584);
or UO_927 (O_927,N_8469,N_8811);
nor UO_928 (O_928,N_8723,N_8490);
or UO_929 (O_929,N_8358,N_9591);
and UO_930 (O_930,N_8378,N_8266);
or UO_931 (O_931,N_9106,N_8024);
nand UO_932 (O_932,N_8985,N_8385);
nand UO_933 (O_933,N_8938,N_8796);
and UO_934 (O_934,N_8287,N_8351);
or UO_935 (O_935,N_8859,N_9415);
nor UO_936 (O_936,N_8390,N_9700);
nand UO_937 (O_937,N_8033,N_8650);
or UO_938 (O_938,N_8883,N_8718);
nand UO_939 (O_939,N_8066,N_8722);
and UO_940 (O_940,N_9903,N_9187);
nor UO_941 (O_941,N_8361,N_9329);
nor UO_942 (O_942,N_9518,N_8709);
nor UO_943 (O_943,N_8341,N_9602);
nor UO_944 (O_944,N_9040,N_9341);
nand UO_945 (O_945,N_9465,N_8804);
or UO_946 (O_946,N_8975,N_8533);
and UO_947 (O_947,N_8766,N_9357);
nand UO_948 (O_948,N_9876,N_9013);
nor UO_949 (O_949,N_8042,N_8194);
and UO_950 (O_950,N_8501,N_9939);
and UO_951 (O_951,N_9643,N_8759);
nand UO_952 (O_952,N_9763,N_8707);
nor UO_953 (O_953,N_8992,N_8595);
and UO_954 (O_954,N_8577,N_9926);
and UO_955 (O_955,N_8733,N_8095);
or UO_956 (O_956,N_9790,N_8699);
nor UO_957 (O_957,N_9808,N_8339);
or UO_958 (O_958,N_8130,N_9010);
nor UO_959 (O_959,N_8173,N_8435);
or UO_960 (O_960,N_8030,N_9717);
and UO_961 (O_961,N_9697,N_8866);
nand UO_962 (O_962,N_8396,N_9402);
or UO_963 (O_963,N_9346,N_9091);
nor UO_964 (O_964,N_8514,N_8245);
nand UO_965 (O_965,N_9240,N_9548);
and UO_966 (O_966,N_8798,N_8198);
and UO_967 (O_967,N_8678,N_8652);
or UO_968 (O_968,N_9483,N_8166);
and UO_969 (O_969,N_9992,N_9950);
or UO_970 (O_970,N_8706,N_9477);
nor UO_971 (O_971,N_8032,N_9444);
nand UO_972 (O_972,N_9327,N_9113);
and UO_973 (O_973,N_9772,N_9375);
and UO_974 (O_974,N_8305,N_8384);
or UO_975 (O_975,N_9140,N_9961);
or UO_976 (O_976,N_8833,N_9001);
nor UO_977 (O_977,N_9471,N_9907);
nand UO_978 (O_978,N_8180,N_8793);
nor UO_979 (O_979,N_9127,N_9671);
or UO_980 (O_980,N_8623,N_9272);
and UO_981 (O_981,N_8754,N_8502);
and UO_982 (O_982,N_9999,N_9647);
or UO_983 (O_983,N_8493,N_8773);
or UO_984 (O_984,N_8438,N_8892);
nor UO_985 (O_985,N_8086,N_8054);
or UO_986 (O_986,N_8346,N_9535);
xnor UO_987 (O_987,N_8240,N_9938);
or UO_988 (O_988,N_9893,N_9681);
and UO_989 (O_989,N_9751,N_9534);
nor UO_990 (O_990,N_9599,N_9838);
or UO_991 (O_991,N_9585,N_9025);
or UO_992 (O_992,N_8439,N_8075);
nand UO_993 (O_993,N_9094,N_8738);
or UO_994 (O_994,N_8249,N_8875);
nand UO_995 (O_995,N_8103,N_9078);
or UO_996 (O_996,N_8023,N_9887);
nand UO_997 (O_997,N_9080,N_8306);
nand UO_998 (O_998,N_9168,N_9558);
or UO_999 (O_999,N_8431,N_9590);
and UO_1000 (O_1000,N_9114,N_8801);
nand UO_1001 (O_1001,N_9235,N_9457);
or UO_1002 (O_1002,N_8654,N_9286);
or UO_1003 (O_1003,N_8928,N_8037);
and UO_1004 (O_1004,N_9640,N_9064);
nor UO_1005 (O_1005,N_8076,N_8779);
nor UO_1006 (O_1006,N_8591,N_9659);
nor UO_1007 (O_1007,N_8093,N_9409);
or UO_1008 (O_1008,N_8103,N_8244);
nand UO_1009 (O_1009,N_8903,N_8047);
nor UO_1010 (O_1010,N_9481,N_8183);
or UO_1011 (O_1011,N_8360,N_9436);
nand UO_1012 (O_1012,N_8745,N_8686);
nand UO_1013 (O_1013,N_9089,N_8359);
nand UO_1014 (O_1014,N_8155,N_9151);
nand UO_1015 (O_1015,N_9800,N_8683);
nor UO_1016 (O_1016,N_8317,N_8255);
and UO_1017 (O_1017,N_9441,N_8882);
and UO_1018 (O_1018,N_9766,N_9916);
or UO_1019 (O_1019,N_9771,N_9714);
and UO_1020 (O_1020,N_8969,N_8925);
nor UO_1021 (O_1021,N_8094,N_8306);
nand UO_1022 (O_1022,N_8839,N_8565);
or UO_1023 (O_1023,N_8784,N_8536);
nor UO_1024 (O_1024,N_9881,N_8543);
or UO_1025 (O_1025,N_9051,N_9178);
nor UO_1026 (O_1026,N_8403,N_9180);
and UO_1027 (O_1027,N_9500,N_8609);
nand UO_1028 (O_1028,N_8153,N_9179);
or UO_1029 (O_1029,N_8968,N_8462);
nor UO_1030 (O_1030,N_9215,N_9439);
or UO_1031 (O_1031,N_8678,N_9446);
or UO_1032 (O_1032,N_8887,N_8056);
nand UO_1033 (O_1033,N_9118,N_9473);
and UO_1034 (O_1034,N_9273,N_9811);
or UO_1035 (O_1035,N_8001,N_8177);
or UO_1036 (O_1036,N_8007,N_8564);
nand UO_1037 (O_1037,N_8913,N_8076);
nor UO_1038 (O_1038,N_9207,N_9720);
nor UO_1039 (O_1039,N_8439,N_9380);
or UO_1040 (O_1040,N_9206,N_9531);
or UO_1041 (O_1041,N_8351,N_8318);
nand UO_1042 (O_1042,N_9874,N_8405);
nand UO_1043 (O_1043,N_8668,N_9665);
and UO_1044 (O_1044,N_8990,N_9752);
nor UO_1045 (O_1045,N_9325,N_9267);
nor UO_1046 (O_1046,N_9113,N_9486);
nor UO_1047 (O_1047,N_8076,N_9114);
or UO_1048 (O_1048,N_8929,N_9873);
nor UO_1049 (O_1049,N_9569,N_8636);
and UO_1050 (O_1050,N_8595,N_8855);
nand UO_1051 (O_1051,N_9681,N_8033);
or UO_1052 (O_1052,N_9085,N_8140);
or UO_1053 (O_1053,N_8175,N_8415);
or UO_1054 (O_1054,N_9808,N_8027);
and UO_1055 (O_1055,N_9853,N_8709);
nor UO_1056 (O_1056,N_9470,N_9283);
or UO_1057 (O_1057,N_8551,N_9232);
or UO_1058 (O_1058,N_8430,N_9346);
and UO_1059 (O_1059,N_8581,N_8507);
or UO_1060 (O_1060,N_8190,N_9958);
nand UO_1061 (O_1061,N_9014,N_9401);
and UO_1062 (O_1062,N_9687,N_9539);
or UO_1063 (O_1063,N_8322,N_8202);
nand UO_1064 (O_1064,N_9880,N_9733);
and UO_1065 (O_1065,N_8859,N_8277);
or UO_1066 (O_1066,N_8896,N_9403);
and UO_1067 (O_1067,N_9455,N_8896);
or UO_1068 (O_1068,N_8142,N_9755);
or UO_1069 (O_1069,N_9199,N_9499);
or UO_1070 (O_1070,N_9012,N_8887);
nand UO_1071 (O_1071,N_9823,N_9639);
nand UO_1072 (O_1072,N_8126,N_9555);
and UO_1073 (O_1073,N_9190,N_8755);
and UO_1074 (O_1074,N_9591,N_9260);
and UO_1075 (O_1075,N_8832,N_8228);
nor UO_1076 (O_1076,N_8843,N_8102);
nor UO_1077 (O_1077,N_8211,N_9451);
or UO_1078 (O_1078,N_9617,N_8414);
or UO_1079 (O_1079,N_9819,N_8891);
or UO_1080 (O_1080,N_8714,N_9445);
nand UO_1081 (O_1081,N_8977,N_8380);
nor UO_1082 (O_1082,N_8182,N_9792);
nand UO_1083 (O_1083,N_9136,N_9687);
nand UO_1084 (O_1084,N_9470,N_8559);
nor UO_1085 (O_1085,N_8716,N_9323);
and UO_1086 (O_1086,N_9676,N_8750);
nor UO_1087 (O_1087,N_8569,N_9427);
nor UO_1088 (O_1088,N_9394,N_9699);
nand UO_1089 (O_1089,N_8226,N_9634);
nand UO_1090 (O_1090,N_8668,N_9875);
or UO_1091 (O_1091,N_8880,N_8164);
nor UO_1092 (O_1092,N_8354,N_9654);
nand UO_1093 (O_1093,N_9118,N_8647);
nor UO_1094 (O_1094,N_9890,N_9085);
or UO_1095 (O_1095,N_9378,N_9782);
nand UO_1096 (O_1096,N_9253,N_8060);
nor UO_1097 (O_1097,N_9799,N_8726);
nand UO_1098 (O_1098,N_8689,N_8209);
and UO_1099 (O_1099,N_9585,N_9930);
and UO_1100 (O_1100,N_8768,N_8248);
or UO_1101 (O_1101,N_9980,N_8861);
and UO_1102 (O_1102,N_9552,N_9073);
or UO_1103 (O_1103,N_9108,N_9643);
or UO_1104 (O_1104,N_9503,N_9034);
nand UO_1105 (O_1105,N_9715,N_8390);
or UO_1106 (O_1106,N_9260,N_9922);
nor UO_1107 (O_1107,N_9937,N_8002);
nand UO_1108 (O_1108,N_8163,N_8982);
or UO_1109 (O_1109,N_8345,N_9791);
or UO_1110 (O_1110,N_8253,N_8804);
nor UO_1111 (O_1111,N_8127,N_8133);
nor UO_1112 (O_1112,N_9931,N_8238);
or UO_1113 (O_1113,N_9045,N_9995);
nor UO_1114 (O_1114,N_9906,N_8136);
nand UO_1115 (O_1115,N_9655,N_8952);
nor UO_1116 (O_1116,N_9113,N_8998);
and UO_1117 (O_1117,N_8425,N_8424);
nor UO_1118 (O_1118,N_8621,N_9467);
nor UO_1119 (O_1119,N_9754,N_9532);
nor UO_1120 (O_1120,N_9256,N_8596);
and UO_1121 (O_1121,N_9574,N_9825);
nor UO_1122 (O_1122,N_9538,N_8335);
nor UO_1123 (O_1123,N_9733,N_9431);
nand UO_1124 (O_1124,N_8303,N_9402);
and UO_1125 (O_1125,N_9611,N_8281);
nand UO_1126 (O_1126,N_9834,N_8143);
nor UO_1127 (O_1127,N_9185,N_8960);
and UO_1128 (O_1128,N_8461,N_8234);
and UO_1129 (O_1129,N_8046,N_8483);
and UO_1130 (O_1130,N_9578,N_9646);
nand UO_1131 (O_1131,N_8631,N_8915);
or UO_1132 (O_1132,N_9198,N_9854);
nor UO_1133 (O_1133,N_9072,N_9056);
and UO_1134 (O_1134,N_8370,N_9424);
nand UO_1135 (O_1135,N_8924,N_8683);
and UO_1136 (O_1136,N_9704,N_9178);
or UO_1137 (O_1137,N_9454,N_8777);
nor UO_1138 (O_1138,N_8855,N_9339);
nand UO_1139 (O_1139,N_8921,N_8818);
nand UO_1140 (O_1140,N_9165,N_8343);
and UO_1141 (O_1141,N_8699,N_9580);
nand UO_1142 (O_1142,N_8074,N_9620);
nor UO_1143 (O_1143,N_8592,N_9184);
nor UO_1144 (O_1144,N_9790,N_9637);
or UO_1145 (O_1145,N_8179,N_9601);
nor UO_1146 (O_1146,N_9870,N_8383);
and UO_1147 (O_1147,N_8339,N_9798);
and UO_1148 (O_1148,N_8645,N_9445);
nor UO_1149 (O_1149,N_8449,N_8398);
nor UO_1150 (O_1150,N_8440,N_8875);
nor UO_1151 (O_1151,N_9887,N_8712);
or UO_1152 (O_1152,N_9698,N_8335);
or UO_1153 (O_1153,N_9986,N_8262);
nand UO_1154 (O_1154,N_9666,N_8142);
or UO_1155 (O_1155,N_9880,N_8643);
or UO_1156 (O_1156,N_9592,N_9394);
nor UO_1157 (O_1157,N_8830,N_9346);
and UO_1158 (O_1158,N_9199,N_8623);
or UO_1159 (O_1159,N_9327,N_9642);
nand UO_1160 (O_1160,N_9191,N_9449);
nor UO_1161 (O_1161,N_9978,N_9908);
nor UO_1162 (O_1162,N_9174,N_9811);
and UO_1163 (O_1163,N_8428,N_8678);
and UO_1164 (O_1164,N_9165,N_9502);
and UO_1165 (O_1165,N_9878,N_8378);
or UO_1166 (O_1166,N_8830,N_9381);
and UO_1167 (O_1167,N_8963,N_9483);
nor UO_1168 (O_1168,N_9264,N_8254);
or UO_1169 (O_1169,N_9973,N_9807);
or UO_1170 (O_1170,N_9674,N_8801);
nand UO_1171 (O_1171,N_8050,N_8609);
nor UO_1172 (O_1172,N_8577,N_8343);
nand UO_1173 (O_1173,N_8713,N_8684);
and UO_1174 (O_1174,N_9715,N_8052);
nor UO_1175 (O_1175,N_8054,N_8120);
and UO_1176 (O_1176,N_8480,N_8744);
nor UO_1177 (O_1177,N_9943,N_8570);
and UO_1178 (O_1178,N_8810,N_9130);
or UO_1179 (O_1179,N_8111,N_9991);
or UO_1180 (O_1180,N_9594,N_9959);
or UO_1181 (O_1181,N_9538,N_8668);
nor UO_1182 (O_1182,N_8921,N_9036);
nand UO_1183 (O_1183,N_8427,N_9606);
or UO_1184 (O_1184,N_9258,N_9266);
or UO_1185 (O_1185,N_8013,N_9157);
or UO_1186 (O_1186,N_9143,N_9832);
or UO_1187 (O_1187,N_8087,N_9761);
or UO_1188 (O_1188,N_8361,N_8277);
and UO_1189 (O_1189,N_8032,N_8341);
and UO_1190 (O_1190,N_8792,N_8669);
xnor UO_1191 (O_1191,N_9051,N_8052);
nand UO_1192 (O_1192,N_9503,N_8783);
and UO_1193 (O_1193,N_8901,N_9816);
or UO_1194 (O_1194,N_9548,N_8818);
nor UO_1195 (O_1195,N_8364,N_8172);
nor UO_1196 (O_1196,N_9226,N_9295);
nand UO_1197 (O_1197,N_9783,N_9136);
or UO_1198 (O_1198,N_9667,N_9984);
or UO_1199 (O_1199,N_9429,N_8967);
nor UO_1200 (O_1200,N_9821,N_8058);
and UO_1201 (O_1201,N_9495,N_8501);
or UO_1202 (O_1202,N_9974,N_8453);
or UO_1203 (O_1203,N_8196,N_8992);
nand UO_1204 (O_1204,N_8650,N_9664);
nand UO_1205 (O_1205,N_9235,N_8493);
or UO_1206 (O_1206,N_9059,N_9294);
or UO_1207 (O_1207,N_9104,N_8516);
and UO_1208 (O_1208,N_9962,N_8967);
and UO_1209 (O_1209,N_9041,N_8800);
and UO_1210 (O_1210,N_8435,N_9501);
or UO_1211 (O_1211,N_9803,N_9136);
and UO_1212 (O_1212,N_8389,N_9051);
or UO_1213 (O_1213,N_8986,N_8380);
nand UO_1214 (O_1214,N_9941,N_8993);
or UO_1215 (O_1215,N_8709,N_9034);
nor UO_1216 (O_1216,N_9938,N_8702);
or UO_1217 (O_1217,N_9728,N_8982);
nor UO_1218 (O_1218,N_8988,N_9470);
nor UO_1219 (O_1219,N_8068,N_9633);
nand UO_1220 (O_1220,N_8951,N_9508);
nand UO_1221 (O_1221,N_8732,N_8577);
nor UO_1222 (O_1222,N_8774,N_8428);
nand UO_1223 (O_1223,N_8663,N_8341);
nor UO_1224 (O_1224,N_9696,N_9157);
nand UO_1225 (O_1225,N_8786,N_9159);
nor UO_1226 (O_1226,N_8020,N_9130);
or UO_1227 (O_1227,N_9640,N_9699);
nor UO_1228 (O_1228,N_9526,N_9194);
nor UO_1229 (O_1229,N_8944,N_8174);
and UO_1230 (O_1230,N_8832,N_9412);
xnor UO_1231 (O_1231,N_9226,N_8857);
nand UO_1232 (O_1232,N_8710,N_9919);
nand UO_1233 (O_1233,N_8386,N_8955);
and UO_1234 (O_1234,N_8127,N_9049);
nor UO_1235 (O_1235,N_9256,N_9020);
nand UO_1236 (O_1236,N_8338,N_8808);
nor UO_1237 (O_1237,N_8650,N_8165);
nor UO_1238 (O_1238,N_9511,N_9958);
or UO_1239 (O_1239,N_8803,N_8175);
and UO_1240 (O_1240,N_9342,N_8657);
nor UO_1241 (O_1241,N_9351,N_9989);
and UO_1242 (O_1242,N_8426,N_8347);
and UO_1243 (O_1243,N_9645,N_9829);
or UO_1244 (O_1244,N_9498,N_9282);
nand UO_1245 (O_1245,N_8501,N_8678);
and UO_1246 (O_1246,N_8548,N_9451);
or UO_1247 (O_1247,N_9736,N_9941);
nand UO_1248 (O_1248,N_9576,N_9859);
nand UO_1249 (O_1249,N_8078,N_9197);
nor UO_1250 (O_1250,N_8444,N_9948);
or UO_1251 (O_1251,N_9983,N_8511);
nor UO_1252 (O_1252,N_8783,N_9381);
and UO_1253 (O_1253,N_8683,N_9804);
or UO_1254 (O_1254,N_9265,N_8305);
or UO_1255 (O_1255,N_8557,N_9464);
nor UO_1256 (O_1256,N_9046,N_8812);
and UO_1257 (O_1257,N_9932,N_9625);
nor UO_1258 (O_1258,N_9191,N_8094);
nand UO_1259 (O_1259,N_8750,N_9911);
or UO_1260 (O_1260,N_8963,N_8650);
nand UO_1261 (O_1261,N_9418,N_9196);
and UO_1262 (O_1262,N_8935,N_8831);
nand UO_1263 (O_1263,N_8572,N_8536);
or UO_1264 (O_1264,N_8275,N_8495);
nor UO_1265 (O_1265,N_9715,N_9157);
and UO_1266 (O_1266,N_9847,N_9707);
nor UO_1267 (O_1267,N_9503,N_9700);
and UO_1268 (O_1268,N_8077,N_9720);
nand UO_1269 (O_1269,N_9939,N_8593);
nor UO_1270 (O_1270,N_9526,N_8562);
and UO_1271 (O_1271,N_9200,N_9191);
nand UO_1272 (O_1272,N_8465,N_9859);
or UO_1273 (O_1273,N_8162,N_9559);
and UO_1274 (O_1274,N_8562,N_9209);
or UO_1275 (O_1275,N_9254,N_9721);
nor UO_1276 (O_1276,N_8181,N_9832);
nor UO_1277 (O_1277,N_9938,N_8635);
nand UO_1278 (O_1278,N_9221,N_8978);
nor UO_1279 (O_1279,N_9413,N_8551);
and UO_1280 (O_1280,N_8694,N_8535);
and UO_1281 (O_1281,N_9533,N_9499);
nor UO_1282 (O_1282,N_9675,N_8807);
nor UO_1283 (O_1283,N_8358,N_9046);
and UO_1284 (O_1284,N_9654,N_8961);
or UO_1285 (O_1285,N_9941,N_9425);
or UO_1286 (O_1286,N_9292,N_9990);
nand UO_1287 (O_1287,N_8503,N_8515);
or UO_1288 (O_1288,N_8553,N_9393);
nand UO_1289 (O_1289,N_8789,N_9177);
xor UO_1290 (O_1290,N_8916,N_9448);
and UO_1291 (O_1291,N_9029,N_8138);
nor UO_1292 (O_1292,N_8368,N_8539);
nor UO_1293 (O_1293,N_9617,N_8718);
or UO_1294 (O_1294,N_8184,N_9505);
nor UO_1295 (O_1295,N_8142,N_9864);
or UO_1296 (O_1296,N_9814,N_8897);
nand UO_1297 (O_1297,N_8379,N_8838);
and UO_1298 (O_1298,N_8842,N_9500);
nor UO_1299 (O_1299,N_8371,N_9131);
nand UO_1300 (O_1300,N_9509,N_9951);
nand UO_1301 (O_1301,N_8002,N_8209);
and UO_1302 (O_1302,N_9400,N_8008);
and UO_1303 (O_1303,N_8206,N_9975);
nor UO_1304 (O_1304,N_8438,N_8916);
nor UO_1305 (O_1305,N_8340,N_8677);
nor UO_1306 (O_1306,N_8485,N_9429);
or UO_1307 (O_1307,N_8023,N_8070);
nand UO_1308 (O_1308,N_9194,N_8954);
or UO_1309 (O_1309,N_8765,N_8360);
nor UO_1310 (O_1310,N_9331,N_8433);
nor UO_1311 (O_1311,N_9515,N_9192);
nor UO_1312 (O_1312,N_8820,N_8893);
nand UO_1313 (O_1313,N_8102,N_9555);
nor UO_1314 (O_1314,N_9692,N_9412);
and UO_1315 (O_1315,N_9209,N_9833);
and UO_1316 (O_1316,N_9782,N_8460);
nand UO_1317 (O_1317,N_8307,N_9345);
nor UO_1318 (O_1318,N_8408,N_9581);
xnor UO_1319 (O_1319,N_8392,N_9944);
or UO_1320 (O_1320,N_8789,N_8315);
and UO_1321 (O_1321,N_9321,N_9728);
nor UO_1322 (O_1322,N_9472,N_8080);
nand UO_1323 (O_1323,N_9562,N_8387);
and UO_1324 (O_1324,N_8007,N_8000);
or UO_1325 (O_1325,N_9069,N_9216);
nor UO_1326 (O_1326,N_8536,N_9675);
and UO_1327 (O_1327,N_9155,N_8693);
nor UO_1328 (O_1328,N_8863,N_8798);
nand UO_1329 (O_1329,N_9450,N_8714);
and UO_1330 (O_1330,N_8119,N_8066);
nand UO_1331 (O_1331,N_9368,N_9399);
and UO_1332 (O_1332,N_8777,N_9386);
nand UO_1333 (O_1333,N_9309,N_9131);
nand UO_1334 (O_1334,N_8672,N_9991);
and UO_1335 (O_1335,N_8799,N_9440);
or UO_1336 (O_1336,N_8471,N_8030);
nor UO_1337 (O_1337,N_9990,N_9389);
and UO_1338 (O_1338,N_9009,N_8065);
nor UO_1339 (O_1339,N_8238,N_8052);
nand UO_1340 (O_1340,N_8464,N_8025);
or UO_1341 (O_1341,N_8809,N_8711);
nor UO_1342 (O_1342,N_8900,N_9952);
nand UO_1343 (O_1343,N_9102,N_9896);
or UO_1344 (O_1344,N_8515,N_9218);
nand UO_1345 (O_1345,N_8529,N_8669);
nand UO_1346 (O_1346,N_9653,N_9521);
nand UO_1347 (O_1347,N_8489,N_9812);
or UO_1348 (O_1348,N_9360,N_8536);
nor UO_1349 (O_1349,N_9600,N_9618);
nand UO_1350 (O_1350,N_8836,N_8867);
nand UO_1351 (O_1351,N_8608,N_9494);
and UO_1352 (O_1352,N_8218,N_8238);
nor UO_1353 (O_1353,N_9233,N_9457);
nand UO_1354 (O_1354,N_9331,N_9014);
or UO_1355 (O_1355,N_9931,N_8588);
and UO_1356 (O_1356,N_9906,N_8813);
and UO_1357 (O_1357,N_8562,N_9433);
and UO_1358 (O_1358,N_8049,N_9034);
nand UO_1359 (O_1359,N_9594,N_9053);
or UO_1360 (O_1360,N_9052,N_8152);
and UO_1361 (O_1361,N_8444,N_8826);
nor UO_1362 (O_1362,N_8673,N_9033);
xor UO_1363 (O_1363,N_9556,N_8617);
nand UO_1364 (O_1364,N_8819,N_8668);
or UO_1365 (O_1365,N_8313,N_8785);
or UO_1366 (O_1366,N_9256,N_9547);
or UO_1367 (O_1367,N_8280,N_8216);
and UO_1368 (O_1368,N_9791,N_9572);
nor UO_1369 (O_1369,N_8257,N_8610);
and UO_1370 (O_1370,N_8737,N_9867);
and UO_1371 (O_1371,N_8572,N_9780);
nand UO_1372 (O_1372,N_8806,N_8066);
or UO_1373 (O_1373,N_8894,N_8296);
nand UO_1374 (O_1374,N_8306,N_8271);
nand UO_1375 (O_1375,N_9052,N_8610);
and UO_1376 (O_1376,N_8557,N_9038);
nor UO_1377 (O_1377,N_8887,N_8910);
nand UO_1378 (O_1378,N_8529,N_8190);
and UO_1379 (O_1379,N_9595,N_8332);
or UO_1380 (O_1380,N_8858,N_8874);
or UO_1381 (O_1381,N_8919,N_8825);
nor UO_1382 (O_1382,N_9380,N_9506);
and UO_1383 (O_1383,N_8359,N_9175);
nand UO_1384 (O_1384,N_9678,N_9594);
or UO_1385 (O_1385,N_8567,N_8278);
nand UO_1386 (O_1386,N_8119,N_9246);
nor UO_1387 (O_1387,N_8225,N_8975);
nor UO_1388 (O_1388,N_9387,N_8415);
or UO_1389 (O_1389,N_9065,N_9164);
nand UO_1390 (O_1390,N_9278,N_9242);
nor UO_1391 (O_1391,N_9342,N_8541);
nand UO_1392 (O_1392,N_8800,N_9176);
or UO_1393 (O_1393,N_8617,N_8632);
and UO_1394 (O_1394,N_8603,N_8337);
nand UO_1395 (O_1395,N_9794,N_9347);
and UO_1396 (O_1396,N_8024,N_9074);
nor UO_1397 (O_1397,N_8465,N_8243);
and UO_1398 (O_1398,N_8574,N_8143);
and UO_1399 (O_1399,N_8930,N_9939);
nor UO_1400 (O_1400,N_8889,N_8326);
nor UO_1401 (O_1401,N_9425,N_9347);
nand UO_1402 (O_1402,N_8581,N_9064);
or UO_1403 (O_1403,N_8631,N_9600);
and UO_1404 (O_1404,N_8658,N_8159);
and UO_1405 (O_1405,N_9512,N_8448);
nand UO_1406 (O_1406,N_8175,N_9874);
and UO_1407 (O_1407,N_9380,N_9507);
and UO_1408 (O_1408,N_9665,N_8935);
xnor UO_1409 (O_1409,N_8775,N_8772);
or UO_1410 (O_1410,N_8100,N_9796);
and UO_1411 (O_1411,N_8232,N_8445);
and UO_1412 (O_1412,N_9637,N_8116);
or UO_1413 (O_1413,N_9281,N_9267);
and UO_1414 (O_1414,N_8244,N_9508);
nor UO_1415 (O_1415,N_9719,N_8633);
xnor UO_1416 (O_1416,N_9729,N_8913);
and UO_1417 (O_1417,N_8959,N_9603);
nand UO_1418 (O_1418,N_9889,N_8436);
or UO_1419 (O_1419,N_8311,N_8596);
and UO_1420 (O_1420,N_8468,N_8662);
or UO_1421 (O_1421,N_8373,N_8737);
nor UO_1422 (O_1422,N_9655,N_8779);
nand UO_1423 (O_1423,N_8667,N_8303);
or UO_1424 (O_1424,N_8735,N_8515);
nand UO_1425 (O_1425,N_8486,N_9030);
and UO_1426 (O_1426,N_9105,N_9709);
nor UO_1427 (O_1427,N_8098,N_9390);
and UO_1428 (O_1428,N_8322,N_8030);
nand UO_1429 (O_1429,N_8253,N_9172);
nand UO_1430 (O_1430,N_8483,N_8978);
and UO_1431 (O_1431,N_9564,N_9585);
nand UO_1432 (O_1432,N_8130,N_9824);
or UO_1433 (O_1433,N_9509,N_8780);
or UO_1434 (O_1434,N_9912,N_8838);
and UO_1435 (O_1435,N_9779,N_9361);
nand UO_1436 (O_1436,N_8515,N_8336);
or UO_1437 (O_1437,N_8327,N_8804);
nor UO_1438 (O_1438,N_8657,N_9672);
or UO_1439 (O_1439,N_9332,N_8490);
nor UO_1440 (O_1440,N_8297,N_9344);
or UO_1441 (O_1441,N_8718,N_8049);
and UO_1442 (O_1442,N_8725,N_8056);
or UO_1443 (O_1443,N_9197,N_9768);
or UO_1444 (O_1444,N_8421,N_8840);
nand UO_1445 (O_1445,N_8945,N_9538);
and UO_1446 (O_1446,N_9882,N_8496);
nand UO_1447 (O_1447,N_9950,N_8524);
nor UO_1448 (O_1448,N_8808,N_9030);
nor UO_1449 (O_1449,N_8764,N_9698);
or UO_1450 (O_1450,N_8924,N_9148);
and UO_1451 (O_1451,N_8746,N_8053);
nand UO_1452 (O_1452,N_8122,N_8841);
and UO_1453 (O_1453,N_8122,N_9854);
nand UO_1454 (O_1454,N_8465,N_9834);
nor UO_1455 (O_1455,N_8541,N_9071);
nor UO_1456 (O_1456,N_9607,N_8883);
or UO_1457 (O_1457,N_8167,N_9684);
and UO_1458 (O_1458,N_8092,N_8030);
and UO_1459 (O_1459,N_9426,N_9622);
nor UO_1460 (O_1460,N_9419,N_8599);
or UO_1461 (O_1461,N_8856,N_8164);
or UO_1462 (O_1462,N_8902,N_9460);
and UO_1463 (O_1463,N_9055,N_8408);
nor UO_1464 (O_1464,N_9285,N_8891);
nor UO_1465 (O_1465,N_9560,N_8037);
or UO_1466 (O_1466,N_8844,N_9693);
nor UO_1467 (O_1467,N_9936,N_9115);
and UO_1468 (O_1468,N_8735,N_8864);
nor UO_1469 (O_1469,N_9087,N_8149);
nor UO_1470 (O_1470,N_9442,N_9276);
and UO_1471 (O_1471,N_9837,N_8625);
nand UO_1472 (O_1472,N_8870,N_8145);
and UO_1473 (O_1473,N_8841,N_9513);
nand UO_1474 (O_1474,N_8968,N_9038);
and UO_1475 (O_1475,N_8396,N_8965);
or UO_1476 (O_1476,N_9657,N_9040);
or UO_1477 (O_1477,N_9303,N_9271);
and UO_1478 (O_1478,N_9518,N_9138);
and UO_1479 (O_1479,N_8785,N_9677);
nor UO_1480 (O_1480,N_9119,N_9447);
or UO_1481 (O_1481,N_8512,N_9140);
nand UO_1482 (O_1482,N_8757,N_8618);
nor UO_1483 (O_1483,N_8384,N_8902);
nor UO_1484 (O_1484,N_8560,N_9681);
nor UO_1485 (O_1485,N_8196,N_8202);
nand UO_1486 (O_1486,N_9069,N_9081);
or UO_1487 (O_1487,N_9364,N_9374);
nor UO_1488 (O_1488,N_9166,N_8396);
nor UO_1489 (O_1489,N_8052,N_9847);
or UO_1490 (O_1490,N_9291,N_8616);
and UO_1491 (O_1491,N_9719,N_9069);
nor UO_1492 (O_1492,N_9445,N_9617);
or UO_1493 (O_1493,N_9050,N_8644);
nand UO_1494 (O_1494,N_9245,N_9744);
and UO_1495 (O_1495,N_9710,N_9215);
nor UO_1496 (O_1496,N_9125,N_9324);
or UO_1497 (O_1497,N_8080,N_8010);
and UO_1498 (O_1498,N_8338,N_8296);
or UO_1499 (O_1499,N_9116,N_8212);
endmodule