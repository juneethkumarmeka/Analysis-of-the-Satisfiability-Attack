module basic_1000_10000_1500_10_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_474,In_451);
nor U1 (N_1,In_150,In_869);
xnor U2 (N_2,In_859,In_639);
xnor U3 (N_3,In_970,In_50);
xnor U4 (N_4,In_117,In_473);
nor U5 (N_5,In_865,In_858);
or U6 (N_6,In_59,In_571);
or U7 (N_7,In_308,In_90);
or U8 (N_8,In_259,In_65);
nor U9 (N_9,In_875,In_387);
or U10 (N_10,In_876,In_0);
or U11 (N_11,In_882,In_977);
nand U12 (N_12,In_362,In_357);
or U13 (N_13,In_825,In_124);
nand U14 (N_14,In_167,In_763);
nand U15 (N_15,In_670,In_930);
nor U16 (N_16,In_266,In_126);
or U17 (N_17,In_247,In_191);
or U18 (N_18,In_132,In_91);
nand U19 (N_19,In_181,In_727);
nand U20 (N_20,In_155,In_919);
or U21 (N_21,In_598,In_234);
nor U22 (N_22,In_256,In_146);
nand U23 (N_23,In_114,In_99);
nor U24 (N_24,In_341,In_228);
xor U25 (N_25,In_276,In_540);
nand U26 (N_26,In_136,In_866);
nand U27 (N_27,In_425,In_106);
and U28 (N_28,In_547,In_394);
or U29 (N_29,In_567,In_609);
nor U30 (N_30,In_775,In_189);
nor U31 (N_31,In_856,In_129);
and U32 (N_32,In_310,In_364);
nor U33 (N_33,In_732,In_834);
xor U34 (N_34,In_820,In_695);
nand U35 (N_35,In_261,In_360);
or U36 (N_36,In_384,In_439);
nand U37 (N_37,In_583,In_996);
or U38 (N_38,In_511,In_229);
nor U39 (N_39,In_239,In_885);
and U40 (N_40,In_741,In_306);
and U41 (N_41,In_765,In_333);
nor U42 (N_42,In_494,In_46);
and U43 (N_43,In_322,In_340);
and U44 (N_44,In_734,In_161);
nor U45 (N_45,In_270,In_7);
nor U46 (N_46,In_211,In_339);
nand U47 (N_47,In_331,In_397);
and U48 (N_48,In_319,In_575);
nand U49 (N_49,In_900,In_554);
nor U50 (N_50,In_512,In_610);
nor U51 (N_51,In_49,In_243);
nand U52 (N_52,In_915,In_354);
nand U53 (N_53,In_180,In_534);
nor U54 (N_54,In_258,In_574);
and U55 (N_55,In_173,In_216);
or U56 (N_56,In_221,In_315);
nor U57 (N_57,In_367,In_215);
and U58 (N_58,In_537,In_469);
and U59 (N_59,In_570,In_93);
nor U60 (N_60,In_72,In_892);
nand U61 (N_61,In_186,In_1);
nand U62 (N_62,In_110,In_486);
xnor U63 (N_63,In_946,In_391);
nor U64 (N_64,In_11,In_896);
nand U65 (N_65,In_751,In_926);
nor U66 (N_66,In_768,In_895);
and U67 (N_67,In_159,In_585);
nor U68 (N_68,In_304,In_950);
nor U69 (N_69,In_939,In_351);
xnor U70 (N_70,In_48,In_648);
nand U71 (N_71,In_918,In_388);
and U72 (N_72,In_293,In_368);
and U73 (N_73,In_720,In_395);
and U74 (N_74,In_36,In_974);
nand U75 (N_75,In_767,In_785);
nor U76 (N_76,In_416,In_699);
or U77 (N_77,In_23,In_448);
nor U78 (N_78,In_249,In_497);
nand U79 (N_79,In_994,In_576);
nor U80 (N_80,In_78,In_112);
and U81 (N_81,In_881,In_353);
or U82 (N_82,In_645,In_927);
nor U83 (N_83,In_418,In_894);
xnor U84 (N_84,In_764,In_281);
nand U85 (N_85,In_466,In_849);
nor U86 (N_86,In_685,In_361);
xnor U87 (N_87,In_641,In_27);
nor U88 (N_88,In_62,In_912);
nand U89 (N_89,In_246,In_454);
or U90 (N_90,In_325,In_985);
and U91 (N_91,In_171,In_156);
nand U92 (N_92,In_484,In_737);
or U93 (N_93,In_203,In_967);
nor U94 (N_94,In_210,In_123);
nor U95 (N_95,In_908,In_43);
nand U96 (N_96,In_682,In_613);
or U97 (N_97,In_412,In_477);
nor U98 (N_98,In_470,In_952);
and U99 (N_99,In_515,In_519);
or U100 (N_100,In_868,In_64);
or U101 (N_101,In_476,In_461);
or U102 (N_102,In_546,In_483);
or U103 (N_103,In_482,In_651);
and U104 (N_104,In_642,In_224);
nand U105 (N_105,In_53,In_703);
and U106 (N_106,In_716,In_819);
nand U107 (N_107,In_843,In_817);
nand U108 (N_108,In_860,In_627);
or U109 (N_109,In_640,In_20);
and U110 (N_110,In_260,In_45);
nor U111 (N_111,In_710,In_671);
or U112 (N_112,In_424,In_431);
nand U113 (N_113,In_52,In_141);
or U114 (N_114,In_182,In_678);
nand U115 (N_115,In_564,In_521);
nor U116 (N_116,In_986,In_214);
or U117 (N_117,In_997,In_905);
or U118 (N_118,In_691,In_760);
or U119 (N_119,In_271,In_717);
nand U120 (N_120,In_404,In_343);
nand U121 (N_121,In_558,In_85);
and U122 (N_122,In_586,In_984);
or U123 (N_123,In_969,In_55);
nor U124 (N_124,In_749,In_272);
nand U125 (N_125,In_995,In_514);
or U126 (N_126,In_793,In_233);
nor U127 (N_127,In_545,In_97);
and U128 (N_128,In_795,In_76);
and U129 (N_129,In_375,In_163);
and U130 (N_130,In_369,In_536);
or U131 (N_131,In_807,In_621);
nor U132 (N_132,In_355,In_693);
nand U133 (N_133,In_157,In_430);
and U134 (N_134,In_383,In_619);
or U135 (N_135,In_565,In_955);
nor U136 (N_136,In_836,In_581);
nand U137 (N_137,In_615,In_411);
or U138 (N_138,In_30,In_127);
xnor U139 (N_139,In_426,In_176);
xnor U140 (N_140,In_646,In_206);
xnor U141 (N_141,In_195,In_965);
xor U142 (N_142,In_573,In_551);
nor U143 (N_143,In_240,In_471);
nand U144 (N_144,In_659,In_874);
and U145 (N_145,In_104,In_89);
nor U146 (N_146,In_287,In_312);
xor U147 (N_147,In_971,In_634);
nand U148 (N_148,In_294,In_465);
and U149 (N_149,In_614,In_596);
or U150 (N_150,In_457,In_956);
xor U151 (N_151,In_878,In_916);
and U152 (N_152,In_787,In_638);
and U153 (N_153,In_135,In_872);
nor U154 (N_154,In_406,In_120);
or U155 (N_155,In_784,In_501);
xor U156 (N_156,In_830,In_92);
nand U157 (N_157,In_962,In_376);
nor U158 (N_158,In_917,In_747);
nor U159 (N_159,In_602,In_718);
xor U160 (N_160,In_263,In_160);
nand U161 (N_161,In_326,In_495);
or U162 (N_162,In_844,In_746);
nand U163 (N_163,In_972,In_169);
nand U164 (N_164,In_623,In_944);
and U165 (N_165,In_380,In_405);
and U166 (N_166,In_608,In_831);
or U167 (N_167,In_202,In_697);
or U168 (N_168,In_788,In_102);
or U169 (N_169,In_840,In_218);
and U170 (N_170,In_667,In_673);
nor U171 (N_171,In_480,In_278);
nor U172 (N_172,In_21,In_624);
xor U173 (N_173,In_329,In_599);
or U174 (N_174,In_232,In_442);
nand U175 (N_175,In_879,In_337);
nand U176 (N_176,In_550,In_696);
nand U177 (N_177,In_715,In_108);
nor U178 (N_178,In_957,In_744);
and U179 (N_179,In_643,In_561);
nor U180 (N_180,In_488,In_655);
xor U181 (N_181,In_147,In_101);
nor U182 (N_182,In_725,In_154);
or U183 (N_183,In_230,In_222);
and U184 (N_184,In_818,In_739);
nor U185 (N_185,In_264,In_556);
xor U186 (N_186,In_225,In_100);
nor U187 (N_187,In_566,In_274);
nand U188 (N_188,In_724,In_37);
xnor U189 (N_189,In_137,In_863);
xor U190 (N_190,In_372,In_538);
nand U191 (N_191,In_6,In_933);
or U192 (N_192,In_653,In_47);
and U193 (N_193,In_604,In_932);
nor U194 (N_194,In_183,In_428);
and U195 (N_195,In_806,In_209);
and U196 (N_196,In_557,In_398);
nand U197 (N_197,In_292,In_140);
nand U198 (N_198,In_686,In_403);
xnor U199 (N_199,In_657,In_75);
and U200 (N_200,In_899,In_832);
nand U201 (N_201,In_177,In_267);
nand U202 (N_202,In_904,In_95);
nand U203 (N_203,In_936,In_630);
and U204 (N_204,In_420,In_527);
nor U205 (N_205,In_752,In_683);
or U206 (N_206,In_890,In_253);
or U207 (N_207,In_756,In_204);
and U208 (N_208,In_505,In_804);
or U209 (N_209,In_948,In_188);
and U210 (N_210,In_794,In_980);
nand U211 (N_211,In_897,In_589);
nor U212 (N_212,In_422,In_689);
nand U213 (N_213,In_198,In_982);
and U214 (N_214,In_450,In_553);
or U215 (N_215,In_63,In_783);
nand U216 (N_216,In_94,In_711);
nand U217 (N_217,In_838,In_433);
or U218 (N_218,In_786,In_814);
nand U219 (N_219,In_929,In_719);
and U220 (N_220,In_620,In_200);
or U221 (N_221,In_907,In_219);
and U222 (N_222,In_616,In_635);
nor U223 (N_223,In_77,In_286);
and U224 (N_224,In_330,In_170);
nand U225 (N_225,In_166,In_297);
and U226 (N_226,In_130,In_38);
or U227 (N_227,In_409,In_883);
and U228 (N_228,In_694,In_288);
nor U229 (N_229,In_805,In_845);
or U230 (N_230,In_880,In_867);
nand U231 (N_231,In_712,In_138);
nor U232 (N_232,In_73,In_728);
and U233 (N_233,In_318,In_766);
and U234 (N_234,In_745,In_810);
or U235 (N_235,In_321,In_975);
nand U236 (N_236,In_777,In_220);
or U237 (N_237,In_432,In_365);
nor U238 (N_238,In_812,In_870);
nor U239 (N_239,In_194,In_663);
nand U240 (N_240,In_781,In_612);
xor U241 (N_241,In_601,In_298);
xor U242 (N_242,In_174,In_208);
and U243 (N_243,In_945,In_305);
nand U244 (N_244,In_371,In_808);
nor U245 (N_245,In_61,In_611);
or U246 (N_246,In_713,In_96);
or U247 (N_247,In_662,In_31);
xor U248 (N_248,In_603,In_893);
xnor U249 (N_249,In_801,In_410);
nor U250 (N_250,In_937,In_226);
nand U251 (N_251,In_668,In_498);
nor U252 (N_252,In_563,In_798);
nand U253 (N_253,In_593,In_847);
nand U254 (N_254,In_823,In_647);
nand U255 (N_255,In_66,In_217);
xor U256 (N_256,In_778,In_921);
and U257 (N_257,In_854,In_453);
or U258 (N_258,In_821,In_987);
and U259 (N_259,In_600,In_503);
and U260 (N_260,In_753,In_769);
xor U261 (N_261,In_569,In_485);
and U262 (N_262,In_931,In_207);
nor U263 (N_263,In_607,In_731);
nand U264 (N_264,In_58,In_676);
xor U265 (N_265,In_508,In_345);
nand U266 (N_266,In_153,In_625);
nand U267 (N_267,In_344,In_109);
or U268 (N_268,In_197,In_891);
nand U269 (N_269,In_743,In_733);
and U270 (N_270,In_782,In_80);
nor U271 (N_271,In_86,In_489);
nor U272 (N_272,In_184,In_456);
nand U273 (N_273,In_938,In_913);
nand U274 (N_274,In_780,In_530);
and U275 (N_275,In_327,In_871);
or U276 (N_276,In_903,In_981);
or U277 (N_277,In_920,In_317);
or U278 (N_278,In_579,In_235);
nand U279 (N_279,In_506,In_636);
nor U280 (N_280,In_148,In_618);
nand U281 (N_281,In_953,In_12);
nand U282 (N_282,In_835,In_444);
or U283 (N_283,In_923,In_520);
and U284 (N_284,In_963,In_726);
nor U285 (N_285,In_708,In_359);
and U286 (N_286,In_60,In_824);
and U287 (N_287,In_487,In_386);
or U288 (N_288,In_650,In_320);
nand U289 (N_289,In_684,In_669);
nor U290 (N_290,In_257,In_706);
nor U291 (N_291,In_179,In_594);
xnor U292 (N_292,In_158,In_791);
or U293 (N_293,In_18,In_951);
nand U294 (N_294,In_978,In_789);
nor U295 (N_295,In_468,In_231);
or U296 (N_296,In_853,In_901);
nor U297 (N_297,In_107,In_35);
or U298 (N_298,In_29,In_679);
nand U299 (N_299,In_842,In_850);
or U300 (N_300,In_750,In_828);
and U301 (N_301,In_943,In_307);
nor U302 (N_302,In_187,In_139);
or U303 (N_303,In_415,In_666);
or U304 (N_304,In_988,In_370);
nor U305 (N_305,In_71,In_934);
nand U306 (N_306,In_690,In_419);
or U307 (N_307,In_526,In_111);
xor U308 (N_308,In_884,In_976);
or U309 (N_309,In_34,In_4);
nand U310 (N_310,In_452,In_698);
and U311 (N_311,In_151,In_723);
nor U312 (N_312,In_434,In_479);
nor U313 (N_313,In_525,In_507);
or U314 (N_314,In_242,In_909);
and U315 (N_315,In_449,In_423);
xnor U316 (N_316,In_128,In_709);
or U317 (N_317,In_990,In_389);
nor U318 (N_318,In_363,In_629);
nand U319 (N_319,In_762,In_770);
nand U320 (N_320,In_280,In_300);
and U321 (N_321,In_236,In_83);
nand U322 (N_322,In_478,In_522);
and U323 (N_323,In_378,In_803);
nor U324 (N_324,In_660,In_16);
and U325 (N_325,In_533,In_82);
nor U326 (N_326,In_774,In_911);
nor U327 (N_327,In_730,In_999);
and U328 (N_328,In_374,In_134);
nor U329 (N_329,In_622,In_989);
nor U330 (N_330,In_87,In_324);
nor U331 (N_331,In_886,In_888);
xnor U332 (N_332,In_959,In_437);
nand U333 (N_333,In_144,In_721);
nand U334 (N_334,In_382,In_39);
or U335 (N_335,In_119,In_458);
nand U336 (N_336,In_3,In_510);
and U337 (N_337,In_175,In_69);
and U338 (N_338,In_941,In_857);
nand U339 (N_339,In_539,In_516);
xnor U340 (N_340,In_414,In_637);
and U341 (N_341,In_771,In_649);
nor U342 (N_342,In_961,In_284);
nor U343 (N_343,In_88,In_311);
nand U344 (N_344,In_346,In_509);
nand U345 (N_345,In_25,In_314);
and U346 (N_346,In_966,In_262);
and U347 (N_347,In_56,In_654);
nor U348 (N_348,In_595,In_532);
nor U349 (N_349,In_125,In_998);
nand U350 (N_350,In_692,In_658);
and U351 (N_351,In_42,In_675);
nor U352 (N_352,In_687,In_942);
and U353 (N_353,In_289,In_283);
or U354 (N_354,In_446,In_5);
or U355 (N_355,In_493,In_544);
and U356 (N_356,In_295,In_922);
nand U357 (N_357,In_290,In_250);
xnor U358 (N_358,In_877,In_736);
xnor U359 (N_359,In_273,In_811);
or U360 (N_360,In_67,In_702);
nand U361 (N_361,In_592,In_626);
or U362 (N_362,In_902,In_949);
xor U363 (N_363,In_122,In_652);
nand U364 (N_364,In_336,In_185);
and U365 (N_365,In_51,In_460);
and U366 (N_366,In_190,In_254);
and U367 (N_367,In_162,In_542);
nand U368 (N_368,In_664,In_392);
nor U369 (N_369,In_816,In_269);
or U370 (N_370,In_568,In_906);
and U371 (N_371,In_445,In_688);
or U372 (N_372,In_168,In_864);
xnor U373 (N_373,In_531,In_779);
or U374 (N_374,In_705,In_24);
or U375 (N_375,In_960,In_9);
and U376 (N_376,In_381,In_268);
and U377 (N_377,In_947,In_591);
nor U378 (N_378,In_455,In_848);
or U379 (N_379,In_928,In_584);
or U380 (N_380,In_562,In_342);
xor U381 (N_381,In_606,In_81);
nor U382 (N_382,In_41,In_681);
and U383 (N_383,In_26,In_390);
and U384 (N_384,In_898,In_152);
nand U385 (N_385,In_84,In_757);
or U386 (N_386,In_761,In_373);
xnor U387 (N_387,In_914,In_707);
or U388 (N_388,In_172,In_924);
and U389 (N_389,In_227,In_265);
nor U390 (N_390,In_396,In_577);
and U391 (N_391,In_98,In_958);
and U392 (N_392,In_491,In_964);
nor U393 (N_393,In_285,In_983);
and U394 (N_394,In_677,In_131);
or U395 (N_395,In_889,In_335);
xor U396 (N_396,In_349,In_772);
nor U397 (N_397,In_303,In_925);
nor U398 (N_398,In_358,In_524);
and U399 (N_399,In_193,In_490);
and U400 (N_400,In_427,In_587);
or U401 (N_401,In_113,In_837);
nor U402 (N_402,In_441,In_582);
nand U403 (N_403,In_323,In_887);
nand U404 (N_404,In_115,In_475);
and U405 (N_405,In_499,In_103);
and U406 (N_406,In_644,In_28);
nor U407 (N_407,In_301,In_393);
nor U408 (N_408,In_873,In_377);
or U409 (N_409,In_993,In_199);
and U410 (N_410,In_776,In_133);
nand U411 (N_411,In_523,In_54);
xnor U412 (N_412,In_633,In_991);
nand U413 (N_413,In_597,In_245);
nand U414 (N_414,In_758,In_438);
xnor U415 (N_415,In_447,In_348);
nor U416 (N_416,In_464,In_588);
or U417 (N_417,In_379,In_401);
or U418 (N_418,In_502,In_839);
xnor U419 (N_419,In_628,In_316);
xor U420 (N_420,In_296,In_70);
nor U421 (N_421,In_738,In_201);
and U422 (N_422,In_15,In_17);
xor U423 (N_423,In_529,In_467);
or U424 (N_424,In_631,In_237);
or U425 (N_425,In_385,In_347);
and U426 (N_426,In_861,In_33);
or U427 (N_427,In_541,In_833);
nor U428 (N_428,In_813,In_742);
nand U429 (N_429,In_19,In_178);
nand U430 (N_430,In_145,In_338);
and U431 (N_431,In_462,In_313);
or U432 (N_432,In_790,In_279);
and U433 (N_433,In_472,In_255);
nand U434 (N_434,In_238,In_862);
nor U435 (N_435,In_149,In_759);
nand U436 (N_436,In_164,In_299);
nor U437 (N_437,In_407,In_754);
nand U438 (N_438,In_755,In_500);
nand U439 (N_439,In_8,In_578);
and U440 (N_440,In_735,In_142);
nor U441 (N_441,In_535,In_617);
xnor U442 (N_442,In_661,In_822);
xor U443 (N_443,In_632,In_350);
nor U444 (N_444,In_74,In_252);
and U445 (N_445,In_192,In_665);
and U446 (N_446,In_674,In_435);
or U447 (N_447,In_729,In_552);
nor U448 (N_448,In_118,In_796);
nor U449 (N_449,In_443,In_559);
nand U450 (N_450,In_244,In_399);
nor U451 (N_451,In_973,In_459);
or U452 (N_452,In_165,In_400);
or U453 (N_453,In_543,In_421);
nor U454 (N_454,In_44,In_792);
or U455 (N_455,In_829,In_413);
nand U456 (N_456,In_463,In_196);
and U457 (N_457,In_809,In_302);
nand U458 (N_458,In_704,In_57);
nand U459 (N_459,In_121,In_797);
and U460 (N_460,In_440,In_672);
and U461 (N_461,In_496,In_143);
and U462 (N_462,In_366,In_408);
nor U463 (N_463,In_528,In_251);
nand U464 (N_464,In_940,In_802);
or U465 (N_465,In_701,In_846);
nand U466 (N_466,In_827,In_205);
nand U467 (N_467,In_2,In_555);
nand U468 (N_468,In_13,In_572);
and U469 (N_469,In_277,In_590);
nor U470 (N_470,In_800,In_700);
or U471 (N_471,In_841,In_212);
nor U472 (N_472,In_328,In_815);
nor U473 (N_473,In_605,In_40);
xnor U474 (N_474,In_352,In_248);
and U475 (N_475,In_356,In_680);
and U476 (N_476,In_748,In_968);
or U477 (N_477,In_22,In_213);
nor U478 (N_478,In_517,In_282);
and U479 (N_479,In_402,In_504);
and U480 (N_480,In_417,In_773);
nor U481 (N_481,In_241,In_935);
nor U482 (N_482,In_332,In_275);
or U483 (N_483,In_334,In_580);
xor U484 (N_484,In_429,In_309);
and U485 (N_485,In_992,In_492);
nand U486 (N_486,In_954,In_436);
nor U487 (N_487,In_105,In_518);
or U488 (N_488,In_223,In_116);
nor U489 (N_489,In_10,In_852);
nor U490 (N_490,In_291,In_979);
nand U491 (N_491,In_549,In_851);
or U492 (N_492,In_513,In_79);
and U493 (N_493,In_481,In_656);
nand U494 (N_494,In_722,In_855);
or U495 (N_495,In_799,In_826);
nand U496 (N_496,In_560,In_714);
nand U497 (N_497,In_910,In_14);
nor U498 (N_498,In_68,In_740);
and U499 (N_499,In_32,In_548);
and U500 (N_500,In_377,In_737);
and U501 (N_501,In_376,In_919);
or U502 (N_502,In_586,In_851);
or U503 (N_503,In_850,In_796);
nor U504 (N_504,In_368,In_445);
or U505 (N_505,In_812,In_605);
xnor U506 (N_506,In_733,In_372);
nand U507 (N_507,In_731,In_444);
and U508 (N_508,In_241,In_169);
or U509 (N_509,In_730,In_160);
and U510 (N_510,In_930,In_713);
nand U511 (N_511,In_351,In_153);
nor U512 (N_512,In_749,In_601);
nor U513 (N_513,In_495,In_601);
and U514 (N_514,In_915,In_474);
nor U515 (N_515,In_76,In_552);
and U516 (N_516,In_192,In_723);
nor U517 (N_517,In_397,In_584);
nand U518 (N_518,In_758,In_261);
nand U519 (N_519,In_713,In_3);
xor U520 (N_520,In_312,In_150);
nand U521 (N_521,In_599,In_756);
and U522 (N_522,In_517,In_915);
and U523 (N_523,In_522,In_32);
nand U524 (N_524,In_687,In_115);
xor U525 (N_525,In_25,In_394);
nor U526 (N_526,In_610,In_360);
xor U527 (N_527,In_281,In_289);
or U528 (N_528,In_31,In_987);
nand U529 (N_529,In_499,In_27);
and U530 (N_530,In_43,In_111);
nand U531 (N_531,In_558,In_802);
or U532 (N_532,In_916,In_142);
and U533 (N_533,In_631,In_106);
and U534 (N_534,In_217,In_49);
nor U535 (N_535,In_93,In_711);
xnor U536 (N_536,In_606,In_361);
and U537 (N_537,In_455,In_811);
and U538 (N_538,In_291,In_176);
xnor U539 (N_539,In_23,In_52);
nand U540 (N_540,In_150,In_41);
nor U541 (N_541,In_138,In_115);
nor U542 (N_542,In_293,In_983);
nor U543 (N_543,In_926,In_275);
or U544 (N_544,In_183,In_85);
nor U545 (N_545,In_589,In_506);
and U546 (N_546,In_355,In_869);
xor U547 (N_547,In_399,In_709);
nor U548 (N_548,In_899,In_283);
or U549 (N_549,In_942,In_283);
nand U550 (N_550,In_634,In_920);
nor U551 (N_551,In_145,In_761);
nor U552 (N_552,In_829,In_723);
nor U553 (N_553,In_471,In_57);
and U554 (N_554,In_367,In_294);
nor U555 (N_555,In_434,In_867);
nor U556 (N_556,In_465,In_476);
nor U557 (N_557,In_580,In_261);
or U558 (N_558,In_834,In_137);
or U559 (N_559,In_311,In_347);
nor U560 (N_560,In_363,In_659);
nor U561 (N_561,In_840,In_948);
nand U562 (N_562,In_641,In_139);
nor U563 (N_563,In_174,In_171);
xnor U564 (N_564,In_172,In_419);
nor U565 (N_565,In_219,In_14);
and U566 (N_566,In_737,In_733);
nand U567 (N_567,In_456,In_482);
nand U568 (N_568,In_837,In_438);
nand U569 (N_569,In_505,In_830);
or U570 (N_570,In_743,In_295);
and U571 (N_571,In_139,In_597);
or U572 (N_572,In_283,In_297);
or U573 (N_573,In_966,In_46);
or U574 (N_574,In_207,In_17);
and U575 (N_575,In_912,In_741);
or U576 (N_576,In_315,In_855);
and U577 (N_577,In_695,In_421);
nor U578 (N_578,In_125,In_631);
and U579 (N_579,In_462,In_415);
and U580 (N_580,In_783,In_508);
nor U581 (N_581,In_815,In_671);
xor U582 (N_582,In_419,In_970);
nor U583 (N_583,In_319,In_526);
and U584 (N_584,In_812,In_765);
and U585 (N_585,In_883,In_591);
nand U586 (N_586,In_315,In_542);
xnor U587 (N_587,In_578,In_601);
or U588 (N_588,In_212,In_355);
or U589 (N_589,In_896,In_804);
nand U590 (N_590,In_376,In_710);
nand U591 (N_591,In_697,In_380);
or U592 (N_592,In_236,In_902);
or U593 (N_593,In_865,In_293);
nand U594 (N_594,In_494,In_547);
nand U595 (N_595,In_664,In_361);
and U596 (N_596,In_500,In_225);
nand U597 (N_597,In_807,In_76);
nand U598 (N_598,In_901,In_385);
or U599 (N_599,In_15,In_833);
and U600 (N_600,In_822,In_883);
nor U601 (N_601,In_504,In_503);
nand U602 (N_602,In_896,In_259);
or U603 (N_603,In_528,In_26);
nand U604 (N_604,In_126,In_872);
or U605 (N_605,In_162,In_139);
or U606 (N_606,In_36,In_714);
or U607 (N_607,In_320,In_911);
nor U608 (N_608,In_134,In_931);
xor U609 (N_609,In_763,In_408);
nand U610 (N_610,In_898,In_536);
xnor U611 (N_611,In_623,In_888);
and U612 (N_612,In_638,In_708);
and U613 (N_613,In_851,In_114);
nor U614 (N_614,In_365,In_949);
nand U615 (N_615,In_721,In_628);
nand U616 (N_616,In_885,In_148);
nand U617 (N_617,In_225,In_641);
xor U618 (N_618,In_148,In_727);
or U619 (N_619,In_662,In_190);
nand U620 (N_620,In_618,In_915);
or U621 (N_621,In_26,In_236);
nor U622 (N_622,In_897,In_476);
nand U623 (N_623,In_52,In_273);
xnor U624 (N_624,In_169,In_906);
nor U625 (N_625,In_217,In_512);
nor U626 (N_626,In_653,In_380);
and U627 (N_627,In_438,In_72);
nor U628 (N_628,In_194,In_427);
or U629 (N_629,In_481,In_547);
nand U630 (N_630,In_319,In_356);
and U631 (N_631,In_949,In_612);
or U632 (N_632,In_714,In_602);
or U633 (N_633,In_580,In_231);
nor U634 (N_634,In_625,In_842);
or U635 (N_635,In_514,In_482);
nand U636 (N_636,In_746,In_476);
nor U637 (N_637,In_370,In_432);
and U638 (N_638,In_389,In_523);
nor U639 (N_639,In_646,In_107);
nand U640 (N_640,In_867,In_97);
nor U641 (N_641,In_861,In_509);
and U642 (N_642,In_182,In_393);
nand U643 (N_643,In_461,In_83);
nor U644 (N_644,In_746,In_929);
or U645 (N_645,In_442,In_576);
and U646 (N_646,In_527,In_878);
nor U647 (N_647,In_103,In_765);
xor U648 (N_648,In_869,In_416);
nor U649 (N_649,In_45,In_556);
or U650 (N_650,In_877,In_713);
nand U651 (N_651,In_609,In_255);
and U652 (N_652,In_749,In_697);
nand U653 (N_653,In_219,In_250);
nand U654 (N_654,In_600,In_320);
nor U655 (N_655,In_489,In_619);
and U656 (N_656,In_748,In_835);
and U657 (N_657,In_131,In_519);
and U658 (N_658,In_250,In_952);
or U659 (N_659,In_191,In_608);
nor U660 (N_660,In_260,In_240);
xnor U661 (N_661,In_866,In_411);
xor U662 (N_662,In_793,In_178);
or U663 (N_663,In_569,In_551);
or U664 (N_664,In_484,In_811);
nor U665 (N_665,In_356,In_402);
and U666 (N_666,In_349,In_881);
or U667 (N_667,In_452,In_322);
or U668 (N_668,In_851,In_635);
or U669 (N_669,In_961,In_736);
nor U670 (N_670,In_722,In_169);
or U671 (N_671,In_971,In_979);
nand U672 (N_672,In_745,In_841);
and U673 (N_673,In_90,In_735);
nand U674 (N_674,In_89,In_792);
nor U675 (N_675,In_788,In_561);
nor U676 (N_676,In_9,In_478);
or U677 (N_677,In_222,In_630);
and U678 (N_678,In_42,In_28);
xor U679 (N_679,In_603,In_160);
and U680 (N_680,In_37,In_431);
and U681 (N_681,In_804,In_15);
or U682 (N_682,In_254,In_179);
or U683 (N_683,In_64,In_351);
or U684 (N_684,In_415,In_606);
or U685 (N_685,In_991,In_23);
and U686 (N_686,In_278,In_685);
and U687 (N_687,In_524,In_576);
xor U688 (N_688,In_172,In_64);
or U689 (N_689,In_922,In_766);
or U690 (N_690,In_220,In_898);
and U691 (N_691,In_530,In_402);
nand U692 (N_692,In_766,In_928);
nand U693 (N_693,In_161,In_659);
xnor U694 (N_694,In_505,In_92);
and U695 (N_695,In_210,In_659);
or U696 (N_696,In_278,In_34);
nand U697 (N_697,In_18,In_229);
nand U698 (N_698,In_863,In_451);
and U699 (N_699,In_93,In_743);
and U700 (N_700,In_488,In_826);
and U701 (N_701,In_420,In_717);
and U702 (N_702,In_136,In_950);
and U703 (N_703,In_716,In_634);
nand U704 (N_704,In_881,In_203);
xor U705 (N_705,In_456,In_285);
nand U706 (N_706,In_715,In_122);
nor U707 (N_707,In_551,In_496);
nor U708 (N_708,In_292,In_775);
and U709 (N_709,In_285,In_770);
or U710 (N_710,In_524,In_646);
and U711 (N_711,In_717,In_529);
nor U712 (N_712,In_815,In_522);
nor U713 (N_713,In_819,In_150);
nor U714 (N_714,In_922,In_993);
or U715 (N_715,In_557,In_259);
or U716 (N_716,In_314,In_489);
nand U717 (N_717,In_405,In_479);
nor U718 (N_718,In_588,In_471);
nand U719 (N_719,In_302,In_368);
and U720 (N_720,In_306,In_345);
or U721 (N_721,In_607,In_217);
nand U722 (N_722,In_992,In_458);
nand U723 (N_723,In_696,In_492);
or U724 (N_724,In_611,In_247);
nor U725 (N_725,In_719,In_956);
or U726 (N_726,In_262,In_893);
and U727 (N_727,In_59,In_371);
xor U728 (N_728,In_492,In_196);
and U729 (N_729,In_146,In_100);
nor U730 (N_730,In_178,In_509);
and U731 (N_731,In_675,In_446);
nand U732 (N_732,In_537,In_751);
nor U733 (N_733,In_831,In_826);
nand U734 (N_734,In_215,In_617);
nand U735 (N_735,In_622,In_7);
and U736 (N_736,In_212,In_486);
nand U737 (N_737,In_223,In_433);
and U738 (N_738,In_404,In_521);
nor U739 (N_739,In_412,In_863);
nand U740 (N_740,In_966,In_957);
nand U741 (N_741,In_813,In_711);
nor U742 (N_742,In_615,In_699);
and U743 (N_743,In_852,In_112);
and U744 (N_744,In_251,In_415);
and U745 (N_745,In_276,In_680);
nor U746 (N_746,In_853,In_703);
xor U747 (N_747,In_22,In_767);
nand U748 (N_748,In_163,In_532);
nor U749 (N_749,In_918,In_392);
and U750 (N_750,In_719,In_367);
nand U751 (N_751,In_245,In_359);
and U752 (N_752,In_974,In_440);
nand U753 (N_753,In_254,In_200);
and U754 (N_754,In_749,In_282);
xnor U755 (N_755,In_434,In_792);
and U756 (N_756,In_320,In_309);
and U757 (N_757,In_8,In_514);
nor U758 (N_758,In_118,In_155);
nand U759 (N_759,In_100,In_119);
and U760 (N_760,In_627,In_5);
nand U761 (N_761,In_421,In_72);
or U762 (N_762,In_101,In_968);
and U763 (N_763,In_848,In_899);
or U764 (N_764,In_351,In_755);
nor U765 (N_765,In_416,In_331);
nand U766 (N_766,In_673,In_744);
nor U767 (N_767,In_223,In_77);
nor U768 (N_768,In_26,In_329);
or U769 (N_769,In_158,In_284);
xnor U770 (N_770,In_369,In_294);
and U771 (N_771,In_489,In_784);
nand U772 (N_772,In_854,In_157);
nor U773 (N_773,In_389,In_160);
or U774 (N_774,In_137,In_390);
nand U775 (N_775,In_479,In_236);
or U776 (N_776,In_656,In_298);
xnor U777 (N_777,In_318,In_787);
or U778 (N_778,In_565,In_78);
and U779 (N_779,In_461,In_144);
and U780 (N_780,In_804,In_178);
nand U781 (N_781,In_934,In_565);
and U782 (N_782,In_416,In_206);
nand U783 (N_783,In_996,In_736);
or U784 (N_784,In_739,In_287);
nand U785 (N_785,In_543,In_793);
and U786 (N_786,In_125,In_301);
or U787 (N_787,In_220,In_582);
nor U788 (N_788,In_486,In_191);
nor U789 (N_789,In_91,In_550);
nor U790 (N_790,In_345,In_718);
and U791 (N_791,In_898,In_79);
nand U792 (N_792,In_577,In_862);
nand U793 (N_793,In_427,In_735);
nor U794 (N_794,In_569,In_159);
or U795 (N_795,In_571,In_922);
nor U796 (N_796,In_654,In_988);
or U797 (N_797,In_971,In_884);
xnor U798 (N_798,In_280,In_450);
and U799 (N_799,In_552,In_797);
and U800 (N_800,In_221,In_346);
nand U801 (N_801,In_547,In_562);
nor U802 (N_802,In_110,In_321);
nand U803 (N_803,In_745,In_640);
or U804 (N_804,In_397,In_69);
and U805 (N_805,In_689,In_178);
or U806 (N_806,In_473,In_348);
nor U807 (N_807,In_924,In_605);
or U808 (N_808,In_859,In_267);
xor U809 (N_809,In_858,In_147);
nor U810 (N_810,In_238,In_62);
nand U811 (N_811,In_137,In_284);
nor U812 (N_812,In_213,In_545);
and U813 (N_813,In_676,In_44);
nor U814 (N_814,In_236,In_461);
and U815 (N_815,In_250,In_807);
or U816 (N_816,In_788,In_802);
nor U817 (N_817,In_338,In_652);
nand U818 (N_818,In_263,In_596);
or U819 (N_819,In_271,In_227);
and U820 (N_820,In_921,In_895);
xnor U821 (N_821,In_82,In_475);
and U822 (N_822,In_243,In_656);
nand U823 (N_823,In_396,In_946);
and U824 (N_824,In_909,In_819);
nand U825 (N_825,In_97,In_868);
nor U826 (N_826,In_812,In_262);
nor U827 (N_827,In_294,In_844);
and U828 (N_828,In_824,In_738);
or U829 (N_829,In_907,In_422);
nor U830 (N_830,In_44,In_723);
nand U831 (N_831,In_159,In_397);
nand U832 (N_832,In_312,In_99);
xnor U833 (N_833,In_954,In_283);
xnor U834 (N_834,In_884,In_684);
xor U835 (N_835,In_822,In_252);
or U836 (N_836,In_116,In_710);
nor U837 (N_837,In_7,In_693);
or U838 (N_838,In_724,In_261);
nor U839 (N_839,In_741,In_294);
nor U840 (N_840,In_579,In_92);
nand U841 (N_841,In_988,In_987);
xor U842 (N_842,In_742,In_595);
or U843 (N_843,In_334,In_636);
nor U844 (N_844,In_55,In_198);
and U845 (N_845,In_621,In_768);
nand U846 (N_846,In_339,In_497);
or U847 (N_847,In_210,In_862);
or U848 (N_848,In_384,In_529);
and U849 (N_849,In_586,In_877);
or U850 (N_850,In_220,In_103);
or U851 (N_851,In_519,In_584);
nand U852 (N_852,In_732,In_910);
or U853 (N_853,In_506,In_806);
nand U854 (N_854,In_798,In_292);
or U855 (N_855,In_561,In_766);
xor U856 (N_856,In_883,In_789);
and U857 (N_857,In_838,In_260);
and U858 (N_858,In_525,In_359);
nand U859 (N_859,In_980,In_824);
and U860 (N_860,In_892,In_666);
or U861 (N_861,In_662,In_532);
nor U862 (N_862,In_673,In_363);
nor U863 (N_863,In_888,In_35);
nor U864 (N_864,In_522,In_168);
nand U865 (N_865,In_562,In_99);
and U866 (N_866,In_659,In_550);
and U867 (N_867,In_471,In_669);
or U868 (N_868,In_481,In_486);
nor U869 (N_869,In_327,In_630);
nor U870 (N_870,In_332,In_579);
and U871 (N_871,In_74,In_911);
nand U872 (N_872,In_987,In_649);
nor U873 (N_873,In_948,In_175);
and U874 (N_874,In_984,In_231);
and U875 (N_875,In_957,In_849);
nand U876 (N_876,In_152,In_420);
nand U877 (N_877,In_272,In_212);
nand U878 (N_878,In_43,In_666);
nor U879 (N_879,In_784,In_214);
and U880 (N_880,In_308,In_905);
nor U881 (N_881,In_264,In_262);
or U882 (N_882,In_16,In_163);
nand U883 (N_883,In_522,In_692);
nor U884 (N_884,In_518,In_158);
nor U885 (N_885,In_749,In_377);
or U886 (N_886,In_438,In_493);
and U887 (N_887,In_367,In_448);
and U888 (N_888,In_249,In_804);
or U889 (N_889,In_808,In_380);
nor U890 (N_890,In_264,In_896);
or U891 (N_891,In_867,In_35);
xnor U892 (N_892,In_323,In_969);
xnor U893 (N_893,In_707,In_490);
xor U894 (N_894,In_555,In_185);
nand U895 (N_895,In_749,In_190);
and U896 (N_896,In_544,In_7);
or U897 (N_897,In_21,In_354);
nand U898 (N_898,In_143,In_623);
nand U899 (N_899,In_543,In_209);
and U900 (N_900,In_444,In_215);
nor U901 (N_901,In_848,In_675);
nor U902 (N_902,In_870,In_319);
nor U903 (N_903,In_676,In_340);
nand U904 (N_904,In_84,In_653);
xnor U905 (N_905,In_221,In_200);
nor U906 (N_906,In_277,In_682);
or U907 (N_907,In_726,In_181);
nand U908 (N_908,In_138,In_680);
xnor U909 (N_909,In_652,In_500);
nor U910 (N_910,In_358,In_817);
nor U911 (N_911,In_175,In_571);
or U912 (N_912,In_462,In_603);
and U913 (N_913,In_405,In_818);
and U914 (N_914,In_565,In_24);
xnor U915 (N_915,In_59,In_435);
or U916 (N_916,In_690,In_150);
nor U917 (N_917,In_712,In_779);
or U918 (N_918,In_125,In_487);
or U919 (N_919,In_235,In_419);
and U920 (N_920,In_622,In_656);
nor U921 (N_921,In_196,In_982);
or U922 (N_922,In_285,In_561);
nor U923 (N_923,In_269,In_844);
or U924 (N_924,In_152,In_907);
nand U925 (N_925,In_529,In_172);
and U926 (N_926,In_560,In_267);
and U927 (N_927,In_364,In_472);
nor U928 (N_928,In_470,In_587);
nor U929 (N_929,In_303,In_154);
or U930 (N_930,In_415,In_225);
nor U931 (N_931,In_138,In_930);
nor U932 (N_932,In_914,In_474);
nand U933 (N_933,In_938,In_871);
xnor U934 (N_934,In_163,In_25);
and U935 (N_935,In_932,In_8);
nor U936 (N_936,In_981,In_306);
nor U937 (N_937,In_919,In_965);
or U938 (N_938,In_618,In_703);
nand U939 (N_939,In_181,In_135);
or U940 (N_940,In_163,In_693);
nand U941 (N_941,In_0,In_288);
nand U942 (N_942,In_733,In_934);
nor U943 (N_943,In_277,In_70);
or U944 (N_944,In_933,In_174);
nand U945 (N_945,In_404,In_744);
nand U946 (N_946,In_456,In_844);
nor U947 (N_947,In_913,In_698);
and U948 (N_948,In_291,In_838);
or U949 (N_949,In_597,In_228);
and U950 (N_950,In_110,In_319);
and U951 (N_951,In_275,In_303);
nor U952 (N_952,In_148,In_628);
and U953 (N_953,In_614,In_804);
or U954 (N_954,In_572,In_464);
or U955 (N_955,In_466,In_667);
nor U956 (N_956,In_567,In_945);
nand U957 (N_957,In_505,In_513);
and U958 (N_958,In_871,In_581);
nand U959 (N_959,In_142,In_710);
or U960 (N_960,In_86,In_571);
xor U961 (N_961,In_764,In_527);
and U962 (N_962,In_776,In_695);
nand U963 (N_963,In_582,In_949);
and U964 (N_964,In_379,In_767);
or U965 (N_965,In_837,In_990);
or U966 (N_966,In_754,In_182);
nor U967 (N_967,In_454,In_927);
and U968 (N_968,In_307,In_155);
nand U969 (N_969,In_818,In_202);
or U970 (N_970,In_964,In_812);
nor U971 (N_971,In_983,In_227);
and U972 (N_972,In_997,In_322);
and U973 (N_973,In_465,In_715);
nand U974 (N_974,In_784,In_14);
nand U975 (N_975,In_44,In_193);
and U976 (N_976,In_446,In_115);
nor U977 (N_977,In_252,In_373);
or U978 (N_978,In_593,In_728);
nor U979 (N_979,In_938,In_13);
xnor U980 (N_980,In_21,In_916);
and U981 (N_981,In_28,In_996);
and U982 (N_982,In_871,In_788);
nor U983 (N_983,In_24,In_736);
and U984 (N_984,In_2,In_938);
nor U985 (N_985,In_318,In_260);
xnor U986 (N_986,In_698,In_126);
and U987 (N_987,In_683,In_707);
and U988 (N_988,In_866,In_233);
xor U989 (N_989,In_418,In_151);
nand U990 (N_990,In_421,In_655);
nand U991 (N_991,In_634,In_40);
nor U992 (N_992,In_545,In_347);
nor U993 (N_993,In_378,In_671);
nor U994 (N_994,In_597,In_594);
xnor U995 (N_995,In_970,In_238);
and U996 (N_996,In_486,In_798);
nor U997 (N_997,In_221,In_445);
and U998 (N_998,In_584,In_177);
and U999 (N_999,In_547,In_808);
xor U1000 (N_1000,N_494,N_727);
xnor U1001 (N_1001,N_760,N_543);
or U1002 (N_1002,N_608,N_163);
and U1003 (N_1003,N_409,N_707);
or U1004 (N_1004,N_769,N_264);
or U1005 (N_1005,N_911,N_174);
or U1006 (N_1006,N_213,N_555);
nand U1007 (N_1007,N_94,N_445);
nor U1008 (N_1008,N_741,N_528);
nor U1009 (N_1009,N_466,N_438);
or U1010 (N_1010,N_255,N_340);
xnor U1011 (N_1011,N_927,N_449);
or U1012 (N_1012,N_522,N_57);
and U1013 (N_1013,N_969,N_617);
nand U1014 (N_1014,N_881,N_566);
nor U1015 (N_1015,N_754,N_38);
nor U1016 (N_1016,N_204,N_259);
xnor U1017 (N_1017,N_496,N_670);
or U1018 (N_1018,N_530,N_159);
nor U1019 (N_1019,N_41,N_498);
nor U1020 (N_1020,N_432,N_840);
nand U1021 (N_1021,N_958,N_776);
xnor U1022 (N_1022,N_730,N_33);
nand U1023 (N_1023,N_268,N_448);
nand U1024 (N_1024,N_74,N_281);
xor U1025 (N_1025,N_913,N_86);
nand U1026 (N_1026,N_215,N_651);
nand U1027 (N_1027,N_362,N_85);
xor U1028 (N_1028,N_361,N_283);
or U1029 (N_1029,N_368,N_737);
or U1030 (N_1030,N_818,N_938);
nand U1031 (N_1031,N_965,N_602);
or U1032 (N_1032,N_747,N_66);
and U1033 (N_1033,N_526,N_887);
or U1034 (N_1034,N_841,N_547);
or U1035 (N_1035,N_946,N_2);
nor U1036 (N_1036,N_604,N_620);
nand U1037 (N_1037,N_400,N_132);
nand U1038 (N_1038,N_549,N_857);
or U1039 (N_1039,N_854,N_676);
xnor U1040 (N_1040,N_332,N_93);
xor U1041 (N_1041,N_369,N_842);
nand U1042 (N_1042,N_856,N_299);
nor U1043 (N_1043,N_349,N_901);
and U1044 (N_1044,N_762,N_492);
nand U1045 (N_1045,N_551,N_247);
and U1046 (N_1046,N_452,N_790);
and U1047 (N_1047,N_487,N_750);
and U1048 (N_1048,N_151,N_673);
nand U1049 (N_1049,N_5,N_387);
nor U1050 (N_1050,N_891,N_815);
or U1051 (N_1051,N_282,N_154);
nor U1052 (N_1052,N_210,N_296);
or U1053 (N_1053,N_457,N_11);
nand U1054 (N_1054,N_874,N_529);
and U1055 (N_1055,N_755,N_257);
and U1056 (N_1056,N_334,N_718);
or U1057 (N_1057,N_469,N_434);
xor U1058 (N_1058,N_675,N_150);
and U1059 (N_1059,N_404,N_574);
and U1060 (N_1060,N_502,N_298);
xnor U1061 (N_1061,N_272,N_258);
nand U1062 (N_1062,N_781,N_644);
or U1063 (N_1063,N_288,N_73);
xnor U1064 (N_1064,N_343,N_793);
and U1065 (N_1065,N_831,N_43);
and U1066 (N_1066,N_293,N_879);
xor U1067 (N_1067,N_801,N_926);
or U1068 (N_1068,N_811,N_626);
nor U1069 (N_1069,N_735,N_906);
and U1070 (N_1070,N_907,N_472);
and U1071 (N_1071,N_714,N_647);
nor U1072 (N_1072,N_637,N_702);
nor U1073 (N_1073,N_389,N_843);
and U1074 (N_1074,N_925,N_55);
nor U1075 (N_1075,N_836,N_796);
and U1076 (N_1076,N_46,N_991);
and U1077 (N_1077,N_511,N_423);
nor U1078 (N_1078,N_351,N_412);
and U1079 (N_1079,N_367,N_286);
or U1080 (N_1080,N_59,N_32);
nand U1081 (N_1081,N_540,N_273);
and U1082 (N_1082,N_768,N_83);
xor U1083 (N_1083,N_375,N_613);
and U1084 (N_1084,N_701,N_194);
or U1085 (N_1085,N_786,N_700);
or U1086 (N_1086,N_648,N_106);
nand U1087 (N_1087,N_200,N_744);
nor U1088 (N_1088,N_669,N_234);
nand U1089 (N_1089,N_847,N_439);
and U1090 (N_1090,N_348,N_309);
or U1091 (N_1091,N_704,N_712);
nand U1092 (N_1092,N_554,N_482);
nand U1093 (N_1093,N_591,N_139);
or U1094 (N_1094,N_437,N_941);
nor U1095 (N_1095,N_483,N_471);
nand U1096 (N_1096,N_695,N_899);
or U1097 (N_1097,N_756,N_201);
nand U1098 (N_1098,N_825,N_81);
xor U1099 (N_1099,N_671,N_516);
nor U1100 (N_1100,N_640,N_870);
or U1101 (N_1101,N_816,N_307);
and U1102 (N_1102,N_238,N_277);
xor U1103 (N_1103,N_972,N_416);
nor U1104 (N_1104,N_377,N_433);
nand U1105 (N_1105,N_632,N_560);
or U1106 (N_1106,N_886,N_500);
or U1107 (N_1107,N_686,N_563);
and U1108 (N_1108,N_582,N_183);
and U1109 (N_1109,N_82,N_550);
nor U1110 (N_1110,N_719,N_198);
or U1111 (N_1111,N_365,N_544);
nor U1112 (N_1112,N_845,N_758);
nand U1113 (N_1113,N_14,N_628);
nand U1114 (N_1114,N_725,N_752);
nor U1115 (N_1115,N_363,N_239);
and U1116 (N_1116,N_7,N_493);
nand U1117 (N_1117,N_785,N_65);
nor U1118 (N_1118,N_230,N_397);
and U1119 (N_1119,N_723,N_173);
and U1120 (N_1120,N_470,N_577);
and U1121 (N_1121,N_28,N_948);
and U1122 (N_1122,N_520,N_778);
or U1123 (N_1123,N_146,N_622);
nor U1124 (N_1124,N_917,N_128);
xnor U1125 (N_1125,N_13,N_848);
nand U1126 (N_1126,N_40,N_625);
nand U1127 (N_1127,N_463,N_844);
nand U1128 (N_1128,N_42,N_971);
or U1129 (N_1129,N_592,N_101);
nand U1130 (N_1130,N_383,N_461);
and U1131 (N_1131,N_152,N_681);
or U1132 (N_1132,N_133,N_656);
nand U1133 (N_1133,N_692,N_325);
xnor U1134 (N_1134,N_262,N_54);
nand U1135 (N_1135,N_192,N_571);
xor U1136 (N_1136,N_413,N_237);
nand U1137 (N_1137,N_871,N_980);
nand U1138 (N_1138,N_666,N_863);
or U1139 (N_1139,N_484,N_63);
xor U1140 (N_1140,N_175,N_889);
nand U1141 (N_1141,N_379,N_552);
and U1142 (N_1142,N_524,N_638);
or U1143 (N_1143,N_978,N_578);
or U1144 (N_1144,N_398,N_372);
xnor U1145 (N_1145,N_355,N_267);
and U1146 (N_1146,N_422,N_459);
xnor U1147 (N_1147,N_19,N_519);
or U1148 (N_1148,N_318,N_542);
nor U1149 (N_1149,N_885,N_214);
nor U1150 (N_1150,N_820,N_580);
nor U1151 (N_1151,N_224,N_548);
or U1152 (N_1152,N_127,N_961);
or U1153 (N_1153,N_557,N_491);
or U1154 (N_1154,N_505,N_269);
nor U1155 (N_1155,N_664,N_629);
xnor U1156 (N_1156,N_882,N_593);
nor U1157 (N_1157,N_738,N_960);
or U1158 (N_1158,N_77,N_4);
and U1159 (N_1159,N_957,N_301);
nor U1160 (N_1160,N_933,N_266);
or U1161 (N_1161,N_35,N_849);
nand U1162 (N_1162,N_350,N_833);
nand U1163 (N_1163,N_428,N_3);
nor U1164 (N_1164,N_444,N_804);
and U1165 (N_1165,N_187,N_859);
nor U1166 (N_1166,N_410,N_561);
or U1167 (N_1167,N_34,N_805);
or U1168 (N_1168,N_535,N_248);
nand U1169 (N_1169,N_431,N_462);
and U1170 (N_1170,N_323,N_953);
or U1171 (N_1171,N_691,N_109);
xnor U1172 (N_1172,N_211,N_839);
and U1173 (N_1173,N_601,N_921);
or U1174 (N_1174,N_373,N_244);
or U1175 (N_1175,N_955,N_188);
nand U1176 (N_1176,N_536,N_830);
and U1177 (N_1177,N_382,N_27);
nor U1178 (N_1178,N_759,N_420);
nor U1179 (N_1179,N_576,N_655);
nand U1180 (N_1180,N_274,N_895);
nor U1181 (N_1181,N_905,N_876);
nand U1182 (N_1182,N_386,N_618);
nor U1183 (N_1183,N_260,N_419);
and U1184 (N_1184,N_384,N_556);
and U1185 (N_1185,N_757,N_477);
xor U1186 (N_1186,N_641,N_104);
nor U1187 (N_1187,N_517,N_454);
or U1188 (N_1188,N_185,N_436);
and U1189 (N_1189,N_120,N_374);
nor U1190 (N_1190,N_732,N_303);
nor U1191 (N_1191,N_986,N_335);
nor U1192 (N_1192,N_407,N_533);
nor U1193 (N_1193,N_440,N_391);
nand U1194 (N_1194,N_84,N_18);
nor U1195 (N_1195,N_406,N_162);
or U1196 (N_1196,N_142,N_645);
or U1197 (N_1197,N_996,N_562);
nand U1198 (N_1198,N_590,N_709);
or U1199 (N_1199,N_579,N_983);
xor U1200 (N_1200,N_292,N_15);
nor U1201 (N_1201,N_534,N_869);
or U1202 (N_1202,N_165,N_791);
nand U1203 (N_1203,N_376,N_861);
and U1204 (N_1204,N_568,N_855);
nor U1205 (N_1205,N_521,N_792);
nand U1206 (N_1206,N_287,N_541);
and U1207 (N_1207,N_923,N_306);
nor U1208 (N_1208,N_963,N_388);
nand U1209 (N_1209,N_71,N_64);
and U1210 (N_1210,N_635,N_261);
nor U1211 (N_1211,N_821,N_974);
and U1212 (N_1212,N_121,N_356);
nand U1213 (N_1213,N_231,N_212);
and U1214 (N_1214,N_789,N_324);
and U1215 (N_1215,N_100,N_873);
xor U1216 (N_1216,N_240,N_176);
nand U1217 (N_1217,N_249,N_17);
xnor U1218 (N_1218,N_243,N_161);
or U1219 (N_1219,N_353,N_624);
or U1220 (N_1220,N_606,N_97);
nand U1221 (N_1221,N_250,N_179);
or U1222 (N_1222,N_587,N_581);
or U1223 (N_1223,N_837,N_39);
nand U1224 (N_1224,N_572,N_236);
or U1225 (N_1225,N_987,N_456);
nand U1226 (N_1226,N_902,N_490);
xnor U1227 (N_1227,N_583,N_141);
nand U1228 (N_1228,N_25,N_443);
nand U1229 (N_1229,N_88,N_924);
and U1230 (N_1230,N_614,N_393);
nor U1231 (N_1231,N_21,N_26);
nand U1232 (N_1232,N_171,N_317);
and U1233 (N_1233,N_829,N_979);
and U1234 (N_1234,N_321,N_326);
nand U1235 (N_1235,N_51,N_415);
nor U1236 (N_1236,N_114,N_525);
nor U1237 (N_1237,N_951,N_310);
nand U1238 (N_1238,N_631,N_867);
and U1239 (N_1239,N_252,N_619);
or U1240 (N_1240,N_731,N_890);
xor U1241 (N_1241,N_235,N_126);
or U1242 (N_1242,N_285,N_743);
xor U1243 (N_1243,N_233,N_610);
or U1244 (N_1244,N_850,N_144);
and U1245 (N_1245,N_706,N_228);
or U1246 (N_1246,N_812,N_220);
or U1247 (N_1247,N_337,N_347);
or U1248 (N_1248,N_797,N_392);
and U1249 (N_1249,N_425,N_649);
nor U1250 (N_1250,N_575,N_328);
nand U1251 (N_1251,N_265,N_111);
and U1252 (N_1252,N_254,N_729);
xor U1253 (N_1253,N_746,N_75);
or U1254 (N_1254,N_209,N_105);
nor U1255 (N_1255,N_358,N_123);
and U1256 (N_1256,N_131,N_92);
and U1257 (N_1257,N_742,N_880);
xor U1258 (N_1258,N_91,N_596);
and U1259 (N_1259,N_920,N_807);
and U1260 (N_1260,N_689,N_380);
nor U1261 (N_1261,N_232,N_672);
and U1262 (N_1262,N_460,N_817);
nand U1263 (N_1263,N_80,N_12);
or U1264 (N_1264,N_767,N_865);
or U1265 (N_1265,N_822,N_523);
or U1266 (N_1266,N_799,N_512);
nor U1267 (N_1267,N_202,N_253);
nor U1268 (N_1268,N_458,N_984);
nand U1269 (N_1269,N_206,N_605);
nor U1270 (N_1270,N_166,N_115);
or U1271 (N_1271,N_720,N_788);
xnor U1272 (N_1272,N_745,N_771);
and U1273 (N_1273,N_682,N_118);
and U1274 (N_1274,N_98,N_584);
nand U1275 (N_1275,N_748,N_721);
nor U1276 (N_1276,N_450,N_506);
xor U1277 (N_1277,N_573,N_129);
xor U1278 (N_1278,N_772,N_661);
and U1279 (N_1279,N_952,N_276);
or U1280 (N_1280,N_931,N_795);
nor U1281 (N_1281,N_783,N_609);
and U1282 (N_1282,N_878,N_975);
or U1283 (N_1283,N_813,N_476);
nand U1284 (N_1284,N_339,N_251);
nand U1285 (N_1285,N_360,N_87);
nand U1286 (N_1286,N_193,N_79);
and U1287 (N_1287,N_153,N_241);
or U1288 (N_1288,N_338,N_346);
or U1289 (N_1289,N_381,N_207);
nor U1290 (N_1290,N_678,N_780);
nor U1291 (N_1291,N_916,N_60);
nand U1292 (N_1292,N_950,N_611);
nor U1293 (N_1293,N_455,N_47);
nor U1294 (N_1294,N_177,N_595);
nor U1295 (N_1295,N_954,N_710);
or U1296 (N_1296,N_515,N_160);
xnor U1297 (N_1297,N_403,N_538);
nand U1298 (N_1298,N_167,N_623);
and U1299 (N_1299,N_504,N_62);
nand U1300 (N_1300,N_427,N_693);
and U1301 (N_1301,N_95,N_134);
nand U1302 (N_1302,N_553,N_909);
nor U1303 (N_1303,N_956,N_819);
xnor U1304 (N_1304,N_157,N_749);
nand U1305 (N_1305,N_872,N_915);
nor U1306 (N_1306,N_586,N_826);
or U1307 (N_1307,N_72,N_378);
and U1308 (N_1308,N_997,N_802);
nand U1309 (N_1309,N_914,N_56);
nor U1310 (N_1310,N_302,N_344);
and U1311 (N_1311,N_329,N_195);
and U1312 (N_1312,N_30,N_703);
nand U1313 (N_1313,N_513,N_858);
xnor U1314 (N_1314,N_441,N_140);
and U1315 (N_1315,N_156,N_1);
nor U1316 (N_1316,N_823,N_945);
nand U1317 (N_1317,N_942,N_774);
xor U1318 (N_1318,N_734,N_654);
xnor U1319 (N_1319,N_447,N_999);
xnor U1320 (N_1320,N_119,N_0);
nor U1321 (N_1321,N_846,N_218);
nand U1322 (N_1322,N_475,N_627);
nand U1323 (N_1323,N_932,N_765);
nor U1324 (N_1324,N_782,N_994);
or U1325 (N_1325,N_621,N_489);
xor U1326 (N_1326,N_495,N_169);
or U1327 (N_1327,N_117,N_108);
nor U1328 (N_1328,N_168,N_37);
or U1329 (N_1329,N_103,N_6);
nand U1330 (N_1330,N_316,N_898);
and U1331 (N_1331,N_53,N_229);
nor U1332 (N_1332,N_478,N_429);
nand U1333 (N_1333,N_770,N_465);
nor U1334 (N_1334,N_507,N_943);
nand U1335 (N_1335,N_677,N_158);
nor U1336 (N_1336,N_311,N_565);
and U1337 (N_1337,N_935,N_834);
and U1338 (N_1338,N_155,N_658);
and U1339 (N_1339,N_866,N_514);
nand U1340 (N_1340,N_308,N_336);
nor U1341 (N_1341,N_903,N_989);
nor U1342 (N_1342,N_205,N_45);
and U1343 (N_1343,N_705,N_52);
and U1344 (N_1344,N_527,N_145);
or U1345 (N_1345,N_68,N_683);
nor U1346 (N_1346,N_739,N_149);
xnor U1347 (N_1347,N_982,N_148);
xor U1348 (N_1348,N_208,N_616);
nor U1349 (N_1349,N_981,N_451);
or U1350 (N_1350,N_518,N_680);
or U1351 (N_1351,N_467,N_305);
and U1352 (N_1352,N_688,N_589);
and U1353 (N_1353,N_357,N_246);
nor U1354 (N_1354,N_877,N_196);
nor U1355 (N_1355,N_414,N_401);
or U1356 (N_1356,N_221,N_814);
or U1357 (N_1357,N_354,N_314);
and U1358 (N_1358,N_832,N_643);
or U1359 (N_1359,N_853,N_291);
or U1360 (N_1360,N_135,N_99);
nor U1361 (N_1361,N_480,N_947);
nor U1362 (N_1362,N_147,N_189);
nand U1363 (N_1363,N_223,N_190);
nor U1364 (N_1364,N_278,N_904);
and U1365 (N_1365,N_405,N_696);
and U1366 (N_1366,N_499,N_949);
nor U1367 (N_1367,N_684,N_722);
nor U1368 (N_1368,N_399,N_182);
nor U1369 (N_1369,N_304,N_934);
nor U1370 (N_1370,N_539,N_559);
or U1371 (N_1371,N_426,N_531);
nor U1372 (N_1372,N_970,N_411);
or U1373 (N_1373,N_275,N_69);
or U1374 (N_1374,N_418,N_612);
and U1375 (N_1375,N_508,N_23);
xor U1376 (N_1376,N_537,N_313);
and U1377 (N_1377,N_633,N_24);
and U1378 (N_1378,N_180,N_315);
or U1379 (N_1379,N_884,N_300);
nor U1380 (N_1380,N_646,N_203);
or U1381 (N_1381,N_888,N_509);
nor U1382 (N_1382,N_713,N_690);
nor U1383 (N_1383,N_922,N_191);
or U1384 (N_1384,N_396,N_715);
and U1385 (N_1385,N_588,N_78);
nor U1386 (N_1386,N_798,N_468);
or U1387 (N_1387,N_615,N_9);
or U1388 (N_1388,N_775,N_779);
nand U1389 (N_1389,N_10,N_665);
or U1390 (N_1390,N_256,N_851);
nand U1391 (N_1391,N_36,N_421);
or U1392 (N_1392,N_137,N_402);
nor U1393 (N_1393,N_116,N_16);
or U1394 (N_1394,N_453,N_44);
and U1395 (N_1395,N_564,N_122);
and U1396 (N_1396,N_226,N_96);
nand U1397 (N_1397,N_630,N_985);
or U1398 (N_1398,N_50,N_810);
nand U1399 (N_1399,N_89,N_394);
nor U1400 (N_1400,N_312,N_22);
xnor U1401 (N_1401,N_634,N_322);
and U1402 (N_1402,N_928,N_446);
xnor U1403 (N_1403,N_352,N_61);
or U1404 (N_1404,N_966,N_501);
nor U1405 (N_1405,N_359,N_716);
nor U1406 (N_1406,N_178,N_333);
nor U1407 (N_1407,N_371,N_603);
and U1408 (N_1408,N_652,N_875);
and U1409 (N_1409,N_919,N_138);
nand U1410 (N_1410,N_699,N_184);
nor U1411 (N_1411,N_740,N_320);
nor U1412 (N_1412,N_893,N_967);
and U1413 (N_1413,N_199,N_319);
or U1414 (N_1414,N_284,N_297);
nand U1415 (N_1415,N_959,N_216);
nand U1416 (N_1416,N_977,N_107);
or U1417 (N_1417,N_327,N_864);
xnor U1418 (N_1418,N_708,N_599);
and U1419 (N_1419,N_366,N_990);
and U1420 (N_1420,N_76,N_70);
nand U1421 (N_1421,N_607,N_242);
and U1422 (N_1422,N_170,N_939);
nand U1423 (N_1423,N_497,N_733);
and U1424 (N_1424,N_197,N_835);
nand U1425 (N_1425,N_892,N_569);
nor U1426 (N_1426,N_806,N_912);
nor U1427 (N_1427,N_546,N_964);
nand U1428 (N_1428,N_58,N_636);
or U1429 (N_1429,N_809,N_222);
nor U1430 (N_1430,N_639,N_364);
nor U1431 (N_1431,N_998,N_385);
nand U1432 (N_1432,N_827,N_289);
nand U1433 (N_1433,N_558,N_164);
and U1434 (N_1434,N_31,N_976);
and U1435 (N_1435,N_667,N_330);
nor U1436 (N_1436,N_736,N_345);
nor U1437 (N_1437,N_883,N_130);
nor U1438 (N_1438,N_724,N_594);
and U1439 (N_1439,N_486,N_424);
nand U1440 (N_1440,N_761,N_408);
and U1441 (N_1441,N_124,N_763);
and U1442 (N_1442,N_918,N_8);
nor U1443 (N_1443,N_280,N_937);
nor U1444 (N_1444,N_217,N_824);
nor U1445 (N_1445,N_936,N_993);
nand U1446 (N_1446,N_598,N_481);
and U1447 (N_1447,N_112,N_270);
xnor U1448 (N_1448,N_642,N_473);
or U1449 (N_1449,N_331,N_181);
xnor U1450 (N_1450,N_464,N_766);
and U1451 (N_1451,N_442,N_370);
and U1452 (N_1452,N_479,N_838);
or U1453 (N_1453,N_787,N_794);
and U1454 (N_1454,N_227,N_697);
nor U1455 (N_1455,N_662,N_125);
nand U1456 (N_1456,N_668,N_245);
or U1457 (N_1457,N_929,N_717);
nor U1458 (N_1458,N_910,N_659);
xor U1459 (N_1459,N_510,N_532);
or U1460 (N_1460,N_435,N_726);
and U1461 (N_1461,N_488,N_940);
nand U1462 (N_1462,N_49,N_570);
or U1463 (N_1463,N_992,N_90);
nor U1464 (N_1464,N_172,N_279);
xor U1465 (N_1465,N_687,N_597);
or U1466 (N_1466,N_930,N_862);
or U1467 (N_1467,N_110,N_962);
and U1468 (N_1468,N_263,N_968);
or U1469 (N_1469,N_868,N_784);
nor U1470 (N_1470,N_600,N_474);
xnor U1471 (N_1471,N_711,N_660);
or U1472 (N_1472,N_67,N_897);
nand U1473 (N_1473,N_225,N_503);
nand U1474 (N_1474,N_585,N_653);
nand U1475 (N_1475,N_29,N_545);
nor U1476 (N_1476,N_808,N_674);
or U1477 (N_1477,N_290,N_698);
or U1478 (N_1478,N_113,N_852);
xnor U1479 (N_1479,N_567,N_764);
or U1480 (N_1480,N_485,N_143);
or U1481 (N_1481,N_430,N_417);
and U1482 (N_1482,N_186,N_136);
nand U1483 (N_1483,N_753,N_803);
and U1484 (N_1484,N_341,N_908);
nor U1485 (N_1485,N_48,N_390);
or U1486 (N_1486,N_860,N_679);
nand U1487 (N_1487,N_342,N_900);
or U1488 (N_1488,N_828,N_751);
or U1489 (N_1489,N_973,N_295);
nor U1490 (N_1490,N_894,N_657);
nor U1491 (N_1491,N_102,N_685);
or U1492 (N_1492,N_663,N_896);
nand U1493 (N_1493,N_773,N_694);
nand U1494 (N_1494,N_995,N_728);
nor U1495 (N_1495,N_800,N_294);
nand U1496 (N_1496,N_944,N_271);
nand U1497 (N_1497,N_219,N_20);
and U1498 (N_1498,N_777,N_395);
or U1499 (N_1499,N_988,N_650);
nor U1500 (N_1500,N_604,N_707);
or U1501 (N_1501,N_258,N_427);
and U1502 (N_1502,N_923,N_187);
or U1503 (N_1503,N_798,N_655);
xor U1504 (N_1504,N_393,N_691);
or U1505 (N_1505,N_689,N_783);
and U1506 (N_1506,N_78,N_969);
and U1507 (N_1507,N_469,N_477);
and U1508 (N_1508,N_571,N_499);
and U1509 (N_1509,N_944,N_390);
xnor U1510 (N_1510,N_367,N_784);
nor U1511 (N_1511,N_965,N_912);
nor U1512 (N_1512,N_677,N_362);
nor U1513 (N_1513,N_336,N_245);
nand U1514 (N_1514,N_2,N_148);
nand U1515 (N_1515,N_524,N_342);
nor U1516 (N_1516,N_230,N_446);
nand U1517 (N_1517,N_730,N_149);
or U1518 (N_1518,N_411,N_29);
nand U1519 (N_1519,N_879,N_85);
nor U1520 (N_1520,N_509,N_400);
nand U1521 (N_1521,N_620,N_572);
xor U1522 (N_1522,N_742,N_604);
and U1523 (N_1523,N_744,N_359);
or U1524 (N_1524,N_610,N_342);
nor U1525 (N_1525,N_414,N_87);
or U1526 (N_1526,N_905,N_746);
nor U1527 (N_1527,N_511,N_778);
nand U1528 (N_1528,N_940,N_818);
xnor U1529 (N_1529,N_486,N_161);
nand U1530 (N_1530,N_530,N_136);
nor U1531 (N_1531,N_261,N_55);
nor U1532 (N_1532,N_23,N_748);
xor U1533 (N_1533,N_223,N_841);
or U1534 (N_1534,N_964,N_775);
nor U1535 (N_1535,N_625,N_493);
and U1536 (N_1536,N_86,N_869);
or U1537 (N_1537,N_162,N_337);
nor U1538 (N_1538,N_858,N_668);
nand U1539 (N_1539,N_500,N_20);
and U1540 (N_1540,N_455,N_557);
and U1541 (N_1541,N_536,N_139);
or U1542 (N_1542,N_322,N_757);
and U1543 (N_1543,N_432,N_169);
nor U1544 (N_1544,N_881,N_701);
and U1545 (N_1545,N_737,N_674);
or U1546 (N_1546,N_720,N_273);
xor U1547 (N_1547,N_824,N_225);
xor U1548 (N_1548,N_481,N_639);
nand U1549 (N_1549,N_466,N_208);
xor U1550 (N_1550,N_638,N_420);
or U1551 (N_1551,N_437,N_470);
nor U1552 (N_1552,N_712,N_367);
and U1553 (N_1553,N_405,N_524);
or U1554 (N_1554,N_516,N_605);
nor U1555 (N_1555,N_501,N_213);
xnor U1556 (N_1556,N_235,N_911);
and U1557 (N_1557,N_633,N_506);
xor U1558 (N_1558,N_21,N_875);
xor U1559 (N_1559,N_34,N_582);
nand U1560 (N_1560,N_676,N_639);
nor U1561 (N_1561,N_954,N_591);
xnor U1562 (N_1562,N_430,N_83);
and U1563 (N_1563,N_39,N_949);
or U1564 (N_1564,N_464,N_427);
and U1565 (N_1565,N_806,N_342);
nor U1566 (N_1566,N_849,N_959);
nor U1567 (N_1567,N_515,N_357);
nor U1568 (N_1568,N_222,N_623);
and U1569 (N_1569,N_672,N_395);
or U1570 (N_1570,N_792,N_632);
xor U1571 (N_1571,N_170,N_259);
or U1572 (N_1572,N_617,N_346);
xor U1573 (N_1573,N_429,N_593);
or U1574 (N_1574,N_360,N_129);
or U1575 (N_1575,N_371,N_562);
and U1576 (N_1576,N_319,N_758);
and U1577 (N_1577,N_974,N_211);
and U1578 (N_1578,N_783,N_711);
or U1579 (N_1579,N_913,N_659);
or U1580 (N_1580,N_411,N_258);
and U1581 (N_1581,N_540,N_740);
nor U1582 (N_1582,N_587,N_718);
or U1583 (N_1583,N_372,N_212);
nor U1584 (N_1584,N_355,N_12);
or U1585 (N_1585,N_774,N_512);
and U1586 (N_1586,N_917,N_151);
or U1587 (N_1587,N_970,N_883);
nand U1588 (N_1588,N_590,N_267);
and U1589 (N_1589,N_271,N_354);
nand U1590 (N_1590,N_53,N_805);
nor U1591 (N_1591,N_879,N_993);
nor U1592 (N_1592,N_352,N_464);
or U1593 (N_1593,N_571,N_924);
and U1594 (N_1594,N_660,N_283);
and U1595 (N_1595,N_649,N_633);
nor U1596 (N_1596,N_539,N_657);
or U1597 (N_1597,N_306,N_998);
nor U1598 (N_1598,N_678,N_307);
nand U1599 (N_1599,N_445,N_574);
or U1600 (N_1600,N_986,N_313);
or U1601 (N_1601,N_595,N_118);
xor U1602 (N_1602,N_128,N_109);
xor U1603 (N_1603,N_220,N_498);
nand U1604 (N_1604,N_281,N_784);
nor U1605 (N_1605,N_229,N_797);
nand U1606 (N_1606,N_801,N_825);
nand U1607 (N_1607,N_329,N_63);
xnor U1608 (N_1608,N_128,N_875);
nor U1609 (N_1609,N_430,N_293);
nand U1610 (N_1610,N_489,N_385);
and U1611 (N_1611,N_383,N_982);
or U1612 (N_1612,N_941,N_83);
or U1613 (N_1613,N_459,N_538);
and U1614 (N_1614,N_949,N_483);
and U1615 (N_1615,N_891,N_747);
nand U1616 (N_1616,N_13,N_212);
and U1617 (N_1617,N_697,N_899);
nand U1618 (N_1618,N_537,N_123);
nor U1619 (N_1619,N_975,N_317);
nand U1620 (N_1620,N_430,N_136);
or U1621 (N_1621,N_39,N_598);
nand U1622 (N_1622,N_190,N_787);
or U1623 (N_1623,N_669,N_755);
xor U1624 (N_1624,N_347,N_869);
or U1625 (N_1625,N_809,N_310);
and U1626 (N_1626,N_598,N_992);
nor U1627 (N_1627,N_585,N_734);
nor U1628 (N_1628,N_669,N_70);
and U1629 (N_1629,N_791,N_663);
nand U1630 (N_1630,N_426,N_548);
and U1631 (N_1631,N_583,N_408);
or U1632 (N_1632,N_785,N_346);
xnor U1633 (N_1633,N_294,N_657);
xnor U1634 (N_1634,N_289,N_67);
and U1635 (N_1635,N_9,N_603);
or U1636 (N_1636,N_154,N_327);
nor U1637 (N_1637,N_583,N_451);
nor U1638 (N_1638,N_892,N_879);
or U1639 (N_1639,N_808,N_910);
or U1640 (N_1640,N_550,N_145);
nor U1641 (N_1641,N_595,N_915);
and U1642 (N_1642,N_908,N_275);
or U1643 (N_1643,N_992,N_873);
nor U1644 (N_1644,N_289,N_799);
nand U1645 (N_1645,N_641,N_725);
or U1646 (N_1646,N_20,N_856);
nor U1647 (N_1647,N_9,N_654);
or U1648 (N_1648,N_851,N_846);
nor U1649 (N_1649,N_332,N_152);
or U1650 (N_1650,N_642,N_916);
or U1651 (N_1651,N_235,N_680);
and U1652 (N_1652,N_300,N_943);
nor U1653 (N_1653,N_295,N_261);
nand U1654 (N_1654,N_398,N_445);
xor U1655 (N_1655,N_780,N_803);
xnor U1656 (N_1656,N_61,N_733);
and U1657 (N_1657,N_470,N_262);
nand U1658 (N_1658,N_93,N_458);
xor U1659 (N_1659,N_630,N_753);
nor U1660 (N_1660,N_389,N_926);
and U1661 (N_1661,N_354,N_903);
xor U1662 (N_1662,N_256,N_142);
and U1663 (N_1663,N_939,N_13);
or U1664 (N_1664,N_225,N_384);
or U1665 (N_1665,N_5,N_285);
xnor U1666 (N_1666,N_493,N_803);
nor U1667 (N_1667,N_728,N_472);
and U1668 (N_1668,N_502,N_147);
and U1669 (N_1669,N_281,N_345);
nor U1670 (N_1670,N_949,N_712);
and U1671 (N_1671,N_504,N_373);
or U1672 (N_1672,N_371,N_415);
nor U1673 (N_1673,N_363,N_880);
nor U1674 (N_1674,N_953,N_311);
xnor U1675 (N_1675,N_990,N_57);
and U1676 (N_1676,N_896,N_538);
and U1677 (N_1677,N_571,N_481);
nand U1678 (N_1678,N_498,N_137);
nand U1679 (N_1679,N_902,N_657);
nand U1680 (N_1680,N_40,N_525);
nor U1681 (N_1681,N_762,N_291);
or U1682 (N_1682,N_495,N_744);
nor U1683 (N_1683,N_173,N_836);
and U1684 (N_1684,N_187,N_939);
and U1685 (N_1685,N_104,N_676);
nand U1686 (N_1686,N_909,N_659);
or U1687 (N_1687,N_626,N_613);
and U1688 (N_1688,N_533,N_357);
nor U1689 (N_1689,N_165,N_964);
and U1690 (N_1690,N_136,N_533);
or U1691 (N_1691,N_234,N_395);
or U1692 (N_1692,N_635,N_480);
nand U1693 (N_1693,N_101,N_636);
or U1694 (N_1694,N_881,N_27);
nand U1695 (N_1695,N_509,N_826);
and U1696 (N_1696,N_769,N_40);
xnor U1697 (N_1697,N_598,N_22);
nand U1698 (N_1698,N_770,N_995);
and U1699 (N_1699,N_166,N_905);
nand U1700 (N_1700,N_73,N_637);
nand U1701 (N_1701,N_371,N_38);
and U1702 (N_1702,N_683,N_832);
and U1703 (N_1703,N_526,N_858);
and U1704 (N_1704,N_198,N_194);
and U1705 (N_1705,N_288,N_341);
or U1706 (N_1706,N_396,N_515);
and U1707 (N_1707,N_955,N_215);
nand U1708 (N_1708,N_898,N_740);
or U1709 (N_1709,N_417,N_285);
nand U1710 (N_1710,N_95,N_84);
or U1711 (N_1711,N_683,N_945);
or U1712 (N_1712,N_41,N_913);
nand U1713 (N_1713,N_388,N_20);
nor U1714 (N_1714,N_14,N_685);
nand U1715 (N_1715,N_550,N_468);
and U1716 (N_1716,N_447,N_915);
nand U1717 (N_1717,N_676,N_828);
nand U1718 (N_1718,N_552,N_194);
nand U1719 (N_1719,N_49,N_974);
nand U1720 (N_1720,N_997,N_46);
and U1721 (N_1721,N_539,N_595);
and U1722 (N_1722,N_341,N_239);
and U1723 (N_1723,N_514,N_280);
nand U1724 (N_1724,N_563,N_411);
and U1725 (N_1725,N_822,N_418);
and U1726 (N_1726,N_358,N_650);
or U1727 (N_1727,N_713,N_191);
or U1728 (N_1728,N_997,N_421);
nand U1729 (N_1729,N_523,N_693);
and U1730 (N_1730,N_217,N_233);
nand U1731 (N_1731,N_873,N_411);
or U1732 (N_1732,N_776,N_828);
nor U1733 (N_1733,N_387,N_235);
xnor U1734 (N_1734,N_974,N_884);
nand U1735 (N_1735,N_765,N_632);
or U1736 (N_1736,N_891,N_657);
nand U1737 (N_1737,N_668,N_44);
nor U1738 (N_1738,N_633,N_469);
and U1739 (N_1739,N_152,N_895);
and U1740 (N_1740,N_859,N_908);
or U1741 (N_1741,N_948,N_317);
nor U1742 (N_1742,N_966,N_646);
or U1743 (N_1743,N_950,N_6);
or U1744 (N_1744,N_460,N_596);
nand U1745 (N_1745,N_695,N_209);
or U1746 (N_1746,N_804,N_725);
and U1747 (N_1747,N_147,N_658);
xor U1748 (N_1748,N_487,N_174);
nor U1749 (N_1749,N_750,N_21);
or U1750 (N_1750,N_186,N_421);
and U1751 (N_1751,N_453,N_501);
nor U1752 (N_1752,N_405,N_185);
or U1753 (N_1753,N_62,N_728);
nand U1754 (N_1754,N_804,N_216);
and U1755 (N_1755,N_160,N_653);
or U1756 (N_1756,N_650,N_206);
xnor U1757 (N_1757,N_668,N_100);
nor U1758 (N_1758,N_26,N_391);
nand U1759 (N_1759,N_507,N_885);
or U1760 (N_1760,N_9,N_349);
nor U1761 (N_1761,N_530,N_535);
nor U1762 (N_1762,N_359,N_198);
or U1763 (N_1763,N_780,N_533);
nor U1764 (N_1764,N_340,N_903);
nor U1765 (N_1765,N_997,N_586);
nor U1766 (N_1766,N_892,N_221);
or U1767 (N_1767,N_285,N_449);
nor U1768 (N_1768,N_627,N_455);
xor U1769 (N_1769,N_885,N_207);
xor U1770 (N_1770,N_256,N_958);
nor U1771 (N_1771,N_9,N_655);
nand U1772 (N_1772,N_947,N_74);
xor U1773 (N_1773,N_606,N_527);
nand U1774 (N_1774,N_553,N_123);
nor U1775 (N_1775,N_291,N_509);
nand U1776 (N_1776,N_751,N_645);
nor U1777 (N_1777,N_418,N_235);
or U1778 (N_1778,N_516,N_142);
nand U1779 (N_1779,N_844,N_87);
nand U1780 (N_1780,N_392,N_319);
xnor U1781 (N_1781,N_385,N_517);
xor U1782 (N_1782,N_623,N_248);
nor U1783 (N_1783,N_908,N_621);
nand U1784 (N_1784,N_839,N_768);
and U1785 (N_1785,N_964,N_606);
and U1786 (N_1786,N_580,N_581);
and U1787 (N_1787,N_54,N_991);
and U1788 (N_1788,N_156,N_851);
and U1789 (N_1789,N_35,N_754);
or U1790 (N_1790,N_81,N_777);
or U1791 (N_1791,N_968,N_789);
or U1792 (N_1792,N_922,N_706);
or U1793 (N_1793,N_772,N_129);
nand U1794 (N_1794,N_599,N_150);
and U1795 (N_1795,N_275,N_634);
nor U1796 (N_1796,N_114,N_911);
nand U1797 (N_1797,N_509,N_307);
nand U1798 (N_1798,N_298,N_177);
or U1799 (N_1799,N_534,N_491);
or U1800 (N_1800,N_228,N_563);
or U1801 (N_1801,N_912,N_777);
xnor U1802 (N_1802,N_325,N_436);
or U1803 (N_1803,N_936,N_995);
or U1804 (N_1804,N_547,N_117);
nand U1805 (N_1805,N_981,N_8);
nand U1806 (N_1806,N_313,N_586);
nand U1807 (N_1807,N_664,N_693);
and U1808 (N_1808,N_104,N_583);
nor U1809 (N_1809,N_290,N_804);
nor U1810 (N_1810,N_970,N_45);
nand U1811 (N_1811,N_222,N_151);
xnor U1812 (N_1812,N_820,N_19);
nand U1813 (N_1813,N_302,N_455);
nand U1814 (N_1814,N_258,N_681);
or U1815 (N_1815,N_229,N_143);
nand U1816 (N_1816,N_536,N_194);
and U1817 (N_1817,N_55,N_612);
xnor U1818 (N_1818,N_34,N_851);
nand U1819 (N_1819,N_683,N_328);
nand U1820 (N_1820,N_764,N_858);
nand U1821 (N_1821,N_589,N_912);
and U1822 (N_1822,N_673,N_38);
xnor U1823 (N_1823,N_355,N_813);
nor U1824 (N_1824,N_660,N_648);
nand U1825 (N_1825,N_162,N_499);
xor U1826 (N_1826,N_917,N_473);
nor U1827 (N_1827,N_2,N_217);
and U1828 (N_1828,N_737,N_890);
and U1829 (N_1829,N_476,N_443);
and U1830 (N_1830,N_661,N_913);
and U1831 (N_1831,N_532,N_727);
or U1832 (N_1832,N_135,N_837);
and U1833 (N_1833,N_93,N_911);
nor U1834 (N_1834,N_611,N_585);
or U1835 (N_1835,N_133,N_721);
nor U1836 (N_1836,N_946,N_653);
nor U1837 (N_1837,N_982,N_673);
nand U1838 (N_1838,N_401,N_830);
or U1839 (N_1839,N_633,N_146);
nor U1840 (N_1840,N_180,N_935);
nand U1841 (N_1841,N_155,N_271);
nor U1842 (N_1842,N_326,N_873);
or U1843 (N_1843,N_212,N_603);
nor U1844 (N_1844,N_427,N_492);
xnor U1845 (N_1845,N_929,N_66);
xnor U1846 (N_1846,N_787,N_392);
or U1847 (N_1847,N_922,N_138);
or U1848 (N_1848,N_129,N_454);
or U1849 (N_1849,N_22,N_311);
nor U1850 (N_1850,N_54,N_924);
nand U1851 (N_1851,N_955,N_878);
and U1852 (N_1852,N_977,N_0);
nor U1853 (N_1853,N_750,N_604);
or U1854 (N_1854,N_732,N_215);
nand U1855 (N_1855,N_298,N_956);
nand U1856 (N_1856,N_226,N_607);
xnor U1857 (N_1857,N_126,N_151);
and U1858 (N_1858,N_954,N_231);
nand U1859 (N_1859,N_663,N_364);
and U1860 (N_1860,N_583,N_849);
nand U1861 (N_1861,N_83,N_668);
xor U1862 (N_1862,N_362,N_114);
and U1863 (N_1863,N_751,N_695);
or U1864 (N_1864,N_619,N_327);
and U1865 (N_1865,N_845,N_858);
nand U1866 (N_1866,N_993,N_624);
and U1867 (N_1867,N_712,N_735);
and U1868 (N_1868,N_48,N_57);
nand U1869 (N_1869,N_814,N_178);
nor U1870 (N_1870,N_140,N_899);
nor U1871 (N_1871,N_2,N_788);
and U1872 (N_1872,N_575,N_459);
nor U1873 (N_1873,N_811,N_413);
xnor U1874 (N_1874,N_247,N_620);
nor U1875 (N_1875,N_979,N_158);
nor U1876 (N_1876,N_855,N_296);
nor U1877 (N_1877,N_520,N_578);
nor U1878 (N_1878,N_44,N_395);
or U1879 (N_1879,N_892,N_47);
nor U1880 (N_1880,N_802,N_821);
and U1881 (N_1881,N_768,N_554);
xor U1882 (N_1882,N_747,N_942);
or U1883 (N_1883,N_993,N_408);
xor U1884 (N_1884,N_163,N_171);
nand U1885 (N_1885,N_67,N_591);
and U1886 (N_1886,N_721,N_841);
or U1887 (N_1887,N_785,N_502);
xor U1888 (N_1888,N_202,N_127);
or U1889 (N_1889,N_180,N_638);
and U1890 (N_1890,N_936,N_852);
or U1891 (N_1891,N_881,N_115);
and U1892 (N_1892,N_272,N_577);
and U1893 (N_1893,N_720,N_526);
nor U1894 (N_1894,N_264,N_416);
and U1895 (N_1895,N_528,N_24);
nor U1896 (N_1896,N_405,N_722);
or U1897 (N_1897,N_453,N_843);
and U1898 (N_1898,N_793,N_306);
xor U1899 (N_1899,N_480,N_446);
nand U1900 (N_1900,N_131,N_545);
xnor U1901 (N_1901,N_721,N_239);
or U1902 (N_1902,N_392,N_69);
nor U1903 (N_1903,N_304,N_796);
and U1904 (N_1904,N_580,N_315);
or U1905 (N_1905,N_230,N_118);
and U1906 (N_1906,N_220,N_853);
and U1907 (N_1907,N_963,N_111);
and U1908 (N_1908,N_835,N_557);
nor U1909 (N_1909,N_185,N_652);
or U1910 (N_1910,N_380,N_409);
or U1911 (N_1911,N_757,N_447);
nor U1912 (N_1912,N_434,N_199);
or U1913 (N_1913,N_564,N_152);
nand U1914 (N_1914,N_29,N_104);
nand U1915 (N_1915,N_685,N_417);
nor U1916 (N_1916,N_423,N_535);
and U1917 (N_1917,N_586,N_129);
and U1918 (N_1918,N_247,N_170);
nor U1919 (N_1919,N_909,N_953);
and U1920 (N_1920,N_209,N_771);
and U1921 (N_1921,N_509,N_934);
or U1922 (N_1922,N_798,N_372);
xor U1923 (N_1923,N_484,N_701);
or U1924 (N_1924,N_824,N_961);
or U1925 (N_1925,N_570,N_522);
or U1926 (N_1926,N_17,N_938);
and U1927 (N_1927,N_578,N_770);
or U1928 (N_1928,N_59,N_498);
or U1929 (N_1929,N_628,N_925);
nand U1930 (N_1930,N_195,N_267);
nor U1931 (N_1931,N_975,N_635);
nand U1932 (N_1932,N_565,N_415);
nand U1933 (N_1933,N_429,N_963);
nand U1934 (N_1934,N_439,N_145);
and U1935 (N_1935,N_776,N_890);
nor U1936 (N_1936,N_89,N_381);
nand U1937 (N_1937,N_701,N_907);
nand U1938 (N_1938,N_613,N_23);
and U1939 (N_1939,N_871,N_525);
nor U1940 (N_1940,N_313,N_798);
or U1941 (N_1941,N_346,N_220);
nand U1942 (N_1942,N_678,N_410);
nand U1943 (N_1943,N_474,N_178);
nor U1944 (N_1944,N_893,N_608);
and U1945 (N_1945,N_182,N_834);
or U1946 (N_1946,N_834,N_777);
nand U1947 (N_1947,N_773,N_676);
or U1948 (N_1948,N_82,N_337);
or U1949 (N_1949,N_916,N_989);
xnor U1950 (N_1950,N_509,N_843);
nor U1951 (N_1951,N_713,N_149);
or U1952 (N_1952,N_741,N_965);
or U1953 (N_1953,N_495,N_564);
nor U1954 (N_1954,N_920,N_756);
and U1955 (N_1955,N_431,N_920);
or U1956 (N_1956,N_30,N_654);
or U1957 (N_1957,N_87,N_961);
or U1958 (N_1958,N_545,N_80);
nor U1959 (N_1959,N_281,N_965);
or U1960 (N_1960,N_257,N_83);
xor U1961 (N_1961,N_401,N_302);
nand U1962 (N_1962,N_329,N_597);
nor U1963 (N_1963,N_735,N_856);
xor U1964 (N_1964,N_832,N_7);
nor U1965 (N_1965,N_148,N_167);
nand U1966 (N_1966,N_303,N_809);
and U1967 (N_1967,N_871,N_547);
nand U1968 (N_1968,N_43,N_556);
nand U1969 (N_1969,N_800,N_454);
xnor U1970 (N_1970,N_399,N_69);
nor U1971 (N_1971,N_613,N_656);
or U1972 (N_1972,N_734,N_763);
or U1973 (N_1973,N_255,N_36);
nand U1974 (N_1974,N_465,N_900);
xor U1975 (N_1975,N_499,N_49);
or U1976 (N_1976,N_494,N_425);
xor U1977 (N_1977,N_876,N_108);
nand U1978 (N_1978,N_244,N_665);
and U1979 (N_1979,N_62,N_92);
nor U1980 (N_1980,N_341,N_635);
and U1981 (N_1981,N_142,N_596);
nand U1982 (N_1982,N_852,N_489);
or U1983 (N_1983,N_812,N_920);
and U1984 (N_1984,N_493,N_738);
or U1985 (N_1985,N_149,N_566);
and U1986 (N_1986,N_790,N_963);
nor U1987 (N_1987,N_313,N_202);
nand U1988 (N_1988,N_563,N_153);
and U1989 (N_1989,N_685,N_846);
nor U1990 (N_1990,N_828,N_236);
nor U1991 (N_1991,N_93,N_436);
or U1992 (N_1992,N_791,N_862);
nor U1993 (N_1993,N_447,N_325);
or U1994 (N_1994,N_168,N_791);
or U1995 (N_1995,N_260,N_569);
nor U1996 (N_1996,N_122,N_384);
and U1997 (N_1997,N_651,N_765);
nand U1998 (N_1998,N_527,N_981);
and U1999 (N_1999,N_881,N_332);
xor U2000 (N_2000,N_1556,N_1991);
and U2001 (N_2001,N_1914,N_1413);
nand U2002 (N_2002,N_1568,N_1963);
or U2003 (N_2003,N_1392,N_1237);
xor U2004 (N_2004,N_1138,N_1211);
nand U2005 (N_2005,N_1449,N_1286);
xor U2006 (N_2006,N_1615,N_1673);
nand U2007 (N_2007,N_1471,N_1669);
or U2008 (N_2008,N_1090,N_1672);
nor U2009 (N_2009,N_1889,N_1185);
or U2010 (N_2010,N_1801,N_1439);
or U2011 (N_2011,N_1637,N_1870);
or U2012 (N_2012,N_1034,N_1872);
and U2013 (N_2013,N_1805,N_1551);
and U2014 (N_2014,N_1245,N_1654);
nand U2015 (N_2015,N_1169,N_1099);
or U2016 (N_2016,N_1937,N_1597);
nor U2017 (N_2017,N_1520,N_1902);
nand U2018 (N_2018,N_1328,N_1311);
or U2019 (N_2019,N_1252,N_1670);
and U2020 (N_2020,N_1083,N_1527);
nor U2021 (N_2021,N_1003,N_1078);
nor U2022 (N_2022,N_1068,N_1592);
nor U2023 (N_2023,N_1072,N_1335);
or U2024 (N_2024,N_1105,N_1277);
or U2025 (N_2025,N_1101,N_1031);
nand U2026 (N_2026,N_1743,N_1194);
or U2027 (N_2027,N_1760,N_1887);
nand U2028 (N_2028,N_1632,N_1084);
and U2029 (N_2029,N_1502,N_1605);
and U2030 (N_2030,N_1524,N_1240);
nand U2031 (N_2031,N_1396,N_1258);
nand U2032 (N_2032,N_1552,N_1585);
and U2033 (N_2033,N_1880,N_1865);
and U2034 (N_2034,N_1994,N_1156);
and U2035 (N_2035,N_1326,N_1466);
nor U2036 (N_2036,N_1726,N_1886);
and U2037 (N_2037,N_1267,N_1111);
and U2038 (N_2038,N_1687,N_1680);
and U2039 (N_2039,N_1975,N_1723);
nand U2040 (N_2040,N_1410,N_1008);
and U2041 (N_2041,N_1787,N_1448);
nand U2042 (N_2042,N_1222,N_1776);
nor U2043 (N_2043,N_1708,N_1565);
or U2044 (N_2044,N_1069,N_1728);
nand U2045 (N_2045,N_1757,N_1122);
and U2046 (N_2046,N_1430,N_1148);
and U2047 (N_2047,N_1528,N_1697);
or U2048 (N_2048,N_1694,N_1955);
nor U2049 (N_2049,N_1231,N_1043);
xor U2050 (N_2050,N_1879,N_1295);
and U2051 (N_2051,N_1229,N_1476);
or U2052 (N_2052,N_1992,N_1184);
nand U2053 (N_2053,N_1517,N_1722);
or U2054 (N_2054,N_1800,N_1186);
xor U2055 (N_2055,N_1192,N_1164);
and U2056 (N_2056,N_1877,N_1956);
nor U2057 (N_2057,N_1265,N_1253);
and U2058 (N_2058,N_1884,N_1584);
or U2059 (N_2059,N_1494,N_1041);
nand U2060 (N_2060,N_1030,N_1998);
xnor U2061 (N_2061,N_1216,N_1049);
nand U2062 (N_2062,N_1289,N_1179);
and U2063 (N_2063,N_1301,N_1193);
and U2064 (N_2064,N_1575,N_1695);
nand U2065 (N_2065,N_1109,N_1067);
and U2066 (N_2066,N_1481,N_1076);
nor U2067 (N_2067,N_1601,N_1491);
nand U2068 (N_2068,N_1214,N_1793);
nand U2069 (N_2069,N_1107,N_1108);
nor U2070 (N_2070,N_1767,N_1054);
and U2071 (N_2071,N_1624,N_1233);
nor U2072 (N_2072,N_1060,N_1735);
nor U2073 (N_2073,N_1098,N_1541);
nor U2074 (N_2074,N_1402,N_1126);
or U2075 (N_2075,N_1540,N_1895);
nor U2076 (N_2076,N_1910,N_1006);
and U2077 (N_2077,N_1748,N_1118);
and U2078 (N_2078,N_1690,N_1503);
nand U2079 (N_2079,N_1951,N_1940);
or U2080 (N_2080,N_1302,N_1828);
or U2081 (N_2081,N_1752,N_1702);
nor U2082 (N_2082,N_1206,N_1273);
and U2083 (N_2083,N_1972,N_1473);
or U2084 (N_2084,N_1939,N_1638);
xor U2085 (N_2085,N_1017,N_1104);
nand U2086 (N_2086,N_1668,N_1871);
nor U2087 (N_2087,N_1275,N_1163);
nor U2088 (N_2088,N_1318,N_1798);
nand U2089 (N_2089,N_1576,N_1778);
nor U2090 (N_2090,N_1603,N_1489);
nor U2091 (N_2091,N_1210,N_1529);
nor U2092 (N_2092,N_1834,N_1139);
or U2093 (N_2093,N_1320,N_1530);
or U2094 (N_2094,N_1047,N_1796);
and U2095 (N_2095,N_1121,N_1911);
nor U2096 (N_2096,N_1634,N_1407);
nor U2097 (N_2097,N_1213,N_1157);
or U2098 (N_2098,N_1200,N_1144);
and U2099 (N_2099,N_1660,N_1720);
and U2100 (N_2100,N_1106,N_1145);
and U2101 (N_2101,N_1095,N_1182);
and U2102 (N_2102,N_1784,N_1094);
or U2103 (N_2103,N_1997,N_1152);
nor U2104 (N_2104,N_1691,N_1881);
or U2105 (N_2105,N_1492,N_1588);
nor U2106 (N_2106,N_1073,N_1897);
and U2107 (N_2107,N_1299,N_1498);
nor U2108 (N_2108,N_1858,N_1838);
and U2109 (N_2109,N_1562,N_1352);
nor U2110 (N_2110,N_1155,N_1025);
or U2111 (N_2111,N_1177,N_1243);
nand U2112 (N_2112,N_1160,N_1933);
or U2113 (N_2113,N_1700,N_1208);
or U2114 (N_2114,N_1052,N_1581);
xor U2115 (N_2115,N_1026,N_1643);
xnor U2116 (N_2116,N_1646,N_1260);
nor U2117 (N_2117,N_1266,N_1633);
nand U2118 (N_2118,N_1433,N_1379);
and U2119 (N_2119,N_1119,N_1709);
nand U2120 (N_2120,N_1401,N_1120);
and U2121 (N_2121,N_1314,N_1075);
nor U2122 (N_2122,N_1679,N_1256);
nand U2123 (N_2123,N_1451,N_1977);
nand U2124 (N_2124,N_1809,N_1554);
nand U2125 (N_2125,N_1522,N_1044);
and U2126 (N_2126,N_1465,N_1436);
or U2127 (N_2127,N_1606,N_1225);
and U2128 (N_2128,N_1876,N_1550);
nand U2129 (N_2129,N_1960,N_1789);
nand U2130 (N_2130,N_1628,N_1322);
or U2131 (N_2131,N_1027,N_1300);
nand U2132 (N_2132,N_1916,N_1346);
nand U2133 (N_2133,N_1427,N_1591);
or U2134 (N_2134,N_1096,N_1404);
xor U2135 (N_2135,N_1719,N_1969);
nor U2136 (N_2136,N_1506,N_1088);
or U2137 (N_2137,N_1467,N_1356);
nand U2138 (N_2138,N_1518,N_1408);
nand U2139 (N_2139,N_1431,N_1059);
nand U2140 (N_2140,N_1390,N_1089);
nand U2141 (N_2141,N_1666,N_1384);
nor U2142 (N_2142,N_1310,N_1345);
nor U2143 (N_2143,N_1202,N_1515);
nor U2144 (N_2144,N_1665,N_1849);
nand U2145 (N_2145,N_1779,N_1365);
or U2146 (N_2146,N_1381,N_1324);
or U2147 (N_2147,N_1747,N_1523);
or U2148 (N_2148,N_1968,N_1901);
xnor U2149 (N_2149,N_1855,N_1617);
xor U2150 (N_2150,N_1713,N_1261);
nand U2151 (N_2151,N_1154,N_1259);
or U2152 (N_2152,N_1715,N_1450);
xor U2153 (N_2153,N_1574,N_1399);
nor U2154 (N_2154,N_1731,N_1526);
nand U2155 (N_2155,N_1899,N_1839);
and U2156 (N_2156,N_1454,N_1029);
xnor U2157 (N_2157,N_1348,N_1819);
nand U2158 (N_2158,N_1387,N_1594);
xnor U2159 (N_2159,N_1452,N_1689);
xor U2160 (N_2160,N_1837,N_1058);
or U2161 (N_2161,N_1903,N_1535);
or U2162 (N_2162,N_1827,N_1740);
or U2163 (N_2163,N_1995,N_1422);
or U2164 (N_2164,N_1547,N_1426);
xnor U2165 (N_2165,N_1024,N_1894);
nor U2166 (N_2166,N_1269,N_1023);
nor U2167 (N_2167,N_1197,N_1678);
or U2168 (N_2168,N_1774,N_1488);
or U2169 (N_2169,N_1630,N_1773);
or U2170 (N_2170,N_1802,N_1781);
and U2171 (N_2171,N_1190,N_1445);
or U2172 (N_2172,N_1463,N_1092);
and U2173 (N_2173,N_1973,N_1768);
nand U2174 (N_2174,N_1948,N_1370);
and U2175 (N_2175,N_1504,N_1274);
nand U2176 (N_2176,N_1223,N_1446);
nor U2177 (N_2177,N_1724,N_1124);
nor U2178 (N_2178,N_1270,N_1170);
nand U2179 (N_2179,N_1389,N_1707);
nand U2180 (N_2180,N_1869,N_1063);
and U2181 (N_2181,N_1055,N_1763);
or U2182 (N_2182,N_1349,N_1005);
nor U2183 (N_2183,N_1593,N_1569);
nor U2184 (N_2184,N_1676,N_1358);
and U2185 (N_2185,N_1864,N_1875);
nor U2186 (N_2186,N_1363,N_1514);
nand U2187 (N_2187,N_1656,N_1685);
nand U2188 (N_2188,N_1579,N_1548);
and U2189 (N_2189,N_1770,N_1361);
nand U2190 (N_2190,N_1856,N_1609);
xor U2191 (N_2191,N_1251,N_1813);
nand U2192 (N_2192,N_1116,N_1854);
nor U2193 (N_2193,N_1683,N_1051);
and U2194 (N_2194,N_1331,N_1555);
nor U2195 (N_2195,N_1979,N_1930);
and U2196 (N_2196,N_1806,N_1571);
nor U2197 (N_2197,N_1946,N_1382);
nand U2198 (N_2198,N_1943,N_1477);
and U2199 (N_2199,N_1868,N_1851);
xnor U2200 (N_2200,N_1674,N_1860);
nor U2201 (N_2201,N_1351,N_1644);
nand U2202 (N_2202,N_1508,N_1079);
nand U2203 (N_2203,N_1961,N_1655);
or U2204 (N_2204,N_1814,N_1925);
or U2205 (N_2205,N_1458,N_1230);
and U2206 (N_2206,N_1965,N_1741);
and U2207 (N_2207,N_1167,N_1783);
and U2208 (N_2208,N_1934,N_1507);
nand U2209 (N_2209,N_1377,N_1519);
and U2210 (N_2210,N_1355,N_1432);
and U2211 (N_2211,N_1171,N_1905);
or U2212 (N_2212,N_1219,N_1172);
or U2213 (N_2213,N_1546,N_1161);
nor U2214 (N_2214,N_1143,N_1406);
or U2215 (N_2215,N_1011,N_1602);
or U2216 (N_2216,N_1647,N_1500);
nor U2217 (N_2217,N_1372,N_1343);
and U2218 (N_2218,N_1195,N_1711);
xnor U2219 (N_2219,N_1996,N_1737);
nand U2220 (N_2220,N_1056,N_1232);
nand U2221 (N_2221,N_1453,N_1703);
nor U2222 (N_2222,N_1915,N_1305);
xor U2223 (N_2223,N_1804,N_1907);
nand U2224 (N_2224,N_1283,N_1811);
nand U2225 (N_2225,N_1766,N_1110);
nand U2226 (N_2226,N_1140,N_1125);
xnor U2227 (N_2227,N_1566,N_1613);
or U2228 (N_2228,N_1599,N_1682);
and U2229 (N_2229,N_1931,N_1873);
nor U2230 (N_2230,N_1021,N_1621);
nor U2231 (N_2231,N_1516,N_1958);
and U2232 (N_2232,N_1196,N_1162);
nand U2233 (N_2233,N_1706,N_1909);
and U2234 (N_2234,N_1714,N_1264);
nor U2235 (N_2235,N_1420,N_1071);
xnor U2236 (N_2236,N_1284,N_1293);
nand U2237 (N_2237,N_1531,N_1288);
and U2238 (N_2238,N_1236,N_1038);
nand U2239 (N_2239,N_1278,N_1241);
nand U2240 (N_2240,N_1521,N_1221);
and U2241 (N_2241,N_1727,N_1572);
nor U2242 (N_2242,N_1501,N_1957);
xor U2243 (N_2243,N_1215,N_1821);
nor U2244 (N_2244,N_1847,N_1619);
nand U2245 (N_2245,N_1191,N_1461);
or U2246 (N_2246,N_1201,N_1165);
xor U2247 (N_2247,N_1829,N_1749);
or U2248 (N_2248,N_1327,N_1850);
or U2249 (N_2249,N_1397,N_1032);
and U2250 (N_2250,N_1564,N_1415);
or U2251 (N_2251,N_1964,N_1559);
nor U2252 (N_2252,N_1984,N_1978);
nor U2253 (N_2253,N_1586,N_1239);
nand U2254 (N_2254,N_1890,N_1701);
and U2255 (N_2255,N_1142,N_1254);
nand U2256 (N_2256,N_1040,N_1962);
or U2257 (N_2257,N_1822,N_1028);
and U2258 (N_2258,N_1388,N_1844);
and U2259 (N_2259,N_1441,N_1205);
nor U2260 (N_2260,N_1831,N_1022);
and U2261 (N_2261,N_1282,N_1938);
and U2262 (N_2262,N_1595,N_1153);
or U2263 (N_2263,N_1020,N_1483);
and U2264 (N_2264,N_1896,N_1730);
nand U2265 (N_2265,N_1539,N_1857);
nor U2266 (N_2266,N_1699,N_1296);
xor U2267 (N_2267,N_1852,N_1612);
or U2268 (N_2268,N_1290,N_1082);
or U2269 (N_2269,N_1651,N_1999);
or U2270 (N_2270,N_1631,N_1967);
xnor U2271 (N_2271,N_1036,N_1893);
nor U2272 (N_2272,N_1671,N_1159);
and U2273 (N_2273,N_1366,N_1537);
and U2274 (N_2274,N_1456,N_1173);
nand U2275 (N_2275,N_1100,N_1070);
or U2276 (N_2276,N_1342,N_1442);
xor U2277 (N_2277,N_1151,N_1587);
and U2278 (N_2278,N_1306,N_1178);
and U2279 (N_2279,N_1563,N_1513);
xnor U2280 (N_2280,N_1980,N_1950);
or U2281 (N_2281,N_1421,N_1340);
and U2282 (N_2282,N_1684,N_1459);
nor U2283 (N_2283,N_1091,N_1443);
nand U2284 (N_2284,N_1490,N_1403);
or U2285 (N_2285,N_1812,N_1657);
or U2286 (N_2286,N_1675,N_1294);
nor U2287 (N_2287,N_1817,N_1220);
or U2288 (N_2288,N_1512,N_1649);
nand U2289 (N_2289,N_1616,N_1457);
nor U2290 (N_2290,N_1622,N_1198);
or U2291 (N_2291,N_1487,N_1014);
and U2292 (N_2292,N_1115,N_1209);
nor U2293 (N_2293,N_1204,N_1097);
nand U2294 (N_2294,N_1117,N_1544);
nor U2295 (N_2295,N_1578,N_1904);
or U2296 (N_2296,N_1478,N_1128);
nand U2297 (N_2297,N_1696,N_1183);
nand U2298 (N_2298,N_1833,N_1046);
or U2299 (N_2299,N_1103,N_1824);
or U2300 (N_2300,N_1988,N_1945);
nand U2301 (N_2301,N_1378,N_1629);
xor U2302 (N_2302,N_1455,N_1888);
or U2303 (N_2303,N_1815,N_1007);
and U2304 (N_2304,N_1661,N_1045);
nor U2305 (N_2305,N_1132,N_1636);
and U2306 (N_2306,N_1228,N_1610);
or U2307 (N_2307,N_1495,N_1212);
nand U2308 (N_2308,N_1836,N_1843);
or U2309 (N_2309,N_1641,N_1600);
nand U2310 (N_2310,N_1199,N_1412);
xor U2311 (N_2311,N_1188,N_1986);
xor U2312 (N_2312,N_1383,N_1368);
or U2313 (N_2313,N_1347,N_1883);
and U2314 (N_2314,N_1042,N_1580);
nand U2315 (N_2315,N_1330,N_1093);
or U2316 (N_2316,N_1064,N_1297);
and U2317 (N_2317,N_1653,N_1010);
nor U2318 (N_2318,N_1435,N_1375);
nor U2319 (N_2319,N_1717,N_1797);
or U2320 (N_2320,N_1891,N_1035);
nor U2321 (N_2321,N_1534,N_1835);
nand U2322 (N_2322,N_1130,N_1405);
and U2323 (N_2323,N_1906,N_1227);
or U2324 (N_2324,N_1648,N_1333);
and U2325 (N_2325,N_1050,N_1536);
and U2326 (N_2326,N_1244,N_1039);
and U2327 (N_2327,N_1848,N_1371);
or U2328 (N_2328,N_1589,N_1218);
or U2329 (N_2329,N_1542,N_1557);
or U2330 (N_2330,N_1423,N_1558);
xnor U2331 (N_2331,N_1733,N_1718);
and U2332 (N_2332,N_1662,N_1015);
nor U2333 (N_2333,N_1898,N_1919);
xnor U2334 (N_2334,N_1102,N_1688);
nand U2335 (N_2335,N_1291,N_1280);
and U2336 (N_2336,N_1048,N_1086);
or U2337 (N_2337,N_1926,N_1560);
nor U2338 (N_2338,N_1739,N_1470);
and U2339 (N_2339,N_1511,N_1496);
or U2340 (N_2340,N_1553,N_1168);
nand U2341 (N_2341,N_1780,N_1983);
nor U2342 (N_2342,N_1181,N_1698);
or U2343 (N_2343,N_1425,N_1892);
nor U2344 (N_2344,N_1364,N_1941);
or U2345 (N_2345,N_1226,N_1842);
or U2346 (N_2346,N_1395,N_1742);
or U2347 (N_2347,N_1002,N_1279);
nor U2348 (N_2348,N_1350,N_1482);
nand U2349 (N_2349,N_1474,N_1065);
and U2350 (N_2350,N_1334,N_1681);
or U2351 (N_2351,N_1922,N_1418);
nand U2352 (N_2352,N_1147,N_1775);
or U2353 (N_2353,N_1137,N_1016);
and U2354 (N_2354,N_1391,N_1317);
and U2355 (N_2355,N_1505,N_1758);
or U2356 (N_2356,N_1133,N_1756);
nand U2357 (N_2357,N_1790,N_1411);
xor U2358 (N_2358,N_1769,N_1863);
or U2359 (N_2359,N_1853,N_1460);
nor U2360 (N_2360,N_1061,N_1549);
nand U2361 (N_2361,N_1583,N_1493);
or U2362 (N_2362,N_1764,N_1645);
and U2363 (N_2363,N_1000,N_1867);
nor U2364 (N_2364,N_1944,N_1927);
nor U2365 (N_2365,N_1971,N_1484);
or U2366 (N_2366,N_1369,N_1820);
and U2367 (N_2367,N_1447,N_1131);
or U2368 (N_2368,N_1792,N_1795);
xnor U2369 (N_2369,N_1928,N_1954);
xor U2370 (N_2370,N_1416,N_1510);
and U2371 (N_2371,N_1429,N_1479);
nand U2372 (N_2372,N_1292,N_1704);
nand U2373 (N_2373,N_1808,N_1913);
nand U2374 (N_2374,N_1625,N_1339);
and U2375 (N_2375,N_1611,N_1596);
nand U2376 (N_2376,N_1235,N_1650);
and U2377 (N_2377,N_1794,N_1745);
nand U2378 (N_2378,N_1755,N_1761);
nor U2379 (N_2379,N_1417,N_1862);
xor U2380 (N_2380,N_1087,N_1917);
nor U2381 (N_2381,N_1362,N_1825);
nor U2382 (N_2382,N_1874,N_1238);
and U2383 (N_2383,N_1658,N_1604);
and U2384 (N_2384,N_1771,N_1062);
or U2385 (N_2385,N_1882,N_1315);
xor U2386 (N_2386,N_1932,N_1693);
or U2387 (N_2387,N_1981,N_1710);
nand U2388 (N_2388,N_1242,N_1246);
xnor U2389 (N_2389,N_1112,N_1263);
or U2390 (N_2390,N_1359,N_1830);
xor U2391 (N_2391,N_1920,N_1725);
nor U2392 (N_2392,N_1398,N_1712);
and U2393 (N_2393,N_1538,N_1248);
nor U2394 (N_2394,N_1791,N_1319);
and U2395 (N_2395,N_1627,N_1545);
and U2396 (N_2396,N_1053,N_1424);
or U2397 (N_2397,N_1912,N_1136);
or U2398 (N_2398,N_1990,N_1386);
nor U2399 (N_2399,N_1705,N_1746);
nand U2400 (N_2400,N_1019,N_1664);
and U2401 (N_2401,N_1271,N_1338);
and U2402 (N_2402,N_1262,N_1440);
nand U2403 (N_2403,N_1176,N_1400);
xnor U2404 (N_2404,N_1772,N_1249);
nor U2405 (N_2405,N_1908,N_1976);
and U2406 (N_2406,N_1736,N_1336);
nand U2407 (N_2407,N_1004,N_1626);
nand U2408 (N_2408,N_1929,N_1750);
and U2409 (N_2409,N_1974,N_1298);
and U2410 (N_2410,N_1543,N_1846);
or U2411 (N_2411,N_1623,N_1360);
and U2412 (N_2412,N_1114,N_1614);
nand U2413 (N_2413,N_1921,N_1826);
or U2414 (N_2414,N_1692,N_1337);
and U2415 (N_2415,N_1759,N_1217);
nor U2416 (N_2416,N_1608,N_1141);
and U2417 (N_2417,N_1485,N_1577);
and U2418 (N_2418,N_1762,N_1033);
xnor U2419 (N_2419,N_1321,N_1303);
xor U2420 (N_2420,N_1085,N_1840);
and U2421 (N_2421,N_1652,N_1942);
and U2422 (N_2422,N_1325,N_1374);
nor U2423 (N_2423,N_1080,N_1618);
nor U2424 (N_2424,N_1642,N_1187);
and U2425 (N_2425,N_1475,N_1127);
xnor U2426 (N_2426,N_1823,N_1716);
or U2427 (N_2427,N_1667,N_1959);
or U2428 (N_2428,N_1532,N_1018);
nor U2429 (N_2429,N_1935,N_1734);
or U2430 (N_2430,N_1437,N_1393);
and U2431 (N_2431,N_1158,N_1859);
nand U2432 (N_2432,N_1367,N_1970);
or U2433 (N_2433,N_1316,N_1861);
and U2434 (N_2434,N_1832,N_1037);
nand U2435 (N_2435,N_1561,N_1567);
xor U2436 (N_2436,N_1257,N_1135);
or U2437 (N_2437,N_1640,N_1376);
and U2438 (N_2438,N_1598,N_1203);
nor U2439 (N_2439,N_1635,N_1786);
nand U2440 (N_2440,N_1738,N_1497);
nand U2441 (N_2441,N_1807,N_1287);
nor U2442 (N_2442,N_1480,N_1953);
xnor U2443 (N_2443,N_1885,N_1799);
nor U2444 (N_2444,N_1509,N_1620);
xor U2445 (N_2445,N_1353,N_1468);
nand U2446 (N_2446,N_1354,N_1918);
xnor U2447 (N_2447,N_1357,N_1134);
and U2448 (N_2448,N_1499,N_1989);
nor U2449 (N_2449,N_1782,N_1841);
or U2450 (N_2450,N_1385,N_1765);
xor U2451 (N_2451,N_1949,N_1234);
or U2452 (N_2452,N_1607,N_1081);
nand U2453 (N_2453,N_1268,N_1472);
nor U2454 (N_2454,N_1309,N_1180);
and U2455 (N_2455,N_1659,N_1985);
or U2456 (N_2456,N_1845,N_1175);
and U2457 (N_2457,N_1123,N_1394);
nor U2458 (N_2458,N_1785,N_1255);
nand U2459 (N_2459,N_1818,N_1753);
or U2460 (N_2460,N_1380,N_1947);
or U2461 (N_2461,N_1729,N_1462);
and U2462 (N_2462,N_1166,N_1066);
nand U2463 (N_2463,N_1582,N_1174);
nand U2464 (N_2464,N_1341,N_1993);
and U2465 (N_2465,N_1009,N_1113);
nand U2466 (N_2466,N_1987,N_1732);
xnor U2467 (N_2467,N_1189,N_1744);
and U2468 (N_2468,N_1866,N_1013);
or U2469 (N_2469,N_1077,N_1329);
nand U2470 (N_2470,N_1677,N_1373);
and U2471 (N_2471,N_1754,N_1878);
and U2472 (N_2472,N_1464,N_1323);
and U2473 (N_2473,N_1307,N_1788);
xnor U2474 (N_2474,N_1001,N_1686);
nand U2475 (N_2475,N_1966,N_1224);
and U2476 (N_2476,N_1923,N_1428);
and U2477 (N_2477,N_1247,N_1074);
and U2478 (N_2478,N_1751,N_1149);
nor U2479 (N_2479,N_1146,N_1272);
xor U2480 (N_2480,N_1469,N_1721);
nand U2481 (N_2481,N_1777,N_1924);
and U2482 (N_2482,N_1525,N_1304);
nor U2483 (N_2483,N_1057,N_1276);
and U2484 (N_2484,N_1639,N_1663);
or U2485 (N_2485,N_1816,N_1982);
and U2486 (N_2486,N_1810,N_1900);
nand U2487 (N_2487,N_1207,N_1313);
nand U2488 (N_2488,N_1952,N_1150);
nor U2489 (N_2489,N_1573,N_1312);
nand U2490 (N_2490,N_1434,N_1570);
or U2491 (N_2491,N_1419,N_1344);
or U2492 (N_2492,N_1332,N_1936);
nand U2493 (N_2493,N_1486,N_1438);
nor U2494 (N_2494,N_1803,N_1409);
and U2495 (N_2495,N_1414,N_1308);
or U2496 (N_2496,N_1285,N_1533);
xnor U2497 (N_2497,N_1590,N_1250);
nand U2498 (N_2498,N_1281,N_1012);
nand U2499 (N_2499,N_1129,N_1444);
nor U2500 (N_2500,N_1721,N_1025);
and U2501 (N_2501,N_1527,N_1219);
and U2502 (N_2502,N_1966,N_1055);
nand U2503 (N_2503,N_1892,N_1306);
and U2504 (N_2504,N_1471,N_1194);
or U2505 (N_2505,N_1949,N_1598);
and U2506 (N_2506,N_1956,N_1431);
nand U2507 (N_2507,N_1951,N_1695);
nand U2508 (N_2508,N_1932,N_1264);
nand U2509 (N_2509,N_1521,N_1756);
xor U2510 (N_2510,N_1504,N_1743);
or U2511 (N_2511,N_1957,N_1271);
or U2512 (N_2512,N_1805,N_1198);
xor U2513 (N_2513,N_1562,N_1600);
nand U2514 (N_2514,N_1766,N_1839);
or U2515 (N_2515,N_1595,N_1977);
and U2516 (N_2516,N_1747,N_1385);
xnor U2517 (N_2517,N_1559,N_1207);
nand U2518 (N_2518,N_1639,N_1794);
and U2519 (N_2519,N_1762,N_1869);
nor U2520 (N_2520,N_1983,N_1004);
and U2521 (N_2521,N_1855,N_1853);
or U2522 (N_2522,N_1990,N_1951);
nand U2523 (N_2523,N_1936,N_1755);
or U2524 (N_2524,N_1845,N_1661);
or U2525 (N_2525,N_1460,N_1907);
or U2526 (N_2526,N_1172,N_1433);
nor U2527 (N_2527,N_1029,N_1204);
and U2528 (N_2528,N_1675,N_1059);
xnor U2529 (N_2529,N_1060,N_1557);
nand U2530 (N_2530,N_1550,N_1662);
nor U2531 (N_2531,N_1646,N_1398);
nand U2532 (N_2532,N_1259,N_1579);
nor U2533 (N_2533,N_1219,N_1970);
and U2534 (N_2534,N_1463,N_1279);
and U2535 (N_2535,N_1536,N_1773);
nor U2536 (N_2536,N_1460,N_1741);
and U2537 (N_2537,N_1116,N_1058);
or U2538 (N_2538,N_1988,N_1899);
and U2539 (N_2539,N_1962,N_1373);
nor U2540 (N_2540,N_1360,N_1599);
or U2541 (N_2541,N_1358,N_1924);
or U2542 (N_2542,N_1645,N_1753);
nand U2543 (N_2543,N_1155,N_1910);
nand U2544 (N_2544,N_1679,N_1095);
and U2545 (N_2545,N_1322,N_1755);
nor U2546 (N_2546,N_1598,N_1505);
nand U2547 (N_2547,N_1226,N_1107);
nor U2548 (N_2548,N_1823,N_1946);
or U2549 (N_2549,N_1404,N_1200);
and U2550 (N_2550,N_1270,N_1958);
or U2551 (N_2551,N_1455,N_1329);
nand U2552 (N_2552,N_1590,N_1635);
nor U2553 (N_2553,N_1860,N_1524);
nand U2554 (N_2554,N_1506,N_1074);
nor U2555 (N_2555,N_1891,N_1724);
nor U2556 (N_2556,N_1461,N_1188);
nor U2557 (N_2557,N_1028,N_1215);
or U2558 (N_2558,N_1960,N_1825);
xor U2559 (N_2559,N_1759,N_1675);
and U2560 (N_2560,N_1640,N_1720);
xor U2561 (N_2561,N_1996,N_1509);
or U2562 (N_2562,N_1973,N_1147);
nor U2563 (N_2563,N_1840,N_1172);
or U2564 (N_2564,N_1339,N_1980);
or U2565 (N_2565,N_1649,N_1306);
nand U2566 (N_2566,N_1848,N_1525);
or U2567 (N_2567,N_1362,N_1983);
or U2568 (N_2568,N_1831,N_1934);
nand U2569 (N_2569,N_1187,N_1997);
and U2570 (N_2570,N_1804,N_1007);
nand U2571 (N_2571,N_1895,N_1805);
and U2572 (N_2572,N_1399,N_1618);
nand U2573 (N_2573,N_1705,N_1033);
xnor U2574 (N_2574,N_1543,N_1941);
nor U2575 (N_2575,N_1527,N_1168);
nor U2576 (N_2576,N_1216,N_1793);
nor U2577 (N_2577,N_1688,N_1534);
and U2578 (N_2578,N_1882,N_1647);
and U2579 (N_2579,N_1523,N_1896);
nor U2580 (N_2580,N_1661,N_1287);
nor U2581 (N_2581,N_1468,N_1883);
or U2582 (N_2582,N_1163,N_1435);
or U2583 (N_2583,N_1285,N_1660);
nand U2584 (N_2584,N_1428,N_1247);
xor U2585 (N_2585,N_1083,N_1340);
nand U2586 (N_2586,N_1007,N_1383);
and U2587 (N_2587,N_1725,N_1367);
or U2588 (N_2588,N_1463,N_1188);
nor U2589 (N_2589,N_1022,N_1537);
and U2590 (N_2590,N_1771,N_1920);
and U2591 (N_2591,N_1199,N_1991);
and U2592 (N_2592,N_1239,N_1625);
and U2593 (N_2593,N_1827,N_1865);
nand U2594 (N_2594,N_1028,N_1140);
nand U2595 (N_2595,N_1417,N_1530);
nand U2596 (N_2596,N_1949,N_1462);
and U2597 (N_2597,N_1010,N_1473);
nor U2598 (N_2598,N_1515,N_1502);
xnor U2599 (N_2599,N_1858,N_1356);
nand U2600 (N_2600,N_1924,N_1164);
or U2601 (N_2601,N_1446,N_1893);
nor U2602 (N_2602,N_1548,N_1613);
nor U2603 (N_2603,N_1740,N_1394);
nand U2604 (N_2604,N_1148,N_1335);
and U2605 (N_2605,N_1487,N_1480);
or U2606 (N_2606,N_1869,N_1603);
nand U2607 (N_2607,N_1051,N_1054);
nor U2608 (N_2608,N_1558,N_1635);
nor U2609 (N_2609,N_1601,N_1819);
or U2610 (N_2610,N_1810,N_1321);
nor U2611 (N_2611,N_1550,N_1392);
and U2612 (N_2612,N_1714,N_1078);
and U2613 (N_2613,N_1621,N_1315);
and U2614 (N_2614,N_1809,N_1549);
xor U2615 (N_2615,N_1036,N_1239);
nand U2616 (N_2616,N_1171,N_1595);
or U2617 (N_2617,N_1237,N_1485);
xor U2618 (N_2618,N_1404,N_1538);
nor U2619 (N_2619,N_1068,N_1892);
nor U2620 (N_2620,N_1274,N_1366);
or U2621 (N_2621,N_1257,N_1198);
and U2622 (N_2622,N_1929,N_1866);
nor U2623 (N_2623,N_1247,N_1736);
or U2624 (N_2624,N_1784,N_1201);
nor U2625 (N_2625,N_1458,N_1486);
nor U2626 (N_2626,N_1806,N_1930);
and U2627 (N_2627,N_1304,N_1209);
nor U2628 (N_2628,N_1386,N_1034);
nand U2629 (N_2629,N_1997,N_1312);
nor U2630 (N_2630,N_1792,N_1037);
nand U2631 (N_2631,N_1691,N_1405);
nor U2632 (N_2632,N_1104,N_1933);
or U2633 (N_2633,N_1916,N_1478);
or U2634 (N_2634,N_1378,N_1215);
nor U2635 (N_2635,N_1606,N_1024);
or U2636 (N_2636,N_1595,N_1401);
nand U2637 (N_2637,N_1520,N_1015);
nor U2638 (N_2638,N_1707,N_1415);
nor U2639 (N_2639,N_1460,N_1919);
xor U2640 (N_2640,N_1070,N_1846);
nor U2641 (N_2641,N_1894,N_1809);
and U2642 (N_2642,N_1787,N_1954);
and U2643 (N_2643,N_1544,N_1212);
nor U2644 (N_2644,N_1463,N_1493);
and U2645 (N_2645,N_1272,N_1526);
nor U2646 (N_2646,N_1554,N_1497);
or U2647 (N_2647,N_1329,N_1710);
or U2648 (N_2648,N_1775,N_1567);
nor U2649 (N_2649,N_1583,N_1693);
and U2650 (N_2650,N_1230,N_1992);
xor U2651 (N_2651,N_1051,N_1580);
nor U2652 (N_2652,N_1105,N_1805);
nor U2653 (N_2653,N_1640,N_1302);
nor U2654 (N_2654,N_1886,N_1062);
nor U2655 (N_2655,N_1549,N_1840);
nor U2656 (N_2656,N_1103,N_1676);
or U2657 (N_2657,N_1104,N_1166);
nand U2658 (N_2658,N_1554,N_1656);
nand U2659 (N_2659,N_1856,N_1163);
or U2660 (N_2660,N_1209,N_1505);
or U2661 (N_2661,N_1295,N_1720);
nor U2662 (N_2662,N_1383,N_1415);
and U2663 (N_2663,N_1247,N_1475);
nor U2664 (N_2664,N_1254,N_1523);
nand U2665 (N_2665,N_1681,N_1505);
nor U2666 (N_2666,N_1333,N_1511);
nand U2667 (N_2667,N_1431,N_1360);
or U2668 (N_2668,N_1443,N_1544);
nor U2669 (N_2669,N_1648,N_1570);
nor U2670 (N_2670,N_1741,N_1020);
or U2671 (N_2671,N_1176,N_1746);
nor U2672 (N_2672,N_1506,N_1684);
nand U2673 (N_2673,N_1435,N_1468);
nor U2674 (N_2674,N_1695,N_1394);
or U2675 (N_2675,N_1786,N_1362);
or U2676 (N_2676,N_1017,N_1663);
nor U2677 (N_2677,N_1622,N_1264);
nor U2678 (N_2678,N_1450,N_1307);
nor U2679 (N_2679,N_1813,N_1079);
or U2680 (N_2680,N_1962,N_1582);
nand U2681 (N_2681,N_1011,N_1819);
or U2682 (N_2682,N_1036,N_1515);
nand U2683 (N_2683,N_1788,N_1390);
or U2684 (N_2684,N_1114,N_1567);
and U2685 (N_2685,N_1064,N_1833);
nand U2686 (N_2686,N_1834,N_1594);
or U2687 (N_2687,N_1899,N_1035);
nand U2688 (N_2688,N_1309,N_1028);
and U2689 (N_2689,N_1649,N_1388);
nand U2690 (N_2690,N_1561,N_1805);
nand U2691 (N_2691,N_1108,N_1519);
nor U2692 (N_2692,N_1980,N_1889);
nand U2693 (N_2693,N_1634,N_1946);
xor U2694 (N_2694,N_1302,N_1522);
xor U2695 (N_2695,N_1973,N_1512);
nand U2696 (N_2696,N_1758,N_1535);
or U2697 (N_2697,N_1714,N_1613);
nand U2698 (N_2698,N_1365,N_1251);
and U2699 (N_2699,N_1742,N_1860);
and U2700 (N_2700,N_1921,N_1058);
or U2701 (N_2701,N_1430,N_1054);
nor U2702 (N_2702,N_1275,N_1160);
xor U2703 (N_2703,N_1386,N_1460);
nand U2704 (N_2704,N_1233,N_1199);
nor U2705 (N_2705,N_1289,N_1417);
or U2706 (N_2706,N_1425,N_1275);
or U2707 (N_2707,N_1525,N_1201);
nand U2708 (N_2708,N_1295,N_1432);
and U2709 (N_2709,N_1962,N_1243);
nand U2710 (N_2710,N_1973,N_1526);
nand U2711 (N_2711,N_1028,N_1015);
and U2712 (N_2712,N_1064,N_1477);
and U2713 (N_2713,N_1693,N_1419);
and U2714 (N_2714,N_1045,N_1708);
xor U2715 (N_2715,N_1291,N_1729);
nor U2716 (N_2716,N_1071,N_1384);
nor U2717 (N_2717,N_1454,N_1006);
or U2718 (N_2718,N_1116,N_1514);
nand U2719 (N_2719,N_1987,N_1845);
and U2720 (N_2720,N_1225,N_1998);
or U2721 (N_2721,N_1905,N_1770);
nor U2722 (N_2722,N_1396,N_1420);
and U2723 (N_2723,N_1892,N_1523);
or U2724 (N_2724,N_1406,N_1683);
or U2725 (N_2725,N_1640,N_1332);
nand U2726 (N_2726,N_1461,N_1823);
and U2727 (N_2727,N_1359,N_1342);
nor U2728 (N_2728,N_1309,N_1203);
nor U2729 (N_2729,N_1255,N_1059);
and U2730 (N_2730,N_1799,N_1354);
nand U2731 (N_2731,N_1811,N_1855);
and U2732 (N_2732,N_1853,N_1492);
and U2733 (N_2733,N_1949,N_1692);
xnor U2734 (N_2734,N_1466,N_1525);
nor U2735 (N_2735,N_1758,N_1695);
nor U2736 (N_2736,N_1703,N_1545);
nand U2737 (N_2737,N_1025,N_1487);
and U2738 (N_2738,N_1293,N_1605);
xor U2739 (N_2739,N_1484,N_1039);
or U2740 (N_2740,N_1938,N_1721);
nor U2741 (N_2741,N_1289,N_1367);
nor U2742 (N_2742,N_1006,N_1771);
nor U2743 (N_2743,N_1932,N_1038);
and U2744 (N_2744,N_1431,N_1185);
xnor U2745 (N_2745,N_1116,N_1787);
and U2746 (N_2746,N_1030,N_1846);
and U2747 (N_2747,N_1015,N_1799);
nand U2748 (N_2748,N_1632,N_1874);
or U2749 (N_2749,N_1003,N_1236);
nor U2750 (N_2750,N_1941,N_1204);
nor U2751 (N_2751,N_1180,N_1670);
xnor U2752 (N_2752,N_1245,N_1994);
and U2753 (N_2753,N_1359,N_1152);
nor U2754 (N_2754,N_1027,N_1367);
nand U2755 (N_2755,N_1515,N_1495);
or U2756 (N_2756,N_1232,N_1616);
xnor U2757 (N_2757,N_1565,N_1278);
nor U2758 (N_2758,N_1729,N_1704);
and U2759 (N_2759,N_1532,N_1749);
nand U2760 (N_2760,N_1006,N_1141);
or U2761 (N_2761,N_1657,N_1468);
nor U2762 (N_2762,N_1436,N_1264);
nand U2763 (N_2763,N_1858,N_1695);
nand U2764 (N_2764,N_1353,N_1411);
and U2765 (N_2765,N_1447,N_1034);
or U2766 (N_2766,N_1785,N_1407);
and U2767 (N_2767,N_1167,N_1486);
nor U2768 (N_2768,N_1955,N_1911);
or U2769 (N_2769,N_1501,N_1057);
nor U2770 (N_2770,N_1301,N_1332);
nor U2771 (N_2771,N_1438,N_1868);
nor U2772 (N_2772,N_1358,N_1147);
nand U2773 (N_2773,N_1381,N_1162);
or U2774 (N_2774,N_1472,N_1252);
or U2775 (N_2775,N_1075,N_1123);
or U2776 (N_2776,N_1658,N_1894);
nand U2777 (N_2777,N_1618,N_1338);
nand U2778 (N_2778,N_1201,N_1781);
nor U2779 (N_2779,N_1239,N_1336);
and U2780 (N_2780,N_1512,N_1564);
or U2781 (N_2781,N_1868,N_1654);
nand U2782 (N_2782,N_1850,N_1282);
or U2783 (N_2783,N_1642,N_1031);
nand U2784 (N_2784,N_1458,N_1280);
and U2785 (N_2785,N_1811,N_1988);
nor U2786 (N_2786,N_1501,N_1972);
nor U2787 (N_2787,N_1479,N_1426);
nand U2788 (N_2788,N_1090,N_1689);
nor U2789 (N_2789,N_1302,N_1222);
or U2790 (N_2790,N_1099,N_1052);
and U2791 (N_2791,N_1425,N_1573);
and U2792 (N_2792,N_1637,N_1438);
and U2793 (N_2793,N_1812,N_1269);
nand U2794 (N_2794,N_1685,N_1259);
and U2795 (N_2795,N_1646,N_1106);
nor U2796 (N_2796,N_1949,N_1396);
and U2797 (N_2797,N_1806,N_1607);
nand U2798 (N_2798,N_1156,N_1595);
nor U2799 (N_2799,N_1222,N_1960);
xor U2800 (N_2800,N_1909,N_1797);
or U2801 (N_2801,N_1925,N_1613);
nor U2802 (N_2802,N_1407,N_1366);
and U2803 (N_2803,N_1919,N_1384);
or U2804 (N_2804,N_1241,N_1447);
or U2805 (N_2805,N_1666,N_1070);
nor U2806 (N_2806,N_1533,N_1002);
nand U2807 (N_2807,N_1683,N_1704);
nor U2808 (N_2808,N_1874,N_1002);
nor U2809 (N_2809,N_1211,N_1015);
or U2810 (N_2810,N_1216,N_1116);
and U2811 (N_2811,N_1027,N_1436);
or U2812 (N_2812,N_1813,N_1908);
nor U2813 (N_2813,N_1368,N_1009);
nor U2814 (N_2814,N_1558,N_1757);
or U2815 (N_2815,N_1471,N_1293);
nor U2816 (N_2816,N_1009,N_1800);
or U2817 (N_2817,N_1320,N_1637);
nor U2818 (N_2818,N_1176,N_1158);
nor U2819 (N_2819,N_1828,N_1654);
nand U2820 (N_2820,N_1202,N_1714);
xor U2821 (N_2821,N_1934,N_1067);
xor U2822 (N_2822,N_1374,N_1238);
and U2823 (N_2823,N_1299,N_1482);
and U2824 (N_2824,N_1511,N_1249);
nor U2825 (N_2825,N_1554,N_1789);
nor U2826 (N_2826,N_1571,N_1815);
nand U2827 (N_2827,N_1790,N_1255);
and U2828 (N_2828,N_1258,N_1681);
nand U2829 (N_2829,N_1243,N_1045);
nand U2830 (N_2830,N_1235,N_1188);
nor U2831 (N_2831,N_1371,N_1187);
and U2832 (N_2832,N_1483,N_1630);
nand U2833 (N_2833,N_1810,N_1515);
and U2834 (N_2834,N_1511,N_1022);
nand U2835 (N_2835,N_1578,N_1594);
and U2836 (N_2836,N_1110,N_1775);
and U2837 (N_2837,N_1884,N_1406);
and U2838 (N_2838,N_1629,N_1728);
or U2839 (N_2839,N_1305,N_1326);
nand U2840 (N_2840,N_1498,N_1654);
nand U2841 (N_2841,N_1226,N_1033);
nand U2842 (N_2842,N_1051,N_1289);
xnor U2843 (N_2843,N_1945,N_1909);
nand U2844 (N_2844,N_1767,N_1021);
or U2845 (N_2845,N_1006,N_1154);
and U2846 (N_2846,N_1145,N_1296);
or U2847 (N_2847,N_1730,N_1456);
nor U2848 (N_2848,N_1996,N_1058);
nor U2849 (N_2849,N_1714,N_1148);
xor U2850 (N_2850,N_1887,N_1967);
xor U2851 (N_2851,N_1185,N_1847);
nand U2852 (N_2852,N_1333,N_1329);
xor U2853 (N_2853,N_1067,N_1243);
nor U2854 (N_2854,N_1698,N_1448);
nand U2855 (N_2855,N_1086,N_1608);
nand U2856 (N_2856,N_1200,N_1675);
nor U2857 (N_2857,N_1740,N_1387);
nor U2858 (N_2858,N_1344,N_1690);
nor U2859 (N_2859,N_1482,N_1245);
xnor U2860 (N_2860,N_1725,N_1284);
nand U2861 (N_2861,N_1088,N_1702);
or U2862 (N_2862,N_1034,N_1185);
xnor U2863 (N_2863,N_1468,N_1950);
nand U2864 (N_2864,N_1590,N_1199);
or U2865 (N_2865,N_1862,N_1400);
and U2866 (N_2866,N_1320,N_1656);
nor U2867 (N_2867,N_1664,N_1475);
nand U2868 (N_2868,N_1252,N_1243);
and U2869 (N_2869,N_1047,N_1934);
and U2870 (N_2870,N_1582,N_1041);
nor U2871 (N_2871,N_1374,N_1333);
nand U2872 (N_2872,N_1068,N_1375);
nand U2873 (N_2873,N_1241,N_1910);
nand U2874 (N_2874,N_1677,N_1887);
nor U2875 (N_2875,N_1731,N_1705);
xor U2876 (N_2876,N_1502,N_1200);
or U2877 (N_2877,N_1965,N_1086);
nor U2878 (N_2878,N_1483,N_1162);
and U2879 (N_2879,N_1218,N_1232);
or U2880 (N_2880,N_1011,N_1835);
and U2881 (N_2881,N_1573,N_1600);
nand U2882 (N_2882,N_1531,N_1347);
and U2883 (N_2883,N_1183,N_1860);
or U2884 (N_2884,N_1651,N_1774);
or U2885 (N_2885,N_1797,N_1506);
nand U2886 (N_2886,N_1612,N_1935);
nand U2887 (N_2887,N_1567,N_1218);
and U2888 (N_2888,N_1463,N_1534);
nor U2889 (N_2889,N_1318,N_1401);
or U2890 (N_2890,N_1608,N_1808);
and U2891 (N_2891,N_1329,N_1344);
nor U2892 (N_2892,N_1564,N_1487);
and U2893 (N_2893,N_1987,N_1994);
nand U2894 (N_2894,N_1370,N_1192);
nand U2895 (N_2895,N_1482,N_1502);
and U2896 (N_2896,N_1788,N_1254);
nor U2897 (N_2897,N_1599,N_1797);
or U2898 (N_2898,N_1993,N_1070);
nor U2899 (N_2899,N_1267,N_1845);
nand U2900 (N_2900,N_1386,N_1081);
nor U2901 (N_2901,N_1336,N_1976);
or U2902 (N_2902,N_1125,N_1939);
and U2903 (N_2903,N_1208,N_1676);
nand U2904 (N_2904,N_1670,N_1339);
xor U2905 (N_2905,N_1857,N_1594);
nor U2906 (N_2906,N_1679,N_1155);
nand U2907 (N_2907,N_1073,N_1632);
and U2908 (N_2908,N_1644,N_1213);
xnor U2909 (N_2909,N_1938,N_1918);
nand U2910 (N_2910,N_1952,N_1777);
and U2911 (N_2911,N_1408,N_1114);
and U2912 (N_2912,N_1779,N_1562);
xor U2913 (N_2913,N_1462,N_1726);
nor U2914 (N_2914,N_1471,N_1943);
or U2915 (N_2915,N_1948,N_1115);
and U2916 (N_2916,N_1414,N_1692);
and U2917 (N_2917,N_1644,N_1472);
and U2918 (N_2918,N_1278,N_1960);
and U2919 (N_2919,N_1218,N_1684);
xor U2920 (N_2920,N_1749,N_1127);
xnor U2921 (N_2921,N_1914,N_1015);
and U2922 (N_2922,N_1845,N_1342);
and U2923 (N_2923,N_1189,N_1062);
or U2924 (N_2924,N_1164,N_1974);
or U2925 (N_2925,N_1052,N_1685);
and U2926 (N_2926,N_1256,N_1745);
nand U2927 (N_2927,N_1264,N_1581);
nand U2928 (N_2928,N_1168,N_1245);
nor U2929 (N_2929,N_1669,N_1253);
and U2930 (N_2930,N_1548,N_1006);
and U2931 (N_2931,N_1291,N_1860);
nand U2932 (N_2932,N_1670,N_1989);
nor U2933 (N_2933,N_1588,N_1092);
nor U2934 (N_2934,N_1825,N_1416);
or U2935 (N_2935,N_1089,N_1320);
or U2936 (N_2936,N_1944,N_1210);
and U2937 (N_2937,N_1738,N_1012);
xor U2938 (N_2938,N_1144,N_1416);
nor U2939 (N_2939,N_1477,N_1268);
and U2940 (N_2940,N_1543,N_1372);
nor U2941 (N_2941,N_1950,N_1894);
or U2942 (N_2942,N_1838,N_1307);
nor U2943 (N_2943,N_1987,N_1191);
and U2944 (N_2944,N_1013,N_1907);
nand U2945 (N_2945,N_1274,N_1270);
or U2946 (N_2946,N_1296,N_1439);
and U2947 (N_2947,N_1213,N_1567);
nor U2948 (N_2948,N_1558,N_1357);
nand U2949 (N_2949,N_1951,N_1036);
nand U2950 (N_2950,N_1833,N_1366);
xnor U2951 (N_2951,N_1406,N_1769);
and U2952 (N_2952,N_1981,N_1201);
and U2953 (N_2953,N_1672,N_1634);
nand U2954 (N_2954,N_1614,N_1240);
and U2955 (N_2955,N_1943,N_1577);
xnor U2956 (N_2956,N_1987,N_1487);
nor U2957 (N_2957,N_1783,N_1153);
nor U2958 (N_2958,N_1005,N_1347);
or U2959 (N_2959,N_1566,N_1015);
nand U2960 (N_2960,N_1685,N_1417);
and U2961 (N_2961,N_1671,N_1108);
nor U2962 (N_2962,N_1862,N_1586);
or U2963 (N_2963,N_1990,N_1286);
nand U2964 (N_2964,N_1087,N_1731);
xor U2965 (N_2965,N_1460,N_1205);
nor U2966 (N_2966,N_1785,N_1194);
and U2967 (N_2967,N_1623,N_1510);
or U2968 (N_2968,N_1750,N_1023);
xnor U2969 (N_2969,N_1216,N_1178);
nor U2970 (N_2970,N_1432,N_1788);
or U2971 (N_2971,N_1038,N_1750);
or U2972 (N_2972,N_1821,N_1844);
nand U2973 (N_2973,N_1858,N_1536);
and U2974 (N_2974,N_1856,N_1665);
xor U2975 (N_2975,N_1941,N_1673);
nor U2976 (N_2976,N_1913,N_1975);
nand U2977 (N_2977,N_1295,N_1482);
and U2978 (N_2978,N_1777,N_1748);
nor U2979 (N_2979,N_1337,N_1363);
nand U2980 (N_2980,N_1238,N_1869);
nand U2981 (N_2981,N_1862,N_1629);
nand U2982 (N_2982,N_1060,N_1706);
and U2983 (N_2983,N_1896,N_1843);
xnor U2984 (N_2984,N_1984,N_1967);
and U2985 (N_2985,N_1703,N_1115);
nand U2986 (N_2986,N_1922,N_1210);
nor U2987 (N_2987,N_1506,N_1897);
nor U2988 (N_2988,N_1245,N_1266);
nor U2989 (N_2989,N_1334,N_1301);
xnor U2990 (N_2990,N_1932,N_1795);
or U2991 (N_2991,N_1839,N_1461);
nor U2992 (N_2992,N_1476,N_1805);
or U2993 (N_2993,N_1082,N_1021);
nor U2994 (N_2994,N_1068,N_1442);
and U2995 (N_2995,N_1021,N_1493);
and U2996 (N_2996,N_1356,N_1452);
nand U2997 (N_2997,N_1210,N_1590);
nor U2998 (N_2998,N_1451,N_1381);
or U2999 (N_2999,N_1518,N_1671);
and U3000 (N_3000,N_2659,N_2039);
nand U3001 (N_3001,N_2246,N_2450);
nor U3002 (N_3002,N_2379,N_2907);
nand U3003 (N_3003,N_2452,N_2015);
xnor U3004 (N_3004,N_2234,N_2301);
nand U3005 (N_3005,N_2276,N_2519);
or U3006 (N_3006,N_2343,N_2461);
nor U3007 (N_3007,N_2896,N_2462);
and U3008 (N_3008,N_2061,N_2347);
nand U3009 (N_3009,N_2420,N_2767);
nand U3010 (N_3010,N_2367,N_2227);
nand U3011 (N_3011,N_2162,N_2577);
nand U3012 (N_3012,N_2010,N_2311);
and U3013 (N_3013,N_2555,N_2055);
and U3014 (N_3014,N_2840,N_2842);
nand U3015 (N_3015,N_2979,N_2387);
nor U3016 (N_3016,N_2744,N_2786);
and U3017 (N_3017,N_2108,N_2133);
and U3018 (N_3018,N_2600,N_2638);
nor U3019 (N_3019,N_2340,N_2059);
nand U3020 (N_3020,N_2229,N_2371);
and U3021 (N_3021,N_2838,N_2255);
nor U3022 (N_3022,N_2500,N_2874);
and U3023 (N_3023,N_2672,N_2766);
nand U3024 (N_3024,N_2054,N_2797);
nand U3025 (N_3025,N_2892,N_2467);
nor U3026 (N_3026,N_2003,N_2938);
xnor U3027 (N_3027,N_2404,N_2771);
or U3028 (N_3028,N_2448,N_2517);
nor U3029 (N_3029,N_2760,N_2894);
and U3030 (N_3030,N_2913,N_2808);
nor U3031 (N_3031,N_2562,N_2280);
and U3032 (N_3032,N_2705,N_2832);
nor U3033 (N_3033,N_2743,N_2897);
xor U3034 (N_3034,N_2460,N_2273);
xnor U3035 (N_3035,N_2606,N_2558);
or U3036 (N_3036,N_2095,N_2489);
or U3037 (N_3037,N_2851,N_2034);
or U3038 (N_3038,N_2927,N_2485);
nor U3039 (N_3039,N_2663,N_2309);
and U3040 (N_3040,N_2285,N_2709);
nand U3041 (N_3041,N_2695,N_2341);
or U3042 (N_3042,N_2845,N_2998);
and U3043 (N_3043,N_2077,N_2445);
nand U3044 (N_3044,N_2856,N_2936);
nor U3045 (N_3045,N_2608,N_2735);
nand U3046 (N_3046,N_2949,N_2532);
or U3047 (N_3047,N_2660,N_2814);
nand U3048 (N_3048,N_2850,N_2506);
nand U3049 (N_3049,N_2964,N_2066);
or U3050 (N_3050,N_2710,N_2590);
nor U3051 (N_3051,N_2393,N_2935);
or U3052 (N_3052,N_2161,N_2314);
and U3053 (N_3053,N_2711,N_2177);
nor U3054 (N_3054,N_2075,N_2300);
nor U3055 (N_3055,N_2728,N_2362);
or U3056 (N_3056,N_2693,N_2138);
nor U3057 (N_3057,N_2875,N_2466);
nand U3058 (N_3058,N_2376,N_2871);
and U3059 (N_3059,N_2768,N_2505);
nor U3060 (N_3060,N_2333,N_2626);
xnor U3061 (N_3061,N_2566,N_2046);
nor U3062 (N_3062,N_2529,N_2584);
nor U3063 (N_3063,N_2097,N_2407);
or U3064 (N_3064,N_2587,N_2270);
or U3065 (N_3065,N_2205,N_2304);
and U3066 (N_3066,N_2675,N_2086);
or U3067 (N_3067,N_2188,N_2109);
and U3068 (N_3068,N_2206,N_2642);
and U3069 (N_3069,N_2761,N_2245);
xor U3070 (N_3070,N_2495,N_2120);
and U3071 (N_3071,N_2523,N_2960);
or U3072 (N_3072,N_2745,N_2018);
nand U3073 (N_3073,N_2346,N_2547);
nand U3074 (N_3074,N_2794,N_2221);
xnor U3075 (N_3075,N_2516,N_2127);
or U3076 (N_3076,N_2037,N_2342);
and U3077 (N_3077,N_2806,N_2176);
nand U3078 (N_3078,N_2607,N_2546);
or U3079 (N_3079,N_2818,N_2671);
nand U3080 (N_3080,N_2948,N_2282);
xor U3081 (N_3081,N_2873,N_2275);
and U3082 (N_3082,N_2307,N_2480);
and U3083 (N_3083,N_2380,N_2576);
or U3084 (N_3084,N_2396,N_2701);
or U3085 (N_3085,N_2373,N_2315);
or U3086 (N_3086,N_2021,N_2996);
or U3087 (N_3087,N_2030,N_2817);
and U3088 (N_3088,N_2085,N_2852);
nand U3089 (N_3089,N_2464,N_2024);
xnor U3090 (N_3090,N_2919,N_2169);
nand U3091 (N_3091,N_2223,N_2604);
nand U3092 (N_3092,N_2782,N_2289);
and U3093 (N_3093,N_2764,N_2661);
or U3094 (N_3094,N_2906,N_2972);
nor U3095 (N_3095,N_2349,N_2416);
or U3096 (N_3096,N_2385,N_2147);
nor U3097 (N_3097,N_2681,N_2124);
and U3098 (N_3098,N_2488,N_2718);
nor U3099 (N_3099,N_2637,N_2890);
and U3100 (N_3100,N_2830,N_2165);
xor U3101 (N_3101,N_2867,N_2070);
xor U3102 (N_3102,N_2599,N_2081);
and U3103 (N_3103,N_2905,N_2235);
nor U3104 (N_3104,N_2211,N_2345);
or U3105 (N_3105,N_2552,N_2049);
or U3106 (N_3106,N_2820,N_2847);
and U3107 (N_3107,N_2633,N_2719);
or U3108 (N_3108,N_2076,N_2225);
xor U3109 (N_3109,N_2178,N_2277);
nand U3110 (N_3110,N_2550,N_2295);
nand U3111 (N_3111,N_2048,N_2459);
xor U3112 (N_3112,N_2943,N_2478);
or U3113 (N_3113,N_2572,N_2180);
or U3114 (N_3114,N_2813,N_2944);
or U3115 (N_3115,N_2585,N_2252);
or U3116 (N_3116,N_2363,N_2163);
xor U3117 (N_3117,N_2833,N_2332);
or U3118 (N_3118,N_2627,N_2187);
nand U3119 (N_3119,N_2405,N_2296);
xnor U3120 (N_3120,N_2423,N_2792);
nor U3121 (N_3121,N_2412,N_2997);
nand U3122 (N_3122,N_2580,N_2593);
nand U3123 (N_3123,N_2962,N_2511);
nor U3124 (N_3124,N_2402,N_2611);
nand U3125 (N_3125,N_2952,N_2185);
and U3126 (N_3126,N_2539,N_2614);
or U3127 (N_3127,N_2381,N_2911);
nand U3128 (N_3128,N_2917,N_2364);
and U3129 (N_3129,N_2146,N_2053);
nor U3130 (N_3130,N_2266,N_2438);
xnor U3131 (N_3131,N_2561,N_2741);
or U3132 (N_3132,N_2502,N_2248);
or U3133 (N_3133,N_2533,N_2787);
nor U3134 (N_3134,N_2522,N_2953);
nor U3135 (N_3135,N_2189,N_2195);
nand U3136 (N_3136,N_2486,N_2645);
nor U3137 (N_3137,N_2630,N_2411);
nor U3138 (N_3138,N_2099,N_2201);
xor U3139 (N_3139,N_2876,N_2389);
or U3140 (N_3140,N_2019,N_2704);
nand U3141 (N_3141,N_2916,N_2754);
nor U3142 (N_3142,N_2612,N_2586);
or U3143 (N_3143,N_2014,N_2549);
nand U3144 (N_3144,N_2837,N_2094);
nor U3145 (N_3145,N_2560,N_2375);
and U3146 (N_3146,N_2118,N_2141);
nor U3147 (N_3147,N_2135,N_2733);
xor U3148 (N_3148,N_2625,N_2443);
nand U3149 (N_3149,N_2433,N_2765);
or U3150 (N_3150,N_2592,N_2357);
xor U3151 (N_3151,N_2801,N_2702);
nand U3152 (N_3152,N_2676,N_2656);
xor U3153 (N_3153,N_2781,N_2924);
or U3154 (N_3154,N_2134,N_2999);
and U3155 (N_3155,N_2929,N_2976);
nand U3156 (N_3156,N_2057,N_2214);
or U3157 (N_3157,N_2720,N_2531);
or U3158 (N_3158,N_2391,N_2022);
nand U3159 (N_3159,N_2267,N_2629);
xnor U3160 (N_3160,N_2060,N_2634);
or U3161 (N_3161,N_2666,N_2199);
and U3162 (N_3162,N_2064,N_2736);
or U3163 (N_3163,N_2468,N_2058);
nand U3164 (N_3164,N_2993,N_2893);
or U3165 (N_3165,N_2356,N_2481);
nand U3166 (N_3166,N_2687,N_2113);
nand U3167 (N_3167,N_2647,N_2012);
and U3168 (N_3168,N_2888,N_2811);
xnor U3169 (N_3169,N_2975,N_2853);
or U3170 (N_3170,N_2131,N_2145);
nor U3171 (N_3171,N_2330,N_2398);
or U3172 (N_3172,N_2657,N_2017);
or U3173 (N_3173,N_2286,N_2355);
nor U3174 (N_3174,N_2759,N_2716);
nor U3175 (N_3175,N_2040,N_2013);
nor U3176 (N_3176,N_2238,N_2490);
nor U3177 (N_3177,N_2557,N_2703);
nor U3178 (N_3178,N_2940,N_2848);
nor U3179 (N_3179,N_2035,N_2351);
nand U3180 (N_3180,N_2181,N_2653);
nand U3181 (N_3181,N_2100,N_2617);
nor U3182 (N_3182,N_2877,N_2780);
and U3183 (N_3183,N_2966,N_2168);
and U3184 (N_3184,N_2925,N_2762);
and U3185 (N_3185,N_2712,N_2954);
nand U3186 (N_3186,N_2664,N_2827);
and U3187 (N_3187,N_2139,N_2475);
nor U3188 (N_3188,N_2023,N_2191);
nor U3189 (N_3189,N_2928,N_2909);
nor U3190 (N_3190,N_2518,N_2287);
nand U3191 (N_3191,N_2117,N_2903);
nand U3192 (N_3192,N_2153,N_2419);
nand U3193 (N_3193,N_2338,N_2155);
xnor U3194 (N_3194,N_2440,N_2254);
or U3195 (N_3195,N_2209,N_2902);
and U3196 (N_3196,N_2541,N_2707);
xnor U3197 (N_3197,N_2990,N_2912);
or U3198 (N_3198,N_2937,N_2544);
nor U3199 (N_3199,N_2150,N_2470);
and U3200 (N_3200,N_2869,N_2706);
nor U3201 (N_3201,N_2449,N_2096);
nor U3202 (N_3202,N_2669,N_2260);
nand U3203 (N_3203,N_2821,N_2933);
xnor U3204 (N_3204,N_2750,N_2644);
and U3205 (N_3205,N_2497,N_2567);
nand U3206 (N_3206,N_2812,N_2403);
nor U3207 (N_3207,N_2824,N_2878);
nand U3208 (N_3208,N_2788,N_2991);
xnor U3209 (N_3209,N_2620,N_2172);
nor U3210 (N_3210,N_2029,N_2215);
nor U3211 (N_3211,N_2027,N_2261);
and U3212 (N_3212,N_2965,N_2374);
xor U3213 (N_3213,N_2388,N_2854);
and U3214 (N_3214,N_2898,N_2320);
nand U3215 (N_3215,N_2233,N_2978);
nor U3216 (N_3216,N_2425,N_2281);
or U3217 (N_3217,N_2082,N_2294);
nand U3218 (N_3218,N_2746,N_2088);
and U3219 (N_3219,N_2640,N_2006);
and U3220 (N_3220,N_2317,N_2957);
or U3221 (N_3221,N_2756,N_2297);
or U3222 (N_3222,N_2025,N_2526);
and U3223 (N_3223,N_2540,N_2200);
or U3224 (N_3224,N_2000,N_2484);
or U3225 (N_3225,N_2222,N_2390);
and U3226 (N_3226,N_2078,N_2900);
nand U3227 (N_3227,N_2598,N_2779);
and U3228 (N_3228,N_2213,N_2578);
nand U3229 (N_3229,N_2887,N_2011);
or U3230 (N_3230,N_2622,N_2713);
nand U3231 (N_3231,N_2417,N_2968);
or U3232 (N_3232,N_2319,N_2044);
nand U3233 (N_3233,N_2548,N_2646);
nand U3234 (N_3234,N_2239,N_2520);
nor U3235 (N_3235,N_2828,N_2154);
and U3236 (N_3236,N_2510,N_2482);
nand U3237 (N_3237,N_2989,N_2372);
and U3238 (N_3238,N_2302,N_2982);
xnor U3239 (N_3239,N_2588,N_2104);
and U3240 (N_3240,N_2737,N_2184);
or U3241 (N_3241,N_2729,N_2748);
and U3242 (N_3242,N_2446,N_2822);
and U3243 (N_3243,N_2083,N_2202);
and U3244 (N_3244,N_2757,N_2228);
xor U3245 (N_3245,N_2148,N_2730);
nor U3246 (N_3246,N_2959,N_2427);
nor U3247 (N_3247,N_2431,N_2512);
xor U3248 (N_3248,N_2359,N_2524);
nand U3249 (N_3249,N_2501,N_2268);
and U3250 (N_3250,N_2802,N_2435);
or U3251 (N_3251,N_2008,N_2253);
and U3252 (N_3252,N_2399,N_2474);
nand U3253 (N_3253,N_2734,N_2103);
nand U3254 (N_3254,N_2951,N_2236);
and U3255 (N_3255,N_2092,N_2331);
nor U3256 (N_3256,N_2366,N_2090);
nand U3257 (N_3257,N_2908,N_2047);
and U3258 (N_3258,N_2799,N_2721);
nor U3259 (N_3259,N_2891,N_2815);
and U3260 (N_3260,N_2934,N_2441);
and U3261 (N_3261,N_2545,N_2932);
nand U3262 (N_3262,N_2122,N_2093);
and U3263 (N_3263,N_2564,N_2665);
and U3264 (N_3264,N_2860,N_2283);
or U3265 (N_3265,N_2826,N_2969);
nor U3266 (N_3266,N_2983,N_2456);
nor U3267 (N_3267,N_2377,N_2152);
nand U3268 (N_3268,N_2408,N_2955);
nor U3269 (N_3269,N_2472,N_2678);
and U3270 (N_3270,N_2498,N_2256);
nor U3271 (N_3271,N_2192,N_2834);
or U3272 (N_3272,N_2062,N_2328);
nand U3273 (N_3273,N_2559,N_2793);
or U3274 (N_3274,N_2609,N_2308);
nand U3275 (N_3275,N_2946,N_2595);
nor U3276 (N_3276,N_2920,N_2007);
nor U3277 (N_3277,N_2386,N_2068);
nand U3278 (N_3278,N_2487,N_2504);
xor U3279 (N_3279,N_2123,N_2002);
nand U3280 (N_3280,N_2800,N_2084);
xnor U3281 (N_3281,N_2218,N_2310);
nand U3282 (N_3282,N_2984,N_2739);
and U3283 (N_3283,N_2543,N_2112);
or U3284 (N_3284,N_2872,N_2028);
nor U3285 (N_3285,N_2732,N_2325);
nor U3286 (N_3286,N_2740,N_2795);
and U3287 (N_3287,N_2855,N_2571);
xor U3288 (N_3288,N_2409,N_2130);
xor U3289 (N_3289,N_2784,N_2473);
xnor U3290 (N_3290,N_2778,N_2686);
and U3291 (N_3291,N_2265,N_2447);
and U3292 (N_3292,N_2400,N_2079);
xor U3293 (N_3293,N_2167,N_2465);
nand U3294 (N_3294,N_2382,N_2941);
nor U3295 (N_3295,N_2414,N_2785);
xor U3296 (N_3296,N_2031,N_2859);
nor U3297 (N_3297,N_2350,N_2910);
nor U3298 (N_3298,N_2683,N_2080);
or U3299 (N_3299,N_2662,N_2271);
nand U3300 (N_3300,N_2866,N_2881);
nor U3301 (N_3301,N_2336,N_2573);
xnor U3302 (N_3302,N_2263,N_2212);
or U3303 (N_3303,N_2335,N_2536);
nor U3304 (N_3304,N_2643,N_2581);
or U3305 (N_3305,N_2886,N_2884);
nand U3306 (N_3306,N_2752,N_2655);
nor U3307 (N_3307,N_2110,N_2186);
nand U3308 (N_3308,N_2950,N_2776);
nand U3309 (N_3309,N_2243,N_2798);
nor U3310 (N_3310,N_2641,N_2603);
nand U3311 (N_3311,N_2742,N_2995);
nand U3312 (N_3312,N_2810,N_2918);
and U3313 (N_3313,N_2458,N_2160);
and U3314 (N_3314,N_2428,N_2885);
xnor U3315 (N_3315,N_2190,N_2791);
nand U3316 (N_3316,N_2005,N_2981);
and U3317 (N_3317,N_2652,N_2985);
and U3318 (N_3318,N_2437,N_2542);
and U3319 (N_3319,N_2923,N_2136);
and U3320 (N_3320,N_2858,N_2582);
and U3321 (N_3321,N_2065,N_2334);
and U3322 (N_3322,N_2554,N_2224);
or U3323 (N_3323,N_2220,N_2203);
nand U3324 (N_3324,N_2673,N_2444);
or U3325 (N_3325,N_2422,N_2324);
xnor U3326 (N_3326,N_2565,N_2026);
nand U3327 (N_3327,N_2279,N_2537);
nor U3328 (N_3328,N_2326,N_2763);
nand U3329 (N_3329,N_2128,N_2628);
and U3330 (N_3330,N_2074,N_2731);
nand U3331 (N_3331,N_2455,N_2208);
nor U3332 (N_3332,N_2632,N_2312);
nand U3333 (N_3333,N_2570,N_2353);
nand U3334 (N_3334,N_2259,N_2365);
nor U3335 (N_3335,N_2901,N_2668);
nand U3336 (N_3336,N_2288,N_2809);
nor U3337 (N_3337,N_2257,N_2613);
and U3338 (N_3338,N_2973,N_2864);
nand U3339 (N_3339,N_2457,N_2773);
nand U3340 (N_3340,N_2667,N_2463);
or U3341 (N_3341,N_2204,N_2251);
or U3342 (N_3342,N_2922,N_2921);
nor U3343 (N_3343,N_2553,N_2738);
nor U3344 (N_3344,N_2835,N_2111);
nand U3345 (N_3345,N_2749,N_2605);
nor U3346 (N_3346,N_2970,N_2831);
nor U3347 (N_3347,N_2509,N_2020);
nor U3348 (N_3348,N_2726,N_2247);
or U3349 (N_3349,N_2825,N_2072);
nand U3350 (N_3350,N_2383,N_2210);
nor U3351 (N_3351,N_2418,N_2140);
nand U3352 (N_3352,N_2692,N_2839);
or U3353 (N_3353,N_2597,N_2159);
nor U3354 (N_3354,N_2197,N_2685);
nor U3355 (N_3355,N_2945,N_2977);
nor U3356 (N_3356,N_2722,N_2636);
xor U3357 (N_3357,N_2971,N_2395);
and U3358 (N_3358,N_2694,N_2410);
nand U3359 (N_3359,N_2508,N_2525);
nor U3360 (N_3360,N_2994,N_2619);
nor U3361 (N_3361,N_2819,N_2535);
nor U3362 (N_3362,N_2930,N_2471);
nor U3363 (N_3363,N_2514,N_2454);
nand U3364 (N_3364,N_2513,N_2004);
nand U3365 (N_3365,N_2434,N_2250);
nand U3366 (N_3366,N_2615,N_2105);
and U3367 (N_3367,N_2610,N_2045);
nand U3368 (N_3368,N_2337,N_2796);
nand U3369 (N_3369,N_2618,N_2521);
xnor U3370 (N_3370,N_2358,N_2313);
xnor U3371 (N_3371,N_2861,N_2496);
nor U3372 (N_3372,N_2836,N_2469);
xor U3373 (N_3373,N_2352,N_2115);
or U3374 (N_3374,N_2714,N_2050);
and U3375 (N_3375,N_2479,N_2804);
nor U3376 (N_3376,N_2439,N_2631);
and U3377 (N_3377,N_2988,N_2538);
xnor U3378 (N_3378,N_2067,N_2596);
nor U3379 (N_3379,N_2551,N_2098);
nand U3380 (N_3380,N_2616,N_2432);
nand U3381 (N_3381,N_2882,N_2394);
nand U3382 (N_3382,N_2226,N_2194);
and U3383 (N_3383,N_2575,N_2001);
or U3384 (N_3384,N_2149,N_2747);
or U3385 (N_3385,N_2865,N_2717);
or U3386 (N_3386,N_2144,N_2967);
nand U3387 (N_3387,N_2670,N_2016);
and U3388 (N_3388,N_2591,N_2244);
xor U3389 (N_3389,N_2883,N_2689);
and U3390 (N_3390,N_2166,N_2777);
nand U3391 (N_3391,N_2725,N_2579);
nor U3392 (N_3392,N_2413,N_2369);
nand U3393 (N_3393,N_2143,N_2829);
nor U3394 (N_3394,N_2121,N_2298);
or U3395 (N_3395,N_2360,N_2451);
or U3396 (N_3396,N_2574,N_2370);
xor U3397 (N_3397,N_2158,N_2368);
or U3398 (N_3398,N_2175,N_2102);
and U3399 (N_3399,N_2316,N_2174);
nand U3400 (N_3400,N_2769,N_2805);
and U3401 (N_3401,N_2089,N_2624);
and U3402 (N_3402,N_2217,N_2361);
nand U3403 (N_3403,N_2033,N_2401);
and U3404 (N_3404,N_2862,N_2758);
nor U3405 (N_3405,N_2556,N_2684);
or U3406 (N_3406,N_2931,N_2715);
or U3407 (N_3407,N_2503,N_2183);
or U3408 (N_3408,N_2107,N_2327);
nand U3409 (N_3409,N_2568,N_2601);
and U3410 (N_3410,N_2043,N_2216);
or U3411 (N_3411,N_2173,N_2677);
nor U3412 (N_3412,N_2262,N_2880);
and U3413 (N_3413,N_2198,N_2406);
or U3414 (N_3414,N_2230,N_2914);
or U3415 (N_3415,N_2339,N_2106);
and U3416 (N_3416,N_2171,N_2041);
and U3417 (N_3417,N_2698,N_2986);
xor U3418 (N_3418,N_2563,N_2430);
nor U3419 (N_3419,N_2032,N_2322);
and U3420 (N_3420,N_2116,N_2980);
xnor U3421 (N_3421,N_2038,N_2274);
nand U3422 (N_3422,N_2649,N_2291);
nor U3423 (N_3423,N_2042,N_2392);
nand U3424 (N_3424,N_2863,N_2700);
nand U3425 (N_3425,N_2182,N_2240);
and U3426 (N_3426,N_2699,N_2963);
and U3427 (N_3427,N_2772,N_2589);
or U3428 (N_3428,N_2691,N_2528);
nor U3429 (N_3429,N_2242,N_2193);
nor U3430 (N_3430,N_2269,N_2857);
nand U3431 (N_3431,N_2114,N_2009);
nand U3432 (N_3432,N_2690,N_2841);
and U3433 (N_3433,N_2843,N_2823);
and U3434 (N_3434,N_2142,N_2483);
nand U3435 (N_3435,N_2602,N_2290);
nand U3436 (N_3436,N_2284,N_2774);
or U3437 (N_3437,N_2534,N_2491);
nor U3438 (N_3438,N_2219,N_2753);
or U3439 (N_3439,N_2091,N_2623);
and U3440 (N_3440,N_2477,N_2056);
or U3441 (N_3441,N_2429,N_2846);
nand U3442 (N_3442,N_2237,N_2087);
or U3443 (N_3443,N_2807,N_2723);
nor U3444 (N_3444,N_2442,N_2958);
nand U3445 (N_3445,N_2132,N_2415);
nor U3446 (N_3446,N_2530,N_2650);
and U3447 (N_3447,N_2974,N_2870);
or U3448 (N_3448,N_2305,N_2674);
and U3449 (N_3449,N_2119,N_2942);
xnor U3450 (N_3450,N_2476,N_2515);
and U3451 (N_3451,N_2051,N_2299);
nor U3452 (N_3452,N_2895,N_2987);
xnor U3453 (N_3453,N_2790,N_2126);
nand U3454 (N_3454,N_2724,N_2426);
nand U3455 (N_3455,N_2755,N_2680);
and U3456 (N_3456,N_2323,N_2679);
xnor U3457 (N_3457,N_2272,N_2436);
and U3458 (N_3458,N_2232,N_2499);
nor U3459 (N_3459,N_2688,N_2329);
xor U3460 (N_3460,N_2697,N_2621);
and U3461 (N_3461,N_2844,N_2378);
or U3462 (N_3462,N_2635,N_2264);
nand U3463 (N_3463,N_2569,N_2751);
xor U3464 (N_3464,N_2170,N_2292);
or U3465 (N_3465,N_2770,N_2639);
nand U3466 (N_3466,N_2727,N_2179);
and U3467 (N_3467,N_2527,N_2947);
or U3468 (N_3468,N_2354,N_2849);
nand U3469 (N_3469,N_2384,N_2583);
or U3470 (N_3470,N_2073,N_2696);
xnor U3471 (N_3471,N_2293,N_2507);
nor U3472 (N_3472,N_2654,N_2816);
nor U3473 (N_3473,N_2783,N_2493);
and U3474 (N_3474,N_2904,N_2803);
and U3475 (N_3475,N_2879,N_2889);
and U3476 (N_3476,N_2421,N_2129);
nor U3477 (N_3477,N_2992,N_2063);
and U3478 (N_3478,N_2241,N_2069);
or U3479 (N_3479,N_2157,N_2397);
or U3480 (N_3480,N_2151,N_2775);
xnor U3481 (N_3481,N_2789,N_2899);
or U3482 (N_3482,N_2249,N_2961);
nand U3483 (N_3483,N_2926,N_2915);
nor U3484 (N_3484,N_2231,N_2344);
nor U3485 (N_3485,N_2303,N_2071);
nand U3486 (N_3486,N_2318,N_2868);
xor U3487 (N_3487,N_2648,N_2207);
nand U3488 (N_3488,N_2306,N_2956);
nor U3489 (N_3489,N_2651,N_2196);
nand U3490 (N_3490,N_2682,N_2658);
or U3491 (N_3491,N_2321,N_2594);
and U3492 (N_3492,N_2453,N_2278);
nand U3493 (N_3493,N_2348,N_2164);
nor U3494 (N_3494,N_2708,N_2494);
or U3495 (N_3495,N_2137,N_2424);
nand U3496 (N_3496,N_2492,N_2036);
nand U3497 (N_3497,N_2101,N_2052);
or U3498 (N_3498,N_2939,N_2156);
or U3499 (N_3499,N_2125,N_2258);
and U3500 (N_3500,N_2594,N_2468);
and U3501 (N_3501,N_2070,N_2388);
and U3502 (N_3502,N_2228,N_2189);
nand U3503 (N_3503,N_2170,N_2948);
xnor U3504 (N_3504,N_2771,N_2836);
and U3505 (N_3505,N_2996,N_2214);
or U3506 (N_3506,N_2227,N_2199);
or U3507 (N_3507,N_2999,N_2309);
or U3508 (N_3508,N_2863,N_2517);
nand U3509 (N_3509,N_2309,N_2666);
nand U3510 (N_3510,N_2620,N_2664);
or U3511 (N_3511,N_2741,N_2336);
nand U3512 (N_3512,N_2745,N_2045);
and U3513 (N_3513,N_2877,N_2670);
and U3514 (N_3514,N_2474,N_2779);
nor U3515 (N_3515,N_2189,N_2134);
or U3516 (N_3516,N_2930,N_2321);
and U3517 (N_3517,N_2703,N_2502);
or U3518 (N_3518,N_2468,N_2151);
and U3519 (N_3519,N_2706,N_2283);
and U3520 (N_3520,N_2242,N_2037);
nor U3521 (N_3521,N_2567,N_2595);
nand U3522 (N_3522,N_2565,N_2786);
or U3523 (N_3523,N_2121,N_2504);
nand U3524 (N_3524,N_2993,N_2639);
or U3525 (N_3525,N_2589,N_2831);
nand U3526 (N_3526,N_2375,N_2196);
nor U3527 (N_3527,N_2466,N_2788);
and U3528 (N_3528,N_2729,N_2256);
nor U3529 (N_3529,N_2490,N_2207);
or U3530 (N_3530,N_2795,N_2159);
and U3531 (N_3531,N_2892,N_2461);
nor U3532 (N_3532,N_2132,N_2549);
and U3533 (N_3533,N_2605,N_2193);
nor U3534 (N_3534,N_2320,N_2662);
or U3535 (N_3535,N_2383,N_2342);
and U3536 (N_3536,N_2962,N_2286);
nor U3537 (N_3537,N_2345,N_2454);
nor U3538 (N_3538,N_2863,N_2572);
or U3539 (N_3539,N_2901,N_2530);
or U3540 (N_3540,N_2313,N_2676);
or U3541 (N_3541,N_2897,N_2359);
nor U3542 (N_3542,N_2290,N_2940);
or U3543 (N_3543,N_2996,N_2367);
nor U3544 (N_3544,N_2466,N_2707);
nor U3545 (N_3545,N_2190,N_2264);
or U3546 (N_3546,N_2037,N_2045);
nor U3547 (N_3547,N_2187,N_2987);
nor U3548 (N_3548,N_2012,N_2013);
nor U3549 (N_3549,N_2015,N_2283);
or U3550 (N_3550,N_2250,N_2323);
or U3551 (N_3551,N_2798,N_2291);
xnor U3552 (N_3552,N_2041,N_2911);
nor U3553 (N_3553,N_2616,N_2399);
nor U3554 (N_3554,N_2790,N_2791);
and U3555 (N_3555,N_2031,N_2625);
or U3556 (N_3556,N_2150,N_2945);
nand U3557 (N_3557,N_2387,N_2739);
nor U3558 (N_3558,N_2628,N_2007);
xor U3559 (N_3559,N_2826,N_2424);
nor U3560 (N_3560,N_2634,N_2997);
xor U3561 (N_3561,N_2618,N_2361);
nor U3562 (N_3562,N_2558,N_2369);
nand U3563 (N_3563,N_2116,N_2435);
nor U3564 (N_3564,N_2157,N_2330);
or U3565 (N_3565,N_2968,N_2217);
or U3566 (N_3566,N_2427,N_2703);
or U3567 (N_3567,N_2314,N_2037);
and U3568 (N_3568,N_2626,N_2107);
nand U3569 (N_3569,N_2851,N_2254);
nor U3570 (N_3570,N_2275,N_2041);
and U3571 (N_3571,N_2110,N_2048);
or U3572 (N_3572,N_2485,N_2040);
nor U3573 (N_3573,N_2777,N_2419);
or U3574 (N_3574,N_2853,N_2098);
or U3575 (N_3575,N_2689,N_2146);
nand U3576 (N_3576,N_2918,N_2771);
and U3577 (N_3577,N_2159,N_2101);
and U3578 (N_3578,N_2966,N_2167);
xnor U3579 (N_3579,N_2397,N_2278);
nor U3580 (N_3580,N_2381,N_2076);
nand U3581 (N_3581,N_2701,N_2640);
nand U3582 (N_3582,N_2806,N_2377);
xor U3583 (N_3583,N_2565,N_2516);
nor U3584 (N_3584,N_2197,N_2454);
and U3585 (N_3585,N_2385,N_2764);
nand U3586 (N_3586,N_2712,N_2970);
nand U3587 (N_3587,N_2755,N_2926);
or U3588 (N_3588,N_2480,N_2233);
and U3589 (N_3589,N_2653,N_2534);
nand U3590 (N_3590,N_2578,N_2923);
nor U3591 (N_3591,N_2999,N_2055);
nor U3592 (N_3592,N_2228,N_2623);
xor U3593 (N_3593,N_2624,N_2398);
nor U3594 (N_3594,N_2347,N_2948);
nand U3595 (N_3595,N_2934,N_2341);
and U3596 (N_3596,N_2260,N_2306);
xnor U3597 (N_3597,N_2069,N_2106);
xnor U3598 (N_3598,N_2954,N_2251);
and U3599 (N_3599,N_2628,N_2544);
nor U3600 (N_3600,N_2260,N_2280);
nand U3601 (N_3601,N_2061,N_2031);
nor U3602 (N_3602,N_2446,N_2338);
xnor U3603 (N_3603,N_2531,N_2494);
nor U3604 (N_3604,N_2513,N_2592);
nor U3605 (N_3605,N_2564,N_2402);
xnor U3606 (N_3606,N_2370,N_2014);
nor U3607 (N_3607,N_2391,N_2467);
and U3608 (N_3608,N_2129,N_2771);
and U3609 (N_3609,N_2498,N_2016);
nor U3610 (N_3610,N_2357,N_2678);
xor U3611 (N_3611,N_2098,N_2319);
nand U3612 (N_3612,N_2271,N_2132);
and U3613 (N_3613,N_2613,N_2733);
xnor U3614 (N_3614,N_2975,N_2665);
and U3615 (N_3615,N_2467,N_2404);
and U3616 (N_3616,N_2462,N_2648);
nor U3617 (N_3617,N_2670,N_2593);
or U3618 (N_3618,N_2271,N_2068);
xnor U3619 (N_3619,N_2158,N_2787);
or U3620 (N_3620,N_2851,N_2016);
nand U3621 (N_3621,N_2974,N_2299);
nand U3622 (N_3622,N_2308,N_2606);
and U3623 (N_3623,N_2127,N_2277);
or U3624 (N_3624,N_2292,N_2905);
nor U3625 (N_3625,N_2166,N_2121);
or U3626 (N_3626,N_2090,N_2193);
or U3627 (N_3627,N_2787,N_2903);
or U3628 (N_3628,N_2329,N_2359);
nand U3629 (N_3629,N_2783,N_2822);
nor U3630 (N_3630,N_2109,N_2925);
or U3631 (N_3631,N_2196,N_2478);
nor U3632 (N_3632,N_2359,N_2685);
nor U3633 (N_3633,N_2722,N_2887);
nand U3634 (N_3634,N_2079,N_2433);
or U3635 (N_3635,N_2866,N_2697);
and U3636 (N_3636,N_2375,N_2558);
or U3637 (N_3637,N_2671,N_2878);
nor U3638 (N_3638,N_2755,N_2613);
nor U3639 (N_3639,N_2490,N_2289);
and U3640 (N_3640,N_2143,N_2950);
nand U3641 (N_3641,N_2234,N_2829);
nor U3642 (N_3642,N_2785,N_2954);
nand U3643 (N_3643,N_2187,N_2109);
xor U3644 (N_3644,N_2041,N_2876);
xnor U3645 (N_3645,N_2513,N_2102);
or U3646 (N_3646,N_2431,N_2233);
xnor U3647 (N_3647,N_2212,N_2941);
nor U3648 (N_3648,N_2286,N_2670);
nand U3649 (N_3649,N_2202,N_2674);
or U3650 (N_3650,N_2960,N_2135);
nand U3651 (N_3651,N_2186,N_2343);
xor U3652 (N_3652,N_2882,N_2760);
nor U3653 (N_3653,N_2283,N_2775);
or U3654 (N_3654,N_2172,N_2438);
and U3655 (N_3655,N_2664,N_2593);
and U3656 (N_3656,N_2627,N_2138);
xnor U3657 (N_3657,N_2177,N_2577);
nor U3658 (N_3658,N_2376,N_2725);
or U3659 (N_3659,N_2598,N_2092);
or U3660 (N_3660,N_2236,N_2806);
and U3661 (N_3661,N_2965,N_2758);
and U3662 (N_3662,N_2101,N_2181);
nand U3663 (N_3663,N_2289,N_2270);
or U3664 (N_3664,N_2131,N_2423);
xnor U3665 (N_3665,N_2397,N_2314);
xnor U3666 (N_3666,N_2092,N_2464);
or U3667 (N_3667,N_2544,N_2859);
and U3668 (N_3668,N_2961,N_2127);
and U3669 (N_3669,N_2322,N_2402);
nor U3670 (N_3670,N_2398,N_2241);
xor U3671 (N_3671,N_2450,N_2501);
nor U3672 (N_3672,N_2833,N_2368);
nand U3673 (N_3673,N_2218,N_2094);
and U3674 (N_3674,N_2633,N_2021);
nand U3675 (N_3675,N_2627,N_2059);
nor U3676 (N_3676,N_2801,N_2887);
and U3677 (N_3677,N_2797,N_2676);
nand U3678 (N_3678,N_2458,N_2674);
or U3679 (N_3679,N_2363,N_2261);
nand U3680 (N_3680,N_2418,N_2529);
nand U3681 (N_3681,N_2545,N_2227);
nand U3682 (N_3682,N_2886,N_2261);
or U3683 (N_3683,N_2543,N_2582);
and U3684 (N_3684,N_2977,N_2229);
or U3685 (N_3685,N_2927,N_2246);
nand U3686 (N_3686,N_2322,N_2310);
and U3687 (N_3687,N_2875,N_2835);
nor U3688 (N_3688,N_2553,N_2381);
and U3689 (N_3689,N_2779,N_2790);
or U3690 (N_3690,N_2092,N_2854);
and U3691 (N_3691,N_2123,N_2493);
and U3692 (N_3692,N_2568,N_2490);
nand U3693 (N_3693,N_2066,N_2521);
and U3694 (N_3694,N_2689,N_2196);
and U3695 (N_3695,N_2797,N_2900);
nand U3696 (N_3696,N_2287,N_2135);
xor U3697 (N_3697,N_2475,N_2979);
nand U3698 (N_3698,N_2393,N_2787);
and U3699 (N_3699,N_2591,N_2607);
or U3700 (N_3700,N_2349,N_2348);
xor U3701 (N_3701,N_2408,N_2081);
nor U3702 (N_3702,N_2342,N_2208);
and U3703 (N_3703,N_2017,N_2520);
or U3704 (N_3704,N_2098,N_2459);
nor U3705 (N_3705,N_2935,N_2562);
nand U3706 (N_3706,N_2604,N_2317);
nor U3707 (N_3707,N_2697,N_2830);
or U3708 (N_3708,N_2844,N_2616);
and U3709 (N_3709,N_2967,N_2172);
or U3710 (N_3710,N_2198,N_2958);
and U3711 (N_3711,N_2026,N_2104);
nor U3712 (N_3712,N_2577,N_2955);
and U3713 (N_3713,N_2083,N_2228);
nor U3714 (N_3714,N_2313,N_2721);
nand U3715 (N_3715,N_2663,N_2514);
xor U3716 (N_3716,N_2977,N_2926);
and U3717 (N_3717,N_2927,N_2801);
nand U3718 (N_3718,N_2598,N_2625);
and U3719 (N_3719,N_2894,N_2897);
nand U3720 (N_3720,N_2111,N_2232);
and U3721 (N_3721,N_2800,N_2622);
or U3722 (N_3722,N_2158,N_2788);
and U3723 (N_3723,N_2412,N_2988);
and U3724 (N_3724,N_2406,N_2938);
nand U3725 (N_3725,N_2515,N_2952);
nand U3726 (N_3726,N_2223,N_2250);
xor U3727 (N_3727,N_2426,N_2372);
or U3728 (N_3728,N_2301,N_2783);
or U3729 (N_3729,N_2499,N_2273);
nand U3730 (N_3730,N_2180,N_2135);
nor U3731 (N_3731,N_2487,N_2955);
xor U3732 (N_3732,N_2563,N_2797);
nand U3733 (N_3733,N_2349,N_2889);
or U3734 (N_3734,N_2941,N_2336);
nand U3735 (N_3735,N_2874,N_2565);
nand U3736 (N_3736,N_2078,N_2488);
nand U3737 (N_3737,N_2957,N_2196);
nand U3738 (N_3738,N_2156,N_2150);
nand U3739 (N_3739,N_2417,N_2768);
nand U3740 (N_3740,N_2504,N_2197);
nor U3741 (N_3741,N_2346,N_2160);
nand U3742 (N_3742,N_2214,N_2134);
nor U3743 (N_3743,N_2934,N_2558);
nor U3744 (N_3744,N_2824,N_2058);
nand U3745 (N_3745,N_2364,N_2845);
nand U3746 (N_3746,N_2440,N_2377);
nand U3747 (N_3747,N_2449,N_2750);
or U3748 (N_3748,N_2526,N_2633);
and U3749 (N_3749,N_2434,N_2921);
xnor U3750 (N_3750,N_2697,N_2726);
nand U3751 (N_3751,N_2909,N_2637);
nor U3752 (N_3752,N_2429,N_2966);
nor U3753 (N_3753,N_2193,N_2208);
or U3754 (N_3754,N_2876,N_2056);
and U3755 (N_3755,N_2144,N_2023);
and U3756 (N_3756,N_2443,N_2621);
or U3757 (N_3757,N_2259,N_2229);
and U3758 (N_3758,N_2339,N_2523);
nor U3759 (N_3759,N_2288,N_2668);
nor U3760 (N_3760,N_2195,N_2221);
nor U3761 (N_3761,N_2957,N_2030);
nand U3762 (N_3762,N_2656,N_2309);
and U3763 (N_3763,N_2483,N_2888);
nor U3764 (N_3764,N_2489,N_2576);
nand U3765 (N_3765,N_2266,N_2863);
nand U3766 (N_3766,N_2956,N_2423);
and U3767 (N_3767,N_2422,N_2940);
xnor U3768 (N_3768,N_2574,N_2149);
nor U3769 (N_3769,N_2539,N_2496);
nand U3770 (N_3770,N_2612,N_2889);
nand U3771 (N_3771,N_2205,N_2611);
xnor U3772 (N_3772,N_2210,N_2816);
nand U3773 (N_3773,N_2531,N_2231);
and U3774 (N_3774,N_2687,N_2562);
nor U3775 (N_3775,N_2068,N_2570);
nor U3776 (N_3776,N_2768,N_2241);
xnor U3777 (N_3777,N_2445,N_2100);
nor U3778 (N_3778,N_2298,N_2748);
and U3779 (N_3779,N_2014,N_2730);
nand U3780 (N_3780,N_2477,N_2513);
nand U3781 (N_3781,N_2321,N_2021);
nor U3782 (N_3782,N_2115,N_2750);
nor U3783 (N_3783,N_2818,N_2591);
nor U3784 (N_3784,N_2955,N_2610);
and U3785 (N_3785,N_2436,N_2561);
and U3786 (N_3786,N_2195,N_2866);
nand U3787 (N_3787,N_2915,N_2616);
nor U3788 (N_3788,N_2256,N_2089);
nand U3789 (N_3789,N_2217,N_2103);
nor U3790 (N_3790,N_2774,N_2105);
and U3791 (N_3791,N_2148,N_2526);
nand U3792 (N_3792,N_2129,N_2516);
and U3793 (N_3793,N_2116,N_2858);
and U3794 (N_3794,N_2130,N_2362);
nand U3795 (N_3795,N_2567,N_2749);
and U3796 (N_3796,N_2224,N_2566);
nor U3797 (N_3797,N_2659,N_2230);
nor U3798 (N_3798,N_2063,N_2874);
xor U3799 (N_3799,N_2942,N_2958);
or U3800 (N_3800,N_2687,N_2466);
nor U3801 (N_3801,N_2789,N_2455);
nor U3802 (N_3802,N_2849,N_2120);
nor U3803 (N_3803,N_2754,N_2725);
and U3804 (N_3804,N_2201,N_2606);
xnor U3805 (N_3805,N_2517,N_2734);
xor U3806 (N_3806,N_2127,N_2103);
and U3807 (N_3807,N_2185,N_2884);
nor U3808 (N_3808,N_2855,N_2585);
nor U3809 (N_3809,N_2762,N_2392);
and U3810 (N_3810,N_2965,N_2538);
or U3811 (N_3811,N_2996,N_2960);
nor U3812 (N_3812,N_2774,N_2448);
xnor U3813 (N_3813,N_2520,N_2189);
nor U3814 (N_3814,N_2968,N_2272);
xnor U3815 (N_3815,N_2744,N_2537);
xor U3816 (N_3816,N_2352,N_2307);
and U3817 (N_3817,N_2861,N_2071);
nor U3818 (N_3818,N_2335,N_2566);
and U3819 (N_3819,N_2641,N_2622);
or U3820 (N_3820,N_2958,N_2033);
nor U3821 (N_3821,N_2462,N_2348);
nand U3822 (N_3822,N_2097,N_2610);
or U3823 (N_3823,N_2932,N_2605);
nor U3824 (N_3824,N_2607,N_2107);
nor U3825 (N_3825,N_2088,N_2698);
nand U3826 (N_3826,N_2490,N_2119);
or U3827 (N_3827,N_2709,N_2708);
or U3828 (N_3828,N_2346,N_2419);
xor U3829 (N_3829,N_2670,N_2496);
nor U3830 (N_3830,N_2414,N_2314);
nor U3831 (N_3831,N_2494,N_2872);
nand U3832 (N_3832,N_2053,N_2652);
or U3833 (N_3833,N_2786,N_2285);
and U3834 (N_3834,N_2642,N_2825);
or U3835 (N_3835,N_2673,N_2381);
and U3836 (N_3836,N_2335,N_2288);
nor U3837 (N_3837,N_2832,N_2085);
and U3838 (N_3838,N_2503,N_2568);
nor U3839 (N_3839,N_2137,N_2657);
and U3840 (N_3840,N_2536,N_2909);
or U3841 (N_3841,N_2690,N_2936);
xnor U3842 (N_3842,N_2635,N_2482);
nor U3843 (N_3843,N_2727,N_2585);
and U3844 (N_3844,N_2939,N_2646);
and U3845 (N_3845,N_2498,N_2422);
nor U3846 (N_3846,N_2272,N_2720);
or U3847 (N_3847,N_2095,N_2610);
nor U3848 (N_3848,N_2487,N_2970);
nand U3849 (N_3849,N_2674,N_2996);
or U3850 (N_3850,N_2278,N_2952);
nand U3851 (N_3851,N_2751,N_2886);
xor U3852 (N_3852,N_2573,N_2461);
or U3853 (N_3853,N_2102,N_2950);
nand U3854 (N_3854,N_2458,N_2708);
or U3855 (N_3855,N_2722,N_2832);
nand U3856 (N_3856,N_2916,N_2434);
or U3857 (N_3857,N_2198,N_2981);
and U3858 (N_3858,N_2794,N_2791);
nand U3859 (N_3859,N_2285,N_2123);
nand U3860 (N_3860,N_2098,N_2653);
and U3861 (N_3861,N_2669,N_2100);
nor U3862 (N_3862,N_2550,N_2267);
and U3863 (N_3863,N_2369,N_2698);
nand U3864 (N_3864,N_2016,N_2514);
nor U3865 (N_3865,N_2855,N_2966);
xnor U3866 (N_3866,N_2220,N_2044);
or U3867 (N_3867,N_2923,N_2572);
nor U3868 (N_3868,N_2577,N_2416);
nand U3869 (N_3869,N_2531,N_2879);
nand U3870 (N_3870,N_2276,N_2352);
nor U3871 (N_3871,N_2792,N_2372);
or U3872 (N_3872,N_2414,N_2382);
and U3873 (N_3873,N_2664,N_2775);
or U3874 (N_3874,N_2454,N_2809);
nand U3875 (N_3875,N_2892,N_2878);
or U3876 (N_3876,N_2418,N_2542);
nand U3877 (N_3877,N_2394,N_2036);
nand U3878 (N_3878,N_2317,N_2520);
xnor U3879 (N_3879,N_2097,N_2016);
nand U3880 (N_3880,N_2610,N_2359);
nor U3881 (N_3881,N_2769,N_2591);
or U3882 (N_3882,N_2244,N_2344);
and U3883 (N_3883,N_2348,N_2957);
nand U3884 (N_3884,N_2894,N_2112);
nor U3885 (N_3885,N_2808,N_2666);
nor U3886 (N_3886,N_2111,N_2328);
nor U3887 (N_3887,N_2262,N_2559);
and U3888 (N_3888,N_2898,N_2056);
or U3889 (N_3889,N_2827,N_2112);
and U3890 (N_3890,N_2175,N_2035);
nand U3891 (N_3891,N_2422,N_2823);
nor U3892 (N_3892,N_2148,N_2421);
nor U3893 (N_3893,N_2721,N_2247);
nand U3894 (N_3894,N_2954,N_2263);
and U3895 (N_3895,N_2752,N_2460);
and U3896 (N_3896,N_2789,N_2237);
nor U3897 (N_3897,N_2752,N_2700);
nor U3898 (N_3898,N_2027,N_2996);
nand U3899 (N_3899,N_2272,N_2577);
nand U3900 (N_3900,N_2917,N_2306);
nand U3901 (N_3901,N_2053,N_2422);
xor U3902 (N_3902,N_2395,N_2356);
nand U3903 (N_3903,N_2564,N_2703);
and U3904 (N_3904,N_2901,N_2182);
nand U3905 (N_3905,N_2546,N_2989);
nand U3906 (N_3906,N_2048,N_2742);
and U3907 (N_3907,N_2609,N_2894);
or U3908 (N_3908,N_2727,N_2458);
or U3909 (N_3909,N_2951,N_2026);
or U3910 (N_3910,N_2474,N_2246);
or U3911 (N_3911,N_2501,N_2021);
nand U3912 (N_3912,N_2890,N_2648);
nand U3913 (N_3913,N_2806,N_2538);
nor U3914 (N_3914,N_2212,N_2309);
xnor U3915 (N_3915,N_2453,N_2097);
nand U3916 (N_3916,N_2642,N_2773);
or U3917 (N_3917,N_2921,N_2231);
nor U3918 (N_3918,N_2440,N_2048);
and U3919 (N_3919,N_2094,N_2227);
nor U3920 (N_3920,N_2085,N_2562);
and U3921 (N_3921,N_2133,N_2170);
nor U3922 (N_3922,N_2821,N_2039);
and U3923 (N_3923,N_2490,N_2329);
or U3924 (N_3924,N_2773,N_2161);
nor U3925 (N_3925,N_2644,N_2634);
and U3926 (N_3926,N_2852,N_2762);
nand U3927 (N_3927,N_2895,N_2852);
or U3928 (N_3928,N_2934,N_2229);
or U3929 (N_3929,N_2970,N_2995);
nand U3930 (N_3930,N_2132,N_2178);
and U3931 (N_3931,N_2998,N_2934);
nand U3932 (N_3932,N_2833,N_2496);
nand U3933 (N_3933,N_2234,N_2179);
and U3934 (N_3934,N_2085,N_2075);
nand U3935 (N_3935,N_2336,N_2239);
xnor U3936 (N_3936,N_2741,N_2028);
nor U3937 (N_3937,N_2612,N_2142);
and U3938 (N_3938,N_2868,N_2060);
nand U3939 (N_3939,N_2988,N_2363);
or U3940 (N_3940,N_2802,N_2465);
nand U3941 (N_3941,N_2770,N_2456);
nand U3942 (N_3942,N_2387,N_2775);
and U3943 (N_3943,N_2343,N_2002);
and U3944 (N_3944,N_2999,N_2074);
and U3945 (N_3945,N_2065,N_2897);
nand U3946 (N_3946,N_2161,N_2572);
or U3947 (N_3947,N_2233,N_2043);
or U3948 (N_3948,N_2247,N_2653);
xnor U3949 (N_3949,N_2555,N_2759);
and U3950 (N_3950,N_2935,N_2464);
or U3951 (N_3951,N_2213,N_2953);
nand U3952 (N_3952,N_2012,N_2637);
nand U3953 (N_3953,N_2682,N_2415);
or U3954 (N_3954,N_2892,N_2288);
nor U3955 (N_3955,N_2479,N_2165);
xnor U3956 (N_3956,N_2556,N_2331);
xor U3957 (N_3957,N_2407,N_2952);
and U3958 (N_3958,N_2011,N_2772);
and U3959 (N_3959,N_2571,N_2070);
nand U3960 (N_3960,N_2669,N_2169);
xor U3961 (N_3961,N_2343,N_2529);
and U3962 (N_3962,N_2565,N_2655);
and U3963 (N_3963,N_2596,N_2242);
nand U3964 (N_3964,N_2850,N_2513);
xor U3965 (N_3965,N_2277,N_2769);
nor U3966 (N_3966,N_2310,N_2963);
and U3967 (N_3967,N_2322,N_2924);
nand U3968 (N_3968,N_2042,N_2793);
nor U3969 (N_3969,N_2699,N_2094);
and U3970 (N_3970,N_2970,N_2899);
nor U3971 (N_3971,N_2943,N_2899);
xnor U3972 (N_3972,N_2971,N_2734);
nand U3973 (N_3973,N_2325,N_2249);
nor U3974 (N_3974,N_2624,N_2190);
or U3975 (N_3975,N_2886,N_2563);
and U3976 (N_3976,N_2283,N_2769);
and U3977 (N_3977,N_2556,N_2830);
or U3978 (N_3978,N_2572,N_2852);
and U3979 (N_3979,N_2558,N_2009);
and U3980 (N_3980,N_2997,N_2932);
and U3981 (N_3981,N_2234,N_2067);
and U3982 (N_3982,N_2047,N_2108);
nor U3983 (N_3983,N_2605,N_2473);
nand U3984 (N_3984,N_2035,N_2482);
or U3985 (N_3985,N_2486,N_2956);
nand U3986 (N_3986,N_2115,N_2571);
nor U3987 (N_3987,N_2066,N_2644);
and U3988 (N_3988,N_2025,N_2044);
or U3989 (N_3989,N_2501,N_2975);
nor U3990 (N_3990,N_2704,N_2214);
nor U3991 (N_3991,N_2060,N_2877);
nor U3992 (N_3992,N_2249,N_2810);
xnor U3993 (N_3993,N_2870,N_2676);
nand U3994 (N_3994,N_2499,N_2916);
or U3995 (N_3995,N_2334,N_2846);
and U3996 (N_3996,N_2966,N_2498);
and U3997 (N_3997,N_2442,N_2351);
or U3998 (N_3998,N_2235,N_2446);
and U3999 (N_3999,N_2573,N_2795);
or U4000 (N_4000,N_3041,N_3024);
nand U4001 (N_4001,N_3536,N_3188);
nor U4002 (N_4002,N_3470,N_3720);
and U4003 (N_4003,N_3394,N_3737);
or U4004 (N_4004,N_3650,N_3766);
and U4005 (N_4005,N_3408,N_3948);
nor U4006 (N_4006,N_3032,N_3416);
nor U4007 (N_4007,N_3550,N_3980);
or U4008 (N_4008,N_3454,N_3316);
or U4009 (N_4009,N_3712,N_3891);
and U4010 (N_4010,N_3736,N_3722);
nor U4011 (N_4011,N_3468,N_3791);
xor U4012 (N_4012,N_3962,N_3079);
nand U4013 (N_4013,N_3974,N_3977);
or U4014 (N_4014,N_3912,N_3862);
or U4015 (N_4015,N_3352,N_3608);
and U4016 (N_4016,N_3195,N_3793);
nand U4017 (N_4017,N_3543,N_3156);
nor U4018 (N_4018,N_3303,N_3346);
nand U4019 (N_4019,N_3497,N_3214);
and U4020 (N_4020,N_3163,N_3746);
nor U4021 (N_4021,N_3186,N_3095);
and U4022 (N_4022,N_3849,N_3823);
nor U4023 (N_4023,N_3057,N_3771);
and U4024 (N_4024,N_3592,N_3495);
or U4025 (N_4025,N_3784,N_3114);
xnor U4026 (N_4026,N_3060,N_3926);
and U4027 (N_4027,N_3896,N_3358);
or U4028 (N_4028,N_3179,N_3199);
nor U4029 (N_4029,N_3970,N_3317);
nand U4030 (N_4030,N_3196,N_3976);
nor U4031 (N_4031,N_3538,N_3225);
xnor U4032 (N_4032,N_3836,N_3778);
xor U4033 (N_4033,N_3119,N_3143);
xnor U4034 (N_4034,N_3264,N_3773);
nor U4035 (N_4035,N_3724,N_3403);
and U4036 (N_4036,N_3305,N_3049);
or U4037 (N_4037,N_3876,N_3460);
nand U4038 (N_4038,N_3443,N_3966);
nor U4039 (N_4039,N_3578,N_3741);
nand U4040 (N_4040,N_3994,N_3643);
nand U4041 (N_4041,N_3355,N_3230);
nand U4042 (N_4042,N_3031,N_3379);
or U4043 (N_4043,N_3476,N_3703);
nor U4044 (N_4044,N_3788,N_3190);
nor U4045 (N_4045,N_3874,N_3751);
or U4046 (N_4046,N_3187,N_3593);
or U4047 (N_4047,N_3298,N_3721);
nor U4048 (N_4048,N_3957,N_3707);
or U4049 (N_4049,N_3365,N_3708);
nor U4050 (N_4050,N_3135,N_3568);
nor U4051 (N_4051,N_3116,N_3146);
and U4052 (N_4052,N_3294,N_3700);
or U4053 (N_4053,N_3904,N_3235);
nand U4054 (N_4054,N_3684,N_3331);
and U4055 (N_4055,N_3493,N_3640);
nor U4056 (N_4056,N_3945,N_3430);
nand U4057 (N_4057,N_3296,N_3239);
and U4058 (N_4058,N_3292,N_3914);
or U4059 (N_4059,N_3338,N_3870);
nor U4060 (N_4060,N_3269,N_3589);
nand U4061 (N_4061,N_3483,N_3665);
or U4062 (N_4062,N_3867,N_3508);
xor U4063 (N_4063,N_3297,N_3542);
xnor U4064 (N_4064,N_3834,N_3801);
nand U4065 (N_4065,N_3702,N_3813);
and U4066 (N_4066,N_3381,N_3289);
nand U4067 (N_4067,N_3604,N_3133);
and U4068 (N_4068,N_3743,N_3015);
nor U4069 (N_4069,N_3878,N_3623);
nand U4070 (N_4070,N_3065,N_3682);
nor U4071 (N_4071,N_3952,N_3609);
xor U4072 (N_4072,N_3614,N_3789);
or U4073 (N_4073,N_3638,N_3237);
nand U4074 (N_4074,N_3663,N_3221);
and U4075 (N_4075,N_3304,N_3790);
nor U4076 (N_4076,N_3459,N_3653);
xnor U4077 (N_4077,N_3206,N_3005);
nand U4078 (N_4078,N_3404,N_3631);
nor U4079 (N_4079,N_3181,N_3928);
nand U4080 (N_4080,N_3231,N_3137);
nor U4081 (N_4081,N_3101,N_3490);
nand U4082 (N_4082,N_3277,N_3322);
nor U4083 (N_4083,N_3852,N_3262);
nor U4084 (N_4084,N_3740,N_3450);
and U4085 (N_4085,N_3571,N_3530);
nor U4086 (N_4086,N_3913,N_3055);
or U4087 (N_4087,N_3339,N_3559);
nand U4088 (N_4088,N_3350,N_3111);
and U4089 (N_4089,N_3319,N_3566);
or U4090 (N_4090,N_3696,N_3671);
or U4091 (N_4091,N_3535,N_3389);
nor U4092 (N_4092,N_3061,N_3882);
or U4093 (N_4093,N_3633,N_3222);
nor U4094 (N_4094,N_3711,N_3687);
or U4095 (N_4095,N_3035,N_3779);
nand U4096 (N_4096,N_3223,N_3437);
or U4097 (N_4097,N_3556,N_3224);
and U4098 (N_4098,N_3284,N_3036);
nand U4099 (N_4099,N_3523,N_3361);
and U4100 (N_4100,N_3669,N_3924);
nor U4101 (N_4101,N_3360,N_3885);
nand U4102 (N_4102,N_3025,N_3109);
nand U4103 (N_4103,N_3953,N_3622);
and U4104 (N_4104,N_3968,N_3798);
nand U4105 (N_4105,N_3286,N_3817);
nor U4106 (N_4106,N_3792,N_3677);
and U4107 (N_4107,N_3986,N_3735);
or U4108 (N_4108,N_3526,N_3883);
and U4109 (N_4109,N_3548,N_3603);
or U4110 (N_4110,N_3840,N_3400);
nor U4111 (N_4111,N_3866,N_3482);
nor U4112 (N_4112,N_3692,N_3325);
nand U4113 (N_4113,N_3879,N_3983);
nand U4114 (N_4114,N_3255,N_3675);
and U4115 (N_4115,N_3178,N_3585);
nor U4116 (N_4116,N_3673,N_3007);
or U4117 (N_4117,N_3067,N_3254);
nand U4118 (N_4118,N_3978,N_3527);
nor U4119 (N_4119,N_3267,N_3356);
xor U4120 (N_4120,N_3959,N_3227);
nor U4121 (N_4121,N_3198,N_3575);
nor U4122 (N_4122,N_3946,N_3960);
nand U4123 (N_4123,N_3209,N_3118);
or U4124 (N_4124,N_3429,N_3886);
and U4125 (N_4125,N_3348,N_3494);
and U4126 (N_4126,N_3780,N_3828);
and U4127 (N_4127,N_3327,N_3981);
nand U4128 (N_4128,N_3308,N_3742);
and U4129 (N_4129,N_3851,N_3330);
nand U4130 (N_4130,N_3342,N_3969);
or U4131 (N_4131,N_3993,N_3856);
nor U4132 (N_4132,N_3377,N_3996);
or U4133 (N_4133,N_3376,N_3372);
or U4134 (N_4134,N_3438,N_3375);
xnor U4135 (N_4135,N_3475,N_3820);
xor U4136 (N_4136,N_3512,N_3194);
nor U4137 (N_4137,N_3138,N_3120);
or U4138 (N_4138,N_3717,N_3956);
nand U4139 (N_4139,N_3949,N_3326);
or U4140 (N_4140,N_3898,N_3887);
nor U4141 (N_4141,N_3918,N_3806);
and U4142 (N_4142,N_3013,N_3018);
nand U4143 (N_4143,N_3023,N_3825);
xnor U4144 (N_4144,N_3447,N_3162);
xor U4145 (N_4145,N_3905,N_3732);
nor U4146 (N_4146,N_3026,N_3954);
nand U4147 (N_4147,N_3261,N_3576);
nand U4148 (N_4148,N_3260,N_3436);
or U4149 (N_4149,N_3747,N_3599);
and U4150 (N_4150,N_3875,N_3144);
nor U4151 (N_4151,N_3397,N_3009);
or U4152 (N_4152,N_3037,N_3080);
or U4153 (N_4153,N_3110,N_3204);
and U4154 (N_4154,N_3321,N_3985);
nand U4155 (N_4155,N_3749,N_3249);
nand U4156 (N_4156,N_3487,N_3931);
or U4157 (N_4157,N_3469,N_3907);
xnor U4158 (N_4158,N_3300,N_3630);
xnor U4159 (N_4159,N_3177,N_3516);
nand U4160 (N_4160,N_3547,N_3515);
xnor U4161 (N_4161,N_3271,N_3033);
and U4162 (N_4162,N_3822,N_3467);
nor U4163 (N_4163,N_3217,N_3533);
or U4164 (N_4164,N_3226,N_3916);
nor U4165 (N_4165,N_3486,N_3274);
or U4166 (N_4166,N_3987,N_3458);
or U4167 (N_4167,N_3888,N_3920);
or U4168 (N_4168,N_3564,N_3328);
nor U4169 (N_4169,N_3594,N_3510);
or U4170 (N_4170,N_3933,N_3910);
or U4171 (N_4171,N_3621,N_3498);
xnor U4172 (N_4172,N_3121,N_3189);
and U4173 (N_4173,N_3815,N_3810);
and U4174 (N_4174,N_3086,N_3719);
nand U4175 (N_4175,N_3629,N_3734);
nor U4176 (N_4176,N_3058,N_3234);
or U4177 (N_4177,N_3044,N_3975);
nand U4178 (N_4178,N_3809,N_3938);
nand U4179 (N_4179,N_3378,N_3030);
or U4180 (N_4180,N_3581,N_3579);
nand U4181 (N_4181,N_3309,N_3656);
nor U4182 (N_4182,N_3529,N_3169);
nand U4183 (N_4183,N_3580,N_3610);
or U4184 (N_4184,N_3624,N_3074);
nor U4185 (N_4185,N_3582,N_3759);
xor U4186 (N_4186,N_3554,N_3832);
or U4187 (N_4187,N_3117,N_3725);
nor U4188 (N_4188,N_3919,N_3345);
nor U4189 (N_4189,N_3864,N_3423);
nor U4190 (N_4190,N_3710,N_3329);
nand U4191 (N_4191,N_3374,N_3145);
and U4192 (N_4192,N_3944,N_3591);
nand U4193 (N_4193,N_3611,N_3415);
nor U4194 (N_4194,N_3038,N_3858);
or U4195 (N_4195,N_3511,N_3107);
nor U4196 (N_4196,N_3029,N_3521);
nand U4197 (N_4197,N_3739,N_3201);
xnor U4198 (N_4198,N_3503,N_3522);
xor U4199 (N_4199,N_3401,N_3626);
and U4200 (N_4200,N_3392,N_3141);
nand U4201 (N_4201,N_3210,N_3391);
nor U4202 (N_4202,N_3865,N_3203);
nand U4203 (N_4203,N_3006,N_3808);
nand U4204 (N_4204,N_3362,N_3565);
nand U4205 (N_4205,N_3685,N_3011);
nand U4206 (N_4206,N_3370,N_3172);
and U4207 (N_4207,N_3413,N_3995);
and U4208 (N_4208,N_3046,N_3802);
nand U4209 (N_4209,N_3691,N_3218);
nor U4210 (N_4210,N_3432,N_3762);
or U4211 (N_4211,N_3730,N_3113);
or U4212 (N_4212,N_3860,N_3320);
nand U4213 (N_4213,N_3558,N_3909);
and U4214 (N_4214,N_3839,N_3216);
and U4215 (N_4215,N_3380,N_3694);
or U4216 (N_4216,N_3173,N_3704);
and U4217 (N_4217,N_3531,N_3008);
or U4218 (N_4218,N_3777,N_3635);
and U4219 (N_4219,N_3848,N_3388);
nand U4220 (N_4220,N_3314,N_3868);
xor U4221 (N_4221,N_3192,N_3890);
and U4222 (N_4222,N_3315,N_3507);
nand U4223 (N_4223,N_3247,N_3070);
or U4224 (N_4224,N_3229,N_3664);
nand U4225 (N_4225,N_3340,N_3765);
nor U4226 (N_4226,N_3412,N_3324);
and U4227 (N_4227,N_3642,N_3076);
or U4228 (N_4228,N_3040,N_3884);
xor U4229 (N_4229,N_3383,N_3803);
and U4230 (N_4230,N_3182,N_3641);
nor U4231 (N_4231,N_3597,N_3505);
nor U4232 (N_4232,N_3627,N_3131);
xnor U4233 (N_4233,N_3963,N_3606);
nand U4234 (N_4234,N_3857,N_3837);
nand U4235 (N_4235,N_3238,N_3184);
nand U4236 (N_4236,N_3804,N_3628);
nand U4237 (N_4237,N_3989,N_3877);
nor U4238 (N_4238,N_3257,N_3967);
and U4239 (N_4239,N_3104,N_3584);
nor U4240 (N_4240,N_3812,N_3845);
xnor U4241 (N_4241,N_3081,N_3453);
and U4242 (N_4242,N_3427,N_3092);
or U4243 (N_4243,N_3425,N_3048);
xnor U4244 (N_4244,N_3841,N_3831);
nand U4245 (N_4245,N_3426,N_3541);
nor U4246 (N_4246,N_3480,N_3772);
or U4247 (N_4247,N_3134,N_3484);
xnor U4248 (N_4248,N_3716,N_3351);
nor U4249 (N_4249,N_3984,N_3781);
nor U4250 (N_4250,N_3528,N_3513);
nand U4251 (N_4251,N_3418,N_3054);
and U4252 (N_4252,N_3754,N_3814);
and U4253 (N_4253,N_3601,N_3170);
or U4254 (N_4254,N_3228,N_3644);
or U4255 (N_4255,N_3850,N_3807);
nor U4256 (N_4256,N_3272,N_3481);
nand U4257 (N_4257,N_3073,N_3448);
xnor U4258 (N_4258,N_3000,N_3902);
or U4259 (N_4259,N_3667,N_3435);
and U4260 (N_4260,N_3616,N_3941);
nand U4261 (N_4261,N_3233,N_3265);
xor U4262 (N_4262,N_3657,N_3386);
nand U4263 (N_4263,N_3191,N_3028);
nor U4264 (N_4264,N_3563,N_3903);
nor U4265 (N_4265,N_3988,N_3520);
or U4266 (N_4266,N_3514,N_3540);
nand U4267 (N_4267,N_3921,N_3596);
or U4268 (N_4268,N_3075,N_3936);
and U4269 (N_4269,N_3307,N_3087);
and U4270 (N_4270,N_3136,N_3193);
xnor U4271 (N_4271,N_3906,N_3488);
and U4272 (N_4272,N_3615,N_3992);
nor U4273 (N_4273,N_3155,N_3698);
or U4274 (N_4274,N_3973,N_3463);
or U4275 (N_4275,N_3768,N_3441);
and U4276 (N_4276,N_3082,N_3417);
and U4277 (N_4277,N_3706,N_3699);
nor U4278 (N_4278,N_3256,N_3409);
nand U4279 (N_4279,N_3034,N_3112);
xor U4280 (N_4280,N_3053,N_3132);
and U4281 (N_4281,N_3894,N_3525);
xor U4282 (N_4282,N_3276,N_3098);
nor U4283 (N_4283,N_3185,N_3471);
or U4284 (N_4284,N_3153,N_3881);
nand U4285 (N_4285,N_3442,N_3390);
xor U4286 (N_4286,N_3853,N_3537);
nor U4287 (N_4287,N_3124,N_3197);
nor U4288 (N_4288,N_3655,N_3932);
nor U4289 (N_4289,N_3022,N_3129);
nor U4290 (N_4290,N_3019,N_3343);
and U4291 (N_4291,N_3750,N_3501);
nor U4292 (N_4292,N_3420,N_3369);
or U4293 (N_4293,N_3440,N_3998);
nand U4294 (N_4294,N_3477,N_3676);
and U4295 (N_4295,N_3639,N_3752);
nor U4296 (N_4296,N_3180,N_3701);
or U4297 (N_4297,N_3612,N_3697);
nor U4298 (N_4298,N_3253,N_3818);
nand U4299 (N_4299,N_3452,N_3561);
nand U4300 (N_4300,N_3705,N_3336);
and U4301 (N_4301,N_3091,N_3115);
nand U4302 (N_4302,N_3940,N_3679);
or U4303 (N_4303,N_3651,N_3843);
xor U4304 (N_4304,N_3003,N_3782);
nand U4305 (N_4305,N_3499,N_3937);
or U4306 (N_4306,N_3660,N_3646);
and U4307 (N_4307,N_3344,N_3128);
and U4308 (N_4308,N_3819,N_3157);
nor U4309 (N_4309,N_3613,N_3318);
or U4310 (N_4310,N_3895,N_3399);
and U4311 (N_4311,N_3103,N_3293);
nand U4312 (N_4312,N_3562,N_3942);
nand U4313 (N_4313,N_3295,N_3683);
nand U4314 (N_4314,N_3551,N_3174);
and U4315 (N_4315,N_3855,N_3042);
nand U4316 (N_4316,N_3236,N_3245);
or U4317 (N_4317,N_3607,N_3424);
nand U4318 (N_4318,N_3659,N_3270);
and U4319 (N_4319,N_3674,N_3775);
xor U4320 (N_4320,N_3496,N_3573);
xnor U4321 (N_4321,N_3451,N_3414);
nand U4322 (N_4322,N_3072,N_3662);
and U4323 (N_4323,N_3398,N_3979);
nand U4324 (N_4324,N_3359,N_3215);
and U4325 (N_4325,N_3445,N_3268);
nand U4326 (N_4326,N_3213,N_3387);
xnor U4327 (N_4327,N_3760,N_3159);
nor U4328 (N_4328,N_3004,N_3106);
or U4329 (N_4329,N_3310,N_3947);
or U4330 (N_4330,N_3354,N_3583);
xor U4331 (N_4331,N_3829,N_3688);
xor U4332 (N_4332,N_3552,N_3925);
or U4333 (N_4333,N_3456,N_3923);
or U4334 (N_4334,N_3334,N_3786);
nand U4335 (N_4335,N_3462,N_3492);
nor U4336 (N_4336,N_3502,N_3439);
xnor U4337 (N_4337,N_3428,N_3094);
xnor U4338 (N_4338,N_3863,N_3266);
or U4339 (N_4339,N_3431,N_3572);
nor U4340 (N_4340,N_3990,N_3280);
xnor U4341 (N_4341,N_3183,N_3205);
nand U4342 (N_4342,N_3273,N_3002);
xor U4343 (N_4343,N_3333,N_3367);
or U4344 (N_4344,N_3248,N_3748);
nand U4345 (N_4345,N_3411,N_3570);
or U4346 (N_4346,N_3958,N_3835);
nand U4347 (N_4347,N_3200,N_3833);
nor U4348 (N_4348,N_3341,N_3385);
nor U4349 (N_4349,N_3083,N_3062);
or U4350 (N_4350,N_3259,N_3617);
nand U4351 (N_4351,N_3755,N_3577);
and U4352 (N_4352,N_3726,N_3142);
or U4353 (N_4353,N_3744,N_3915);
xor U4354 (N_4354,N_3539,N_3299);
and U4355 (N_4355,N_3084,N_3407);
and U4356 (N_4356,N_3147,N_3433);
nand U4357 (N_4357,N_3100,N_3587);
or U4358 (N_4358,N_3500,N_3244);
xnor U4359 (N_4359,N_3219,N_3595);
and U4360 (N_4360,N_3410,N_3421);
nor U4361 (N_4361,N_3282,N_3893);
nor U4362 (N_4362,N_3518,N_3465);
and U4363 (N_4363,N_3444,N_3371);
nand U4364 (N_4364,N_3930,N_3586);
or U4365 (N_4365,N_3821,N_3123);
nand U4366 (N_4366,N_3243,N_3357);
nand U4367 (N_4367,N_3016,N_3869);
and U4368 (N_4368,N_3108,N_3846);
or U4369 (N_4369,N_3285,N_3939);
and U4370 (N_4370,N_3632,N_3063);
xor U4371 (N_4371,N_3672,N_3769);
nand U4372 (N_4372,N_3288,N_3922);
nand U4373 (N_4373,N_3050,N_3176);
or U4374 (N_4374,N_3043,N_3164);
nand U4375 (N_4375,N_3908,N_3871);
xor U4376 (N_4376,N_3774,N_3020);
nand U4377 (N_4377,N_3689,N_3250);
nor U4378 (N_4378,N_3347,N_3695);
and U4379 (N_4379,N_3620,N_3251);
nand U4380 (N_4380,N_3927,N_3634);
nor U4381 (N_4381,N_3506,N_3045);
or U4382 (N_4382,N_3066,N_3275);
nand U4383 (N_4383,N_3158,N_3715);
and U4384 (N_4384,N_3096,N_3934);
nand U4385 (N_4385,N_3532,N_3287);
nor U4386 (N_4386,N_3306,N_3800);
nor U4387 (N_4387,N_3472,N_3999);
nor U4388 (N_4388,N_3648,N_3899);
and U4389 (N_4389,N_3723,N_3139);
nor U4390 (N_4390,N_3770,N_3010);
or U4391 (N_4391,N_3152,N_3466);
or U4392 (N_4392,N_3207,N_3027);
xor U4393 (N_4393,N_3811,N_3872);
or U4394 (N_4394,N_3382,N_3241);
and U4395 (N_4395,N_3714,N_3733);
or U4396 (N_4396,N_3168,N_3929);
or U4397 (N_4397,N_3099,N_3757);
xor U4398 (N_4398,N_3729,N_3419);
nand U4399 (N_4399,N_3311,N_3171);
xnor U4400 (N_4400,N_3127,N_3368);
and U4401 (N_4401,N_3140,N_3301);
and U4402 (N_4402,N_3151,N_3880);
or U4403 (N_4403,N_3078,N_3125);
or U4404 (N_4404,N_3393,N_3900);
and U4405 (N_4405,N_3056,N_3126);
nor U4406 (N_4406,N_3816,N_3861);
nand U4407 (N_4407,N_3859,N_3738);
or U4408 (N_4408,N_3598,N_3457);
nor U4409 (N_4409,N_3709,N_3645);
nand U4410 (N_4410,N_3557,N_3366);
or U4411 (N_4411,N_3461,N_3524);
and U4412 (N_4412,N_3961,N_3093);
nor U4413 (N_4413,N_3824,N_3489);
nor U4414 (N_4414,N_3105,N_3951);
or U4415 (N_4415,N_3220,N_3728);
nand U4416 (N_4416,N_3312,N_3122);
and U4417 (N_4417,N_3668,N_3731);
or U4418 (N_4418,N_3051,N_3509);
or U4419 (N_4419,N_3102,N_3014);
nand U4420 (N_4420,N_3649,N_3670);
nand U4421 (N_4421,N_3085,N_3291);
nand U4422 (N_4422,N_3889,N_3167);
nand U4423 (N_4423,N_3021,N_3149);
nand U4424 (N_4424,N_3785,N_3263);
nor U4425 (N_4425,N_3545,N_3405);
nand U4426 (N_4426,N_3232,N_3842);
nand U4427 (N_4427,N_3165,N_3847);
nand U4428 (N_4428,N_3797,N_3069);
or U4429 (N_4429,N_3796,N_3549);
nor U4430 (N_4430,N_3246,N_3517);
nor U4431 (N_4431,N_3464,N_3827);
xnor U4432 (N_4432,N_3997,N_3240);
xor U4433 (N_4433,N_3666,N_3965);
xor U4434 (N_4434,N_3658,N_3012);
nand U4435 (N_4435,N_3278,N_3052);
nand U4436 (N_4436,N_3647,N_3560);
xor U4437 (N_4437,N_3150,N_3363);
nor U4438 (N_4438,N_3619,N_3625);
nand U4439 (N_4439,N_3485,N_3059);
or U4440 (N_4440,N_3039,N_3943);
nor U4441 (N_4441,N_3693,N_3097);
or U4442 (N_4442,N_3088,N_3795);
nor U4443 (N_4443,N_3402,N_3718);
nand U4444 (N_4444,N_3555,N_3406);
nand U4445 (N_4445,N_3258,N_3017);
or U4446 (N_4446,N_3600,N_3212);
and U4447 (N_4447,N_3982,N_3950);
xor U4448 (N_4448,N_3713,N_3154);
nand U4449 (N_4449,N_3917,N_3302);
or U4450 (N_4450,N_3636,N_3323);
nand U4451 (N_4451,N_3892,N_3618);
and U4452 (N_4452,N_3148,N_3972);
and U4453 (N_4453,N_3064,N_3290);
xor U4454 (N_4454,N_3242,N_3588);
nand U4455 (N_4455,N_3519,N_3335);
nor U4456 (N_4456,N_3449,N_3776);
or U4457 (N_4457,N_3283,N_3422);
nor U4458 (N_4458,N_3787,N_3089);
or U4459 (N_4459,N_3964,N_3783);
and U4460 (N_4460,N_3794,N_3353);
nand U4461 (N_4461,N_3077,N_3690);
and U4462 (N_4462,N_3544,N_3955);
nor U4463 (N_4463,N_3727,N_3763);
nand U4464 (N_4464,N_3935,N_3473);
nor U4465 (N_4465,N_3686,N_3911);
nand U4466 (N_4466,N_3681,N_3434);
nor U4467 (N_4467,N_3211,N_3838);
and U4468 (N_4468,N_3567,N_3047);
and U4469 (N_4469,N_3395,N_3332);
xor U4470 (N_4470,N_3805,N_3252);
nand U4471 (N_4471,N_3166,N_3826);
or U4472 (N_4472,N_3534,N_3652);
nor U4473 (N_4473,N_3202,N_3001);
xor U4474 (N_4474,N_3479,N_3602);
nor U4475 (N_4475,N_3491,N_3130);
nor U4476 (N_4476,N_3160,N_3071);
and U4477 (N_4477,N_3373,N_3680);
nand U4478 (N_4478,N_3854,N_3637);
nand U4479 (N_4479,N_3767,N_3446);
and U4480 (N_4480,N_3753,N_3175);
and U4481 (N_4481,N_3455,N_3279);
nand U4482 (N_4482,N_3678,N_3971);
or U4483 (N_4483,N_3504,N_3764);
nor U4484 (N_4484,N_3844,N_3281);
nor U4485 (N_4485,N_3396,N_3313);
nand U4486 (N_4486,N_3901,N_3799);
xor U4487 (N_4487,N_3337,N_3569);
and U4488 (N_4488,N_3384,N_3991);
or U4489 (N_4489,N_3873,N_3605);
or U4490 (N_4490,N_3756,N_3090);
nor U4491 (N_4491,N_3590,N_3661);
nand U4492 (N_4492,N_3161,N_3897);
and U4493 (N_4493,N_3474,N_3745);
and U4494 (N_4494,N_3758,N_3654);
nand U4495 (N_4495,N_3553,N_3574);
nor U4496 (N_4496,N_3068,N_3546);
and U4497 (N_4497,N_3208,N_3761);
nor U4498 (N_4498,N_3364,N_3830);
or U4499 (N_4499,N_3349,N_3478);
xor U4500 (N_4500,N_3015,N_3422);
and U4501 (N_4501,N_3157,N_3584);
and U4502 (N_4502,N_3640,N_3310);
or U4503 (N_4503,N_3144,N_3486);
nor U4504 (N_4504,N_3644,N_3636);
nor U4505 (N_4505,N_3959,N_3033);
and U4506 (N_4506,N_3875,N_3977);
or U4507 (N_4507,N_3411,N_3640);
nor U4508 (N_4508,N_3520,N_3036);
nand U4509 (N_4509,N_3197,N_3734);
xor U4510 (N_4510,N_3439,N_3954);
nor U4511 (N_4511,N_3432,N_3347);
and U4512 (N_4512,N_3593,N_3286);
nand U4513 (N_4513,N_3377,N_3801);
and U4514 (N_4514,N_3241,N_3830);
nor U4515 (N_4515,N_3615,N_3299);
xnor U4516 (N_4516,N_3987,N_3246);
nand U4517 (N_4517,N_3270,N_3142);
nor U4518 (N_4518,N_3041,N_3962);
or U4519 (N_4519,N_3051,N_3839);
nand U4520 (N_4520,N_3980,N_3857);
or U4521 (N_4521,N_3173,N_3671);
xor U4522 (N_4522,N_3951,N_3773);
nor U4523 (N_4523,N_3214,N_3350);
or U4524 (N_4524,N_3976,N_3990);
and U4525 (N_4525,N_3157,N_3919);
or U4526 (N_4526,N_3236,N_3195);
nand U4527 (N_4527,N_3791,N_3273);
xor U4528 (N_4528,N_3889,N_3093);
or U4529 (N_4529,N_3257,N_3910);
nand U4530 (N_4530,N_3915,N_3074);
or U4531 (N_4531,N_3303,N_3665);
or U4532 (N_4532,N_3899,N_3643);
nand U4533 (N_4533,N_3347,N_3448);
nor U4534 (N_4534,N_3254,N_3761);
nor U4535 (N_4535,N_3947,N_3955);
and U4536 (N_4536,N_3357,N_3639);
xnor U4537 (N_4537,N_3346,N_3473);
xnor U4538 (N_4538,N_3432,N_3628);
nand U4539 (N_4539,N_3983,N_3047);
nand U4540 (N_4540,N_3446,N_3166);
nor U4541 (N_4541,N_3999,N_3427);
nor U4542 (N_4542,N_3900,N_3605);
nand U4543 (N_4543,N_3173,N_3362);
xnor U4544 (N_4544,N_3696,N_3954);
nor U4545 (N_4545,N_3995,N_3178);
or U4546 (N_4546,N_3977,N_3954);
and U4547 (N_4547,N_3705,N_3765);
and U4548 (N_4548,N_3813,N_3206);
nor U4549 (N_4549,N_3334,N_3534);
nor U4550 (N_4550,N_3841,N_3653);
and U4551 (N_4551,N_3421,N_3765);
or U4552 (N_4552,N_3209,N_3162);
or U4553 (N_4553,N_3550,N_3454);
and U4554 (N_4554,N_3008,N_3940);
or U4555 (N_4555,N_3585,N_3505);
nand U4556 (N_4556,N_3670,N_3569);
nor U4557 (N_4557,N_3275,N_3767);
or U4558 (N_4558,N_3329,N_3891);
xor U4559 (N_4559,N_3308,N_3516);
or U4560 (N_4560,N_3252,N_3448);
or U4561 (N_4561,N_3453,N_3172);
nor U4562 (N_4562,N_3920,N_3822);
nor U4563 (N_4563,N_3911,N_3206);
or U4564 (N_4564,N_3178,N_3264);
and U4565 (N_4565,N_3942,N_3585);
nand U4566 (N_4566,N_3051,N_3728);
nand U4567 (N_4567,N_3661,N_3739);
nor U4568 (N_4568,N_3679,N_3158);
nor U4569 (N_4569,N_3158,N_3958);
nor U4570 (N_4570,N_3912,N_3326);
or U4571 (N_4571,N_3920,N_3763);
and U4572 (N_4572,N_3607,N_3813);
or U4573 (N_4573,N_3354,N_3928);
xor U4574 (N_4574,N_3468,N_3672);
nand U4575 (N_4575,N_3453,N_3756);
nor U4576 (N_4576,N_3381,N_3326);
xor U4577 (N_4577,N_3749,N_3920);
or U4578 (N_4578,N_3761,N_3372);
or U4579 (N_4579,N_3446,N_3549);
and U4580 (N_4580,N_3904,N_3983);
nand U4581 (N_4581,N_3053,N_3183);
nand U4582 (N_4582,N_3438,N_3641);
nor U4583 (N_4583,N_3850,N_3269);
nand U4584 (N_4584,N_3422,N_3064);
and U4585 (N_4585,N_3336,N_3443);
nor U4586 (N_4586,N_3919,N_3703);
and U4587 (N_4587,N_3185,N_3798);
or U4588 (N_4588,N_3802,N_3071);
and U4589 (N_4589,N_3200,N_3081);
or U4590 (N_4590,N_3718,N_3196);
nand U4591 (N_4591,N_3557,N_3840);
nand U4592 (N_4592,N_3518,N_3833);
and U4593 (N_4593,N_3322,N_3359);
nor U4594 (N_4594,N_3019,N_3349);
nand U4595 (N_4595,N_3226,N_3590);
nand U4596 (N_4596,N_3784,N_3502);
nor U4597 (N_4597,N_3324,N_3673);
nor U4598 (N_4598,N_3067,N_3745);
nand U4599 (N_4599,N_3236,N_3750);
nand U4600 (N_4600,N_3915,N_3426);
and U4601 (N_4601,N_3092,N_3978);
xor U4602 (N_4602,N_3792,N_3263);
or U4603 (N_4603,N_3898,N_3177);
nand U4604 (N_4604,N_3230,N_3360);
and U4605 (N_4605,N_3481,N_3835);
and U4606 (N_4606,N_3245,N_3860);
and U4607 (N_4607,N_3031,N_3784);
or U4608 (N_4608,N_3962,N_3300);
nand U4609 (N_4609,N_3307,N_3025);
nor U4610 (N_4610,N_3216,N_3166);
nor U4611 (N_4611,N_3607,N_3247);
nand U4612 (N_4612,N_3272,N_3214);
or U4613 (N_4613,N_3478,N_3582);
nor U4614 (N_4614,N_3861,N_3770);
and U4615 (N_4615,N_3526,N_3753);
or U4616 (N_4616,N_3004,N_3627);
nor U4617 (N_4617,N_3045,N_3725);
nand U4618 (N_4618,N_3777,N_3630);
and U4619 (N_4619,N_3306,N_3017);
or U4620 (N_4620,N_3790,N_3330);
nor U4621 (N_4621,N_3789,N_3109);
and U4622 (N_4622,N_3638,N_3307);
or U4623 (N_4623,N_3807,N_3327);
or U4624 (N_4624,N_3169,N_3254);
nand U4625 (N_4625,N_3956,N_3353);
and U4626 (N_4626,N_3424,N_3935);
or U4627 (N_4627,N_3869,N_3033);
and U4628 (N_4628,N_3068,N_3622);
nand U4629 (N_4629,N_3365,N_3093);
nand U4630 (N_4630,N_3516,N_3975);
xor U4631 (N_4631,N_3988,N_3182);
nand U4632 (N_4632,N_3549,N_3740);
and U4633 (N_4633,N_3138,N_3363);
nand U4634 (N_4634,N_3678,N_3601);
xnor U4635 (N_4635,N_3489,N_3120);
xnor U4636 (N_4636,N_3299,N_3188);
or U4637 (N_4637,N_3314,N_3798);
or U4638 (N_4638,N_3105,N_3363);
or U4639 (N_4639,N_3894,N_3456);
or U4640 (N_4640,N_3515,N_3105);
nand U4641 (N_4641,N_3600,N_3412);
and U4642 (N_4642,N_3692,N_3782);
and U4643 (N_4643,N_3688,N_3294);
nand U4644 (N_4644,N_3047,N_3251);
nand U4645 (N_4645,N_3399,N_3941);
xnor U4646 (N_4646,N_3640,N_3972);
nor U4647 (N_4647,N_3803,N_3673);
nand U4648 (N_4648,N_3070,N_3093);
or U4649 (N_4649,N_3519,N_3503);
and U4650 (N_4650,N_3098,N_3055);
nor U4651 (N_4651,N_3286,N_3926);
and U4652 (N_4652,N_3032,N_3355);
and U4653 (N_4653,N_3304,N_3473);
xnor U4654 (N_4654,N_3241,N_3890);
or U4655 (N_4655,N_3346,N_3164);
xnor U4656 (N_4656,N_3290,N_3252);
nor U4657 (N_4657,N_3664,N_3633);
or U4658 (N_4658,N_3576,N_3102);
and U4659 (N_4659,N_3941,N_3185);
nor U4660 (N_4660,N_3219,N_3720);
nand U4661 (N_4661,N_3131,N_3623);
nand U4662 (N_4662,N_3573,N_3002);
or U4663 (N_4663,N_3454,N_3212);
nor U4664 (N_4664,N_3399,N_3244);
or U4665 (N_4665,N_3619,N_3204);
and U4666 (N_4666,N_3746,N_3166);
and U4667 (N_4667,N_3797,N_3688);
and U4668 (N_4668,N_3477,N_3505);
or U4669 (N_4669,N_3507,N_3390);
nand U4670 (N_4670,N_3450,N_3605);
nand U4671 (N_4671,N_3291,N_3392);
and U4672 (N_4672,N_3709,N_3203);
nor U4673 (N_4673,N_3124,N_3384);
nor U4674 (N_4674,N_3695,N_3451);
nor U4675 (N_4675,N_3263,N_3961);
nor U4676 (N_4676,N_3179,N_3949);
nand U4677 (N_4677,N_3045,N_3526);
or U4678 (N_4678,N_3999,N_3327);
or U4679 (N_4679,N_3205,N_3425);
nand U4680 (N_4680,N_3021,N_3963);
nor U4681 (N_4681,N_3942,N_3786);
nor U4682 (N_4682,N_3128,N_3069);
or U4683 (N_4683,N_3588,N_3885);
or U4684 (N_4684,N_3025,N_3137);
nor U4685 (N_4685,N_3224,N_3575);
xor U4686 (N_4686,N_3390,N_3424);
nor U4687 (N_4687,N_3828,N_3820);
nor U4688 (N_4688,N_3734,N_3296);
and U4689 (N_4689,N_3230,N_3056);
nor U4690 (N_4690,N_3329,N_3086);
and U4691 (N_4691,N_3272,N_3824);
and U4692 (N_4692,N_3733,N_3735);
and U4693 (N_4693,N_3099,N_3534);
nand U4694 (N_4694,N_3043,N_3977);
nor U4695 (N_4695,N_3923,N_3975);
or U4696 (N_4696,N_3030,N_3724);
nand U4697 (N_4697,N_3044,N_3435);
nor U4698 (N_4698,N_3301,N_3778);
or U4699 (N_4699,N_3907,N_3141);
nand U4700 (N_4700,N_3860,N_3583);
or U4701 (N_4701,N_3592,N_3328);
nand U4702 (N_4702,N_3061,N_3099);
xor U4703 (N_4703,N_3024,N_3167);
and U4704 (N_4704,N_3186,N_3732);
nor U4705 (N_4705,N_3934,N_3121);
nor U4706 (N_4706,N_3931,N_3980);
and U4707 (N_4707,N_3961,N_3610);
xnor U4708 (N_4708,N_3364,N_3439);
nand U4709 (N_4709,N_3326,N_3636);
nor U4710 (N_4710,N_3919,N_3846);
nor U4711 (N_4711,N_3868,N_3906);
nor U4712 (N_4712,N_3314,N_3406);
xor U4713 (N_4713,N_3410,N_3795);
or U4714 (N_4714,N_3741,N_3459);
nor U4715 (N_4715,N_3418,N_3604);
nor U4716 (N_4716,N_3938,N_3678);
and U4717 (N_4717,N_3521,N_3159);
nor U4718 (N_4718,N_3859,N_3701);
and U4719 (N_4719,N_3498,N_3871);
nand U4720 (N_4720,N_3098,N_3097);
and U4721 (N_4721,N_3155,N_3720);
nand U4722 (N_4722,N_3747,N_3441);
xor U4723 (N_4723,N_3524,N_3660);
nor U4724 (N_4724,N_3324,N_3267);
nor U4725 (N_4725,N_3886,N_3035);
and U4726 (N_4726,N_3141,N_3290);
xnor U4727 (N_4727,N_3882,N_3651);
or U4728 (N_4728,N_3536,N_3505);
nand U4729 (N_4729,N_3004,N_3158);
xnor U4730 (N_4730,N_3109,N_3580);
xnor U4731 (N_4731,N_3493,N_3611);
and U4732 (N_4732,N_3456,N_3802);
nand U4733 (N_4733,N_3187,N_3755);
or U4734 (N_4734,N_3106,N_3035);
and U4735 (N_4735,N_3301,N_3104);
nand U4736 (N_4736,N_3741,N_3975);
nand U4737 (N_4737,N_3367,N_3443);
nand U4738 (N_4738,N_3829,N_3123);
nand U4739 (N_4739,N_3169,N_3035);
xnor U4740 (N_4740,N_3781,N_3236);
nor U4741 (N_4741,N_3336,N_3205);
nand U4742 (N_4742,N_3001,N_3825);
nand U4743 (N_4743,N_3335,N_3203);
or U4744 (N_4744,N_3312,N_3919);
or U4745 (N_4745,N_3218,N_3859);
or U4746 (N_4746,N_3548,N_3390);
nand U4747 (N_4747,N_3964,N_3091);
nand U4748 (N_4748,N_3583,N_3202);
xor U4749 (N_4749,N_3021,N_3623);
nand U4750 (N_4750,N_3378,N_3610);
nor U4751 (N_4751,N_3569,N_3091);
nand U4752 (N_4752,N_3323,N_3698);
or U4753 (N_4753,N_3383,N_3006);
nand U4754 (N_4754,N_3258,N_3840);
and U4755 (N_4755,N_3891,N_3980);
or U4756 (N_4756,N_3704,N_3477);
nor U4757 (N_4757,N_3185,N_3487);
nor U4758 (N_4758,N_3843,N_3972);
nand U4759 (N_4759,N_3309,N_3026);
xnor U4760 (N_4760,N_3903,N_3072);
nand U4761 (N_4761,N_3798,N_3177);
xnor U4762 (N_4762,N_3961,N_3552);
and U4763 (N_4763,N_3619,N_3259);
or U4764 (N_4764,N_3933,N_3123);
and U4765 (N_4765,N_3563,N_3190);
or U4766 (N_4766,N_3826,N_3693);
nand U4767 (N_4767,N_3213,N_3650);
nand U4768 (N_4768,N_3314,N_3446);
nand U4769 (N_4769,N_3736,N_3715);
xor U4770 (N_4770,N_3380,N_3649);
and U4771 (N_4771,N_3373,N_3875);
nand U4772 (N_4772,N_3785,N_3929);
or U4773 (N_4773,N_3790,N_3643);
or U4774 (N_4774,N_3693,N_3481);
and U4775 (N_4775,N_3742,N_3482);
xor U4776 (N_4776,N_3031,N_3076);
and U4777 (N_4777,N_3959,N_3349);
nor U4778 (N_4778,N_3520,N_3707);
or U4779 (N_4779,N_3102,N_3692);
nor U4780 (N_4780,N_3778,N_3980);
nand U4781 (N_4781,N_3598,N_3535);
and U4782 (N_4782,N_3103,N_3430);
nand U4783 (N_4783,N_3648,N_3121);
and U4784 (N_4784,N_3822,N_3687);
nand U4785 (N_4785,N_3892,N_3328);
nor U4786 (N_4786,N_3959,N_3791);
nor U4787 (N_4787,N_3480,N_3558);
xor U4788 (N_4788,N_3918,N_3834);
and U4789 (N_4789,N_3462,N_3153);
nor U4790 (N_4790,N_3028,N_3893);
and U4791 (N_4791,N_3926,N_3977);
xnor U4792 (N_4792,N_3645,N_3211);
xor U4793 (N_4793,N_3486,N_3716);
or U4794 (N_4794,N_3449,N_3690);
and U4795 (N_4795,N_3230,N_3553);
nand U4796 (N_4796,N_3265,N_3086);
or U4797 (N_4797,N_3639,N_3348);
xor U4798 (N_4798,N_3182,N_3903);
nand U4799 (N_4799,N_3558,N_3438);
or U4800 (N_4800,N_3335,N_3902);
and U4801 (N_4801,N_3709,N_3908);
and U4802 (N_4802,N_3618,N_3129);
nor U4803 (N_4803,N_3043,N_3897);
or U4804 (N_4804,N_3047,N_3135);
or U4805 (N_4805,N_3605,N_3775);
and U4806 (N_4806,N_3097,N_3531);
and U4807 (N_4807,N_3683,N_3017);
nor U4808 (N_4808,N_3413,N_3150);
nor U4809 (N_4809,N_3683,N_3929);
nand U4810 (N_4810,N_3889,N_3555);
and U4811 (N_4811,N_3334,N_3434);
and U4812 (N_4812,N_3990,N_3508);
nor U4813 (N_4813,N_3925,N_3757);
xor U4814 (N_4814,N_3350,N_3491);
nand U4815 (N_4815,N_3357,N_3590);
and U4816 (N_4816,N_3822,N_3532);
and U4817 (N_4817,N_3917,N_3654);
nand U4818 (N_4818,N_3749,N_3881);
and U4819 (N_4819,N_3028,N_3140);
or U4820 (N_4820,N_3093,N_3772);
nor U4821 (N_4821,N_3200,N_3054);
xnor U4822 (N_4822,N_3974,N_3759);
and U4823 (N_4823,N_3321,N_3456);
xnor U4824 (N_4824,N_3591,N_3890);
nor U4825 (N_4825,N_3696,N_3505);
or U4826 (N_4826,N_3430,N_3218);
nand U4827 (N_4827,N_3536,N_3683);
and U4828 (N_4828,N_3586,N_3265);
or U4829 (N_4829,N_3263,N_3335);
nand U4830 (N_4830,N_3424,N_3283);
nand U4831 (N_4831,N_3361,N_3557);
nor U4832 (N_4832,N_3581,N_3033);
nand U4833 (N_4833,N_3137,N_3708);
and U4834 (N_4834,N_3766,N_3969);
nand U4835 (N_4835,N_3029,N_3859);
and U4836 (N_4836,N_3475,N_3458);
nor U4837 (N_4837,N_3830,N_3017);
and U4838 (N_4838,N_3287,N_3399);
and U4839 (N_4839,N_3197,N_3907);
or U4840 (N_4840,N_3681,N_3024);
nand U4841 (N_4841,N_3154,N_3950);
xnor U4842 (N_4842,N_3513,N_3853);
and U4843 (N_4843,N_3049,N_3304);
nand U4844 (N_4844,N_3581,N_3196);
nor U4845 (N_4845,N_3348,N_3635);
and U4846 (N_4846,N_3131,N_3354);
or U4847 (N_4847,N_3718,N_3643);
nand U4848 (N_4848,N_3972,N_3558);
or U4849 (N_4849,N_3806,N_3183);
or U4850 (N_4850,N_3585,N_3896);
nor U4851 (N_4851,N_3280,N_3580);
or U4852 (N_4852,N_3979,N_3030);
nor U4853 (N_4853,N_3024,N_3388);
nor U4854 (N_4854,N_3161,N_3725);
or U4855 (N_4855,N_3929,N_3863);
or U4856 (N_4856,N_3596,N_3035);
and U4857 (N_4857,N_3584,N_3561);
or U4858 (N_4858,N_3036,N_3077);
xnor U4859 (N_4859,N_3211,N_3417);
and U4860 (N_4860,N_3710,N_3461);
and U4861 (N_4861,N_3517,N_3536);
nor U4862 (N_4862,N_3121,N_3020);
xor U4863 (N_4863,N_3175,N_3756);
and U4864 (N_4864,N_3761,N_3779);
nand U4865 (N_4865,N_3179,N_3883);
nand U4866 (N_4866,N_3934,N_3016);
or U4867 (N_4867,N_3593,N_3733);
nand U4868 (N_4868,N_3229,N_3912);
or U4869 (N_4869,N_3260,N_3978);
nand U4870 (N_4870,N_3524,N_3775);
and U4871 (N_4871,N_3258,N_3694);
or U4872 (N_4872,N_3270,N_3339);
nand U4873 (N_4873,N_3063,N_3242);
nand U4874 (N_4874,N_3099,N_3504);
or U4875 (N_4875,N_3876,N_3088);
or U4876 (N_4876,N_3014,N_3814);
and U4877 (N_4877,N_3206,N_3083);
nor U4878 (N_4878,N_3147,N_3434);
nor U4879 (N_4879,N_3843,N_3997);
xnor U4880 (N_4880,N_3911,N_3198);
nand U4881 (N_4881,N_3850,N_3265);
nor U4882 (N_4882,N_3119,N_3755);
and U4883 (N_4883,N_3811,N_3862);
and U4884 (N_4884,N_3218,N_3742);
and U4885 (N_4885,N_3404,N_3490);
xnor U4886 (N_4886,N_3134,N_3436);
nand U4887 (N_4887,N_3018,N_3324);
or U4888 (N_4888,N_3662,N_3309);
and U4889 (N_4889,N_3853,N_3924);
nor U4890 (N_4890,N_3500,N_3334);
or U4891 (N_4891,N_3573,N_3779);
nor U4892 (N_4892,N_3770,N_3638);
or U4893 (N_4893,N_3934,N_3065);
nor U4894 (N_4894,N_3678,N_3734);
and U4895 (N_4895,N_3747,N_3745);
nor U4896 (N_4896,N_3091,N_3679);
nand U4897 (N_4897,N_3879,N_3034);
xnor U4898 (N_4898,N_3131,N_3670);
and U4899 (N_4899,N_3810,N_3134);
nand U4900 (N_4900,N_3798,N_3562);
nor U4901 (N_4901,N_3031,N_3037);
nor U4902 (N_4902,N_3548,N_3125);
or U4903 (N_4903,N_3042,N_3691);
and U4904 (N_4904,N_3873,N_3344);
and U4905 (N_4905,N_3411,N_3396);
and U4906 (N_4906,N_3952,N_3962);
and U4907 (N_4907,N_3491,N_3338);
nor U4908 (N_4908,N_3373,N_3053);
and U4909 (N_4909,N_3225,N_3778);
or U4910 (N_4910,N_3791,N_3871);
or U4911 (N_4911,N_3537,N_3140);
nor U4912 (N_4912,N_3980,N_3850);
or U4913 (N_4913,N_3897,N_3210);
nand U4914 (N_4914,N_3784,N_3779);
nand U4915 (N_4915,N_3834,N_3078);
nor U4916 (N_4916,N_3181,N_3582);
nand U4917 (N_4917,N_3550,N_3669);
xnor U4918 (N_4918,N_3857,N_3658);
nor U4919 (N_4919,N_3587,N_3951);
and U4920 (N_4920,N_3328,N_3412);
and U4921 (N_4921,N_3824,N_3023);
nor U4922 (N_4922,N_3488,N_3145);
and U4923 (N_4923,N_3678,N_3676);
or U4924 (N_4924,N_3739,N_3295);
xnor U4925 (N_4925,N_3657,N_3876);
xnor U4926 (N_4926,N_3958,N_3955);
nand U4927 (N_4927,N_3454,N_3807);
and U4928 (N_4928,N_3608,N_3151);
and U4929 (N_4929,N_3835,N_3798);
nand U4930 (N_4930,N_3562,N_3293);
nand U4931 (N_4931,N_3906,N_3405);
nand U4932 (N_4932,N_3140,N_3307);
or U4933 (N_4933,N_3335,N_3472);
and U4934 (N_4934,N_3175,N_3082);
and U4935 (N_4935,N_3873,N_3352);
nor U4936 (N_4936,N_3371,N_3274);
nand U4937 (N_4937,N_3794,N_3699);
or U4938 (N_4938,N_3102,N_3282);
or U4939 (N_4939,N_3546,N_3041);
nand U4940 (N_4940,N_3423,N_3968);
nand U4941 (N_4941,N_3214,N_3541);
and U4942 (N_4942,N_3550,N_3531);
or U4943 (N_4943,N_3707,N_3220);
nor U4944 (N_4944,N_3872,N_3314);
nand U4945 (N_4945,N_3523,N_3394);
and U4946 (N_4946,N_3712,N_3568);
nand U4947 (N_4947,N_3984,N_3601);
nand U4948 (N_4948,N_3126,N_3297);
or U4949 (N_4949,N_3069,N_3089);
nor U4950 (N_4950,N_3986,N_3274);
nor U4951 (N_4951,N_3994,N_3098);
nand U4952 (N_4952,N_3349,N_3115);
and U4953 (N_4953,N_3942,N_3059);
nand U4954 (N_4954,N_3737,N_3074);
or U4955 (N_4955,N_3185,N_3957);
and U4956 (N_4956,N_3244,N_3290);
and U4957 (N_4957,N_3872,N_3492);
nor U4958 (N_4958,N_3987,N_3152);
xor U4959 (N_4959,N_3804,N_3335);
nand U4960 (N_4960,N_3682,N_3868);
nor U4961 (N_4961,N_3624,N_3689);
or U4962 (N_4962,N_3522,N_3899);
nand U4963 (N_4963,N_3552,N_3968);
xor U4964 (N_4964,N_3093,N_3391);
xor U4965 (N_4965,N_3038,N_3218);
nor U4966 (N_4966,N_3047,N_3330);
nand U4967 (N_4967,N_3035,N_3043);
xnor U4968 (N_4968,N_3047,N_3513);
nor U4969 (N_4969,N_3996,N_3397);
nand U4970 (N_4970,N_3913,N_3553);
or U4971 (N_4971,N_3239,N_3690);
xnor U4972 (N_4972,N_3337,N_3887);
and U4973 (N_4973,N_3958,N_3937);
and U4974 (N_4974,N_3161,N_3849);
xnor U4975 (N_4975,N_3886,N_3439);
nor U4976 (N_4976,N_3289,N_3693);
or U4977 (N_4977,N_3464,N_3079);
nand U4978 (N_4978,N_3861,N_3367);
nor U4979 (N_4979,N_3118,N_3582);
and U4980 (N_4980,N_3634,N_3507);
and U4981 (N_4981,N_3687,N_3941);
nand U4982 (N_4982,N_3811,N_3741);
or U4983 (N_4983,N_3832,N_3193);
or U4984 (N_4984,N_3411,N_3560);
nand U4985 (N_4985,N_3119,N_3864);
nand U4986 (N_4986,N_3317,N_3289);
or U4987 (N_4987,N_3050,N_3939);
nor U4988 (N_4988,N_3962,N_3403);
nor U4989 (N_4989,N_3605,N_3954);
and U4990 (N_4990,N_3481,N_3109);
nand U4991 (N_4991,N_3419,N_3935);
and U4992 (N_4992,N_3377,N_3762);
nor U4993 (N_4993,N_3978,N_3082);
nor U4994 (N_4994,N_3363,N_3980);
nand U4995 (N_4995,N_3863,N_3396);
xnor U4996 (N_4996,N_3474,N_3942);
nor U4997 (N_4997,N_3164,N_3712);
or U4998 (N_4998,N_3930,N_3487);
and U4999 (N_4999,N_3963,N_3361);
nand U5000 (N_5000,N_4031,N_4796);
nand U5001 (N_5001,N_4297,N_4591);
nor U5002 (N_5002,N_4980,N_4434);
xnor U5003 (N_5003,N_4019,N_4476);
xor U5004 (N_5004,N_4793,N_4597);
xnor U5005 (N_5005,N_4770,N_4180);
nor U5006 (N_5006,N_4859,N_4001);
and U5007 (N_5007,N_4798,N_4114);
or U5008 (N_5008,N_4857,N_4893);
nand U5009 (N_5009,N_4659,N_4924);
nand U5010 (N_5010,N_4842,N_4223);
or U5011 (N_5011,N_4200,N_4609);
nand U5012 (N_5012,N_4767,N_4193);
nand U5013 (N_5013,N_4618,N_4566);
nand U5014 (N_5014,N_4478,N_4670);
or U5015 (N_5015,N_4251,N_4643);
nor U5016 (N_5016,N_4804,N_4576);
nor U5017 (N_5017,N_4567,N_4161);
nand U5018 (N_5018,N_4064,N_4726);
nor U5019 (N_5019,N_4951,N_4721);
xor U5020 (N_5020,N_4540,N_4565);
and U5021 (N_5021,N_4153,N_4267);
nor U5022 (N_5022,N_4009,N_4274);
nor U5023 (N_5023,N_4769,N_4886);
nor U5024 (N_5024,N_4282,N_4482);
nor U5025 (N_5025,N_4410,N_4426);
or U5026 (N_5026,N_4712,N_4380);
and U5027 (N_5027,N_4676,N_4499);
and U5028 (N_5028,N_4090,N_4132);
nor U5029 (N_5029,N_4934,N_4967);
xnor U5030 (N_5030,N_4930,N_4062);
nand U5031 (N_5031,N_4950,N_4880);
and U5032 (N_5032,N_4667,N_4133);
and U5033 (N_5033,N_4570,N_4918);
or U5034 (N_5034,N_4559,N_4779);
nand U5035 (N_5035,N_4481,N_4421);
and U5036 (N_5036,N_4878,N_4703);
and U5037 (N_5037,N_4414,N_4104);
and U5038 (N_5038,N_4883,N_4407);
or U5039 (N_5039,N_4965,N_4942);
or U5040 (N_5040,N_4052,N_4530);
nor U5041 (N_5041,N_4357,N_4836);
and U5042 (N_5042,N_4127,N_4868);
and U5043 (N_5043,N_4413,N_4008);
and U5044 (N_5044,N_4821,N_4985);
and U5045 (N_5045,N_4771,N_4665);
nor U5046 (N_5046,N_4018,N_4048);
or U5047 (N_5047,N_4841,N_4017);
nor U5048 (N_5048,N_4870,N_4534);
and U5049 (N_5049,N_4671,N_4376);
nor U5050 (N_5050,N_4863,N_4602);
and U5051 (N_5051,N_4701,N_4990);
xnor U5052 (N_5052,N_4194,N_4473);
nand U5053 (N_5053,N_4864,N_4760);
nor U5054 (N_5054,N_4440,N_4378);
xnor U5055 (N_5055,N_4435,N_4622);
or U5056 (N_5056,N_4190,N_4386);
xor U5057 (N_5057,N_4640,N_4523);
nand U5058 (N_5058,N_4151,N_4642);
xor U5059 (N_5059,N_4139,N_4572);
xnor U5060 (N_5060,N_4011,N_4637);
nor U5061 (N_5061,N_4252,N_4409);
xor U5062 (N_5062,N_4269,N_4869);
nand U5063 (N_5063,N_4500,N_4563);
or U5064 (N_5064,N_4388,N_4368);
nand U5065 (N_5065,N_4292,N_4152);
or U5066 (N_5066,N_4799,N_4862);
nand U5067 (N_5067,N_4734,N_4268);
nand U5068 (N_5068,N_4858,N_4636);
and U5069 (N_5069,N_4957,N_4372);
xnor U5070 (N_5070,N_4955,N_4494);
or U5071 (N_5071,N_4895,N_4660);
xor U5072 (N_5072,N_4257,N_4520);
or U5073 (N_5073,N_4207,N_4234);
nand U5074 (N_5074,N_4055,N_4186);
or U5075 (N_5075,N_4022,N_4201);
nor U5076 (N_5076,N_4109,N_4912);
nand U5077 (N_5077,N_4989,N_4512);
nor U5078 (N_5078,N_4837,N_4333);
nor U5079 (N_5079,N_4184,N_4285);
nand U5080 (N_5080,N_4217,N_4855);
or U5081 (N_5081,N_4811,N_4135);
nor U5082 (N_5082,N_4192,N_4829);
nor U5083 (N_5083,N_4826,N_4488);
nor U5084 (N_5084,N_4405,N_4089);
or U5085 (N_5085,N_4644,N_4277);
and U5086 (N_5086,N_4141,N_4050);
nand U5087 (N_5087,N_4203,N_4938);
or U5088 (N_5088,N_4042,N_4711);
or U5089 (N_5089,N_4971,N_4524);
nor U5090 (N_5090,N_4492,N_4468);
and U5091 (N_5091,N_4732,N_4120);
and U5092 (N_5092,N_4555,N_4016);
and U5093 (N_5093,N_4522,N_4954);
xor U5094 (N_5094,N_4349,N_4899);
xnor U5095 (N_5095,N_4136,N_4801);
nand U5096 (N_5096,N_4126,N_4154);
nand U5097 (N_5097,N_4933,N_4900);
or U5098 (N_5098,N_4849,N_4748);
and U5099 (N_5099,N_4049,N_4281);
or U5100 (N_5100,N_4289,N_4057);
nand U5101 (N_5101,N_4013,N_4731);
and U5102 (N_5102,N_4650,N_4588);
and U5103 (N_5103,N_4974,N_4843);
nand U5104 (N_5104,N_4706,N_4084);
nor U5105 (N_5105,N_4266,N_4309);
nand U5106 (N_5106,N_4400,N_4963);
nor U5107 (N_5107,N_4627,N_4233);
nand U5108 (N_5108,N_4395,N_4002);
or U5109 (N_5109,N_4138,N_4077);
nand U5110 (N_5110,N_4081,N_4078);
or U5111 (N_5111,N_4578,N_4908);
or U5112 (N_5112,N_4010,N_4290);
or U5113 (N_5113,N_4171,N_4792);
nand U5114 (N_5114,N_4324,N_4551);
and U5115 (N_5115,N_4496,N_4382);
nor U5116 (N_5116,N_4928,N_4777);
nand U5117 (N_5117,N_4280,N_4250);
and U5118 (N_5118,N_4514,N_4398);
nor U5119 (N_5119,N_4103,N_4890);
or U5120 (N_5120,N_4575,N_4340);
or U5121 (N_5121,N_4352,N_4105);
nor U5122 (N_5122,N_4874,N_4474);
or U5123 (N_5123,N_4994,N_4003);
and U5124 (N_5124,N_4338,N_4142);
and U5125 (N_5125,N_4937,N_4749);
nor U5126 (N_5126,N_4589,N_4754);
nor U5127 (N_5127,N_4036,N_4891);
or U5128 (N_5128,N_4427,N_4302);
and U5129 (N_5129,N_4833,N_4390);
xnor U5130 (N_5130,N_4176,N_4505);
or U5131 (N_5131,N_4825,N_4614);
or U5132 (N_5132,N_4189,N_4681);
or U5133 (N_5133,N_4704,N_4820);
nor U5134 (N_5134,N_4773,N_4719);
xor U5135 (N_5135,N_4447,N_4237);
nand U5136 (N_5136,N_4592,N_4005);
nand U5137 (N_5137,N_4131,N_4260);
nor U5138 (N_5138,N_4088,N_4802);
nor U5139 (N_5139,N_4023,N_4295);
nand U5140 (N_5140,N_4156,N_4460);
xnor U5141 (N_5141,N_4700,N_4165);
nand U5142 (N_5142,N_4655,N_4781);
or U5143 (N_5143,N_4772,N_4399);
nor U5144 (N_5144,N_4553,N_4691);
nor U5145 (N_5145,N_4724,N_4978);
and U5146 (N_5146,N_4949,N_4271);
or U5147 (N_5147,N_4463,N_4850);
and U5148 (N_5148,N_4483,N_4907);
nor U5149 (N_5149,N_4604,N_4879);
nor U5150 (N_5150,N_4973,N_4255);
nor U5151 (N_5151,N_4672,N_4586);
nor U5152 (N_5152,N_4328,N_4789);
and U5153 (N_5153,N_4606,N_4337);
xor U5154 (N_5154,N_4780,N_4174);
or U5155 (N_5155,N_4199,N_4952);
or U5156 (N_5156,N_4976,N_4525);
or U5157 (N_5157,N_4411,N_4902);
and U5158 (N_5158,N_4355,N_4204);
nand U5159 (N_5159,N_4053,N_4240);
xor U5160 (N_5160,N_4202,N_4068);
nor U5161 (N_5161,N_4144,N_4159);
nor U5162 (N_5162,N_4882,N_4872);
nor U5163 (N_5163,N_4892,N_4574);
or U5164 (N_5164,N_4179,N_4856);
nor U5165 (N_5165,N_4617,N_4818);
or U5166 (N_5166,N_4752,N_4953);
nand U5167 (N_5167,N_4106,N_4344);
or U5168 (N_5168,N_4404,N_4730);
nor U5169 (N_5169,N_4956,N_4243);
nand U5170 (N_5170,N_4867,N_4254);
or U5171 (N_5171,N_4046,N_4554);
and U5172 (N_5172,N_4241,N_4692);
nor U5173 (N_5173,N_4852,N_4526);
and U5174 (N_5174,N_4348,N_4288);
or U5175 (N_5175,N_4887,N_4032);
or U5176 (N_5176,N_4823,N_4226);
and U5177 (N_5177,N_4479,N_4939);
xor U5178 (N_5178,N_4970,N_4745);
and U5179 (N_5179,N_4316,N_4817);
nor U5180 (N_5180,N_4958,N_4806);
or U5181 (N_5181,N_4045,N_4219);
and U5182 (N_5182,N_4230,N_4175);
or U5183 (N_5183,N_4437,N_4325);
nand U5184 (N_5184,N_4270,N_4300);
or U5185 (N_5185,N_4472,N_4747);
xnor U5186 (N_5186,N_4304,N_4264);
or U5187 (N_5187,N_4805,N_4246);
xnor U5188 (N_5188,N_4383,N_4097);
or U5189 (N_5189,N_4163,N_4107);
and U5190 (N_5190,N_4682,N_4082);
and U5191 (N_5191,N_4444,N_4516);
nand U5192 (N_5192,N_4205,N_4750);
nand U5193 (N_5193,N_4718,N_4273);
nor U5194 (N_5194,N_4279,N_4430);
and U5195 (N_5195,N_4007,N_4756);
or U5196 (N_5196,N_4112,N_4312);
or U5197 (N_5197,N_4188,N_4982);
nand U5198 (N_5198,N_4757,N_4788);
nor U5199 (N_5199,N_4423,N_4674);
or U5200 (N_5200,N_4929,N_4058);
nand U5201 (N_5201,N_4532,N_4913);
and U5202 (N_5202,N_4791,N_4884);
or U5203 (N_5203,N_4759,N_4262);
or U5204 (N_5204,N_4558,N_4209);
nand U5205 (N_5205,N_4607,N_4485);
nor U5206 (N_5206,N_4897,N_4275);
nand U5207 (N_5207,N_4827,N_4506);
and U5208 (N_5208,N_4143,N_4925);
nand U5209 (N_5209,N_4379,N_4835);
nand U5210 (N_5210,N_4824,N_4387);
or U5211 (N_5211,N_4322,N_4091);
or U5212 (N_5212,N_4210,N_4157);
nor U5213 (N_5213,N_4299,N_4162);
nor U5214 (N_5214,N_4941,N_4653);
nor U5215 (N_5215,N_4441,N_4809);
xor U5216 (N_5216,N_4278,N_4004);
or U5217 (N_5217,N_4239,N_4198);
nor U5218 (N_5218,N_4697,N_4443);
nand U5219 (N_5219,N_4043,N_4206);
nand U5220 (N_5220,N_4145,N_4917);
and U5221 (N_5221,N_4493,N_4742);
nor U5222 (N_5222,N_4147,N_4124);
xnor U5223 (N_5223,N_4944,N_4393);
or U5224 (N_5224,N_4517,N_4548);
and U5225 (N_5225,N_4354,N_4467);
nand U5226 (N_5226,N_4166,N_4168);
xor U5227 (N_5227,N_4694,N_4940);
nor U5228 (N_5228,N_4029,N_4397);
or U5229 (N_5229,N_4464,N_4220);
xor U5230 (N_5230,N_4647,N_4236);
nor U5231 (N_5231,N_4743,N_4272);
or U5232 (N_5232,N_4012,N_4392);
or U5233 (N_5233,N_4995,N_4716);
and U5234 (N_5234,N_4111,N_4889);
or U5235 (N_5235,N_4537,N_4529);
nand U5236 (N_5236,N_4164,N_4433);
and U5237 (N_5237,N_4999,N_4303);
nor U5238 (N_5238,N_4931,N_4119);
nand U5239 (N_5239,N_4027,N_4471);
and U5240 (N_5240,N_4353,N_4079);
nor U5241 (N_5241,N_4905,N_4966);
nand U5242 (N_5242,N_4214,N_4060);
and U5243 (N_5243,N_4118,N_4881);
or U5244 (N_5244,N_4775,N_4394);
nand U5245 (N_5245,N_4211,N_4177);
nor U5246 (N_5246,N_4581,N_4365);
and U5247 (N_5247,N_4787,N_4396);
and U5248 (N_5248,N_4737,N_4083);
nor U5249 (N_5249,N_4646,N_4436);
or U5250 (N_5250,N_4758,N_4533);
nor U5251 (N_5251,N_4580,N_4448);
nand U5252 (N_5252,N_4696,N_4315);
nand U5253 (N_5253,N_4894,N_4687);
or U5254 (N_5254,N_4632,N_4232);
and U5255 (N_5255,N_4469,N_4866);
and U5256 (N_5256,N_4087,N_4401);
or U5257 (N_5257,N_4334,N_4557);
and U5258 (N_5258,N_4936,N_4373);
nand U5259 (N_5259,N_4006,N_4601);
nor U5260 (N_5260,N_4993,N_4419);
nand U5261 (N_5261,N_4336,N_4705);
nand U5262 (N_5262,N_4511,N_4975);
and U5263 (N_5263,N_4185,N_4782);
nor U5264 (N_5264,N_4321,N_4633);
nor U5265 (N_5265,N_4535,N_4800);
or U5266 (N_5266,N_4661,N_4693);
nand U5267 (N_5267,N_4648,N_4587);
or U5268 (N_5268,N_4389,N_4094);
and U5269 (N_5269,N_4624,N_4668);
nand U5270 (N_5270,N_4717,N_4098);
or U5271 (N_5271,N_4612,N_4794);
nand U5272 (N_5272,N_4461,N_4669);
or U5273 (N_5273,N_4170,N_4495);
or U5274 (N_5274,N_4509,N_4491);
nand U5275 (N_5275,N_4259,N_4834);
xnor U5276 (N_5276,N_4755,N_4997);
or U5277 (N_5277,N_4739,N_4992);
nand U5278 (N_5278,N_4224,N_4428);
or U5279 (N_5279,N_4196,N_4733);
or U5280 (N_5280,N_4616,N_4326);
xor U5281 (N_5281,N_4504,N_4599);
nand U5282 (N_5282,N_4417,N_4631);
nor U5283 (N_5283,N_4183,N_4129);
nor U5284 (N_5284,N_4969,N_4073);
nand U5285 (N_5285,N_4298,N_4656);
or U5286 (N_5286,N_4169,N_4155);
or U5287 (N_5287,N_4695,N_4538);
and U5288 (N_5288,N_4291,N_4412);
nor U5289 (N_5289,N_4685,N_4996);
nor U5290 (N_5290,N_4363,N_4341);
xnor U5291 (N_5291,N_4725,N_4072);
and U5292 (N_5292,N_4329,N_4903);
nand U5293 (N_5293,N_4510,N_4848);
xnor U5294 (N_5294,N_4128,N_4034);
nand U5295 (N_5295,N_4221,N_4960);
nand U5296 (N_5296,N_4351,N_4723);
or U5297 (N_5297,N_4342,N_4984);
nor U5298 (N_5298,N_4446,N_4213);
nand U5299 (N_5299,N_4556,N_4158);
and U5300 (N_5300,N_4408,N_4350);
and U5301 (N_5301,N_4470,N_4873);
nand U5302 (N_5302,N_4021,N_4686);
nand U5303 (N_5303,N_4560,N_4763);
and U5304 (N_5304,N_4358,N_4853);
nor U5305 (N_5305,N_4130,N_4314);
or U5306 (N_5306,N_4331,N_4150);
xnor U5307 (N_5307,N_4590,N_4457);
and U5308 (N_5308,N_4455,N_4449);
or U5309 (N_5309,N_4261,N_4608);
xnor U5310 (N_5310,N_4920,N_4063);
or U5311 (N_5311,N_4783,N_4986);
and U5312 (N_5312,N_4453,N_4070);
or U5313 (N_5313,N_4753,N_4764);
nor U5314 (N_5314,N_4489,N_4317);
nand U5315 (N_5315,N_4635,N_4311);
nand U5316 (N_5316,N_4123,N_4287);
and U5317 (N_5317,N_4335,N_4528);
and U5318 (N_5318,N_4222,N_4117);
xnor U5319 (N_5319,N_4487,N_4876);
and U5320 (N_5320,N_4830,N_4727);
nand U5321 (N_5321,N_4641,N_4085);
nand U5322 (N_5322,N_4962,N_4228);
xor U5323 (N_5323,N_4603,N_4366);
and U5324 (N_5324,N_4294,N_4683);
xnor U5325 (N_5325,N_4662,N_4484);
and U5326 (N_5326,N_4610,N_4545);
and U5327 (N_5327,N_4497,N_4371);
and U5328 (N_5328,N_4466,N_4037);
nand U5329 (N_5329,N_4846,N_4657);
or U5330 (N_5330,N_4306,N_4416);
nand U5331 (N_5331,N_4054,N_4025);
nor U5332 (N_5332,N_4439,N_4066);
xor U5333 (N_5333,N_4702,N_4319);
nor U5334 (N_5334,N_4231,N_4564);
nor U5335 (N_5335,N_4596,N_4486);
xnor U5336 (N_5336,N_4649,N_4968);
or U5337 (N_5337,N_4583,N_4541);
nor U5338 (N_5338,N_4584,N_4921);
nand U5339 (N_5339,N_4218,N_4542);
xor U5340 (N_5340,N_4943,N_4465);
nor U5341 (N_5341,N_4991,N_4673);
and U5342 (N_5342,N_4406,N_4547);
nor U5343 (N_5343,N_4041,N_4896);
nor U5344 (N_5344,N_4579,N_4051);
xor U5345 (N_5345,N_4033,N_4562);
or U5346 (N_5346,N_4816,N_4360);
or U5347 (N_5347,N_4911,N_4323);
or U5348 (N_5348,N_4364,N_4362);
xor U5349 (N_5349,N_4713,N_4741);
nor U5350 (N_5350,N_4605,N_4451);
and U5351 (N_5351,N_4216,N_4527);
xor U5352 (N_5352,N_4919,N_4812);
or U5353 (N_5353,N_4822,N_4075);
and U5354 (N_5354,N_4947,N_4707);
nor U5355 (N_5355,N_4736,N_4698);
nand U5356 (N_5356,N_4518,N_4922);
nor U5357 (N_5357,N_4561,N_4480);
nor U5358 (N_5358,N_4728,N_4663);
nor U5359 (N_5359,N_4838,N_4959);
nand U5360 (N_5360,N_4283,N_4069);
nand U5361 (N_5361,N_4582,N_4310);
nor U5362 (N_5362,N_4502,N_4513);
and U5363 (N_5363,N_4948,N_4910);
or U5364 (N_5364,N_4507,N_4044);
or U5365 (N_5365,N_4296,N_4689);
nand U5366 (N_5366,N_4030,N_4501);
nand U5367 (N_5367,N_4654,N_4071);
or U5368 (N_5368,N_4761,N_4598);
or U5369 (N_5369,N_4710,N_4422);
nor U5370 (N_5370,N_4014,N_4450);
or U5371 (N_5371,N_4593,N_4778);
nor U5372 (N_5372,N_4585,N_4208);
nand U5373 (N_5373,N_4977,N_4102);
nor U5374 (N_5374,N_4462,N_4115);
xor U5375 (N_5375,N_4819,N_4865);
nand U5376 (N_5376,N_4595,N_4785);
nor U5377 (N_5377,N_4861,N_4815);
nor U5378 (N_5378,N_4238,N_4454);
nand U5379 (N_5379,N_4225,N_4629);
nor U5380 (N_5380,N_4840,N_4898);
nand U5381 (N_5381,N_4096,N_4093);
and U5382 (N_5382,N_4242,N_4531);
or U5383 (N_5383,N_4550,N_4620);
nor U5384 (N_5384,N_4490,N_4247);
nand U5385 (N_5385,N_4573,N_4735);
and U5386 (N_5386,N_4442,N_4885);
and U5387 (N_5387,N_4038,N_4935);
and U5388 (N_5388,N_4766,N_4318);
or U5389 (N_5389,N_4926,N_4256);
xor U5390 (N_5390,N_4675,N_4915);
nor U5391 (N_5391,N_4375,N_4330);
nand U5392 (N_5392,N_4092,N_4914);
nand U5393 (N_5393,N_4369,N_4790);
nor U5394 (N_5394,N_4658,N_4181);
nand U5395 (N_5395,N_4113,N_4248);
or U5396 (N_5396,N_4377,N_4797);
nor U5397 (N_5397,N_4020,N_4628);
nor U5398 (N_5398,N_4339,N_4245);
or U5399 (N_5399,N_4768,N_4871);
nand U5400 (N_5400,N_4972,N_4498);
nor U5401 (N_5401,N_4122,N_4086);
or U5402 (N_5402,N_4813,N_4577);
nand U5403 (N_5403,N_4215,N_4458);
and U5404 (N_5404,N_4432,N_4108);
xor U5405 (N_5405,N_4784,N_4539);
or U5406 (N_5406,N_4645,N_4307);
nor U5407 (N_5407,N_4456,N_4172);
and U5408 (N_5408,N_4844,N_4945);
xor U5409 (N_5409,N_4116,N_4998);
and U5410 (N_5410,N_4028,N_4626);
nor U5411 (N_5411,N_4875,N_4195);
nand U5412 (N_5412,N_4751,N_4983);
or U5413 (N_5413,N_4249,N_4080);
or U5414 (N_5414,N_4356,N_4431);
or U5415 (N_5415,N_4946,N_4729);
and U5416 (N_5416,N_4359,N_4074);
and U5417 (N_5417,N_4549,N_4927);
and U5418 (N_5418,N_4026,N_4508);
nand U5419 (N_5419,N_4690,N_4076);
and U5420 (N_5420,N_4543,N_4638);
or U5421 (N_5421,N_4803,N_4167);
nand U5422 (N_5422,N_4452,N_4293);
nor U5423 (N_5423,N_4916,N_4146);
or U5424 (N_5424,N_4125,N_4061);
nor U5425 (N_5425,N_4722,N_4475);
nand U5426 (N_5426,N_4385,N_4056);
nand U5427 (N_5427,N_4634,N_4370);
or U5428 (N_5428,N_4828,N_4229);
nor U5429 (N_5429,N_4765,N_4134);
and U5430 (N_5430,N_4445,N_4615);
and U5431 (N_5431,N_4000,N_4024);
nor U5432 (N_5432,N_4901,N_4039);
and U5433 (N_5433,N_4679,N_4688);
nand U5434 (N_5434,N_4503,N_4301);
or U5435 (N_5435,N_4619,N_4276);
nor U5436 (N_5436,N_4308,N_4227);
and U5437 (N_5437,N_4420,N_4059);
xnor U5438 (N_5438,N_4265,N_4860);
nand U5439 (N_5439,N_4845,N_4932);
nand U5440 (N_5440,N_4391,N_4621);
and U5441 (N_5441,N_4847,N_4140);
nand U5442 (N_5442,N_4040,N_4611);
xor U5443 (N_5443,N_4173,N_4101);
nand U5444 (N_5444,N_4424,N_4015);
nand U5445 (N_5445,N_4149,N_4964);
and U5446 (N_5446,N_4402,N_4384);
nand U5447 (N_5447,N_4568,N_4594);
and U5448 (N_5448,N_4786,N_4418);
or U5449 (N_5449,N_4244,N_4720);
and U5450 (N_5450,N_4988,N_4888);
or U5451 (N_5451,N_4651,N_4212);
xor U5452 (N_5452,N_4699,N_4403);
or U5453 (N_5453,N_4569,N_4345);
nor U5454 (N_5454,N_4664,N_4600);
nor U5455 (N_5455,N_4343,N_4923);
or U5456 (N_5456,N_4178,N_4795);
and U5457 (N_5457,N_4099,N_4361);
nand U5458 (N_5458,N_4906,N_4851);
and U5459 (N_5459,N_4438,N_4776);
nor U5460 (N_5460,N_4459,N_4536);
nand U5461 (N_5461,N_4182,N_4284);
and U5462 (N_5462,N_4327,N_4839);
nor U5463 (N_5463,N_4715,N_4904);
and U5464 (N_5464,N_4807,N_4979);
xnor U5465 (N_5465,N_4429,N_4305);
or U5466 (N_5466,N_4035,N_4810);
xor U5467 (N_5467,N_4762,N_4477);
nand U5468 (N_5468,N_4515,N_4625);
or U5469 (N_5469,N_4740,N_4709);
nor U5470 (N_5470,N_4714,N_4187);
and U5471 (N_5471,N_4415,N_4160);
or U5472 (N_5472,N_4100,N_4552);
nand U5473 (N_5473,N_4095,N_4639);
nor U5474 (N_5474,N_4110,N_4987);
xnor U5475 (N_5475,N_4613,N_4367);
and U5476 (N_5476,N_4381,N_4571);
or U5477 (N_5477,N_4521,N_4744);
nand U5478 (N_5478,N_4877,N_4263);
xnor U5479 (N_5479,N_4738,N_4137);
nor U5480 (N_5480,N_4346,N_4832);
xnor U5481 (N_5481,N_4961,N_4067);
or U5482 (N_5482,N_4630,N_4258);
nor U5483 (N_5483,N_4313,N_4253);
nor U5484 (N_5484,N_4374,N_4623);
and U5485 (N_5485,N_4684,N_4814);
or U5486 (N_5486,N_4680,N_4652);
or U5487 (N_5487,N_4347,N_4121);
nand U5488 (N_5488,N_4286,N_4909);
nor U5489 (N_5489,N_4708,N_4544);
nand U5490 (N_5490,N_4981,N_4546);
or U5491 (N_5491,N_4320,N_4746);
xor U5492 (N_5492,N_4235,N_4677);
or U5493 (N_5493,N_4191,N_4808);
or U5494 (N_5494,N_4425,N_4854);
nand U5495 (N_5495,N_4774,N_4666);
nand U5496 (N_5496,N_4197,N_4047);
or U5497 (N_5497,N_4678,N_4332);
and U5498 (N_5498,N_4519,N_4148);
nor U5499 (N_5499,N_4831,N_4065);
and U5500 (N_5500,N_4173,N_4839);
or U5501 (N_5501,N_4364,N_4413);
nor U5502 (N_5502,N_4552,N_4123);
or U5503 (N_5503,N_4525,N_4533);
nand U5504 (N_5504,N_4573,N_4051);
or U5505 (N_5505,N_4784,N_4464);
nand U5506 (N_5506,N_4499,N_4611);
nor U5507 (N_5507,N_4453,N_4983);
nor U5508 (N_5508,N_4994,N_4711);
nand U5509 (N_5509,N_4977,N_4135);
nor U5510 (N_5510,N_4518,N_4385);
nor U5511 (N_5511,N_4402,N_4025);
nand U5512 (N_5512,N_4013,N_4053);
nand U5513 (N_5513,N_4741,N_4684);
nor U5514 (N_5514,N_4168,N_4570);
xor U5515 (N_5515,N_4046,N_4387);
or U5516 (N_5516,N_4166,N_4931);
nand U5517 (N_5517,N_4371,N_4278);
nand U5518 (N_5518,N_4982,N_4255);
and U5519 (N_5519,N_4779,N_4599);
or U5520 (N_5520,N_4910,N_4840);
nand U5521 (N_5521,N_4822,N_4580);
or U5522 (N_5522,N_4191,N_4485);
nand U5523 (N_5523,N_4788,N_4829);
xnor U5524 (N_5524,N_4416,N_4139);
or U5525 (N_5525,N_4300,N_4163);
and U5526 (N_5526,N_4841,N_4162);
nand U5527 (N_5527,N_4239,N_4514);
nand U5528 (N_5528,N_4243,N_4227);
xor U5529 (N_5529,N_4800,N_4267);
nor U5530 (N_5530,N_4357,N_4554);
and U5531 (N_5531,N_4390,N_4412);
nand U5532 (N_5532,N_4489,N_4220);
and U5533 (N_5533,N_4757,N_4020);
nor U5534 (N_5534,N_4169,N_4518);
or U5535 (N_5535,N_4061,N_4723);
and U5536 (N_5536,N_4300,N_4205);
nor U5537 (N_5537,N_4372,N_4058);
nand U5538 (N_5538,N_4918,N_4452);
and U5539 (N_5539,N_4296,N_4010);
xor U5540 (N_5540,N_4316,N_4821);
nand U5541 (N_5541,N_4125,N_4580);
or U5542 (N_5542,N_4075,N_4688);
and U5543 (N_5543,N_4204,N_4112);
nand U5544 (N_5544,N_4700,N_4121);
xor U5545 (N_5545,N_4948,N_4672);
xor U5546 (N_5546,N_4327,N_4059);
or U5547 (N_5547,N_4099,N_4527);
and U5548 (N_5548,N_4374,N_4337);
nand U5549 (N_5549,N_4172,N_4874);
and U5550 (N_5550,N_4735,N_4201);
and U5551 (N_5551,N_4679,N_4345);
xnor U5552 (N_5552,N_4884,N_4829);
nand U5553 (N_5553,N_4041,N_4292);
or U5554 (N_5554,N_4365,N_4691);
xnor U5555 (N_5555,N_4366,N_4589);
nand U5556 (N_5556,N_4815,N_4812);
nand U5557 (N_5557,N_4919,N_4846);
xor U5558 (N_5558,N_4425,N_4852);
xnor U5559 (N_5559,N_4069,N_4966);
and U5560 (N_5560,N_4703,N_4793);
or U5561 (N_5561,N_4591,N_4731);
or U5562 (N_5562,N_4899,N_4751);
and U5563 (N_5563,N_4865,N_4183);
and U5564 (N_5564,N_4531,N_4938);
and U5565 (N_5565,N_4824,N_4738);
or U5566 (N_5566,N_4168,N_4568);
nand U5567 (N_5567,N_4589,N_4520);
nand U5568 (N_5568,N_4640,N_4886);
and U5569 (N_5569,N_4200,N_4806);
or U5570 (N_5570,N_4036,N_4564);
xor U5571 (N_5571,N_4917,N_4586);
nand U5572 (N_5572,N_4941,N_4789);
and U5573 (N_5573,N_4637,N_4398);
nor U5574 (N_5574,N_4323,N_4119);
and U5575 (N_5575,N_4995,N_4028);
or U5576 (N_5576,N_4535,N_4694);
and U5577 (N_5577,N_4119,N_4711);
and U5578 (N_5578,N_4366,N_4361);
or U5579 (N_5579,N_4666,N_4344);
nor U5580 (N_5580,N_4875,N_4613);
nor U5581 (N_5581,N_4556,N_4309);
or U5582 (N_5582,N_4656,N_4739);
and U5583 (N_5583,N_4930,N_4535);
nand U5584 (N_5584,N_4500,N_4312);
nand U5585 (N_5585,N_4857,N_4237);
xnor U5586 (N_5586,N_4340,N_4726);
and U5587 (N_5587,N_4340,N_4478);
nand U5588 (N_5588,N_4354,N_4104);
xor U5589 (N_5589,N_4884,N_4741);
nor U5590 (N_5590,N_4427,N_4868);
xnor U5591 (N_5591,N_4396,N_4536);
and U5592 (N_5592,N_4312,N_4823);
or U5593 (N_5593,N_4770,N_4133);
and U5594 (N_5594,N_4485,N_4244);
nor U5595 (N_5595,N_4008,N_4547);
nor U5596 (N_5596,N_4232,N_4793);
or U5597 (N_5597,N_4810,N_4933);
nor U5598 (N_5598,N_4548,N_4348);
or U5599 (N_5599,N_4949,N_4893);
nor U5600 (N_5600,N_4978,N_4121);
nand U5601 (N_5601,N_4357,N_4986);
nor U5602 (N_5602,N_4248,N_4230);
or U5603 (N_5603,N_4631,N_4193);
nor U5604 (N_5604,N_4376,N_4948);
and U5605 (N_5605,N_4050,N_4558);
xor U5606 (N_5606,N_4846,N_4204);
nor U5607 (N_5607,N_4146,N_4167);
and U5608 (N_5608,N_4274,N_4168);
or U5609 (N_5609,N_4074,N_4293);
nand U5610 (N_5610,N_4153,N_4352);
nor U5611 (N_5611,N_4718,N_4571);
nand U5612 (N_5612,N_4085,N_4272);
nor U5613 (N_5613,N_4486,N_4375);
or U5614 (N_5614,N_4608,N_4639);
and U5615 (N_5615,N_4537,N_4030);
and U5616 (N_5616,N_4165,N_4248);
nand U5617 (N_5617,N_4140,N_4869);
and U5618 (N_5618,N_4202,N_4415);
nor U5619 (N_5619,N_4328,N_4249);
or U5620 (N_5620,N_4152,N_4681);
nor U5621 (N_5621,N_4522,N_4313);
nor U5622 (N_5622,N_4505,N_4977);
nor U5623 (N_5623,N_4718,N_4208);
and U5624 (N_5624,N_4771,N_4836);
nand U5625 (N_5625,N_4734,N_4893);
and U5626 (N_5626,N_4239,N_4025);
xor U5627 (N_5627,N_4482,N_4311);
nor U5628 (N_5628,N_4611,N_4583);
nand U5629 (N_5629,N_4884,N_4576);
xor U5630 (N_5630,N_4682,N_4670);
and U5631 (N_5631,N_4930,N_4210);
xor U5632 (N_5632,N_4614,N_4905);
or U5633 (N_5633,N_4648,N_4959);
nor U5634 (N_5634,N_4690,N_4975);
xnor U5635 (N_5635,N_4770,N_4264);
or U5636 (N_5636,N_4011,N_4195);
nand U5637 (N_5637,N_4826,N_4874);
nor U5638 (N_5638,N_4155,N_4601);
and U5639 (N_5639,N_4785,N_4033);
xor U5640 (N_5640,N_4202,N_4414);
nor U5641 (N_5641,N_4102,N_4685);
and U5642 (N_5642,N_4743,N_4073);
or U5643 (N_5643,N_4742,N_4527);
nand U5644 (N_5644,N_4925,N_4935);
and U5645 (N_5645,N_4707,N_4607);
nand U5646 (N_5646,N_4485,N_4926);
nand U5647 (N_5647,N_4609,N_4198);
nor U5648 (N_5648,N_4166,N_4520);
and U5649 (N_5649,N_4783,N_4440);
nand U5650 (N_5650,N_4617,N_4705);
xnor U5651 (N_5651,N_4292,N_4682);
or U5652 (N_5652,N_4727,N_4104);
and U5653 (N_5653,N_4259,N_4696);
nand U5654 (N_5654,N_4595,N_4433);
xor U5655 (N_5655,N_4833,N_4519);
nand U5656 (N_5656,N_4370,N_4751);
nand U5657 (N_5657,N_4668,N_4066);
xnor U5658 (N_5658,N_4874,N_4416);
and U5659 (N_5659,N_4521,N_4695);
or U5660 (N_5660,N_4095,N_4019);
or U5661 (N_5661,N_4922,N_4830);
nand U5662 (N_5662,N_4592,N_4781);
or U5663 (N_5663,N_4639,N_4927);
nand U5664 (N_5664,N_4572,N_4424);
nor U5665 (N_5665,N_4737,N_4065);
xor U5666 (N_5666,N_4154,N_4456);
nor U5667 (N_5667,N_4246,N_4897);
nor U5668 (N_5668,N_4877,N_4558);
nand U5669 (N_5669,N_4772,N_4844);
nor U5670 (N_5670,N_4447,N_4470);
nand U5671 (N_5671,N_4106,N_4019);
nor U5672 (N_5672,N_4345,N_4541);
or U5673 (N_5673,N_4552,N_4316);
xor U5674 (N_5674,N_4835,N_4242);
and U5675 (N_5675,N_4534,N_4309);
or U5676 (N_5676,N_4957,N_4617);
nand U5677 (N_5677,N_4496,N_4783);
nor U5678 (N_5678,N_4357,N_4527);
nand U5679 (N_5679,N_4801,N_4470);
or U5680 (N_5680,N_4339,N_4882);
nor U5681 (N_5681,N_4664,N_4917);
xnor U5682 (N_5682,N_4526,N_4234);
xor U5683 (N_5683,N_4708,N_4692);
or U5684 (N_5684,N_4993,N_4862);
or U5685 (N_5685,N_4375,N_4271);
xor U5686 (N_5686,N_4296,N_4744);
nand U5687 (N_5687,N_4924,N_4514);
xor U5688 (N_5688,N_4266,N_4128);
or U5689 (N_5689,N_4676,N_4177);
xor U5690 (N_5690,N_4534,N_4390);
or U5691 (N_5691,N_4188,N_4839);
and U5692 (N_5692,N_4010,N_4181);
or U5693 (N_5693,N_4393,N_4695);
nor U5694 (N_5694,N_4946,N_4575);
nor U5695 (N_5695,N_4776,N_4070);
and U5696 (N_5696,N_4948,N_4481);
nor U5697 (N_5697,N_4963,N_4424);
nor U5698 (N_5698,N_4643,N_4237);
or U5699 (N_5699,N_4843,N_4632);
xor U5700 (N_5700,N_4948,N_4678);
xnor U5701 (N_5701,N_4992,N_4330);
nor U5702 (N_5702,N_4680,N_4199);
and U5703 (N_5703,N_4473,N_4830);
xnor U5704 (N_5704,N_4409,N_4089);
nand U5705 (N_5705,N_4251,N_4747);
or U5706 (N_5706,N_4345,N_4036);
and U5707 (N_5707,N_4456,N_4001);
nand U5708 (N_5708,N_4796,N_4434);
nor U5709 (N_5709,N_4153,N_4569);
nand U5710 (N_5710,N_4637,N_4990);
or U5711 (N_5711,N_4890,N_4938);
nor U5712 (N_5712,N_4139,N_4136);
and U5713 (N_5713,N_4541,N_4977);
and U5714 (N_5714,N_4570,N_4537);
and U5715 (N_5715,N_4312,N_4260);
and U5716 (N_5716,N_4352,N_4217);
and U5717 (N_5717,N_4056,N_4800);
or U5718 (N_5718,N_4876,N_4170);
xnor U5719 (N_5719,N_4987,N_4662);
or U5720 (N_5720,N_4011,N_4196);
and U5721 (N_5721,N_4724,N_4788);
nor U5722 (N_5722,N_4938,N_4639);
or U5723 (N_5723,N_4239,N_4295);
or U5724 (N_5724,N_4828,N_4467);
and U5725 (N_5725,N_4662,N_4051);
and U5726 (N_5726,N_4292,N_4084);
or U5727 (N_5727,N_4493,N_4847);
nor U5728 (N_5728,N_4260,N_4463);
nand U5729 (N_5729,N_4625,N_4899);
or U5730 (N_5730,N_4530,N_4439);
and U5731 (N_5731,N_4214,N_4843);
or U5732 (N_5732,N_4659,N_4824);
and U5733 (N_5733,N_4741,N_4150);
or U5734 (N_5734,N_4139,N_4878);
or U5735 (N_5735,N_4464,N_4947);
and U5736 (N_5736,N_4088,N_4598);
or U5737 (N_5737,N_4228,N_4602);
nor U5738 (N_5738,N_4184,N_4129);
and U5739 (N_5739,N_4220,N_4291);
and U5740 (N_5740,N_4933,N_4110);
or U5741 (N_5741,N_4254,N_4438);
and U5742 (N_5742,N_4888,N_4628);
nor U5743 (N_5743,N_4373,N_4125);
nor U5744 (N_5744,N_4964,N_4366);
nor U5745 (N_5745,N_4364,N_4810);
and U5746 (N_5746,N_4853,N_4191);
nand U5747 (N_5747,N_4154,N_4450);
nor U5748 (N_5748,N_4042,N_4735);
and U5749 (N_5749,N_4242,N_4226);
or U5750 (N_5750,N_4382,N_4981);
and U5751 (N_5751,N_4865,N_4680);
or U5752 (N_5752,N_4837,N_4512);
nand U5753 (N_5753,N_4700,N_4002);
and U5754 (N_5754,N_4200,N_4777);
nor U5755 (N_5755,N_4736,N_4588);
or U5756 (N_5756,N_4453,N_4268);
xnor U5757 (N_5757,N_4116,N_4478);
and U5758 (N_5758,N_4079,N_4486);
nand U5759 (N_5759,N_4713,N_4597);
and U5760 (N_5760,N_4403,N_4484);
nor U5761 (N_5761,N_4556,N_4731);
and U5762 (N_5762,N_4348,N_4535);
nand U5763 (N_5763,N_4217,N_4203);
nand U5764 (N_5764,N_4807,N_4750);
or U5765 (N_5765,N_4497,N_4652);
and U5766 (N_5766,N_4699,N_4356);
and U5767 (N_5767,N_4569,N_4381);
nor U5768 (N_5768,N_4120,N_4044);
nand U5769 (N_5769,N_4833,N_4721);
and U5770 (N_5770,N_4060,N_4437);
xnor U5771 (N_5771,N_4295,N_4215);
and U5772 (N_5772,N_4049,N_4374);
and U5773 (N_5773,N_4009,N_4722);
xor U5774 (N_5774,N_4430,N_4122);
nand U5775 (N_5775,N_4099,N_4924);
nand U5776 (N_5776,N_4400,N_4282);
nand U5777 (N_5777,N_4955,N_4642);
or U5778 (N_5778,N_4095,N_4407);
nor U5779 (N_5779,N_4134,N_4098);
xor U5780 (N_5780,N_4439,N_4726);
nor U5781 (N_5781,N_4706,N_4849);
or U5782 (N_5782,N_4619,N_4566);
or U5783 (N_5783,N_4326,N_4810);
or U5784 (N_5784,N_4199,N_4738);
xnor U5785 (N_5785,N_4307,N_4026);
and U5786 (N_5786,N_4655,N_4896);
and U5787 (N_5787,N_4670,N_4769);
nor U5788 (N_5788,N_4040,N_4179);
nor U5789 (N_5789,N_4217,N_4256);
or U5790 (N_5790,N_4448,N_4809);
or U5791 (N_5791,N_4697,N_4682);
or U5792 (N_5792,N_4317,N_4246);
nor U5793 (N_5793,N_4064,N_4379);
or U5794 (N_5794,N_4375,N_4650);
xor U5795 (N_5795,N_4161,N_4002);
nor U5796 (N_5796,N_4358,N_4238);
or U5797 (N_5797,N_4266,N_4935);
or U5798 (N_5798,N_4195,N_4662);
and U5799 (N_5799,N_4799,N_4978);
nor U5800 (N_5800,N_4948,N_4654);
nand U5801 (N_5801,N_4015,N_4929);
or U5802 (N_5802,N_4642,N_4096);
and U5803 (N_5803,N_4775,N_4150);
and U5804 (N_5804,N_4615,N_4310);
or U5805 (N_5805,N_4840,N_4034);
nand U5806 (N_5806,N_4841,N_4212);
and U5807 (N_5807,N_4780,N_4770);
or U5808 (N_5808,N_4736,N_4271);
or U5809 (N_5809,N_4252,N_4784);
nand U5810 (N_5810,N_4776,N_4479);
or U5811 (N_5811,N_4955,N_4046);
nor U5812 (N_5812,N_4596,N_4593);
nor U5813 (N_5813,N_4451,N_4681);
or U5814 (N_5814,N_4033,N_4401);
nand U5815 (N_5815,N_4136,N_4464);
xnor U5816 (N_5816,N_4197,N_4250);
xor U5817 (N_5817,N_4047,N_4060);
or U5818 (N_5818,N_4686,N_4362);
nor U5819 (N_5819,N_4524,N_4076);
xor U5820 (N_5820,N_4831,N_4833);
and U5821 (N_5821,N_4242,N_4189);
nand U5822 (N_5822,N_4363,N_4255);
nand U5823 (N_5823,N_4809,N_4426);
and U5824 (N_5824,N_4588,N_4822);
nand U5825 (N_5825,N_4923,N_4304);
nor U5826 (N_5826,N_4771,N_4900);
and U5827 (N_5827,N_4445,N_4541);
nor U5828 (N_5828,N_4759,N_4267);
or U5829 (N_5829,N_4115,N_4481);
nor U5830 (N_5830,N_4772,N_4994);
nor U5831 (N_5831,N_4026,N_4330);
and U5832 (N_5832,N_4850,N_4935);
nand U5833 (N_5833,N_4565,N_4502);
nand U5834 (N_5834,N_4546,N_4806);
xnor U5835 (N_5835,N_4233,N_4551);
and U5836 (N_5836,N_4929,N_4426);
nor U5837 (N_5837,N_4366,N_4009);
nor U5838 (N_5838,N_4135,N_4198);
nand U5839 (N_5839,N_4537,N_4930);
nand U5840 (N_5840,N_4860,N_4385);
nor U5841 (N_5841,N_4190,N_4256);
or U5842 (N_5842,N_4004,N_4816);
nand U5843 (N_5843,N_4772,N_4440);
or U5844 (N_5844,N_4031,N_4272);
or U5845 (N_5845,N_4605,N_4539);
nor U5846 (N_5846,N_4942,N_4809);
nand U5847 (N_5847,N_4680,N_4340);
xor U5848 (N_5848,N_4152,N_4538);
or U5849 (N_5849,N_4107,N_4749);
and U5850 (N_5850,N_4741,N_4016);
nand U5851 (N_5851,N_4971,N_4731);
xor U5852 (N_5852,N_4603,N_4654);
and U5853 (N_5853,N_4431,N_4439);
or U5854 (N_5854,N_4094,N_4128);
xor U5855 (N_5855,N_4721,N_4234);
or U5856 (N_5856,N_4013,N_4507);
and U5857 (N_5857,N_4343,N_4345);
and U5858 (N_5858,N_4857,N_4792);
or U5859 (N_5859,N_4342,N_4038);
nor U5860 (N_5860,N_4474,N_4482);
nor U5861 (N_5861,N_4508,N_4612);
nor U5862 (N_5862,N_4201,N_4227);
nand U5863 (N_5863,N_4817,N_4443);
and U5864 (N_5864,N_4940,N_4913);
xor U5865 (N_5865,N_4886,N_4670);
xnor U5866 (N_5866,N_4594,N_4889);
nor U5867 (N_5867,N_4180,N_4725);
or U5868 (N_5868,N_4609,N_4221);
and U5869 (N_5869,N_4658,N_4743);
and U5870 (N_5870,N_4588,N_4707);
nand U5871 (N_5871,N_4117,N_4255);
nor U5872 (N_5872,N_4945,N_4528);
nand U5873 (N_5873,N_4547,N_4064);
and U5874 (N_5874,N_4847,N_4450);
or U5875 (N_5875,N_4597,N_4678);
nand U5876 (N_5876,N_4860,N_4606);
nor U5877 (N_5877,N_4927,N_4812);
or U5878 (N_5878,N_4858,N_4604);
nor U5879 (N_5879,N_4823,N_4514);
or U5880 (N_5880,N_4287,N_4760);
nand U5881 (N_5881,N_4673,N_4807);
and U5882 (N_5882,N_4273,N_4033);
and U5883 (N_5883,N_4242,N_4447);
nor U5884 (N_5884,N_4287,N_4446);
and U5885 (N_5885,N_4184,N_4701);
nand U5886 (N_5886,N_4133,N_4626);
nor U5887 (N_5887,N_4239,N_4789);
and U5888 (N_5888,N_4834,N_4526);
nand U5889 (N_5889,N_4744,N_4020);
or U5890 (N_5890,N_4881,N_4169);
xnor U5891 (N_5891,N_4502,N_4590);
and U5892 (N_5892,N_4422,N_4168);
and U5893 (N_5893,N_4971,N_4738);
nor U5894 (N_5894,N_4004,N_4190);
xnor U5895 (N_5895,N_4558,N_4386);
nor U5896 (N_5896,N_4883,N_4787);
nor U5897 (N_5897,N_4048,N_4753);
and U5898 (N_5898,N_4686,N_4811);
xnor U5899 (N_5899,N_4309,N_4627);
nor U5900 (N_5900,N_4131,N_4265);
nor U5901 (N_5901,N_4709,N_4463);
nand U5902 (N_5902,N_4671,N_4909);
or U5903 (N_5903,N_4156,N_4007);
or U5904 (N_5904,N_4796,N_4192);
nor U5905 (N_5905,N_4797,N_4035);
and U5906 (N_5906,N_4219,N_4304);
or U5907 (N_5907,N_4415,N_4133);
or U5908 (N_5908,N_4820,N_4266);
and U5909 (N_5909,N_4316,N_4521);
nand U5910 (N_5910,N_4760,N_4208);
xor U5911 (N_5911,N_4860,N_4216);
nand U5912 (N_5912,N_4297,N_4244);
and U5913 (N_5913,N_4941,N_4279);
nand U5914 (N_5914,N_4484,N_4429);
or U5915 (N_5915,N_4923,N_4476);
or U5916 (N_5916,N_4883,N_4194);
nand U5917 (N_5917,N_4339,N_4986);
or U5918 (N_5918,N_4290,N_4143);
or U5919 (N_5919,N_4802,N_4434);
nand U5920 (N_5920,N_4458,N_4927);
or U5921 (N_5921,N_4624,N_4143);
nor U5922 (N_5922,N_4121,N_4649);
nor U5923 (N_5923,N_4978,N_4728);
or U5924 (N_5924,N_4827,N_4884);
xor U5925 (N_5925,N_4706,N_4384);
or U5926 (N_5926,N_4086,N_4327);
or U5927 (N_5927,N_4995,N_4554);
nand U5928 (N_5928,N_4360,N_4260);
or U5929 (N_5929,N_4475,N_4009);
nor U5930 (N_5930,N_4204,N_4387);
and U5931 (N_5931,N_4326,N_4292);
nand U5932 (N_5932,N_4644,N_4274);
or U5933 (N_5933,N_4097,N_4680);
or U5934 (N_5934,N_4059,N_4734);
and U5935 (N_5935,N_4783,N_4125);
and U5936 (N_5936,N_4502,N_4832);
or U5937 (N_5937,N_4293,N_4771);
nand U5938 (N_5938,N_4780,N_4184);
or U5939 (N_5939,N_4957,N_4014);
nand U5940 (N_5940,N_4005,N_4058);
nor U5941 (N_5941,N_4529,N_4195);
nor U5942 (N_5942,N_4695,N_4826);
and U5943 (N_5943,N_4900,N_4375);
or U5944 (N_5944,N_4925,N_4005);
nand U5945 (N_5945,N_4627,N_4235);
nand U5946 (N_5946,N_4190,N_4147);
nand U5947 (N_5947,N_4315,N_4818);
nor U5948 (N_5948,N_4362,N_4753);
nand U5949 (N_5949,N_4617,N_4263);
or U5950 (N_5950,N_4764,N_4955);
nand U5951 (N_5951,N_4438,N_4312);
or U5952 (N_5952,N_4738,N_4123);
nand U5953 (N_5953,N_4415,N_4507);
nor U5954 (N_5954,N_4276,N_4007);
and U5955 (N_5955,N_4017,N_4909);
nand U5956 (N_5956,N_4008,N_4033);
nand U5957 (N_5957,N_4768,N_4582);
nor U5958 (N_5958,N_4430,N_4607);
or U5959 (N_5959,N_4626,N_4398);
and U5960 (N_5960,N_4302,N_4251);
nor U5961 (N_5961,N_4472,N_4091);
nor U5962 (N_5962,N_4948,N_4774);
xor U5963 (N_5963,N_4234,N_4016);
nand U5964 (N_5964,N_4611,N_4595);
and U5965 (N_5965,N_4886,N_4388);
and U5966 (N_5966,N_4016,N_4960);
nor U5967 (N_5967,N_4434,N_4341);
nor U5968 (N_5968,N_4710,N_4780);
or U5969 (N_5969,N_4856,N_4602);
nor U5970 (N_5970,N_4349,N_4397);
or U5971 (N_5971,N_4157,N_4999);
nor U5972 (N_5972,N_4076,N_4060);
nand U5973 (N_5973,N_4915,N_4026);
or U5974 (N_5974,N_4620,N_4512);
or U5975 (N_5975,N_4518,N_4793);
or U5976 (N_5976,N_4955,N_4784);
nand U5977 (N_5977,N_4178,N_4676);
and U5978 (N_5978,N_4909,N_4493);
nand U5979 (N_5979,N_4238,N_4270);
and U5980 (N_5980,N_4572,N_4978);
nor U5981 (N_5981,N_4587,N_4749);
or U5982 (N_5982,N_4573,N_4238);
and U5983 (N_5983,N_4526,N_4840);
nand U5984 (N_5984,N_4937,N_4857);
nor U5985 (N_5985,N_4444,N_4184);
and U5986 (N_5986,N_4488,N_4762);
and U5987 (N_5987,N_4094,N_4878);
xnor U5988 (N_5988,N_4787,N_4518);
nor U5989 (N_5989,N_4043,N_4654);
and U5990 (N_5990,N_4440,N_4060);
or U5991 (N_5991,N_4447,N_4584);
nand U5992 (N_5992,N_4248,N_4714);
nor U5993 (N_5993,N_4329,N_4689);
nor U5994 (N_5994,N_4095,N_4973);
and U5995 (N_5995,N_4905,N_4627);
or U5996 (N_5996,N_4815,N_4835);
and U5997 (N_5997,N_4130,N_4363);
nand U5998 (N_5998,N_4964,N_4036);
or U5999 (N_5999,N_4346,N_4541);
or U6000 (N_6000,N_5202,N_5752);
nor U6001 (N_6001,N_5015,N_5271);
and U6002 (N_6002,N_5769,N_5732);
xor U6003 (N_6003,N_5276,N_5108);
or U6004 (N_6004,N_5505,N_5217);
nor U6005 (N_6005,N_5790,N_5864);
nand U6006 (N_6006,N_5126,N_5510);
xor U6007 (N_6007,N_5266,N_5008);
nand U6008 (N_6008,N_5262,N_5423);
and U6009 (N_6009,N_5645,N_5796);
nor U6010 (N_6010,N_5178,N_5983);
nor U6011 (N_6011,N_5048,N_5502);
nor U6012 (N_6012,N_5414,N_5124);
or U6013 (N_6013,N_5894,N_5936);
or U6014 (N_6014,N_5078,N_5285);
nor U6015 (N_6015,N_5735,N_5294);
nand U6016 (N_6016,N_5397,N_5680);
and U6017 (N_6017,N_5258,N_5069);
nand U6018 (N_6018,N_5558,N_5738);
nor U6019 (N_6019,N_5062,N_5213);
or U6020 (N_6020,N_5125,N_5961);
nor U6021 (N_6021,N_5185,N_5274);
or U6022 (N_6022,N_5902,N_5569);
nand U6023 (N_6023,N_5838,N_5798);
nor U6024 (N_6024,N_5599,N_5167);
or U6025 (N_6025,N_5565,N_5683);
or U6026 (N_6026,N_5956,N_5340);
nand U6027 (N_6027,N_5914,N_5483);
xor U6028 (N_6028,N_5550,N_5834);
xnor U6029 (N_6029,N_5836,N_5288);
and U6030 (N_6030,N_5652,N_5718);
or U6031 (N_6031,N_5165,N_5189);
and U6032 (N_6032,N_5139,N_5454);
nand U6033 (N_6033,N_5153,N_5416);
or U6034 (N_6034,N_5968,N_5360);
nand U6035 (N_6035,N_5351,N_5622);
nor U6036 (N_6036,N_5916,N_5321);
and U6037 (N_6037,N_5694,N_5417);
nor U6038 (N_6038,N_5230,N_5614);
nand U6039 (N_6039,N_5155,N_5150);
or U6040 (N_6040,N_5160,N_5282);
or U6041 (N_6041,N_5715,N_5755);
nor U6042 (N_6042,N_5335,N_5609);
and U6043 (N_6043,N_5898,N_5758);
nand U6044 (N_6044,N_5116,N_5862);
and U6045 (N_6045,N_5813,N_5883);
or U6046 (N_6046,N_5456,N_5601);
and U6047 (N_6047,N_5990,N_5513);
nor U6048 (N_6048,N_5053,N_5032);
or U6049 (N_6049,N_5603,N_5042);
nand U6050 (N_6050,N_5237,N_5491);
or U6051 (N_6051,N_5016,N_5224);
nor U6052 (N_6052,N_5998,N_5257);
and U6053 (N_6053,N_5296,N_5413);
and U6054 (N_6054,N_5842,N_5904);
xor U6055 (N_6055,N_5049,N_5889);
nor U6056 (N_6056,N_5566,N_5159);
and U6057 (N_6057,N_5547,N_5887);
nor U6058 (N_6058,N_5602,N_5358);
or U6059 (N_6059,N_5175,N_5372);
and U6060 (N_6060,N_5587,N_5176);
xnor U6061 (N_6061,N_5563,N_5831);
nor U6062 (N_6062,N_5516,N_5468);
or U6063 (N_6063,N_5844,N_5597);
xor U6064 (N_6064,N_5627,N_5791);
nor U6065 (N_6065,N_5545,N_5070);
or U6066 (N_6066,N_5264,N_5763);
nand U6067 (N_6067,N_5367,N_5024);
nor U6068 (N_6068,N_5621,N_5462);
xnor U6069 (N_6069,N_5691,N_5700);
nand U6070 (N_6070,N_5331,N_5992);
and U6071 (N_6071,N_5072,N_5435);
or U6072 (N_6072,N_5112,N_5648);
nor U6073 (N_6073,N_5338,N_5754);
and U6074 (N_6074,N_5444,N_5706);
nor U6075 (N_6075,N_5507,N_5439);
nand U6076 (N_6076,N_5649,N_5089);
and U6077 (N_6077,N_5682,N_5473);
nor U6078 (N_6078,N_5390,N_5580);
nor U6079 (N_6079,N_5865,N_5559);
nor U6080 (N_6080,N_5337,N_5501);
or U6081 (N_6081,N_5084,N_5747);
and U6082 (N_6082,N_5114,N_5945);
or U6083 (N_6083,N_5030,N_5544);
nor U6084 (N_6084,N_5477,N_5370);
and U6085 (N_6085,N_5302,N_5971);
or U6086 (N_6086,N_5161,N_5443);
or U6087 (N_6087,N_5759,N_5846);
nor U6088 (N_6088,N_5820,N_5994);
nor U6089 (N_6089,N_5774,N_5673);
nand U6090 (N_6090,N_5654,N_5240);
nand U6091 (N_6091,N_5293,N_5490);
or U6092 (N_6092,N_5907,N_5970);
nand U6093 (N_6093,N_5981,N_5623);
nand U6094 (N_6094,N_5256,N_5832);
nor U6095 (N_6095,N_5695,N_5822);
nor U6096 (N_6096,N_5385,N_5440);
nor U6097 (N_6097,N_5381,N_5849);
nor U6098 (N_6098,N_5221,N_5085);
and U6099 (N_6099,N_5146,N_5812);
and U6100 (N_6100,N_5380,N_5805);
or U6101 (N_6101,N_5847,N_5204);
nor U6102 (N_6102,N_5869,N_5951);
and U6103 (N_6103,N_5325,N_5102);
xnor U6104 (N_6104,N_5690,N_5060);
nor U6105 (N_6105,N_5203,N_5273);
nor U6106 (N_6106,N_5814,N_5918);
or U6107 (N_6107,N_5944,N_5960);
or U6108 (N_6108,N_5263,N_5553);
and U6109 (N_6109,N_5729,N_5934);
and U6110 (N_6110,N_5811,N_5641);
nand U6111 (N_6111,N_5679,N_5574);
and U6112 (N_6112,N_5923,N_5073);
and U6113 (N_6113,N_5929,N_5753);
or U6114 (N_6114,N_5198,N_5947);
or U6115 (N_6115,N_5527,N_5383);
xnor U6116 (N_6116,N_5770,N_5295);
nor U6117 (N_6117,N_5942,N_5526);
nor U6118 (N_6118,N_5626,N_5216);
or U6119 (N_6119,N_5967,N_5669);
nand U6120 (N_6120,N_5333,N_5142);
and U6121 (N_6121,N_5304,N_5637);
nor U6122 (N_6122,N_5064,N_5453);
or U6123 (N_6123,N_5434,N_5620);
and U6124 (N_6124,N_5817,N_5267);
or U6125 (N_6125,N_5474,N_5003);
nand U6126 (N_6126,N_5315,N_5644);
nor U6127 (N_6127,N_5661,N_5861);
or U6128 (N_6128,N_5253,N_5011);
nand U6129 (N_6129,N_5006,N_5152);
nand U6130 (N_6130,N_5249,N_5895);
or U6131 (N_6131,N_5464,N_5816);
or U6132 (N_6132,N_5797,N_5026);
xor U6133 (N_6133,N_5038,N_5875);
nor U6134 (N_6134,N_5134,N_5903);
nor U6135 (N_6135,N_5876,N_5455);
nor U6136 (N_6136,N_5215,N_5299);
nand U6137 (N_6137,N_5672,N_5191);
and U6138 (N_6138,N_5879,N_5306);
nor U6139 (N_6139,N_5818,N_5481);
nand U6140 (N_6140,N_5972,N_5854);
and U6141 (N_6141,N_5398,N_5147);
or U6142 (N_6142,N_5166,N_5128);
or U6143 (N_6143,N_5183,N_5686);
or U6144 (N_6144,N_5487,N_5292);
nor U6145 (N_6145,N_5827,N_5105);
nand U6146 (N_6146,N_5259,N_5446);
nor U6147 (N_6147,N_5873,N_5789);
or U6148 (N_6148,N_5538,N_5039);
nand U6149 (N_6149,N_5077,N_5478);
nor U6150 (N_6150,N_5629,N_5855);
nand U6151 (N_6151,N_5872,N_5802);
or U6152 (N_6152,N_5792,N_5938);
nor U6153 (N_6153,N_5303,N_5449);
and U6154 (N_6154,N_5200,N_5721);
xor U6155 (N_6155,N_5562,N_5014);
or U6156 (N_6156,N_5190,N_5308);
or U6157 (N_6157,N_5788,N_5157);
nand U6158 (N_6158,N_5371,N_5726);
and U6159 (N_6159,N_5619,N_5036);
and U6160 (N_6160,N_5209,N_5823);
or U6161 (N_6161,N_5226,N_5137);
nand U6162 (N_6162,N_5332,N_5833);
and U6163 (N_6163,N_5095,N_5924);
nand U6164 (N_6164,N_5618,N_5127);
nor U6165 (N_6165,N_5821,N_5133);
nand U6166 (N_6166,N_5368,N_5988);
nand U6167 (N_6167,N_5714,N_5437);
and U6168 (N_6168,N_5859,N_5999);
or U6169 (N_6169,N_5570,N_5841);
and U6170 (N_6170,N_5762,N_5467);
nor U6171 (N_6171,N_5132,N_5551);
and U6172 (N_6172,N_5596,N_5197);
xnor U6173 (N_6173,N_5965,N_5906);
and U6174 (N_6174,N_5395,N_5734);
or U6175 (N_6175,N_5799,N_5674);
or U6176 (N_6176,N_5935,N_5109);
and U6177 (N_6177,N_5098,N_5377);
nand U6178 (N_6178,N_5756,N_5366);
xnor U6179 (N_6179,N_5031,N_5640);
xor U6180 (N_6180,N_5279,N_5436);
nor U6181 (N_6181,N_5460,N_5013);
nand U6182 (N_6182,N_5853,N_5701);
or U6183 (N_6183,N_5079,N_5671);
xor U6184 (N_6184,N_5930,N_5451);
and U6185 (N_6185,N_5291,N_5245);
nand U6186 (N_6186,N_5548,N_5374);
or U6187 (N_6187,N_5007,N_5472);
and U6188 (N_6188,N_5466,N_5919);
nor U6189 (N_6189,N_5503,N_5040);
nand U6190 (N_6190,N_5019,N_5184);
nor U6191 (N_6191,N_5524,N_5731);
nor U6192 (N_6192,N_5611,N_5705);
and U6193 (N_6193,N_5409,N_5432);
and U6194 (N_6194,N_5815,N_5996);
xor U6195 (N_6195,N_5037,N_5681);
or U6196 (N_6196,N_5359,N_5350);
nor U6197 (N_6197,N_5154,N_5412);
and U6198 (N_6198,N_5653,N_5430);
nor U6199 (N_6199,N_5606,N_5092);
and U6200 (N_6200,N_5239,N_5136);
nor U6201 (N_6201,N_5195,N_5891);
or U6202 (N_6202,N_5585,N_5260);
and U6203 (N_6203,N_5969,N_5751);
nand U6204 (N_6204,N_5452,N_5741);
or U6205 (N_6205,N_5989,N_5497);
nand U6206 (N_6206,N_5174,N_5808);
or U6207 (N_6207,N_5022,N_5584);
nand U6208 (N_6208,N_5055,N_5532);
or U6209 (N_6209,N_5170,N_5206);
nor U6210 (N_6210,N_5415,N_5075);
or U6211 (N_6211,N_5591,N_5948);
and U6212 (N_6212,N_5489,N_5984);
and U6213 (N_6213,N_5693,N_5687);
or U6214 (N_6214,N_5535,N_5512);
nor U6215 (N_6215,N_5608,N_5579);
and U6216 (N_6216,N_5913,N_5362);
and U6217 (N_6217,N_5399,N_5225);
nand U6218 (N_6218,N_5987,N_5678);
nor U6219 (N_6219,N_5486,N_5405);
nor U6220 (N_6220,N_5047,N_5275);
xor U6221 (N_6221,N_5312,N_5921);
and U6222 (N_6222,N_5378,N_5712);
nor U6223 (N_6223,N_5051,N_5012);
or U6224 (N_6224,N_5773,N_5530);
nand U6225 (N_6225,N_5056,N_5511);
nand U6226 (N_6226,N_5401,N_5061);
or U6227 (N_6227,N_5534,N_5809);
or U6228 (N_6228,N_5316,N_5283);
nand U6229 (N_6229,N_5779,N_5218);
or U6230 (N_6230,N_5748,N_5991);
or U6231 (N_6231,N_5342,N_5193);
or U6232 (N_6232,N_5800,N_5556);
or U6233 (N_6233,N_5871,N_5954);
or U6234 (N_6234,N_5976,N_5063);
nor U6235 (N_6235,N_5442,N_5625);
nor U6236 (N_6236,N_5711,N_5471);
nor U6237 (N_6237,N_5171,N_5247);
nand U6238 (N_6238,N_5708,N_5707);
or U6239 (N_6239,N_5552,N_5313);
and U6240 (N_6240,N_5113,N_5665);
nand U6241 (N_6241,N_5568,N_5910);
nor U6242 (N_6242,N_5586,N_5717);
xnor U6243 (N_6243,N_5349,N_5392);
nand U6244 (N_6244,N_5144,N_5476);
or U6245 (N_6245,N_5341,N_5244);
or U6246 (N_6246,N_5959,N_5784);
nand U6247 (N_6247,N_5946,N_5433);
and U6248 (N_6248,N_5120,N_5713);
and U6249 (N_6249,N_5777,N_5517);
or U6250 (N_6250,N_5973,N_5254);
or U6251 (N_6251,N_5963,N_5506);
nand U6252 (N_6252,N_5172,N_5234);
nor U6253 (N_6253,N_5484,N_5839);
and U6254 (N_6254,N_5575,N_5101);
nand U6255 (N_6255,N_5091,N_5870);
nand U6256 (N_6256,N_5287,N_5050);
nand U6257 (N_6257,N_5962,N_5749);
nor U6258 (N_6258,N_5199,N_5148);
nor U6259 (N_6259,N_5280,N_5179);
and U6260 (N_6260,N_5843,N_5564);
and U6261 (N_6261,N_5458,N_5365);
and U6262 (N_6262,N_5323,N_5353);
and U6263 (N_6263,N_5314,N_5896);
or U6264 (N_6264,N_5448,N_5785);
nor U6265 (N_6265,N_5529,N_5957);
nand U6266 (N_6266,N_5094,N_5986);
nand U6267 (N_6267,N_5787,N_5310);
xnor U6268 (N_6268,N_5186,N_5241);
xor U6269 (N_6269,N_5235,N_5760);
and U6270 (N_6270,N_5743,N_5555);
nand U6271 (N_6271,N_5744,N_5656);
nand U6272 (N_6272,N_5400,N_5252);
or U6273 (N_6273,N_5793,N_5666);
or U6274 (N_6274,N_5428,N_5985);
and U6275 (N_6275,N_5858,N_5523);
nand U6276 (N_6276,N_5525,N_5837);
nand U6277 (N_6277,N_5950,N_5382);
or U6278 (N_6278,N_5236,N_5958);
or U6279 (N_6279,N_5210,N_5806);
and U6280 (N_6280,N_5496,N_5508);
xnor U6281 (N_6281,N_5086,N_5182);
or U6282 (N_6282,N_5018,N_5131);
nand U6283 (N_6283,N_5495,N_5781);
and U6284 (N_6284,N_5357,N_5117);
xnor U6285 (N_6285,N_5001,N_5519);
or U6286 (N_6286,N_5255,N_5647);
nor U6287 (N_6287,N_5461,N_5121);
nor U6288 (N_6288,N_5169,N_5531);
nor U6289 (N_6289,N_5670,N_5498);
and U6290 (N_6290,N_5703,N_5677);
nor U6291 (N_6291,N_5766,N_5201);
and U6292 (N_6292,N_5940,N_5364);
nor U6293 (N_6293,N_5141,N_5388);
xor U6294 (N_6294,N_5933,N_5347);
nor U6295 (N_6295,N_5068,N_5156);
and U6296 (N_6296,N_5162,N_5727);
nor U6297 (N_6297,N_5445,N_5188);
xnor U6298 (N_6298,N_5422,N_5345);
xor U6299 (N_6299,N_5764,N_5192);
nand U6300 (N_6300,N_5305,N_5309);
and U6301 (N_6301,N_5881,N_5475);
nand U6302 (N_6302,N_5868,N_5856);
nor U6303 (N_6303,N_5557,N_5297);
or U6304 (N_6304,N_5181,N_5630);
or U6305 (N_6305,N_5593,N_5023);
xnor U6306 (N_6306,N_5598,N_5664);
and U6307 (N_6307,N_5689,N_5803);
xor U6308 (N_6308,N_5343,N_5403);
nor U6309 (N_6309,N_5915,N_5533);
nand U6310 (N_6310,N_5561,N_5901);
nand U6311 (N_6311,N_5927,N_5583);
nand U6312 (N_6312,N_5373,N_5804);
nor U6313 (N_6313,N_5232,N_5615);
nor U6314 (N_6314,N_5922,N_5667);
nand U6315 (N_6315,N_5576,N_5344);
nor U6316 (N_6316,N_5096,N_5493);
nand U6317 (N_6317,N_5431,N_5725);
and U6318 (N_6318,N_5830,N_5088);
or U6319 (N_6319,N_5326,N_5977);
or U6320 (N_6320,N_5046,N_5021);
or U6321 (N_6321,N_5499,N_5905);
xnor U6322 (N_6322,N_5421,N_5082);
nor U6323 (N_6323,N_5238,N_5867);
and U6324 (N_6324,N_5740,N_5278);
nand U6325 (N_6325,N_5354,N_5801);
or U6326 (N_6326,N_5389,N_5509);
nor U6327 (N_6327,N_5638,N_5767);
xnor U6328 (N_6328,N_5780,N_5187);
nand U6329 (N_6329,N_5227,N_5650);
nand U6330 (N_6330,N_5066,N_5076);
nand U6331 (N_6331,N_5613,N_5911);
nand U6332 (N_6332,N_5250,N_5407);
and U6333 (N_6333,N_5352,N_5418);
nand U6334 (N_6334,N_5723,N_5716);
nand U6335 (N_6335,N_5514,N_5194);
nor U6336 (N_6336,N_5540,N_5457);
nor U6337 (N_6337,N_5857,N_5272);
and U6338 (N_6338,N_5581,N_5783);
xor U6339 (N_6339,N_5692,N_5974);
nand U6340 (N_6340,N_5658,N_5745);
or U6341 (N_6341,N_5328,N_5301);
nor U6342 (N_6342,N_5546,N_5835);
and U6343 (N_6343,N_5000,N_5135);
nor U6344 (N_6344,N_5242,N_5982);
nor U6345 (N_6345,N_5010,N_5450);
or U6346 (N_6346,N_5233,N_5363);
nor U6347 (N_6347,N_5899,N_5852);
nor U6348 (N_6348,N_5775,N_5577);
or U6349 (N_6349,N_5387,N_5330);
nor U6350 (N_6350,N_5828,N_5427);
or U6351 (N_6351,N_5746,N_5663);
or U6352 (N_6352,N_5396,N_5408);
nand U6353 (N_6353,N_5494,N_5097);
nand U6354 (N_6354,N_5284,N_5543);
or U6355 (N_6355,N_5196,N_5027);
nor U6356 (N_6356,N_5628,N_5029);
nor U6357 (N_6357,N_5582,N_5251);
nand U6358 (N_6358,N_5324,N_5860);
nor U6359 (N_6359,N_5697,N_5688);
nor U6360 (N_6360,N_5877,N_5229);
or U6361 (N_6361,N_5020,N_5207);
nand U6362 (N_6362,N_5885,N_5052);
or U6363 (N_6363,N_5979,N_5765);
and U6364 (N_6364,N_5208,N_5660);
nor U6365 (N_6365,N_5463,N_5057);
and U6366 (N_6366,N_5728,N_5261);
nor U6367 (N_6367,N_5786,N_5702);
and U6368 (N_6368,N_5528,N_5426);
xor U6369 (N_6369,N_5866,N_5104);
and U6370 (N_6370,N_5676,N_5110);
xnor U6371 (N_6371,N_5739,N_5459);
nand U6372 (N_6372,N_5002,N_5168);
nor U6373 (N_6373,N_5925,N_5058);
nor U6374 (N_6374,N_5518,N_5699);
and U6375 (N_6375,N_5319,N_5953);
nor U6376 (N_6376,N_5140,N_5639);
nand U6377 (N_6377,N_5268,N_5897);
nor U6378 (N_6378,N_5908,N_5632);
or U6379 (N_6379,N_5311,N_5537);
or U6380 (N_6380,N_5067,N_5163);
nand U6381 (N_6381,N_5033,N_5900);
nor U6382 (N_6382,N_5662,N_5975);
nand U6383 (N_6383,N_5643,N_5485);
nor U6384 (N_6384,N_5219,N_5668);
nor U6385 (N_6385,N_5384,N_5009);
or U6386 (N_6386,N_5005,N_5411);
nand U6387 (N_6387,N_5522,N_5997);
xnor U6388 (N_6388,N_5317,N_5926);
xor U6389 (N_6389,N_5704,N_5243);
or U6390 (N_6390,N_5177,N_5882);
nand U6391 (N_6391,N_5920,N_5419);
nor U6392 (N_6392,N_5980,N_5778);
and U6393 (N_6393,N_5329,N_5750);
or U6394 (N_6394,N_5893,N_5955);
or U6395 (N_6395,N_5761,N_5685);
nor U6396 (N_6396,N_5824,N_5214);
nand U6397 (N_6397,N_5772,N_5736);
nand U6398 (N_6398,N_5059,N_5265);
nand U6399 (N_6399,N_5145,N_5205);
or U6400 (N_6400,N_5479,N_5572);
nand U6401 (N_6401,N_5949,N_5826);
nand U6402 (N_6402,N_5369,N_5932);
or U6403 (N_6403,N_5151,N_5093);
nand U6404 (N_6404,N_5480,N_5406);
and U6405 (N_6405,N_5404,N_5807);
or U6406 (N_6406,N_5318,N_5129);
nand U6407 (N_6407,N_5684,N_5829);
xor U6408 (N_6408,N_5617,N_5709);
xnor U6409 (N_6409,N_5521,N_5863);
or U6410 (N_6410,N_5710,N_5592);
nor U6411 (N_6411,N_5071,N_5567);
and U6412 (N_6412,N_5720,N_5542);
nor U6413 (N_6413,N_5825,N_5118);
or U6414 (N_6414,N_5044,N_5111);
and U6415 (N_6415,N_5536,N_5604);
nor U6416 (N_6416,N_5447,N_5361);
nand U6417 (N_6417,N_5103,N_5375);
and U6418 (N_6418,N_5635,N_5724);
nor U6419 (N_6419,N_5886,N_5890);
xor U6420 (N_6420,N_5616,N_5554);
or U6421 (N_6421,N_5045,N_5300);
nor U6422 (N_6422,N_5099,N_5659);
or U6423 (N_6423,N_5211,N_5269);
nand U6424 (N_6424,N_5090,N_5122);
and U6425 (N_6425,N_5081,N_5878);
or U6426 (N_6426,N_5376,N_5322);
nand U6427 (N_6427,N_5348,N_5470);
nor U6428 (N_6428,N_5771,N_5884);
or U6429 (N_6429,N_5675,N_5850);
nand U6430 (N_6430,N_5539,N_5336);
nand U6431 (N_6431,N_5130,N_5386);
xor U6432 (N_6432,N_5054,N_5143);
and U6433 (N_6433,N_5607,N_5429);
or U6434 (N_6434,N_5424,N_5290);
nand U6435 (N_6435,N_5943,N_5655);
nand U6436 (N_6436,N_5874,N_5776);
nor U6437 (N_6437,N_5931,N_5327);
nor U6438 (N_6438,N_5065,N_5100);
nor U6439 (N_6439,N_5115,N_5636);
or U6440 (N_6440,N_5173,N_5588);
and U6441 (N_6441,N_5119,N_5952);
or U6442 (N_6442,N_5610,N_5624);
nor U6443 (N_6443,N_5590,N_5356);
nand U6444 (N_6444,N_5482,N_5393);
and U6445 (N_6445,N_5041,N_5851);
nand U6446 (N_6446,N_5107,N_5560);
xor U6447 (N_6447,N_5488,N_5083);
xnor U6448 (N_6448,N_5917,N_5289);
nand U6449 (N_6449,N_5541,N_5425);
and U6450 (N_6450,N_5420,N_5220);
or U6451 (N_6451,N_5504,N_5270);
or U6452 (N_6452,N_5087,N_5978);
nor U6453 (N_6453,N_5594,N_5379);
nor U6454 (N_6454,N_5355,N_5909);
nand U6455 (N_6455,N_5228,N_5307);
nand U6456 (N_6456,N_5035,N_5605);
and U6457 (N_6457,N_5722,N_5231);
nor U6458 (N_6458,N_5515,N_5768);
or U6459 (N_6459,N_5025,N_5646);
or U6460 (N_6460,N_5346,N_5149);
nor U6461 (N_6461,N_5246,N_5123);
nor U6462 (N_6462,N_5657,N_5964);
nor U6463 (N_6463,N_5441,N_5028);
or U6464 (N_6464,N_5595,N_5438);
and U6465 (N_6465,N_5391,N_5469);
xnor U6466 (N_6466,N_5248,N_5600);
nand U6467 (N_6467,N_5017,N_5402);
nor U6468 (N_6468,N_5043,N_5819);
nor U6469 (N_6469,N_5223,N_5939);
nand U6470 (N_6470,N_5840,N_5730);
nand U6471 (N_6471,N_5286,N_5719);
nand U6472 (N_6472,N_5880,N_5612);
or U6473 (N_6473,N_5888,N_5394);
xnor U6474 (N_6474,N_5737,N_5848);
xnor U6475 (N_6475,N_5698,N_5794);
nand U6476 (N_6476,N_5281,N_5573);
nor U6477 (N_6477,N_5810,N_5912);
or U6478 (N_6478,N_5633,N_5549);
or U6479 (N_6479,N_5757,N_5164);
or U6480 (N_6480,N_5571,N_5500);
or U6481 (N_6481,N_5520,N_5180);
or U6482 (N_6482,N_5320,N_5642);
nand U6483 (N_6483,N_5993,N_5106);
and U6484 (N_6484,N_5004,N_5892);
nor U6485 (N_6485,N_5410,N_5222);
or U6486 (N_6486,N_5733,N_5334);
and U6487 (N_6487,N_5651,N_5212);
and U6488 (N_6488,N_5465,N_5034);
xor U6489 (N_6489,N_5845,N_5589);
nor U6490 (N_6490,N_5339,N_5795);
or U6491 (N_6491,N_5578,N_5937);
nand U6492 (N_6492,N_5074,N_5492);
nor U6493 (N_6493,N_5782,N_5158);
xor U6494 (N_6494,N_5138,N_5742);
nand U6495 (N_6495,N_5696,N_5298);
or U6496 (N_6496,N_5277,N_5080);
nor U6497 (N_6497,N_5634,N_5966);
nor U6498 (N_6498,N_5928,N_5995);
xnor U6499 (N_6499,N_5941,N_5631);
and U6500 (N_6500,N_5422,N_5133);
or U6501 (N_6501,N_5690,N_5314);
xnor U6502 (N_6502,N_5709,N_5151);
and U6503 (N_6503,N_5997,N_5325);
nand U6504 (N_6504,N_5128,N_5969);
and U6505 (N_6505,N_5403,N_5814);
nor U6506 (N_6506,N_5605,N_5870);
nor U6507 (N_6507,N_5237,N_5019);
nand U6508 (N_6508,N_5915,N_5119);
nand U6509 (N_6509,N_5728,N_5081);
and U6510 (N_6510,N_5137,N_5312);
and U6511 (N_6511,N_5449,N_5085);
and U6512 (N_6512,N_5940,N_5285);
nor U6513 (N_6513,N_5678,N_5593);
nand U6514 (N_6514,N_5667,N_5647);
and U6515 (N_6515,N_5480,N_5681);
and U6516 (N_6516,N_5438,N_5211);
or U6517 (N_6517,N_5498,N_5136);
or U6518 (N_6518,N_5638,N_5615);
nand U6519 (N_6519,N_5430,N_5435);
and U6520 (N_6520,N_5945,N_5373);
and U6521 (N_6521,N_5893,N_5342);
and U6522 (N_6522,N_5078,N_5110);
nor U6523 (N_6523,N_5294,N_5313);
nor U6524 (N_6524,N_5784,N_5558);
nand U6525 (N_6525,N_5695,N_5843);
or U6526 (N_6526,N_5544,N_5309);
nor U6527 (N_6527,N_5614,N_5980);
xnor U6528 (N_6528,N_5210,N_5112);
and U6529 (N_6529,N_5043,N_5087);
and U6530 (N_6530,N_5897,N_5828);
or U6531 (N_6531,N_5470,N_5765);
xnor U6532 (N_6532,N_5263,N_5113);
or U6533 (N_6533,N_5553,N_5637);
or U6534 (N_6534,N_5025,N_5194);
and U6535 (N_6535,N_5925,N_5651);
nand U6536 (N_6536,N_5492,N_5437);
nand U6537 (N_6537,N_5520,N_5005);
nand U6538 (N_6538,N_5879,N_5954);
or U6539 (N_6539,N_5493,N_5655);
or U6540 (N_6540,N_5619,N_5485);
nand U6541 (N_6541,N_5016,N_5027);
nand U6542 (N_6542,N_5330,N_5730);
and U6543 (N_6543,N_5293,N_5096);
nor U6544 (N_6544,N_5832,N_5326);
nor U6545 (N_6545,N_5645,N_5499);
or U6546 (N_6546,N_5125,N_5134);
nand U6547 (N_6547,N_5623,N_5303);
nand U6548 (N_6548,N_5379,N_5500);
nor U6549 (N_6549,N_5277,N_5134);
and U6550 (N_6550,N_5590,N_5856);
nand U6551 (N_6551,N_5036,N_5688);
or U6552 (N_6552,N_5837,N_5398);
nor U6553 (N_6553,N_5489,N_5433);
and U6554 (N_6554,N_5969,N_5795);
nor U6555 (N_6555,N_5742,N_5637);
nand U6556 (N_6556,N_5572,N_5757);
nor U6557 (N_6557,N_5915,N_5606);
and U6558 (N_6558,N_5070,N_5204);
and U6559 (N_6559,N_5008,N_5582);
or U6560 (N_6560,N_5932,N_5607);
and U6561 (N_6561,N_5625,N_5800);
nand U6562 (N_6562,N_5459,N_5341);
or U6563 (N_6563,N_5926,N_5504);
nor U6564 (N_6564,N_5771,N_5165);
and U6565 (N_6565,N_5250,N_5076);
or U6566 (N_6566,N_5727,N_5601);
or U6567 (N_6567,N_5814,N_5511);
nor U6568 (N_6568,N_5301,N_5937);
or U6569 (N_6569,N_5157,N_5016);
nand U6570 (N_6570,N_5906,N_5748);
or U6571 (N_6571,N_5654,N_5605);
or U6572 (N_6572,N_5454,N_5468);
and U6573 (N_6573,N_5226,N_5646);
or U6574 (N_6574,N_5643,N_5351);
nor U6575 (N_6575,N_5452,N_5845);
and U6576 (N_6576,N_5968,N_5673);
or U6577 (N_6577,N_5222,N_5753);
and U6578 (N_6578,N_5232,N_5660);
xnor U6579 (N_6579,N_5499,N_5897);
xor U6580 (N_6580,N_5696,N_5907);
or U6581 (N_6581,N_5744,N_5117);
or U6582 (N_6582,N_5021,N_5350);
nor U6583 (N_6583,N_5042,N_5180);
nor U6584 (N_6584,N_5073,N_5579);
nand U6585 (N_6585,N_5909,N_5444);
nand U6586 (N_6586,N_5059,N_5611);
or U6587 (N_6587,N_5169,N_5813);
xnor U6588 (N_6588,N_5206,N_5408);
or U6589 (N_6589,N_5219,N_5036);
or U6590 (N_6590,N_5171,N_5868);
and U6591 (N_6591,N_5031,N_5191);
or U6592 (N_6592,N_5290,N_5169);
or U6593 (N_6593,N_5994,N_5696);
xor U6594 (N_6594,N_5433,N_5299);
or U6595 (N_6595,N_5357,N_5570);
nand U6596 (N_6596,N_5675,N_5710);
nor U6597 (N_6597,N_5591,N_5802);
nand U6598 (N_6598,N_5433,N_5189);
nor U6599 (N_6599,N_5221,N_5923);
xnor U6600 (N_6600,N_5815,N_5008);
nand U6601 (N_6601,N_5074,N_5863);
nand U6602 (N_6602,N_5051,N_5869);
nor U6603 (N_6603,N_5632,N_5291);
nand U6604 (N_6604,N_5132,N_5062);
and U6605 (N_6605,N_5929,N_5223);
nor U6606 (N_6606,N_5033,N_5125);
and U6607 (N_6607,N_5471,N_5324);
and U6608 (N_6608,N_5850,N_5660);
or U6609 (N_6609,N_5910,N_5206);
xor U6610 (N_6610,N_5256,N_5084);
nor U6611 (N_6611,N_5791,N_5555);
nand U6612 (N_6612,N_5065,N_5399);
or U6613 (N_6613,N_5766,N_5439);
or U6614 (N_6614,N_5514,N_5134);
or U6615 (N_6615,N_5052,N_5182);
nor U6616 (N_6616,N_5804,N_5426);
and U6617 (N_6617,N_5161,N_5639);
xor U6618 (N_6618,N_5299,N_5383);
nor U6619 (N_6619,N_5910,N_5853);
nand U6620 (N_6620,N_5716,N_5013);
nor U6621 (N_6621,N_5725,N_5874);
and U6622 (N_6622,N_5303,N_5647);
and U6623 (N_6623,N_5283,N_5724);
and U6624 (N_6624,N_5425,N_5101);
and U6625 (N_6625,N_5999,N_5121);
or U6626 (N_6626,N_5840,N_5168);
or U6627 (N_6627,N_5511,N_5338);
and U6628 (N_6628,N_5058,N_5185);
or U6629 (N_6629,N_5693,N_5597);
nand U6630 (N_6630,N_5837,N_5083);
nand U6631 (N_6631,N_5801,N_5083);
nand U6632 (N_6632,N_5413,N_5056);
nand U6633 (N_6633,N_5189,N_5158);
xor U6634 (N_6634,N_5476,N_5557);
nor U6635 (N_6635,N_5219,N_5279);
or U6636 (N_6636,N_5994,N_5658);
nor U6637 (N_6637,N_5157,N_5453);
nand U6638 (N_6638,N_5278,N_5336);
or U6639 (N_6639,N_5207,N_5595);
nor U6640 (N_6640,N_5100,N_5596);
nand U6641 (N_6641,N_5060,N_5416);
and U6642 (N_6642,N_5430,N_5355);
and U6643 (N_6643,N_5685,N_5045);
nor U6644 (N_6644,N_5453,N_5095);
nor U6645 (N_6645,N_5172,N_5355);
or U6646 (N_6646,N_5386,N_5315);
nand U6647 (N_6647,N_5422,N_5665);
or U6648 (N_6648,N_5285,N_5647);
nand U6649 (N_6649,N_5164,N_5671);
xor U6650 (N_6650,N_5916,N_5360);
nor U6651 (N_6651,N_5500,N_5508);
or U6652 (N_6652,N_5331,N_5441);
and U6653 (N_6653,N_5409,N_5977);
nor U6654 (N_6654,N_5484,N_5627);
and U6655 (N_6655,N_5747,N_5231);
and U6656 (N_6656,N_5369,N_5959);
or U6657 (N_6657,N_5689,N_5930);
or U6658 (N_6658,N_5125,N_5313);
or U6659 (N_6659,N_5778,N_5744);
nor U6660 (N_6660,N_5645,N_5042);
nand U6661 (N_6661,N_5293,N_5655);
or U6662 (N_6662,N_5477,N_5707);
nor U6663 (N_6663,N_5371,N_5000);
nand U6664 (N_6664,N_5551,N_5742);
xnor U6665 (N_6665,N_5631,N_5141);
and U6666 (N_6666,N_5829,N_5084);
or U6667 (N_6667,N_5702,N_5593);
or U6668 (N_6668,N_5562,N_5524);
nand U6669 (N_6669,N_5112,N_5786);
nor U6670 (N_6670,N_5477,N_5317);
or U6671 (N_6671,N_5852,N_5448);
or U6672 (N_6672,N_5115,N_5787);
nor U6673 (N_6673,N_5829,N_5187);
nand U6674 (N_6674,N_5820,N_5075);
nor U6675 (N_6675,N_5557,N_5290);
nand U6676 (N_6676,N_5316,N_5397);
xor U6677 (N_6677,N_5720,N_5075);
nand U6678 (N_6678,N_5536,N_5829);
and U6679 (N_6679,N_5306,N_5831);
nand U6680 (N_6680,N_5140,N_5179);
or U6681 (N_6681,N_5741,N_5775);
and U6682 (N_6682,N_5027,N_5662);
nand U6683 (N_6683,N_5443,N_5944);
and U6684 (N_6684,N_5935,N_5650);
or U6685 (N_6685,N_5314,N_5310);
nor U6686 (N_6686,N_5981,N_5508);
and U6687 (N_6687,N_5243,N_5065);
or U6688 (N_6688,N_5042,N_5713);
and U6689 (N_6689,N_5410,N_5690);
nand U6690 (N_6690,N_5014,N_5356);
nor U6691 (N_6691,N_5974,N_5272);
xnor U6692 (N_6692,N_5908,N_5787);
xnor U6693 (N_6693,N_5830,N_5484);
or U6694 (N_6694,N_5946,N_5548);
or U6695 (N_6695,N_5897,N_5669);
nand U6696 (N_6696,N_5181,N_5764);
or U6697 (N_6697,N_5832,N_5192);
nand U6698 (N_6698,N_5839,N_5467);
or U6699 (N_6699,N_5103,N_5372);
xnor U6700 (N_6700,N_5736,N_5064);
or U6701 (N_6701,N_5605,N_5885);
nor U6702 (N_6702,N_5353,N_5503);
nand U6703 (N_6703,N_5463,N_5823);
nand U6704 (N_6704,N_5204,N_5599);
xnor U6705 (N_6705,N_5561,N_5646);
nor U6706 (N_6706,N_5822,N_5130);
or U6707 (N_6707,N_5513,N_5459);
and U6708 (N_6708,N_5704,N_5449);
or U6709 (N_6709,N_5396,N_5074);
and U6710 (N_6710,N_5918,N_5014);
nand U6711 (N_6711,N_5455,N_5477);
and U6712 (N_6712,N_5922,N_5438);
nor U6713 (N_6713,N_5951,N_5511);
and U6714 (N_6714,N_5832,N_5743);
nor U6715 (N_6715,N_5974,N_5019);
and U6716 (N_6716,N_5160,N_5465);
nand U6717 (N_6717,N_5954,N_5044);
xnor U6718 (N_6718,N_5313,N_5923);
nor U6719 (N_6719,N_5997,N_5821);
nor U6720 (N_6720,N_5090,N_5356);
or U6721 (N_6721,N_5085,N_5347);
nand U6722 (N_6722,N_5902,N_5022);
nand U6723 (N_6723,N_5548,N_5146);
and U6724 (N_6724,N_5114,N_5250);
nor U6725 (N_6725,N_5370,N_5710);
nor U6726 (N_6726,N_5366,N_5734);
nand U6727 (N_6727,N_5603,N_5848);
and U6728 (N_6728,N_5367,N_5747);
nand U6729 (N_6729,N_5074,N_5760);
and U6730 (N_6730,N_5876,N_5014);
nand U6731 (N_6731,N_5900,N_5377);
and U6732 (N_6732,N_5800,N_5531);
xor U6733 (N_6733,N_5533,N_5051);
nor U6734 (N_6734,N_5397,N_5698);
nor U6735 (N_6735,N_5204,N_5263);
nand U6736 (N_6736,N_5136,N_5684);
nand U6737 (N_6737,N_5247,N_5942);
nor U6738 (N_6738,N_5594,N_5011);
and U6739 (N_6739,N_5632,N_5085);
nand U6740 (N_6740,N_5494,N_5856);
nand U6741 (N_6741,N_5907,N_5463);
and U6742 (N_6742,N_5928,N_5915);
nor U6743 (N_6743,N_5646,N_5218);
xnor U6744 (N_6744,N_5861,N_5620);
and U6745 (N_6745,N_5644,N_5601);
or U6746 (N_6746,N_5030,N_5436);
nand U6747 (N_6747,N_5325,N_5224);
and U6748 (N_6748,N_5381,N_5015);
and U6749 (N_6749,N_5921,N_5550);
or U6750 (N_6750,N_5156,N_5561);
nor U6751 (N_6751,N_5711,N_5917);
nand U6752 (N_6752,N_5331,N_5330);
or U6753 (N_6753,N_5166,N_5463);
xor U6754 (N_6754,N_5325,N_5971);
nand U6755 (N_6755,N_5797,N_5652);
or U6756 (N_6756,N_5325,N_5206);
nor U6757 (N_6757,N_5013,N_5541);
nor U6758 (N_6758,N_5256,N_5692);
nor U6759 (N_6759,N_5222,N_5546);
nor U6760 (N_6760,N_5948,N_5955);
or U6761 (N_6761,N_5452,N_5076);
and U6762 (N_6762,N_5032,N_5810);
or U6763 (N_6763,N_5415,N_5479);
nor U6764 (N_6764,N_5111,N_5739);
and U6765 (N_6765,N_5433,N_5093);
nand U6766 (N_6766,N_5306,N_5531);
and U6767 (N_6767,N_5772,N_5727);
or U6768 (N_6768,N_5144,N_5384);
nand U6769 (N_6769,N_5506,N_5586);
or U6770 (N_6770,N_5211,N_5197);
nand U6771 (N_6771,N_5157,N_5622);
nand U6772 (N_6772,N_5820,N_5114);
nand U6773 (N_6773,N_5130,N_5697);
nor U6774 (N_6774,N_5027,N_5836);
nand U6775 (N_6775,N_5410,N_5102);
nand U6776 (N_6776,N_5074,N_5942);
xor U6777 (N_6777,N_5070,N_5901);
and U6778 (N_6778,N_5888,N_5061);
nand U6779 (N_6779,N_5604,N_5157);
nand U6780 (N_6780,N_5679,N_5343);
nor U6781 (N_6781,N_5185,N_5038);
xor U6782 (N_6782,N_5774,N_5152);
and U6783 (N_6783,N_5076,N_5486);
nand U6784 (N_6784,N_5755,N_5370);
and U6785 (N_6785,N_5381,N_5891);
or U6786 (N_6786,N_5781,N_5866);
and U6787 (N_6787,N_5658,N_5408);
xnor U6788 (N_6788,N_5967,N_5758);
and U6789 (N_6789,N_5477,N_5552);
or U6790 (N_6790,N_5046,N_5254);
nor U6791 (N_6791,N_5370,N_5564);
nand U6792 (N_6792,N_5254,N_5039);
and U6793 (N_6793,N_5602,N_5981);
nand U6794 (N_6794,N_5106,N_5145);
and U6795 (N_6795,N_5540,N_5914);
or U6796 (N_6796,N_5035,N_5943);
nand U6797 (N_6797,N_5088,N_5489);
nor U6798 (N_6798,N_5744,N_5016);
nand U6799 (N_6799,N_5482,N_5431);
nand U6800 (N_6800,N_5378,N_5692);
nand U6801 (N_6801,N_5729,N_5267);
xor U6802 (N_6802,N_5891,N_5909);
nand U6803 (N_6803,N_5076,N_5007);
nand U6804 (N_6804,N_5373,N_5782);
or U6805 (N_6805,N_5020,N_5390);
nand U6806 (N_6806,N_5825,N_5646);
and U6807 (N_6807,N_5615,N_5618);
nor U6808 (N_6808,N_5788,N_5169);
or U6809 (N_6809,N_5434,N_5184);
and U6810 (N_6810,N_5073,N_5377);
nand U6811 (N_6811,N_5689,N_5404);
or U6812 (N_6812,N_5808,N_5852);
nand U6813 (N_6813,N_5524,N_5092);
nand U6814 (N_6814,N_5594,N_5825);
and U6815 (N_6815,N_5949,N_5772);
nand U6816 (N_6816,N_5629,N_5031);
nor U6817 (N_6817,N_5825,N_5470);
nand U6818 (N_6818,N_5309,N_5019);
nand U6819 (N_6819,N_5888,N_5173);
xor U6820 (N_6820,N_5345,N_5193);
nand U6821 (N_6821,N_5463,N_5559);
nand U6822 (N_6822,N_5106,N_5672);
xor U6823 (N_6823,N_5986,N_5067);
nor U6824 (N_6824,N_5723,N_5601);
nor U6825 (N_6825,N_5573,N_5945);
and U6826 (N_6826,N_5597,N_5205);
or U6827 (N_6827,N_5111,N_5094);
nand U6828 (N_6828,N_5788,N_5174);
xor U6829 (N_6829,N_5596,N_5939);
xor U6830 (N_6830,N_5221,N_5926);
nor U6831 (N_6831,N_5431,N_5483);
or U6832 (N_6832,N_5020,N_5383);
and U6833 (N_6833,N_5525,N_5756);
or U6834 (N_6834,N_5835,N_5396);
nor U6835 (N_6835,N_5187,N_5675);
xnor U6836 (N_6836,N_5882,N_5840);
and U6837 (N_6837,N_5397,N_5621);
nand U6838 (N_6838,N_5622,N_5765);
xor U6839 (N_6839,N_5482,N_5864);
or U6840 (N_6840,N_5950,N_5071);
or U6841 (N_6841,N_5203,N_5514);
nor U6842 (N_6842,N_5442,N_5661);
nand U6843 (N_6843,N_5706,N_5103);
nor U6844 (N_6844,N_5241,N_5420);
nand U6845 (N_6845,N_5661,N_5667);
nor U6846 (N_6846,N_5985,N_5490);
or U6847 (N_6847,N_5214,N_5699);
and U6848 (N_6848,N_5771,N_5500);
nor U6849 (N_6849,N_5426,N_5762);
nor U6850 (N_6850,N_5893,N_5599);
nand U6851 (N_6851,N_5696,N_5338);
and U6852 (N_6852,N_5280,N_5097);
or U6853 (N_6853,N_5340,N_5487);
nor U6854 (N_6854,N_5295,N_5572);
nor U6855 (N_6855,N_5242,N_5786);
nand U6856 (N_6856,N_5374,N_5825);
xnor U6857 (N_6857,N_5517,N_5919);
and U6858 (N_6858,N_5859,N_5643);
xor U6859 (N_6859,N_5579,N_5209);
or U6860 (N_6860,N_5639,N_5841);
nor U6861 (N_6861,N_5981,N_5570);
or U6862 (N_6862,N_5297,N_5342);
and U6863 (N_6863,N_5411,N_5374);
nor U6864 (N_6864,N_5819,N_5788);
and U6865 (N_6865,N_5915,N_5175);
and U6866 (N_6866,N_5342,N_5183);
or U6867 (N_6867,N_5377,N_5193);
and U6868 (N_6868,N_5920,N_5571);
xnor U6869 (N_6869,N_5917,N_5964);
and U6870 (N_6870,N_5991,N_5385);
or U6871 (N_6871,N_5206,N_5890);
nand U6872 (N_6872,N_5568,N_5637);
nand U6873 (N_6873,N_5372,N_5853);
and U6874 (N_6874,N_5819,N_5589);
and U6875 (N_6875,N_5728,N_5215);
xnor U6876 (N_6876,N_5754,N_5714);
nand U6877 (N_6877,N_5960,N_5733);
xor U6878 (N_6878,N_5301,N_5041);
and U6879 (N_6879,N_5966,N_5432);
or U6880 (N_6880,N_5728,N_5823);
or U6881 (N_6881,N_5519,N_5091);
and U6882 (N_6882,N_5017,N_5717);
nand U6883 (N_6883,N_5269,N_5685);
and U6884 (N_6884,N_5624,N_5071);
nor U6885 (N_6885,N_5620,N_5651);
nor U6886 (N_6886,N_5354,N_5202);
nor U6887 (N_6887,N_5111,N_5710);
and U6888 (N_6888,N_5003,N_5940);
and U6889 (N_6889,N_5886,N_5687);
xnor U6890 (N_6890,N_5406,N_5337);
and U6891 (N_6891,N_5559,N_5163);
and U6892 (N_6892,N_5594,N_5202);
or U6893 (N_6893,N_5341,N_5601);
and U6894 (N_6894,N_5109,N_5785);
or U6895 (N_6895,N_5487,N_5767);
nand U6896 (N_6896,N_5028,N_5763);
nor U6897 (N_6897,N_5277,N_5358);
nand U6898 (N_6898,N_5126,N_5653);
nor U6899 (N_6899,N_5367,N_5611);
nor U6900 (N_6900,N_5780,N_5718);
or U6901 (N_6901,N_5208,N_5279);
and U6902 (N_6902,N_5701,N_5916);
or U6903 (N_6903,N_5789,N_5403);
nand U6904 (N_6904,N_5601,N_5745);
nand U6905 (N_6905,N_5215,N_5279);
or U6906 (N_6906,N_5028,N_5450);
nor U6907 (N_6907,N_5165,N_5913);
nor U6908 (N_6908,N_5598,N_5350);
nor U6909 (N_6909,N_5427,N_5196);
nand U6910 (N_6910,N_5935,N_5531);
or U6911 (N_6911,N_5494,N_5705);
and U6912 (N_6912,N_5583,N_5918);
and U6913 (N_6913,N_5598,N_5919);
nand U6914 (N_6914,N_5818,N_5598);
or U6915 (N_6915,N_5431,N_5950);
or U6916 (N_6916,N_5415,N_5371);
nand U6917 (N_6917,N_5248,N_5927);
xnor U6918 (N_6918,N_5918,N_5685);
and U6919 (N_6919,N_5001,N_5856);
nor U6920 (N_6920,N_5252,N_5418);
or U6921 (N_6921,N_5468,N_5819);
xnor U6922 (N_6922,N_5169,N_5040);
nor U6923 (N_6923,N_5463,N_5266);
or U6924 (N_6924,N_5274,N_5654);
nor U6925 (N_6925,N_5573,N_5008);
and U6926 (N_6926,N_5116,N_5625);
nor U6927 (N_6927,N_5431,N_5963);
and U6928 (N_6928,N_5944,N_5145);
or U6929 (N_6929,N_5250,N_5935);
and U6930 (N_6930,N_5385,N_5078);
and U6931 (N_6931,N_5915,N_5553);
nand U6932 (N_6932,N_5399,N_5387);
xor U6933 (N_6933,N_5009,N_5595);
and U6934 (N_6934,N_5198,N_5544);
nand U6935 (N_6935,N_5764,N_5188);
nor U6936 (N_6936,N_5368,N_5097);
or U6937 (N_6937,N_5489,N_5107);
xor U6938 (N_6938,N_5992,N_5286);
xor U6939 (N_6939,N_5461,N_5806);
nor U6940 (N_6940,N_5907,N_5025);
nor U6941 (N_6941,N_5460,N_5269);
or U6942 (N_6942,N_5337,N_5975);
or U6943 (N_6943,N_5114,N_5733);
and U6944 (N_6944,N_5643,N_5068);
xnor U6945 (N_6945,N_5560,N_5799);
or U6946 (N_6946,N_5908,N_5676);
nand U6947 (N_6947,N_5085,N_5712);
or U6948 (N_6948,N_5077,N_5005);
nor U6949 (N_6949,N_5343,N_5175);
nor U6950 (N_6950,N_5910,N_5605);
nand U6951 (N_6951,N_5088,N_5310);
nor U6952 (N_6952,N_5038,N_5996);
or U6953 (N_6953,N_5337,N_5395);
nand U6954 (N_6954,N_5533,N_5682);
and U6955 (N_6955,N_5994,N_5977);
nor U6956 (N_6956,N_5434,N_5203);
and U6957 (N_6957,N_5436,N_5415);
and U6958 (N_6958,N_5642,N_5438);
nor U6959 (N_6959,N_5800,N_5115);
or U6960 (N_6960,N_5252,N_5557);
nand U6961 (N_6961,N_5568,N_5935);
nor U6962 (N_6962,N_5365,N_5109);
nand U6963 (N_6963,N_5091,N_5543);
and U6964 (N_6964,N_5029,N_5945);
and U6965 (N_6965,N_5246,N_5015);
nor U6966 (N_6966,N_5371,N_5813);
nor U6967 (N_6967,N_5496,N_5841);
or U6968 (N_6968,N_5616,N_5942);
or U6969 (N_6969,N_5978,N_5054);
nand U6970 (N_6970,N_5442,N_5428);
nor U6971 (N_6971,N_5707,N_5457);
xor U6972 (N_6972,N_5093,N_5162);
or U6973 (N_6973,N_5139,N_5460);
nor U6974 (N_6974,N_5634,N_5302);
nand U6975 (N_6975,N_5111,N_5340);
and U6976 (N_6976,N_5241,N_5541);
or U6977 (N_6977,N_5008,N_5343);
and U6978 (N_6978,N_5166,N_5314);
xor U6979 (N_6979,N_5415,N_5585);
or U6980 (N_6980,N_5564,N_5771);
nor U6981 (N_6981,N_5331,N_5724);
or U6982 (N_6982,N_5325,N_5958);
nor U6983 (N_6983,N_5216,N_5594);
nand U6984 (N_6984,N_5284,N_5573);
nand U6985 (N_6985,N_5739,N_5026);
xor U6986 (N_6986,N_5036,N_5404);
nand U6987 (N_6987,N_5284,N_5382);
xnor U6988 (N_6988,N_5600,N_5717);
nand U6989 (N_6989,N_5047,N_5330);
and U6990 (N_6990,N_5980,N_5369);
nand U6991 (N_6991,N_5167,N_5372);
or U6992 (N_6992,N_5709,N_5592);
and U6993 (N_6993,N_5184,N_5402);
nand U6994 (N_6994,N_5186,N_5191);
or U6995 (N_6995,N_5456,N_5921);
xor U6996 (N_6996,N_5097,N_5475);
or U6997 (N_6997,N_5649,N_5321);
and U6998 (N_6998,N_5415,N_5472);
nand U6999 (N_6999,N_5145,N_5344);
nor U7000 (N_7000,N_6747,N_6491);
nor U7001 (N_7001,N_6307,N_6639);
or U7002 (N_7002,N_6276,N_6489);
and U7003 (N_7003,N_6928,N_6001);
xnor U7004 (N_7004,N_6107,N_6341);
nor U7005 (N_7005,N_6227,N_6630);
nand U7006 (N_7006,N_6859,N_6025);
or U7007 (N_7007,N_6569,N_6159);
nand U7008 (N_7008,N_6999,N_6775);
nor U7009 (N_7009,N_6452,N_6918);
nor U7010 (N_7010,N_6469,N_6779);
or U7011 (N_7011,N_6059,N_6576);
nand U7012 (N_7012,N_6397,N_6670);
and U7013 (N_7013,N_6182,N_6427);
and U7014 (N_7014,N_6231,N_6363);
xnor U7015 (N_7015,N_6915,N_6819);
nor U7016 (N_7016,N_6888,N_6386);
nand U7017 (N_7017,N_6834,N_6590);
and U7018 (N_7018,N_6479,N_6215);
nand U7019 (N_7019,N_6753,N_6607);
or U7020 (N_7020,N_6718,N_6869);
nor U7021 (N_7021,N_6253,N_6330);
nor U7022 (N_7022,N_6632,N_6580);
nor U7023 (N_7023,N_6306,N_6143);
and U7024 (N_7024,N_6631,N_6514);
or U7025 (N_7025,N_6780,N_6765);
and U7026 (N_7026,N_6290,N_6114);
nor U7027 (N_7027,N_6179,N_6511);
or U7028 (N_7028,N_6816,N_6743);
or U7029 (N_7029,N_6536,N_6190);
nor U7030 (N_7030,N_6558,N_6681);
nor U7031 (N_7031,N_6833,N_6594);
and U7032 (N_7032,N_6380,N_6548);
nor U7033 (N_7033,N_6012,N_6252);
nor U7034 (N_7034,N_6907,N_6428);
and U7035 (N_7035,N_6930,N_6887);
and U7036 (N_7036,N_6156,N_6298);
or U7037 (N_7037,N_6521,N_6959);
or U7038 (N_7038,N_6537,N_6690);
xor U7039 (N_7039,N_6510,N_6993);
nor U7040 (N_7040,N_6618,N_6198);
or U7041 (N_7041,N_6901,N_6409);
nor U7042 (N_7042,N_6531,N_6850);
or U7043 (N_7043,N_6754,N_6002);
and U7044 (N_7044,N_6599,N_6097);
and U7045 (N_7045,N_6167,N_6440);
nor U7046 (N_7046,N_6328,N_6103);
and U7047 (N_7047,N_6449,N_6144);
and U7048 (N_7048,N_6369,N_6324);
nand U7049 (N_7049,N_6540,N_6291);
nor U7050 (N_7050,N_6476,N_6702);
nor U7051 (N_7051,N_6318,N_6154);
or U7052 (N_7052,N_6044,N_6446);
nor U7053 (N_7053,N_6111,N_6422);
nor U7054 (N_7054,N_6908,N_6662);
and U7055 (N_7055,N_6211,N_6858);
and U7056 (N_7056,N_6501,N_6798);
nor U7057 (N_7057,N_6278,N_6948);
and U7058 (N_7058,N_6042,N_6867);
nor U7059 (N_7059,N_6795,N_6561);
nor U7060 (N_7060,N_6498,N_6832);
nand U7061 (N_7061,N_6596,N_6021);
nor U7062 (N_7062,N_6756,N_6193);
nand U7063 (N_7063,N_6367,N_6106);
nor U7064 (N_7064,N_6050,N_6934);
xor U7065 (N_7065,N_6016,N_6168);
nand U7066 (N_7066,N_6040,N_6643);
xnor U7067 (N_7067,N_6235,N_6383);
or U7068 (N_7068,N_6192,N_6708);
and U7069 (N_7069,N_6712,N_6588);
and U7070 (N_7070,N_6882,N_6396);
nor U7071 (N_7071,N_6509,N_6185);
or U7072 (N_7072,N_6433,N_6308);
or U7073 (N_7073,N_6410,N_6861);
and U7074 (N_7074,N_6385,N_6462);
xor U7075 (N_7075,N_6529,N_6188);
nor U7076 (N_7076,N_6853,N_6085);
nand U7077 (N_7077,N_6007,N_6246);
xnor U7078 (N_7078,N_6605,N_6089);
nand U7079 (N_7079,N_6372,N_6474);
xnor U7080 (N_7080,N_6401,N_6657);
nand U7081 (N_7081,N_6723,N_6357);
and U7082 (N_7082,N_6968,N_6541);
and U7083 (N_7083,N_6266,N_6609);
nor U7084 (N_7084,N_6953,N_6319);
nor U7085 (N_7085,N_6137,N_6333);
or U7086 (N_7086,N_6829,N_6448);
or U7087 (N_7087,N_6186,N_6418);
and U7088 (N_7088,N_6988,N_6384);
nand U7089 (N_7089,N_6742,N_6438);
nand U7090 (N_7090,N_6560,N_6998);
or U7091 (N_7091,N_6792,N_6623);
nand U7092 (N_7092,N_6148,N_6904);
and U7093 (N_7093,N_6563,N_6480);
and U7094 (N_7094,N_6698,N_6459);
and U7095 (N_7095,N_6081,N_6502);
and U7096 (N_7096,N_6967,N_6553);
and U7097 (N_7097,N_6975,N_6054);
and U7098 (N_7098,N_6844,N_6098);
nor U7099 (N_7099,N_6647,N_6169);
nor U7100 (N_7100,N_6600,N_6077);
or U7101 (N_7101,N_6304,N_6910);
or U7102 (N_7102,N_6807,N_6732);
or U7103 (N_7103,N_6682,N_6450);
nand U7104 (N_7104,N_6269,N_6736);
xor U7105 (N_7105,N_6245,N_6105);
nand U7106 (N_7106,N_6676,N_6404);
and U7107 (N_7107,N_6272,N_6950);
nor U7108 (N_7108,N_6302,N_6472);
xnor U7109 (N_7109,N_6031,N_6104);
nor U7110 (N_7110,N_6991,N_6320);
or U7111 (N_7111,N_6322,N_6769);
or U7112 (N_7112,N_6897,N_6287);
and U7113 (N_7113,N_6666,N_6359);
or U7114 (N_7114,N_6203,N_6321);
or U7115 (N_7115,N_6108,N_6225);
or U7116 (N_7116,N_6247,N_6109);
nor U7117 (N_7117,N_6067,N_6880);
and U7118 (N_7118,N_6947,N_6872);
nor U7119 (N_7119,N_6575,N_6274);
and U7120 (N_7120,N_6585,N_6513);
nand U7121 (N_7121,N_6977,N_6425);
or U7122 (N_7122,N_6160,N_6564);
and U7123 (N_7123,N_6808,N_6899);
nor U7124 (N_7124,N_6492,N_6379);
or U7125 (N_7125,N_6648,N_6006);
nand U7126 (N_7126,N_6499,N_6815);
nor U7127 (N_7127,N_6823,N_6431);
nor U7128 (N_7128,N_6522,N_6751);
and U7129 (N_7129,N_6113,N_6554);
nand U7130 (N_7130,N_6229,N_6207);
nor U7131 (N_7131,N_6292,N_6763);
nor U7132 (N_7132,N_6752,N_6789);
nor U7133 (N_7133,N_6738,N_6473);
and U7134 (N_7134,N_6348,N_6084);
nor U7135 (N_7135,N_6778,N_6705);
nand U7136 (N_7136,N_6351,N_6400);
or U7137 (N_7137,N_6912,N_6932);
nor U7138 (N_7138,N_6584,N_6494);
nor U7139 (N_7139,N_6342,N_6072);
nor U7140 (N_7140,N_6875,N_6679);
or U7141 (N_7141,N_6000,N_6056);
xnor U7142 (N_7142,N_6771,N_6281);
nor U7143 (N_7143,N_6957,N_6528);
nor U7144 (N_7144,N_6123,N_6255);
nand U7145 (N_7145,N_6195,N_6260);
or U7146 (N_7146,N_6525,N_6399);
or U7147 (N_7147,N_6885,N_6060);
xnor U7148 (N_7148,N_6956,N_6865);
nor U7149 (N_7149,N_6080,N_6533);
nor U7150 (N_7150,N_6301,N_6187);
nand U7151 (N_7151,N_6430,N_6376);
nand U7152 (N_7152,N_6254,N_6543);
nand U7153 (N_7153,N_6100,N_6724);
nor U7154 (N_7154,N_6295,N_6750);
nor U7155 (N_7155,N_6735,N_6746);
nand U7156 (N_7156,N_6699,N_6674);
xnor U7157 (N_7157,N_6809,N_6094);
or U7158 (N_7158,N_6261,N_6545);
nand U7159 (N_7159,N_6730,N_6866);
or U7160 (N_7160,N_6256,N_6625);
or U7161 (N_7161,N_6960,N_6652);
or U7162 (N_7162,N_6530,N_6366);
nand U7163 (N_7163,N_6748,N_6610);
or U7164 (N_7164,N_6691,N_6797);
nor U7165 (N_7165,N_6764,N_6390);
nor U7166 (N_7166,N_6370,N_6936);
xnor U7167 (N_7167,N_6248,N_6571);
nor U7168 (N_7168,N_6183,N_6411);
and U7169 (N_7169,N_6398,N_6675);
xnor U7170 (N_7170,N_6938,N_6920);
nor U7171 (N_7171,N_6707,N_6194);
or U7172 (N_7172,N_6943,N_6635);
or U7173 (N_7173,N_6737,N_6202);
nand U7174 (N_7174,N_6275,N_6009);
and U7175 (N_7175,N_6228,N_6079);
xor U7176 (N_7176,N_6672,N_6568);
nor U7177 (N_7177,N_6268,N_6622);
nor U7178 (N_7178,N_6878,N_6534);
nand U7179 (N_7179,N_6589,N_6236);
and U7180 (N_7180,N_6488,N_6884);
nand U7181 (N_7181,N_6152,N_6919);
nand U7182 (N_7182,N_6461,N_6812);
xnor U7183 (N_7183,N_6762,N_6843);
xor U7184 (N_7184,N_6835,N_6958);
or U7185 (N_7185,N_6346,N_6034);
nand U7186 (N_7186,N_6983,N_6606);
and U7187 (N_7187,N_6353,N_6023);
and U7188 (N_7188,N_6005,N_6371);
or U7189 (N_7189,N_6744,N_6969);
nand U7190 (N_7190,N_6896,N_6971);
or U7191 (N_7191,N_6995,N_6329);
xor U7192 (N_7192,N_6118,N_6165);
nand U7193 (N_7193,N_6313,N_6454);
or U7194 (N_7194,N_6112,N_6134);
xor U7195 (N_7195,N_6490,N_6004);
nand U7196 (N_7196,N_6593,N_6601);
xor U7197 (N_7197,N_6556,N_6683);
xnor U7198 (N_7198,N_6781,N_6810);
or U7199 (N_7199,N_6890,N_6616);
nor U7200 (N_7200,N_6264,N_6458);
xnor U7201 (N_7201,N_6519,N_6020);
nand U7202 (N_7202,N_6503,N_6693);
nor U7203 (N_7203,N_6538,N_6138);
or U7204 (N_7204,N_6049,N_6455);
nand U7205 (N_7205,N_6980,N_6344);
nor U7206 (N_7206,N_6760,N_6848);
and U7207 (N_7207,N_6602,N_6877);
nand U7208 (N_7208,N_6745,N_6030);
nor U7209 (N_7209,N_6382,N_6061);
nor U7210 (N_7210,N_6913,N_6240);
or U7211 (N_7211,N_6035,N_6841);
and U7212 (N_7212,N_6713,N_6994);
or U7213 (N_7213,N_6239,N_6767);
or U7214 (N_7214,N_6046,N_6559);
nor U7215 (N_7215,N_6706,N_6787);
nand U7216 (N_7216,N_6740,N_6273);
nand U7217 (N_7217,N_6925,N_6209);
or U7218 (N_7218,N_6770,N_6963);
or U7219 (N_7219,N_6258,N_6587);
or U7220 (N_7220,N_6064,N_6136);
nor U7221 (N_7221,N_6505,N_6336);
nor U7222 (N_7222,N_6687,N_6378);
or U7223 (N_7223,N_6902,N_6206);
and U7224 (N_7224,N_6684,N_6347);
and U7225 (N_7225,N_6870,N_6626);
or U7226 (N_7226,N_6524,N_6331);
nor U7227 (N_7227,N_6377,N_6813);
nand U7228 (N_7228,N_6364,N_6102);
and U7229 (N_7229,N_6128,N_6715);
xnor U7230 (N_7230,N_6220,N_6052);
nand U7231 (N_7231,N_6267,N_6442);
nor U7232 (N_7232,N_6900,N_6387);
and U7233 (N_7233,N_6555,N_6695);
and U7234 (N_7234,N_6677,N_6126);
or U7235 (N_7235,N_6921,N_6470);
or U7236 (N_7236,N_6285,N_6297);
nand U7237 (N_7237,N_6145,N_6613);
or U7238 (N_7238,N_6286,N_6181);
nand U7239 (N_7239,N_6226,N_6727);
and U7240 (N_7240,N_6218,N_6250);
xnor U7241 (N_7241,N_6817,N_6392);
nand U7242 (N_7242,N_6339,N_6170);
xnor U7243 (N_7243,N_6277,N_6360);
nand U7244 (N_7244,N_6842,N_6484);
nor U7245 (N_7245,N_6132,N_6766);
or U7246 (N_7246,N_6628,N_6774);
or U7247 (N_7247,N_6703,N_6173);
or U7248 (N_7248,N_6840,N_6660);
nand U7249 (N_7249,N_6851,N_6375);
and U7250 (N_7250,N_6697,N_6311);
nor U7251 (N_7251,N_6493,N_6496);
or U7252 (N_7252,N_6653,N_6008);
nor U7253 (N_7253,N_6638,N_6349);
or U7254 (N_7254,N_6180,N_6076);
or U7255 (N_7255,N_6233,N_6037);
and U7256 (N_7256,N_6784,N_6903);
nand U7257 (N_7257,N_6146,N_6916);
nand U7258 (N_7258,N_6946,N_6063);
xor U7259 (N_7259,N_6471,N_6191);
nand U7260 (N_7260,N_6133,N_6365);
and U7261 (N_7261,N_6673,N_6722);
nor U7262 (N_7262,N_6828,N_6634);
nand U7263 (N_7263,N_6550,N_6846);
nor U7264 (N_7264,N_6725,N_6728);
nand U7265 (N_7265,N_6806,N_6964);
xnor U7266 (N_7266,N_6654,N_6586);
nor U7267 (N_7267,N_6891,N_6871);
nor U7268 (N_7268,N_6694,N_6656);
or U7269 (N_7269,N_6700,N_6482);
and U7270 (N_7270,N_6283,N_6243);
or U7271 (N_7271,N_6820,N_6939);
and U7272 (N_7272,N_6954,N_6032);
or U7273 (N_7273,N_6139,N_6314);
or U7274 (N_7274,N_6873,N_6827);
nand U7275 (N_7275,N_6130,N_6047);
and U7276 (N_7276,N_6800,N_6895);
or U7277 (N_7277,N_6803,N_6926);
nor U7278 (N_7278,N_6949,N_6931);
or U7279 (N_7279,N_6014,N_6280);
and U7280 (N_7280,N_6270,N_6062);
or U7281 (N_7281,N_6583,N_6624);
or U7282 (N_7282,N_6345,N_6189);
xnor U7283 (N_7283,N_6312,N_6051);
xor U7284 (N_7284,N_6847,N_6640);
or U7285 (N_7285,N_6573,N_6979);
nor U7286 (N_7286,N_6069,N_6201);
nand U7287 (N_7287,N_6855,N_6577);
nand U7288 (N_7288,N_6874,N_6412);
or U7289 (N_7289,N_6726,N_6523);
or U7290 (N_7290,N_6238,N_6804);
nand U7291 (N_7291,N_6029,N_6826);
and U7292 (N_7292,N_6883,N_6512);
nand U7293 (N_7293,N_6124,N_6557);
nor U7294 (N_7294,N_6300,N_6417);
and U7295 (N_7295,N_6839,N_6017);
and U7296 (N_7296,N_6974,N_6845);
nand U7297 (N_7297,N_6068,N_6922);
nand U7298 (N_7298,N_6714,N_6213);
or U7299 (N_7299,N_6335,N_6175);
nor U7300 (N_7300,N_6027,N_6811);
nor U7301 (N_7301,N_6095,N_6777);
or U7302 (N_7302,N_6090,N_6038);
nor U7303 (N_7303,N_6337,N_6821);
nand U7304 (N_7304,N_6216,N_6093);
nand U7305 (N_7305,N_6592,N_6197);
xnor U7306 (N_7306,N_6944,N_6432);
or U7307 (N_7307,N_6793,N_6232);
or U7308 (N_7308,N_6177,N_6414);
nand U7309 (N_7309,N_6026,N_6096);
or U7310 (N_7310,N_6794,N_6039);
nor U7311 (N_7311,N_6429,N_6539);
xor U7312 (N_7312,N_6403,N_6444);
and U7313 (N_7313,N_6305,N_6658);
and U7314 (N_7314,N_6970,N_6955);
nor U7315 (N_7315,N_6951,N_6437);
nor U7316 (N_7316,N_6696,N_6504);
nor U7317 (N_7317,N_6508,N_6244);
and U7318 (N_7318,N_6172,N_6129);
nor U7319 (N_7319,N_6914,N_6552);
and U7320 (N_7320,N_6310,N_6234);
nor U7321 (N_7321,N_6487,N_6315);
nor U7322 (N_7322,N_6140,N_6117);
xor U7323 (N_7323,N_6099,N_6436);
and U7324 (N_7324,N_6636,N_6535);
or U7325 (N_7325,N_6898,N_6831);
nor U7326 (N_7326,N_6786,N_6485);
and U7327 (N_7327,N_6719,N_6518);
nand U7328 (N_7328,N_6729,N_6393);
nand U7329 (N_7329,N_6434,N_6710);
or U7330 (N_7330,N_6597,N_6174);
nor U7331 (N_7331,N_6987,N_6716);
nor U7332 (N_7332,N_6516,N_6468);
nor U7333 (N_7333,N_6120,N_6478);
nand U7334 (N_7334,N_6391,N_6671);
nor U7335 (N_7335,N_6619,N_6196);
and U7336 (N_7336,N_6617,N_6200);
nor U7337 (N_7337,N_6070,N_6155);
nand U7338 (N_7338,N_6688,N_6296);
nor U7339 (N_7339,N_6927,N_6435);
nand U7340 (N_7340,N_6802,N_6356);
and U7341 (N_7341,N_6720,N_6092);
nor U7342 (N_7342,N_6520,N_6158);
nand U7343 (N_7343,N_6121,N_6645);
nor U7344 (N_7344,N_6340,N_6066);
nand U7345 (N_7345,N_6241,N_6733);
nand U7346 (N_7346,N_6591,N_6612);
or U7347 (N_7347,N_6416,N_6326);
nand U7348 (N_7348,N_6598,N_6909);
and U7349 (N_7349,N_6783,N_6151);
nor U7350 (N_7350,N_6003,N_6028);
nand U7351 (N_7351,N_6426,N_6734);
nand U7352 (N_7352,N_6407,N_6776);
or U7353 (N_7353,N_6395,N_6966);
nor U7354 (N_7354,N_6611,N_6952);
and U7355 (N_7355,N_6731,N_6447);
xor U7356 (N_7356,N_6415,N_6667);
or U7357 (N_7357,N_6814,N_6082);
and U7358 (N_7358,N_6940,N_6796);
and U7359 (N_7359,N_6864,N_6976);
or U7360 (N_7360,N_6857,N_6973);
nand U7361 (N_7361,N_6057,N_6053);
xor U7362 (N_7362,N_6757,N_6036);
and U7363 (N_7363,N_6838,N_6608);
or U7364 (N_7364,N_6782,N_6544);
or U7365 (N_7365,N_6204,N_6354);
or U7366 (N_7366,N_6373,N_6701);
or U7367 (N_7367,N_6071,N_6149);
or U7368 (N_7368,N_6506,N_6650);
nor U7369 (N_7369,N_6486,N_6852);
nor U7370 (N_7370,N_6289,N_6222);
or U7371 (N_7371,N_6646,N_6578);
or U7372 (N_7372,N_6570,N_6581);
nor U7373 (N_7373,N_6551,N_6299);
or U7374 (N_7374,N_6157,N_6905);
nand U7375 (N_7375,N_6221,N_6879);
nor U7376 (N_7376,N_6282,N_6374);
nand U7377 (N_7377,N_6445,N_6889);
nor U7378 (N_7378,N_6574,N_6721);
nand U7379 (N_7379,N_6131,N_6352);
nand U7380 (N_7380,N_6279,N_6739);
or U7381 (N_7381,N_6924,N_6451);
nand U7382 (N_7382,N_6125,N_6637);
xnor U7383 (N_7383,N_6547,N_6214);
and U7384 (N_7384,N_6615,N_6515);
nand U7385 (N_7385,N_6649,N_6961);
and U7386 (N_7386,N_6361,N_6633);
nand U7387 (N_7387,N_6704,N_6122);
nand U7388 (N_7388,N_6223,N_6992);
or U7389 (N_7389,N_6937,N_6162);
and U7390 (N_7390,N_6074,N_6199);
nand U7391 (N_7391,N_6978,N_6565);
nand U7392 (N_7392,N_6692,N_6680);
nor U7393 (N_7393,N_6881,N_6772);
or U7394 (N_7394,N_6982,N_6171);
nor U7395 (N_7395,N_6265,N_6024);
nor U7396 (N_7396,N_6837,N_6466);
or U7397 (N_7397,N_6423,N_6166);
nor U7398 (N_7398,N_6685,N_6224);
or U7399 (N_7399,N_6424,N_6665);
xor U7400 (N_7400,N_6086,N_6309);
or U7401 (N_7401,N_6962,N_6262);
or U7402 (N_7402,N_6825,N_6711);
and U7403 (N_7403,N_6799,N_6621);
and U7404 (N_7404,N_6164,N_6284);
or U7405 (N_7405,N_6655,N_6065);
nand U7406 (N_7406,N_6388,N_6603);
and U7407 (N_7407,N_6303,N_6010);
nand U7408 (N_7408,N_6893,N_6500);
or U7409 (N_7409,N_6453,N_6562);
and U7410 (N_7410,N_6582,N_6989);
nor U7411 (N_7411,N_6087,N_6460);
nor U7412 (N_7412,N_6790,N_6542);
nor U7413 (N_7413,N_6986,N_6439);
and U7414 (N_7414,N_6237,N_6421);
nor U7415 (N_7415,N_6116,N_6150);
or U7416 (N_7416,N_6849,N_6294);
or U7417 (N_7417,N_6664,N_6022);
and U7418 (N_7418,N_6058,N_6788);
or U7419 (N_7419,N_6323,N_6184);
nor U7420 (N_7420,N_6251,N_6101);
or U7421 (N_7421,N_6886,N_6443);
nand U7422 (N_7422,N_6717,N_6856);
or U7423 (N_7423,N_6018,N_6317);
and U7424 (N_7424,N_6011,N_6801);
and U7425 (N_7425,N_6642,N_6205);
nand U7426 (N_7426,N_6507,N_6257);
nor U7427 (N_7427,N_6293,N_6091);
and U7428 (N_7428,N_6818,N_6567);
nor U7429 (N_7429,N_6997,N_6115);
or U7430 (N_7430,N_6495,N_6629);
and U7431 (N_7431,N_6259,N_6768);
nor U7432 (N_7432,N_6013,N_6045);
and U7433 (N_7433,N_6127,N_6678);
nand U7434 (N_7434,N_6135,N_6892);
nand U7435 (N_7435,N_6863,N_6791);
nand U7436 (N_7436,N_6475,N_6941);
and U7437 (N_7437,N_6394,N_6627);
nor U7438 (N_7438,N_6644,N_6981);
nor U7439 (N_7439,N_6595,N_6659);
nor U7440 (N_7440,N_6338,N_6942);
and U7441 (N_7441,N_6332,N_6327);
or U7442 (N_7442,N_6935,N_6517);
nor U7443 (N_7443,N_6406,N_6860);
nand U7444 (N_7444,N_6483,N_6441);
xnor U7445 (N_7445,N_6405,N_6210);
xor U7446 (N_7446,N_6078,N_6830);
nand U7447 (N_7447,N_6316,N_6355);
nand U7448 (N_7448,N_6457,N_6343);
or U7449 (N_7449,N_6463,N_6984);
nor U7450 (N_7450,N_6996,N_6041);
nand U7451 (N_7451,N_6153,N_6350);
or U7452 (N_7452,N_6669,N_6668);
nor U7453 (N_7453,N_6358,N_6073);
or U7454 (N_7454,N_6985,N_6119);
nand U7455 (N_7455,N_6288,N_6990);
xnor U7456 (N_7456,N_6161,N_6141);
xor U7457 (N_7457,N_6972,N_6945);
or U7458 (N_7458,N_6325,N_6212);
and U7459 (N_7459,N_6249,N_6755);
nor U7460 (N_7460,N_6526,N_6334);
nand U7461 (N_7461,N_6911,N_6689);
nand U7462 (N_7462,N_6477,N_6402);
or U7463 (N_7463,N_6362,N_6773);
nand U7464 (N_7464,N_6083,N_6230);
or U7465 (N_7465,N_6651,N_6758);
nor U7466 (N_7466,N_6686,N_6894);
and U7467 (N_7467,N_6604,N_6532);
or U7468 (N_7468,N_6420,N_6043);
or U7469 (N_7469,N_6497,N_6868);
or U7470 (N_7470,N_6033,N_6933);
and U7471 (N_7471,N_6527,N_6048);
nand U7472 (N_7472,N_6465,N_6271);
nor U7473 (N_7473,N_6389,N_6709);
nand U7474 (N_7474,N_6055,N_6759);
nor U7475 (N_7475,N_6176,N_6876);
and U7476 (N_7476,N_6242,N_6219);
nor U7477 (N_7477,N_6614,N_6419);
nor U7478 (N_7478,N_6088,N_6408);
and U7479 (N_7479,N_6854,N_6208);
nand U7480 (N_7480,N_6163,N_6368);
nand U7481 (N_7481,N_6749,N_6467);
or U7482 (N_7482,N_6805,N_6761);
and U7483 (N_7483,N_6142,N_6549);
nand U7484 (N_7484,N_6110,N_6263);
nor U7485 (N_7485,N_6906,N_6178);
nand U7486 (N_7486,N_6381,N_6579);
or U7487 (N_7487,N_6464,N_6824);
nand U7488 (N_7488,N_6572,N_6413);
and U7489 (N_7489,N_6663,N_6217);
or U7490 (N_7490,N_6929,N_6641);
and U7491 (N_7491,N_6566,N_6917);
and U7492 (N_7492,N_6456,N_6836);
nor U7493 (N_7493,N_6923,N_6546);
nand U7494 (N_7494,N_6741,N_6147);
or U7495 (N_7495,N_6862,N_6661);
nor U7496 (N_7496,N_6620,N_6822);
xor U7497 (N_7497,N_6075,N_6015);
or U7498 (N_7498,N_6481,N_6019);
xor U7499 (N_7499,N_6785,N_6965);
nand U7500 (N_7500,N_6623,N_6055);
or U7501 (N_7501,N_6279,N_6574);
or U7502 (N_7502,N_6657,N_6181);
and U7503 (N_7503,N_6770,N_6213);
nor U7504 (N_7504,N_6360,N_6581);
nand U7505 (N_7505,N_6346,N_6794);
nand U7506 (N_7506,N_6373,N_6215);
nand U7507 (N_7507,N_6318,N_6484);
and U7508 (N_7508,N_6538,N_6961);
nor U7509 (N_7509,N_6840,N_6341);
nand U7510 (N_7510,N_6425,N_6333);
or U7511 (N_7511,N_6021,N_6292);
and U7512 (N_7512,N_6898,N_6917);
and U7513 (N_7513,N_6004,N_6839);
or U7514 (N_7514,N_6358,N_6322);
xor U7515 (N_7515,N_6711,N_6598);
nor U7516 (N_7516,N_6767,N_6171);
nor U7517 (N_7517,N_6222,N_6931);
or U7518 (N_7518,N_6724,N_6102);
and U7519 (N_7519,N_6654,N_6411);
nand U7520 (N_7520,N_6677,N_6140);
or U7521 (N_7521,N_6156,N_6466);
and U7522 (N_7522,N_6825,N_6154);
and U7523 (N_7523,N_6579,N_6914);
nand U7524 (N_7524,N_6327,N_6028);
nand U7525 (N_7525,N_6328,N_6574);
nor U7526 (N_7526,N_6239,N_6050);
or U7527 (N_7527,N_6422,N_6482);
nor U7528 (N_7528,N_6921,N_6093);
and U7529 (N_7529,N_6021,N_6840);
nand U7530 (N_7530,N_6208,N_6367);
and U7531 (N_7531,N_6354,N_6870);
nand U7532 (N_7532,N_6930,N_6052);
and U7533 (N_7533,N_6730,N_6311);
nor U7534 (N_7534,N_6600,N_6310);
nand U7535 (N_7535,N_6568,N_6909);
or U7536 (N_7536,N_6583,N_6519);
nand U7537 (N_7537,N_6208,N_6037);
or U7538 (N_7538,N_6154,N_6275);
nor U7539 (N_7539,N_6459,N_6859);
or U7540 (N_7540,N_6755,N_6131);
nand U7541 (N_7541,N_6590,N_6332);
nor U7542 (N_7542,N_6816,N_6832);
nor U7543 (N_7543,N_6079,N_6515);
nand U7544 (N_7544,N_6617,N_6284);
or U7545 (N_7545,N_6888,N_6434);
and U7546 (N_7546,N_6059,N_6022);
nor U7547 (N_7547,N_6125,N_6300);
xnor U7548 (N_7548,N_6554,N_6153);
or U7549 (N_7549,N_6887,N_6329);
or U7550 (N_7550,N_6102,N_6215);
and U7551 (N_7551,N_6794,N_6567);
or U7552 (N_7552,N_6906,N_6808);
and U7553 (N_7553,N_6999,N_6384);
or U7554 (N_7554,N_6980,N_6521);
nor U7555 (N_7555,N_6467,N_6162);
xor U7556 (N_7556,N_6622,N_6165);
nand U7557 (N_7557,N_6953,N_6989);
nor U7558 (N_7558,N_6041,N_6040);
nand U7559 (N_7559,N_6181,N_6185);
or U7560 (N_7560,N_6610,N_6760);
nor U7561 (N_7561,N_6797,N_6341);
xor U7562 (N_7562,N_6131,N_6285);
nor U7563 (N_7563,N_6574,N_6975);
nor U7564 (N_7564,N_6480,N_6133);
or U7565 (N_7565,N_6497,N_6336);
and U7566 (N_7566,N_6508,N_6065);
nor U7567 (N_7567,N_6504,N_6245);
or U7568 (N_7568,N_6934,N_6859);
or U7569 (N_7569,N_6609,N_6202);
or U7570 (N_7570,N_6437,N_6761);
and U7571 (N_7571,N_6064,N_6530);
nand U7572 (N_7572,N_6397,N_6038);
and U7573 (N_7573,N_6780,N_6347);
nand U7574 (N_7574,N_6594,N_6931);
or U7575 (N_7575,N_6854,N_6966);
nor U7576 (N_7576,N_6641,N_6208);
nand U7577 (N_7577,N_6308,N_6486);
and U7578 (N_7578,N_6896,N_6631);
xnor U7579 (N_7579,N_6737,N_6853);
xnor U7580 (N_7580,N_6945,N_6915);
nor U7581 (N_7581,N_6133,N_6818);
or U7582 (N_7582,N_6990,N_6530);
nor U7583 (N_7583,N_6789,N_6311);
or U7584 (N_7584,N_6315,N_6126);
xor U7585 (N_7585,N_6681,N_6147);
xnor U7586 (N_7586,N_6362,N_6720);
xor U7587 (N_7587,N_6442,N_6707);
and U7588 (N_7588,N_6036,N_6138);
nor U7589 (N_7589,N_6933,N_6487);
nand U7590 (N_7590,N_6623,N_6132);
and U7591 (N_7591,N_6344,N_6672);
nor U7592 (N_7592,N_6608,N_6475);
and U7593 (N_7593,N_6604,N_6373);
nor U7594 (N_7594,N_6781,N_6426);
nand U7595 (N_7595,N_6027,N_6712);
xor U7596 (N_7596,N_6873,N_6847);
nor U7597 (N_7597,N_6213,N_6377);
and U7598 (N_7598,N_6405,N_6052);
or U7599 (N_7599,N_6534,N_6817);
nand U7600 (N_7600,N_6391,N_6907);
nand U7601 (N_7601,N_6871,N_6777);
nor U7602 (N_7602,N_6046,N_6346);
and U7603 (N_7603,N_6856,N_6143);
nand U7604 (N_7604,N_6147,N_6756);
nor U7605 (N_7605,N_6629,N_6510);
or U7606 (N_7606,N_6151,N_6280);
xnor U7607 (N_7607,N_6621,N_6953);
nand U7608 (N_7608,N_6373,N_6075);
and U7609 (N_7609,N_6112,N_6227);
nor U7610 (N_7610,N_6756,N_6179);
or U7611 (N_7611,N_6276,N_6528);
and U7612 (N_7612,N_6748,N_6702);
nor U7613 (N_7613,N_6680,N_6867);
or U7614 (N_7614,N_6129,N_6379);
nor U7615 (N_7615,N_6889,N_6407);
and U7616 (N_7616,N_6456,N_6012);
nor U7617 (N_7617,N_6374,N_6837);
or U7618 (N_7618,N_6206,N_6665);
nand U7619 (N_7619,N_6731,N_6214);
and U7620 (N_7620,N_6408,N_6197);
nor U7621 (N_7621,N_6531,N_6545);
or U7622 (N_7622,N_6939,N_6704);
nor U7623 (N_7623,N_6035,N_6292);
and U7624 (N_7624,N_6361,N_6605);
or U7625 (N_7625,N_6008,N_6042);
nor U7626 (N_7626,N_6557,N_6249);
and U7627 (N_7627,N_6573,N_6626);
or U7628 (N_7628,N_6603,N_6856);
or U7629 (N_7629,N_6476,N_6522);
and U7630 (N_7630,N_6597,N_6659);
or U7631 (N_7631,N_6665,N_6501);
nor U7632 (N_7632,N_6206,N_6501);
nand U7633 (N_7633,N_6430,N_6591);
or U7634 (N_7634,N_6692,N_6995);
nor U7635 (N_7635,N_6444,N_6941);
nand U7636 (N_7636,N_6029,N_6708);
nand U7637 (N_7637,N_6300,N_6269);
or U7638 (N_7638,N_6313,N_6650);
nand U7639 (N_7639,N_6563,N_6048);
nand U7640 (N_7640,N_6907,N_6092);
or U7641 (N_7641,N_6084,N_6451);
or U7642 (N_7642,N_6334,N_6431);
and U7643 (N_7643,N_6558,N_6321);
or U7644 (N_7644,N_6496,N_6926);
and U7645 (N_7645,N_6984,N_6580);
nor U7646 (N_7646,N_6777,N_6023);
and U7647 (N_7647,N_6668,N_6108);
or U7648 (N_7648,N_6362,N_6572);
nand U7649 (N_7649,N_6106,N_6728);
nand U7650 (N_7650,N_6288,N_6035);
or U7651 (N_7651,N_6818,N_6360);
or U7652 (N_7652,N_6516,N_6798);
or U7653 (N_7653,N_6469,N_6675);
nor U7654 (N_7654,N_6491,N_6978);
nand U7655 (N_7655,N_6414,N_6127);
or U7656 (N_7656,N_6513,N_6660);
and U7657 (N_7657,N_6858,N_6292);
and U7658 (N_7658,N_6315,N_6116);
nand U7659 (N_7659,N_6089,N_6266);
nor U7660 (N_7660,N_6872,N_6671);
nand U7661 (N_7661,N_6606,N_6884);
nor U7662 (N_7662,N_6870,N_6908);
or U7663 (N_7663,N_6516,N_6551);
nand U7664 (N_7664,N_6679,N_6026);
nor U7665 (N_7665,N_6386,N_6950);
nor U7666 (N_7666,N_6664,N_6563);
or U7667 (N_7667,N_6840,N_6459);
nor U7668 (N_7668,N_6977,N_6220);
nand U7669 (N_7669,N_6306,N_6327);
and U7670 (N_7670,N_6457,N_6054);
nand U7671 (N_7671,N_6451,N_6798);
nor U7672 (N_7672,N_6489,N_6236);
xnor U7673 (N_7673,N_6789,N_6602);
nand U7674 (N_7674,N_6244,N_6790);
nand U7675 (N_7675,N_6505,N_6973);
or U7676 (N_7676,N_6721,N_6875);
nand U7677 (N_7677,N_6475,N_6060);
and U7678 (N_7678,N_6644,N_6278);
xnor U7679 (N_7679,N_6985,N_6036);
or U7680 (N_7680,N_6445,N_6443);
and U7681 (N_7681,N_6101,N_6474);
nand U7682 (N_7682,N_6469,N_6507);
and U7683 (N_7683,N_6062,N_6362);
xor U7684 (N_7684,N_6994,N_6024);
and U7685 (N_7685,N_6593,N_6397);
xnor U7686 (N_7686,N_6808,N_6989);
or U7687 (N_7687,N_6252,N_6113);
nand U7688 (N_7688,N_6009,N_6040);
nand U7689 (N_7689,N_6616,N_6057);
or U7690 (N_7690,N_6030,N_6981);
or U7691 (N_7691,N_6411,N_6994);
nand U7692 (N_7692,N_6953,N_6649);
nor U7693 (N_7693,N_6604,N_6378);
nor U7694 (N_7694,N_6256,N_6802);
nor U7695 (N_7695,N_6230,N_6410);
nand U7696 (N_7696,N_6082,N_6608);
nand U7697 (N_7697,N_6236,N_6242);
nor U7698 (N_7698,N_6233,N_6017);
nor U7699 (N_7699,N_6637,N_6429);
or U7700 (N_7700,N_6773,N_6403);
nor U7701 (N_7701,N_6279,N_6138);
or U7702 (N_7702,N_6788,N_6025);
nand U7703 (N_7703,N_6062,N_6906);
nor U7704 (N_7704,N_6281,N_6206);
or U7705 (N_7705,N_6643,N_6257);
or U7706 (N_7706,N_6532,N_6814);
xor U7707 (N_7707,N_6623,N_6219);
nand U7708 (N_7708,N_6792,N_6277);
xnor U7709 (N_7709,N_6787,N_6728);
or U7710 (N_7710,N_6559,N_6657);
nor U7711 (N_7711,N_6918,N_6366);
or U7712 (N_7712,N_6649,N_6586);
nand U7713 (N_7713,N_6305,N_6422);
xor U7714 (N_7714,N_6161,N_6171);
or U7715 (N_7715,N_6221,N_6875);
or U7716 (N_7716,N_6076,N_6737);
nor U7717 (N_7717,N_6849,N_6724);
or U7718 (N_7718,N_6053,N_6172);
nand U7719 (N_7719,N_6575,N_6038);
and U7720 (N_7720,N_6117,N_6163);
nand U7721 (N_7721,N_6640,N_6022);
nor U7722 (N_7722,N_6324,N_6417);
or U7723 (N_7723,N_6638,N_6858);
and U7724 (N_7724,N_6347,N_6281);
or U7725 (N_7725,N_6214,N_6865);
or U7726 (N_7726,N_6375,N_6767);
nor U7727 (N_7727,N_6811,N_6418);
nor U7728 (N_7728,N_6271,N_6153);
and U7729 (N_7729,N_6677,N_6991);
and U7730 (N_7730,N_6633,N_6551);
and U7731 (N_7731,N_6664,N_6740);
or U7732 (N_7732,N_6678,N_6810);
or U7733 (N_7733,N_6593,N_6327);
nor U7734 (N_7734,N_6624,N_6282);
or U7735 (N_7735,N_6070,N_6950);
xor U7736 (N_7736,N_6404,N_6502);
xnor U7737 (N_7737,N_6314,N_6808);
nand U7738 (N_7738,N_6011,N_6473);
nor U7739 (N_7739,N_6008,N_6378);
or U7740 (N_7740,N_6393,N_6494);
nor U7741 (N_7741,N_6265,N_6768);
nor U7742 (N_7742,N_6839,N_6618);
nor U7743 (N_7743,N_6152,N_6763);
and U7744 (N_7744,N_6484,N_6382);
or U7745 (N_7745,N_6385,N_6931);
xor U7746 (N_7746,N_6193,N_6310);
nor U7747 (N_7747,N_6734,N_6442);
nand U7748 (N_7748,N_6930,N_6683);
nor U7749 (N_7749,N_6155,N_6397);
and U7750 (N_7750,N_6179,N_6554);
nand U7751 (N_7751,N_6647,N_6435);
and U7752 (N_7752,N_6104,N_6622);
nand U7753 (N_7753,N_6294,N_6511);
and U7754 (N_7754,N_6292,N_6108);
or U7755 (N_7755,N_6729,N_6659);
nand U7756 (N_7756,N_6240,N_6740);
and U7757 (N_7757,N_6430,N_6792);
nand U7758 (N_7758,N_6965,N_6171);
nor U7759 (N_7759,N_6291,N_6226);
or U7760 (N_7760,N_6714,N_6026);
xor U7761 (N_7761,N_6383,N_6575);
nand U7762 (N_7762,N_6843,N_6945);
nand U7763 (N_7763,N_6058,N_6308);
and U7764 (N_7764,N_6630,N_6625);
or U7765 (N_7765,N_6295,N_6321);
or U7766 (N_7766,N_6475,N_6777);
nor U7767 (N_7767,N_6339,N_6626);
nand U7768 (N_7768,N_6684,N_6880);
and U7769 (N_7769,N_6568,N_6014);
nand U7770 (N_7770,N_6456,N_6736);
and U7771 (N_7771,N_6035,N_6537);
and U7772 (N_7772,N_6088,N_6740);
nand U7773 (N_7773,N_6272,N_6610);
and U7774 (N_7774,N_6581,N_6565);
nand U7775 (N_7775,N_6936,N_6245);
nor U7776 (N_7776,N_6481,N_6120);
nand U7777 (N_7777,N_6040,N_6265);
and U7778 (N_7778,N_6566,N_6148);
nor U7779 (N_7779,N_6986,N_6124);
nand U7780 (N_7780,N_6866,N_6298);
nand U7781 (N_7781,N_6822,N_6305);
nor U7782 (N_7782,N_6657,N_6728);
nor U7783 (N_7783,N_6381,N_6374);
xor U7784 (N_7784,N_6944,N_6619);
and U7785 (N_7785,N_6295,N_6602);
or U7786 (N_7786,N_6660,N_6843);
and U7787 (N_7787,N_6704,N_6725);
and U7788 (N_7788,N_6483,N_6444);
nand U7789 (N_7789,N_6075,N_6541);
nand U7790 (N_7790,N_6597,N_6082);
or U7791 (N_7791,N_6486,N_6445);
and U7792 (N_7792,N_6630,N_6879);
or U7793 (N_7793,N_6730,N_6786);
xor U7794 (N_7794,N_6731,N_6144);
nand U7795 (N_7795,N_6898,N_6275);
xor U7796 (N_7796,N_6273,N_6361);
nor U7797 (N_7797,N_6228,N_6475);
and U7798 (N_7798,N_6500,N_6827);
nand U7799 (N_7799,N_6268,N_6293);
nand U7800 (N_7800,N_6738,N_6825);
or U7801 (N_7801,N_6871,N_6518);
or U7802 (N_7802,N_6004,N_6695);
and U7803 (N_7803,N_6819,N_6223);
nor U7804 (N_7804,N_6780,N_6181);
and U7805 (N_7805,N_6250,N_6475);
and U7806 (N_7806,N_6985,N_6808);
nor U7807 (N_7807,N_6094,N_6922);
or U7808 (N_7808,N_6953,N_6930);
or U7809 (N_7809,N_6701,N_6049);
or U7810 (N_7810,N_6632,N_6833);
nand U7811 (N_7811,N_6923,N_6255);
and U7812 (N_7812,N_6883,N_6911);
xor U7813 (N_7813,N_6307,N_6768);
nor U7814 (N_7814,N_6592,N_6736);
nand U7815 (N_7815,N_6213,N_6437);
nand U7816 (N_7816,N_6512,N_6555);
nand U7817 (N_7817,N_6844,N_6818);
and U7818 (N_7818,N_6719,N_6090);
and U7819 (N_7819,N_6938,N_6895);
xor U7820 (N_7820,N_6219,N_6101);
nor U7821 (N_7821,N_6845,N_6684);
or U7822 (N_7822,N_6181,N_6041);
or U7823 (N_7823,N_6128,N_6180);
and U7824 (N_7824,N_6658,N_6712);
nor U7825 (N_7825,N_6105,N_6692);
or U7826 (N_7826,N_6710,N_6939);
nor U7827 (N_7827,N_6454,N_6639);
and U7828 (N_7828,N_6836,N_6665);
nor U7829 (N_7829,N_6468,N_6895);
or U7830 (N_7830,N_6498,N_6686);
and U7831 (N_7831,N_6783,N_6651);
nor U7832 (N_7832,N_6616,N_6946);
nand U7833 (N_7833,N_6175,N_6198);
xnor U7834 (N_7834,N_6296,N_6791);
and U7835 (N_7835,N_6629,N_6792);
nand U7836 (N_7836,N_6817,N_6822);
xor U7837 (N_7837,N_6029,N_6022);
and U7838 (N_7838,N_6351,N_6204);
nand U7839 (N_7839,N_6820,N_6198);
or U7840 (N_7840,N_6303,N_6241);
nor U7841 (N_7841,N_6300,N_6653);
nand U7842 (N_7842,N_6100,N_6997);
nand U7843 (N_7843,N_6224,N_6112);
and U7844 (N_7844,N_6301,N_6356);
nor U7845 (N_7845,N_6712,N_6641);
and U7846 (N_7846,N_6136,N_6537);
xor U7847 (N_7847,N_6660,N_6964);
xnor U7848 (N_7848,N_6336,N_6349);
and U7849 (N_7849,N_6341,N_6849);
or U7850 (N_7850,N_6024,N_6529);
or U7851 (N_7851,N_6503,N_6741);
nand U7852 (N_7852,N_6239,N_6261);
nor U7853 (N_7853,N_6312,N_6418);
or U7854 (N_7854,N_6339,N_6254);
and U7855 (N_7855,N_6154,N_6150);
nand U7856 (N_7856,N_6235,N_6460);
nor U7857 (N_7857,N_6185,N_6475);
or U7858 (N_7858,N_6216,N_6382);
nand U7859 (N_7859,N_6331,N_6064);
nor U7860 (N_7860,N_6839,N_6826);
or U7861 (N_7861,N_6102,N_6134);
or U7862 (N_7862,N_6991,N_6016);
nor U7863 (N_7863,N_6669,N_6907);
nor U7864 (N_7864,N_6141,N_6204);
nand U7865 (N_7865,N_6608,N_6194);
xor U7866 (N_7866,N_6468,N_6987);
xnor U7867 (N_7867,N_6567,N_6521);
or U7868 (N_7868,N_6606,N_6020);
nor U7869 (N_7869,N_6549,N_6863);
and U7870 (N_7870,N_6339,N_6570);
or U7871 (N_7871,N_6786,N_6812);
nand U7872 (N_7872,N_6369,N_6374);
and U7873 (N_7873,N_6979,N_6549);
nand U7874 (N_7874,N_6160,N_6906);
nor U7875 (N_7875,N_6251,N_6655);
or U7876 (N_7876,N_6250,N_6090);
nand U7877 (N_7877,N_6319,N_6628);
or U7878 (N_7878,N_6766,N_6448);
xnor U7879 (N_7879,N_6513,N_6200);
or U7880 (N_7880,N_6175,N_6131);
and U7881 (N_7881,N_6611,N_6588);
nor U7882 (N_7882,N_6641,N_6161);
xnor U7883 (N_7883,N_6465,N_6235);
nand U7884 (N_7884,N_6021,N_6200);
nor U7885 (N_7885,N_6782,N_6382);
or U7886 (N_7886,N_6792,N_6085);
and U7887 (N_7887,N_6184,N_6665);
or U7888 (N_7888,N_6979,N_6108);
and U7889 (N_7889,N_6241,N_6560);
xor U7890 (N_7890,N_6280,N_6204);
or U7891 (N_7891,N_6957,N_6153);
xnor U7892 (N_7892,N_6915,N_6636);
xor U7893 (N_7893,N_6814,N_6249);
nand U7894 (N_7894,N_6142,N_6672);
xor U7895 (N_7895,N_6570,N_6970);
and U7896 (N_7896,N_6848,N_6107);
or U7897 (N_7897,N_6481,N_6672);
nand U7898 (N_7898,N_6329,N_6353);
nand U7899 (N_7899,N_6717,N_6315);
and U7900 (N_7900,N_6110,N_6354);
or U7901 (N_7901,N_6552,N_6157);
nor U7902 (N_7902,N_6838,N_6809);
nor U7903 (N_7903,N_6612,N_6613);
nor U7904 (N_7904,N_6063,N_6492);
nand U7905 (N_7905,N_6024,N_6001);
xnor U7906 (N_7906,N_6562,N_6626);
nand U7907 (N_7907,N_6152,N_6507);
nor U7908 (N_7908,N_6486,N_6065);
nor U7909 (N_7909,N_6608,N_6158);
or U7910 (N_7910,N_6288,N_6153);
and U7911 (N_7911,N_6645,N_6658);
nor U7912 (N_7912,N_6451,N_6353);
nor U7913 (N_7913,N_6228,N_6714);
nor U7914 (N_7914,N_6226,N_6361);
nand U7915 (N_7915,N_6052,N_6206);
nor U7916 (N_7916,N_6026,N_6394);
nand U7917 (N_7917,N_6113,N_6972);
nand U7918 (N_7918,N_6398,N_6117);
and U7919 (N_7919,N_6290,N_6768);
nor U7920 (N_7920,N_6869,N_6231);
nor U7921 (N_7921,N_6753,N_6330);
and U7922 (N_7922,N_6725,N_6038);
and U7923 (N_7923,N_6904,N_6814);
or U7924 (N_7924,N_6199,N_6187);
nand U7925 (N_7925,N_6438,N_6646);
and U7926 (N_7926,N_6345,N_6014);
xnor U7927 (N_7927,N_6606,N_6832);
nor U7928 (N_7928,N_6495,N_6215);
nand U7929 (N_7929,N_6053,N_6111);
or U7930 (N_7930,N_6877,N_6360);
nand U7931 (N_7931,N_6349,N_6522);
or U7932 (N_7932,N_6513,N_6592);
and U7933 (N_7933,N_6370,N_6000);
and U7934 (N_7934,N_6045,N_6893);
nor U7935 (N_7935,N_6127,N_6520);
or U7936 (N_7936,N_6748,N_6458);
nor U7937 (N_7937,N_6245,N_6775);
or U7938 (N_7938,N_6155,N_6588);
and U7939 (N_7939,N_6994,N_6906);
nor U7940 (N_7940,N_6350,N_6135);
and U7941 (N_7941,N_6236,N_6339);
nor U7942 (N_7942,N_6491,N_6512);
nor U7943 (N_7943,N_6457,N_6842);
or U7944 (N_7944,N_6870,N_6490);
or U7945 (N_7945,N_6288,N_6416);
or U7946 (N_7946,N_6780,N_6486);
or U7947 (N_7947,N_6711,N_6536);
or U7948 (N_7948,N_6250,N_6455);
and U7949 (N_7949,N_6332,N_6589);
xnor U7950 (N_7950,N_6664,N_6219);
or U7951 (N_7951,N_6563,N_6333);
nand U7952 (N_7952,N_6767,N_6411);
nand U7953 (N_7953,N_6762,N_6123);
or U7954 (N_7954,N_6394,N_6899);
nor U7955 (N_7955,N_6842,N_6433);
or U7956 (N_7956,N_6542,N_6005);
nor U7957 (N_7957,N_6053,N_6568);
nor U7958 (N_7958,N_6476,N_6556);
and U7959 (N_7959,N_6397,N_6903);
and U7960 (N_7960,N_6045,N_6140);
nand U7961 (N_7961,N_6099,N_6970);
xnor U7962 (N_7962,N_6052,N_6036);
or U7963 (N_7963,N_6847,N_6438);
nor U7964 (N_7964,N_6830,N_6712);
or U7965 (N_7965,N_6535,N_6416);
or U7966 (N_7966,N_6004,N_6477);
nor U7967 (N_7967,N_6719,N_6736);
or U7968 (N_7968,N_6278,N_6153);
nor U7969 (N_7969,N_6160,N_6676);
or U7970 (N_7970,N_6515,N_6686);
nand U7971 (N_7971,N_6044,N_6160);
nor U7972 (N_7972,N_6143,N_6344);
or U7973 (N_7973,N_6195,N_6154);
or U7974 (N_7974,N_6494,N_6025);
and U7975 (N_7975,N_6911,N_6491);
or U7976 (N_7976,N_6199,N_6532);
nand U7977 (N_7977,N_6572,N_6491);
and U7978 (N_7978,N_6722,N_6211);
nor U7979 (N_7979,N_6758,N_6490);
nor U7980 (N_7980,N_6244,N_6243);
nand U7981 (N_7981,N_6102,N_6485);
nor U7982 (N_7982,N_6131,N_6007);
xor U7983 (N_7983,N_6420,N_6486);
or U7984 (N_7984,N_6827,N_6366);
nand U7985 (N_7985,N_6767,N_6494);
nand U7986 (N_7986,N_6124,N_6783);
and U7987 (N_7987,N_6201,N_6510);
and U7988 (N_7988,N_6996,N_6892);
xor U7989 (N_7989,N_6505,N_6035);
nand U7990 (N_7990,N_6195,N_6037);
xor U7991 (N_7991,N_6513,N_6917);
xor U7992 (N_7992,N_6319,N_6945);
or U7993 (N_7993,N_6703,N_6983);
and U7994 (N_7994,N_6968,N_6870);
nand U7995 (N_7995,N_6732,N_6627);
or U7996 (N_7996,N_6231,N_6900);
and U7997 (N_7997,N_6115,N_6592);
and U7998 (N_7998,N_6869,N_6017);
nor U7999 (N_7999,N_6179,N_6309);
nor U8000 (N_8000,N_7620,N_7067);
or U8001 (N_8001,N_7233,N_7205);
and U8002 (N_8002,N_7771,N_7898);
nor U8003 (N_8003,N_7585,N_7519);
nand U8004 (N_8004,N_7170,N_7389);
nor U8005 (N_8005,N_7655,N_7195);
and U8006 (N_8006,N_7449,N_7154);
and U8007 (N_8007,N_7095,N_7946);
or U8008 (N_8008,N_7662,N_7610);
nand U8009 (N_8009,N_7457,N_7561);
or U8010 (N_8010,N_7715,N_7252);
or U8011 (N_8011,N_7129,N_7162);
nor U8012 (N_8012,N_7375,N_7717);
nand U8013 (N_8013,N_7007,N_7214);
or U8014 (N_8014,N_7918,N_7684);
or U8015 (N_8015,N_7035,N_7444);
nor U8016 (N_8016,N_7520,N_7969);
and U8017 (N_8017,N_7299,N_7703);
nand U8018 (N_8018,N_7454,N_7658);
and U8019 (N_8019,N_7335,N_7704);
or U8020 (N_8020,N_7612,N_7452);
or U8021 (N_8021,N_7223,N_7880);
and U8022 (N_8022,N_7671,N_7025);
nor U8023 (N_8023,N_7075,N_7408);
nand U8024 (N_8024,N_7152,N_7925);
xnor U8025 (N_8025,N_7575,N_7398);
nand U8026 (N_8026,N_7827,N_7243);
nand U8027 (N_8027,N_7222,N_7697);
xnor U8028 (N_8028,N_7015,N_7748);
nor U8029 (N_8029,N_7582,N_7884);
nand U8030 (N_8030,N_7388,N_7857);
nand U8031 (N_8031,N_7694,N_7669);
xnor U8032 (N_8032,N_7426,N_7167);
and U8033 (N_8033,N_7951,N_7163);
nand U8034 (N_8034,N_7189,N_7732);
xnor U8035 (N_8035,N_7467,N_7029);
xnor U8036 (N_8036,N_7374,N_7183);
nor U8037 (N_8037,N_7063,N_7401);
nand U8038 (N_8038,N_7562,N_7654);
nand U8039 (N_8039,N_7216,N_7586);
or U8040 (N_8040,N_7746,N_7212);
and U8041 (N_8041,N_7573,N_7279);
nand U8042 (N_8042,N_7229,N_7307);
or U8043 (N_8043,N_7310,N_7415);
and U8044 (N_8044,N_7413,N_7277);
and U8045 (N_8045,N_7339,N_7574);
nor U8046 (N_8046,N_7498,N_7967);
xor U8047 (N_8047,N_7066,N_7423);
and U8048 (N_8048,N_7246,N_7634);
nand U8049 (N_8049,N_7799,N_7466);
nor U8050 (N_8050,N_7316,N_7802);
or U8051 (N_8051,N_7357,N_7461);
nor U8052 (N_8052,N_7440,N_7087);
xnor U8053 (N_8053,N_7819,N_7058);
nand U8054 (N_8054,N_7679,N_7270);
and U8055 (N_8055,N_7230,N_7200);
nand U8056 (N_8056,N_7783,N_7708);
nand U8057 (N_8057,N_7173,N_7462);
and U8058 (N_8058,N_7516,N_7930);
nand U8059 (N_8059,N_7014,N_7098);
and U8060 (N_8060,N_7139,N_7022);
or U8061 (N_8061,N_7936,N_7053);
and U8062 (N_8062,N_7455,N_7278);
nor U8063 (N_8063,N_7425,N_7240);
and U8064 (N_8064,N_7912,N_7852);
and U8065 (N_8065,N_7084,N_7554);
and U8066 (N_8066,N_7446,N_7097);
or U8067 (N_8067,N_7101,N_7241);
nor U8068 (N_8068,N_7903,N_7393);
nor U8069 (N_8069,N_7009,N_7529);
and U8070 (N_8070,N_7823,N_7821);
or U8071 (N_8071,N_7938,N_7759);
and U8072 (N_8072,N_7418,N_7504);
nor U8073 (N_8073,N_7020,N_7537);
nor U8074 (N_8074,N_7650,N_7992);
or U8075 (N_8075,N_7292,N_7735);
nor U8076 (N_8076,N_7138,N_7714);
nand U8077 (N_8077,N_7400,N_7550);
or U8078 (N_8078,N_7798,N_7756);
or U8079 (N_8079,N_7631,N_7136);
and U8080 (N_8080,N_7244,N_7795);
or U8081 (N_8081,N_7890,N_7604);
xnor U8082 (N_8082,N_7849,N_7813);
and U8083 (N_8083,N_7153,N_7206);
nand U8084 (N_8084,N_7940,N_7439);
nand U8085 (N_8085,N_7709,N_7851);
nor U8086 (N_8086,N_7286,N_7038);
nand U8087 (N_8087,N_7046,N_7738);
nor U8088 (N_8088,N_7869,N_7338);
or U8089 (N_8089,N_7227,N_7909);
nand U8090 (N_8090,N_7594,N_7830);
or U8091 (N_8091,N_7961,N_7028);
nor U8092 (N_8092,N_7970,N_7803);
or U8093 (N_8093,N_7993,N_7282);
and U8094 (N_8094,N_7826,N_7469);
xor U8095 (N_8095,N_7488,N_7831);
and U8096 (N_8096,N_7668,N_7172);
nand U8097 (N_8097,N_7623,N_7531);
or U8098 (N_8098,N_7683,N_7928);
nor U8099 (N_8099,N_7239,N_7253);
nor U8100 (N_8100,N_7257,N_7117);
nand U8101 (N_8101,N_7944,N_7350);
or U8102 (N_8102,N_7559,N_7192);
nand U8103 (N_8103,N_7770,N_7601);
and U8104 (N_8104,N_7924,N_7718);
xor U8105 (N_8105,N_7361,N_7474);
or U8106 (N_8106,N_7571,N_7442);
nor U8107 (N_8107,N_7207,N_7451);
nand U8108 (N_8108,N_7533,N_7532);
nor U8109 (N_8109,N_7228,N_7273);
nand U8110 (N_8110,N_7690,N_7952);
nor U8111 (N_8111,N_7850,N_7731);
xnor U8112 (N_8112,N_7224,N_7329);
nand U8113 (N_8113,N_7313,N_7337);
and U8114 (N_8114,N_7921,N_7419);
and U8115 (N_8115,N_7185,N_7635);
nand U8116 (N_8116,N_7569,N_7838);
or U8117 (N_8117,N_7094,N_7584);
nand U8118 (N_8118,N_7019,N_7589);
and U8119 (N_8119,N_7365,N_7816);
xnor U8120 (N_8120,N_7932,N_7905);
nor U8121 (N_8121,N_7927,N_7876);
and U8122 (N_8122,N_7232,N_7399);
and U8123 (N_8123,N_7283,N_7373);
nor U8124 (N_8124,N_7395,N_7051);
nand U8125 (N_8125,N_7054,N_7633);
or U8126 (N_8126,N_7079,N_7006);
nand U8127 (N_8127,N_7591,N_7236);
nand U8128 (N_8128,N_7215,N_7080);
or U8129 (N_8129,N_7264,N_7954);
nor U8130 (N_8130,N_7476,N_7203);
xor U8131 (N_8131,N_7701,N_7037);
nand U8132 (N_8132,N_7693,N_7722);
and U8133 (N_8133,N_7651,N_7837);
and U8134 (N_8134,N_7602,N_7652);
nor U8135 (N_8135,N_7753,N_7359);
or U8136 (N_8136,N_7017,N_7674);
and U8137 (N_8137,N_7560,N_7113);
nor U8138 (N_8138,N_7985,N_7441);
xor U8139 (N_8139,N_7894,N_7456);
nand U8140 (N_8140,N_7854,N_7371);
nand U8141 (N_8141,N_7306,N_7887);
and U8142 (N_8142,N_7742,N_7839);
nor U8143 (N_8143,N_7551,N_7832);
or U8144 (N_8144,N_7406,N_7128);
or U8145 (N_8145,N_7209,N_7906);
nor U8146 (N_8146,N_7500,N_7546);
or U8147 (N_8147,N_7515,N_7011);
nand U8148 (N_8148,N_7809,N_7260);
xor U8149 (N_8149,N_7323,N_7119);
nor U8150 (N_8150,N_7123,N_7778);
and U8151 (N_8151,N_7979,N_7131);
and U8152 (N_8152,N_7645,N_7625);
and U8153 (N_8153,N_7489,N_7998);
nand U8154 (N_8154,N_7547,N_7424);
and U8155 (N_8155,N_7380,N_7583);
nand U8156 (N_8156,N_7397,N_7872);
nor U8157 (N_8157,N_7013,N_7508);
nand U8158 (N_8158,N_7590,N_7176);
nand U8159 (N_8159,N_7100,N_7293);
nor U8160 (N_8160,N_7268,N_7737);
nand U8161 (N_8161,N_7390,N_7699);
nand U8162 (N_8162,N_7367,N_7787);
nand U8163 (N_8163,N_7042,N_7453);
and U8164 (N_8164,N_7682,N_7065);
and U8165 (N_8165,N_7405,N_7002);
nor U8166 (N_8166,N_7160,N_7866);
nand U8167 (N_8167,N_7739,N_7311);
nor U8168 (N_8168,N_7910,N_7353);
or U8169 (N_8169,N_7638,N_7664);
or U8170 (N_8170,N_7641,N_7956);
nand U8171 (N_8171,N_7609,N_7934);
nand U8172 (N_8172,N_7070,N_7143);
nor U8173 (N_8173,N_7522,N_7345);
or U8174 (N_8174,N_7475,N_7146);
nand U8175 (N_8175,N_7259,N_7768);
nand U8176 (N_8176,N_7685,N_7317);
nand U8177 (N_8177,N_7719,N_7812);
nand U8178 (N_8178,N_7542,N_7071);
or U8179 (N_8179,N_7501,N_7964);
nor U8180 (N_8180,N_7741,N_7555);
or U8181 (N_8181,N_7549,N_7191);
nand U8182 (N_8182,N_7363,N_7607);
nor U8183 (N_8183,N_7174,N_7328);
or U8184 (N_8184,N_7412,N_7284);
xnor U8185 (N_8185,N_7465,N_7868);
and U8186 (N_8186,N_7125,N_7657);
or U8187 (N_8187,N_7057,N_7744);
or U8188 (N_8188,N_7908,N_7618);
nand U8189 (N_8189,N_7793,N_7566);
xor U8190 (N_8190,N_7073,N_7644);
nor U8191 (N_8191,N_7960,N_7939);
and U8192 (N_8192,N_7841,N_7580);
and U8193 (N_8193,N_7369,N_7261);
and U8194 (N_8194,N_7751,N_7164);
or U8195 (N_8195,N_7889,N_7289);
or U8196 (N_8196,N_7696,N_7613);
nand U8197 (N_8197,N_7687,N_7962);
and U8198 (N_8198,N_7106,N_7496);
nor U8199 (N_8199,N_7161,N_7341);
xor U8200 (N_8200,N_7061,N_7179);
and U8201 (N_8201,N_7312,N_7196);
xnor U8202 (N_8202,N_7178,N_7221);
and U8203 (N_8203,N_7304,N_7581);
and U8204 (N_8204,N_7991,N_7198);
nor U8205 (N_8205,N_7151,N_7409);
or U8206 (N_8206,N_7303,N_7211);
or U8207 (N_8207,N_7135,N_7484);
xor U8208 (N_8208,N_7104,N_7729);
xnor U8209 (N_8209,N_7391,N_7362);
or U8210 (N_8210,N_7647,N_7616);
and U8211 (N_8211,N_7743,N_7309);
nor U8212 (N_8212,N_7472,N_7570);
or U8213 (N_8213,N_7319,N_7976);
and U8214 (N_8214,N_7263,N_7110);
nor U8215 (N_8215,N_7443,N_7430);
nor U8216 (N_8216,N_7606,N_7855);
or U8217 (N_8217,N_7226,N_7049);
nor U8218 (N_8218,N_7186,N_7235);
and U8219 (N_8219,N_7349,N_7072);
or U8220 (N_8220,N_7346,N_7245);
nand U8221 (N_8221,N_7711,N_7957);
nor U8222 (N_8222,N_7535,N_7291);
nor U8223 (N_8223,N_7997,N_7929);
or U8224 (N_8224,N_7220,N_7420);
nand U8225 (N_8225,N_7911,N_7392);
or U8226 (N_8226,N_7473,N_7158);
nor U8227 (N_8227,N_7495,N_7450);
nor U8228 (N_8228,N_7864,N_7706);
and U8229 (N_8229,N_7807,N_7190);
and U8230 (N_8230,N_7937,N_7916);
and U8231 (N_8231,N_7863,N_7681);
nor U8232 (N_8232,N_7315,N_7112);
or U8233 (N_8233,N_7434,N_7386);
or U8234 (N_8234,N_7695,N_7765);
nor U8235 (N_8235,N_7217,N_7619);
nand U8236 (N_8236,N_7394,N_7530);
nor U8237 (N_8237,N_7790,N_7817);
or U8238 (N_8238,N_7920,N_7527);
or U8239 (N_8239,N_7935,N_7132);
nand U8240 (N_8240,N_7672,N_7250);
nor U8241 (N_8241,N_7130,N_7897);
xnor U8242 (N_8242,N_7210,N_7707);
nor U8243 (N_8243,N_7432,N_7758);
nand U8244 (N_8244,N_7092,N_7843);
and U8245 (N_8245,N_7358,N_7077);
nand U8246 (N_8246,N_7387,N_7248);
xnor U8247 (N_8247,N_7596,N_7081);
or U8248 (N_8248,N_7971,N_7325);
nand U8249 (N_8249,N_7494,N_7523);
and U8250 (N_8250,N_7579,N_7538);
nor U8251 (N_8251,N_7105,N_7789);
nor U8252 (N_8252,N_7567,N_7989);
nor U8253 (N_8253,N_7822,N_7806);
and U8254 (N_8254,N_7421,N_7902);
or U8255 (N_8255,N_7667,N_7385);
nor U8256 (N_8256,N_7725,N_7481);
nand U8257 (N_8257,N_7564,N_7086);
nand U8258 (N_8258,N_7507,N_7984);
or U8259 (N_8259,N_7521,N_7640);
and U8260 (N_8260,N_7900,N_7274);
or U8261 (N_8261,N_7008,N_7673);
nor U8262 (N_8262,N_7977,N_7942);
nand U8263 (N_8263,N_7755,N_7797);
nand U8264 (N_8264,N_7656,N_7525);
nor U8265 (N_8265,N_7676,N_7487);
nand U8266 (N_8266,N_7485,N_7320);
or U8267 (N_8267,N_7513,N_7121);
and U8268 (N_8268,N_7847,N_7052);
nor U8269 (N_8269,N_7262,N_7727);
nand U8270 (N_8270,N_7776,N_7680);
or U8271 (N_8271,N_7834,N_7041);
nor U8272 (N_8272,N_7111,N_7760);
nor U8273 (N_8273,N_7572,N_7692);
or U8274 (N_8274,N_7414,N_7490);
nor U8275 (N_8275,N_7477,N_7251);
nor U8276 (N_8276,N_7318,N_7347);
nand U8277 (N_8277,N_7933,N_7901);
nand U8278 (N_8278,N_7553,N_7980);
nor U8279 (N_8279,N_7828,N_7314);
xnor U8280 (N_8280,N_7763,N_7360);
or U8281 (N_8281,N_7899,N_7871);
or U8282 (N_8282,N_7438,N_7342);
and U8283 (N_8283,N_7886,N_7630);
nor U8284 (N_8284,N_7913,N_7588);
nor U8285 (N_8285,N_7782,N_7503);
or U8286 (N_8286,N_7914,N_7091);
nor U8287 (N_8287,N_7417,N_7429);
and U8288 (N_8288,N_7608,N_7180);
xor U8289 (N_8289,N_7800,N_7445);
nor U8290 (N_8290,N_7747,N_7234);
xnor U8291 (N_8291,N_7033,N_7599);
nor U8292 (N_8292,N_7950,N_7032);
or U8293 (N_8293,N_7730,N_7344);
or U8294 (N_8294,N_7305,N_7885);
nor U8295 (N_8295,N_7724,N_7090);
and U8296 (N_8296,N_7552,N_7159);
and U8297 (N_8297,N_7356,N_7096);
nand U8298 (N_8298,N_7332,N_7825);
and U8299 (N_8299,N_7670,N_7941);
nor U8300 (N_8300,N_7265,N_7773);
nor U8301 (N_8301,N_7848,N_7781);
or U8302 (N_8302,N_7749,N_7578);
nor U8303 (N_8303,N_7736,N_7486);
and U8304 (N_8304,N_7811,N_7126);
or U8305 (N_8305,N_7459,N_7285);
or U8306 (N_8306,N_7171,N_7779);
and U8307 (N_8307,N_7416,N_7115);
or U8308 (N_8308,N_7840,N_7557);
and U8309 (N_8309,N_7888,N_7045);
nor U8310 (N_8310,N_7231,N_7431);
nor U8311 (N_8311,N_7348,N_7202);
nand U8312 (N_8312,N_7904,N_7829);
nor U8313 (N_8313,N_7947,N_7102);
nand U8314 (N_8314,N_7255,N_7861);
and U8315 (N_8315,N_7512,N_7322);
or U8316 (N_8316,N_7030,N_7169);
or U8317 (N_8317,N_7517,N_7024);
nand U8318 (N_8318,N_7534,N_7506);
nor U8319 (N_8319,N_7114,N_7577);
xnor U8320 (N_8320,N_7463,N_7468);
nor U8321 (N_8321,N_7368,N_7437);
and U8322 (N_8322,N_7615,N_7915);
nor U8323 (N_8323,N_7204,N_7187);
xnor U8324 (N_8324,N_7858,N_7376);
and U8325 (N_8325,N_7127,N_7044);
or U8326 (N_8326,N_7786,N_7108);
nor U8327 (N_8327,N_7099,N_7769);
or U8328 (N_8328,N_7624,N_7675);
and U8329 (N_8329,N_7815,N_7056);
nand U8330 (N_8330,N_7791,N_7981);
or U8331 (N_8331,N_7726,N_7945);
and U8332 (N_8332,N_7213,N_7378);
xnor U8333 (N_8333,N_7048,N_7540);
xnor U8334 (N_8334,N_7458,N_7565);
nand U8335 (N_8335,N_7201,N_7777);
and U8336 (N_8336,N_7986,N_7844);
or U8337 (N_8337,N_7188,N_7012);
or U8338 (N_8338,N_7059,N_7275);
nor U8339 (N_8339,N_7614,N_7592);
or U8340 (N_8340,N_7563,N_7384);
nand U8341 (N_8341,N_7034,N_7688);
nor U8342 (N_8342,N_7973,N_7772);
nand U8343 (N_8343,N_7193,N_7321);
nand U8344 (N_8344,N_7931,N_7788);
or U8345 (N_8345,N_7874,N_7785);
and U8346 (N_8346,N_7109,N_7740);
and U8347 (N_8347,N_7780,N_7340);
nand U8348 (N_8348,N_7600,N_7556);
nor U8349 (N_8349,N_7974,N_7301);
nor U8350 (N_8350,N_7107,N_7155);
nand U8351 (N_8351,N_7483,N_7471);
nand U8352 (N_8352,N_7018,N_7089);
and U8353 (N_8353,N_7595,N_7805);
nor U8354 (N_8354,N_7611,N_7147);
or U8355 (N_8355,N_7666,N_7082);
nand U8356 (N_8356,N_7088,N_7000);
xor U8357 (N_8357,N_7764,N_7218);
nand U8358 (N_8358,N_7448,N_7853);
and U8359 (N_8359,N_7403,N_7558);
and U8360 (N_8360,N_7966,N_7678);
and U8361 (N_8361,N_7258,N_7050);
and U8362 (N_8362,N_7539,N_7728);
or U8363 (N_8363,N_7882,N_7156);
or U8364 (N_8364,N_7796,N_7083);
nand U8365 (N_8365,N_7404,N_7761);
and U8366 (N_8366,N_7004,N_7518);
and U8367 (N_8367,N_7120,N_7297);
or U8368 (N_8368,N_7548,N_7288);
or U8369 (N_8369,N_7686,N_7766);
and U8370 (N_8370,N_7237,N_7794);
and U8371 (N_8371,N_7482,N_7895);
nand U8372 (N_8372,N_7355,N_7269);
nor U8373 (N_8373,N_7140,N_7435);
and U8374 (N_8374,N_7846,N_7383);
nor U8375 (N_8375,N_7597,N_7295);
or U8376 (N_8376,N_7988,N_7122);
nand U8377 (N_8377,N_7302,N_7639);
or U8378 (N_8378,N_7272,N_7010);
nand U8379 (N_8379,N_7326,N_7150);
and U8380 (N_8380,N_7856,N_7661);
or U8381 (N_8381,N_7478,N_7382);
xor U8382 (N_8382,N_7784,N_7116);
nor U8383 (N_8383,N_7464,N_7721);
and U8384 (N_8384,N_7959,N_7750);
and U8385 (N_8385,N_7076,N_7493);
or U8386 (N_8386,N_7824,N_7923);
or U8387 (N_8387,N_7331,N_7433);
or U8388 (N_8388,N_7137,N_7300);
nor U8389 (N_8389,N_7402,N_7949);
xnor U8390 (N_8390,N_7509,N_7963);
and U8391 (N_8391,N_7396,N_7814);
nor U8392 (N_8392,N_7298,N_7175);
or U8393 (N_8393,N_7660,N_7142);
or U8394 (N_8394,N_7536,N_7505);
nand U8395 (N_8395,N_7256,N_7955);
and U8396 (N_8396,N_7877,N_7039);
nor U8397 (N_8397,N_7343,N_7208);
and U8398 (N_8398,N_7165,N_7064);
or U8399 (N_8399,N_7713,N_7643);
nand U8400 (N_8400,N_7975,N_7665);
nand U8401 (N_8401,N_7637,N_7896);
and U8402 (N_8402,N_7677,N_7407);
and U8403 (N_8403,N_7965,N_7948);
and U8404 (N_8404,N_7526,N_7103);
or U8405 (N_8405,N_7524,N_7712);
and U8406 (N_8406,N_7999,N_7266);
and U8407 (N_8407,N_7290,N_7276);
or U8408 (N_8408,N_7447,N_7922);
xnor U8409 (N_8409,N_7026,N_7238);
and U8410 (N_8410,N_7649,N_7182);
and U8411 (N_8411,N_7514,N_7626);
xnor U8412 (N_8412,N_7069,N_7249);
nand U8413 (N_8413,N_7281,N_7436);
nand U8414 (N_8414,N_7568,N_7541);
nor U8415 (N_8415,N_7497,N_7628);
nand U8416 (N_8416,N_7808,N_7324);
nor U8417 (N_8417,N_7733,N_7296);
nand U8418 (N_8418,N_7544,N_7003);
and U8419 (N_8419,N_7757,N_7381);
nor U8420 (N_8420,N_7953,N_7411);
nand U8421 (N_8421,N_7804,N_7280);
and U8422 (N_8422,N_7702,N_7491);
nand U8423 (N_8423,N_7219,N_7181);
and U8424 (N_8424,N_7754,N_7124);
and U8425 (N_8425,N_7197,N_7642);
and U8426 (N_8426,N_7351,N_7716);
and U8427 (N_8427,N_7184,N_7605);
and U8428 (N_8428,N_7873,N_7333);
and U8429 (N_8429,N_7168,N_7775);
xnor U8430 (N_8430,N_7134,N_7422);
nor U8431 (N_8431,N_7698,N_7859);
or U8432 (N_8432,N_7528,N_7366);
nor U8433 (N_8433,N_7078,N_7074);
or U8434 (N_8434,N_7502,N_7801);
or U8435 (N_8435,N_7372,N_7720);
and U8436 (N_8436,N_7752,N_7043);
nand U8437 (N_8437,N_7767,N_7603);
nor U8438 (N_8438,N_7689,N_7917);
nor U8439 (N_8439,N_7133,N_7040);
or U8440 (N_8440,N_7646,N_7379);
or U8441 (N_8441,N_7354,N_7627);
and U8442 (N_8442,N_7427,N_7867);
or U8443 (N_8443,N_7648,N_7845);
or U8444 (N_8444,N_7177,N_7835);
or U8445 (N_8445,N_7617,N_7470);
xnor U8446 (N_8446,N_7023,N_7016);
nand U8447 (N_8447,N_7294,N_7144);
or U8448 (N_8448,N_7621,N_7149);
nor U8449 (N_8449,N_7968,N_7943);
and U8450 (N_8450,N_7878,N_7576);
nand U8451 (N_8451,N_7199,N_7891);
nor U8452 (N_8452,N_7148,N_7242);
or U8453 (N_8453,N_7005,N_7141);
or U8454 (N_8454,N_7330,N_7166);
nand U8455 (N_8455,N_7511,N_7870);
nor U8456 (N_8456,N_7479,N_7875);
nand U8457 (N_8457,N_7700,N_7062);
nor U8458 (N_8458,N_7545,N_7990);
nor U8459 (N_8459,N_7893,N_7865);
nor U8460 (N_8460,N_7267,N_7972);
or U8461 (N_8461,N_7792,N_7410);
or U8462 (N_8462,N_7145,N_7892);
nor U8463 (N_8463,N_7587,N_7833);
and U8464 (N_8464,N_7036,N_7810);
nand U8465 (N_8465,N_7068,N_7593);
nand U8466 (N_8466,N_7254,N_7862);
xor U8467 (N_8467,N_7774,N_7659);
and U8468 (N_8468,N_7031,N_7836);
and U8469 (N_8469,N_7926,N_7636);
xor U8470 (N_8470,N_7653,N_7987);
nor U8471 (N_8471,N_7994,N_7364);
nand U8472 (N_8472,N_7047,N_7978);
and U8473 (N_8473,N_7705,N_7598);
xor U8474 (N_8474,N_7499,N_7710);
nand U8475 (N_8475,N_7996,N_7428);
nand U8476 (N_8476,N_7271,N_7958);
xor U8477 (N_8477,N_7093,N_7881);
or U8478 (N_8478,N_7860,N_7287);
nand U8479 (N_8479,N_7629,N_7883);
xnor U8480 (N_8480,N_7622,N_7842);
or U8481 (N_8481,N_7510,N_7691);
nor U8482 (N_8482,N_7907,N_7370);
nor U8483 (N_8483,N_7327,N_7480);
and U8484 (N_8484,N_7820,N_7157);
or U8485 (N_8485,N_7995,N_7460);
and U8486 (N_8486,N_7543,N_7352);
nand U8487 (N_8487,N_7118,N_7492);
xnor U8488 (N_8488,N_7334,N_7632);
xnor U8489 (N_8489,N_7308,N_7194);
or U8490 (N_8490,N_7247,N_7001);
nand U8491 (N_8491,N_7021,N_7377);
or U8492 (N_8492,N_7085,N_7818);
xnor U8493 (N_8493,N_7663,N_7762);
nand U8494 (N_8494,N_7734,N_7055);
or U8495 (N_8495,N_7919,N_7745);
nor U8496 (N_8496,N_7027,N_7225);
or U8497 (N_8497,N_7060,N_7723);
nand U8498 (N_8498,N_7983,N_7879);
or U8499 (N_8499,N_7336,N_7982);
xnor U8500 (N_8500,N_7832,N_7315);
or U8501 (N_8501,N_7950,N_7946);
or U8502 (N_8502,N_7988,N_7347);
nand U8503 (N_8503,N_7688,N_7916);
nor U8504 (N_8504,N_7633,N_7218);
or U8505 (N_8505,N_7115,N_7846);
nor U8506 (N_8506,N_7836,N_7035);
nor U8507 (N_8507,N_7564,N_7819);
or U8508 (N_8508,N_7245,N_7992);
nor U8509 (N_8509,N_7467,N_7813);
xnor U8510 (N_8510,N_7818,N_7737);
nor U8511 (N_8511,N_7812,N_7500);
nand U8512 (N_8512,N_7262,N_7489);
nand U8513 (N_8513,N_7483,N_7170);
or U8514 (N_8514,N_7650,N_7848);
and U8515 (N_8515,N_7544,N_7434);
nand U8516 (N_8516,N_7620,N_7807);
and U8517 (N_8517,N_7105,N_7193);
nor U8518 (N_8518,N_7062,N_7786);
nand U8519 (N_8519,N_7318,N_7265);
nor U8520 (N_8520,N_7767,N_7223);
nor U8521 (N_8521,N_7298,N_7284);
nor U8522 (N_8522,N_7838,N_7017);
or U8523 (N_8523,N_7794,N_7095);
or U8524 (N_8524,N_7501,N_7252);
nand U8525 (N_8525,N_7696,N_7632);
and U8526 (N_8526,N_7304,N_7758);
nand U8527 (N_8527,N_7838,N_7822);
nor U8528 (N_8528,N_7862,N_7367);
and U8529 (N_8529,N_7334,N_7593);
xnor U8530 (N_8530,N_7375,N_7733);
and U8531 (N_8531,N_7524,N_7348);
and U8532 (N_8532,N_7366,N_7263);
or U8533 (N_8533,N_7966,N_7013);
nor U8534 (N_8534,N_7715,N_7374);
nor U8535 (N_8535,N_7050,N_7125);
and U8536 (N_8536,N_7458,N_7387);
and U8537 (N_8537,N_7858,N_7394);
nor U8538 (N_8538,N_7522,N_7250);
nor U8539 (N_8539,N_7504,N_7411);
nand U8540 (N_8540,N_7174,N_7514);
nor U8541 (N_8541,N_7959,N_7391);
or U8542 (N_8542,N_7781,N_7709);
or U8543 (N_8543,N_7800,N_7787);
and U8544 (N_8544,N_7673,N_7866);
and U8545 (N_8545,N_7863,N_7673);
nor U8546 (N_8546,N_7074,N_7719);
and U8547 (N_8547,N_7084,N_7099);
nor U8548 (N_8548,N_7561,N_7787);
or U8549 (N_8549,N_7178,N_7762);
and U8550 (N_8550,N_7042,N_7799);
or U8551 (N_8551,N_7545,N_7939);
nor U8552 (N_8552,N_7700,N_7626);
and U8553 (N_8553,N_7516,N_7974);
and U8554 (N_8554,N_7950,N_7757);
and U8555 (N_8555,N_7855,N_7804);
nand U8556 (N_8556,N_7290,N_7910);
nand U8557 (N_8557,N_7697,N_7054);
nand U8558 (N_8558,N_7692,N_7192);
or U8559 (N_8559,N_7555,N_7528);
nand U8560 (N_8560,N_7221,N_7919);
or U8561 (N_8561,N_7014,N_7660);
nand U8562 (N_8562,N_7500,N_7964);
nor U8563 (N_8563,N_7063,N_7630);
nand U8564 (N_8564,N_7748,N_7395);
and U8565 (N_8565,N_7504,N_7371);
and U8566 (N_8566,N_7993,N_7768);
or U8567 (N_8567,N_7130,N_7797);
nand U8568 (N_8568,N_7508,N_7835);
or U8569 (N_8569,N_7688,N_7412);
and U8570 (N_8570,N_7662,N_7265);
nor U8571 (N_8571,N_7264,N_7395);
nand U8572 (N_8572,N_7688,N_7741);
and U8573 (N_8573,N_7991,N_7982);
xnor U8574 (N_8574,N_7104,N_7098);
and U8575 (N_8575,N_7564,N_7612);
or U8576 (N_8576,N_7703,N_7523);
xnor U8577 (N_8577,N_7356,N_7798);
xor U8578 (N_8578,N_7763,N_7907);
xnor U8579 (N_8579,N_7989,N_7448);
and U8580 (N_8580,N_7164,N_7267);
nand U8581 (N_8581,N_7038,N_7296);
and U8582 (N_8582,N_7423,N_7947);
or U8583 (N_8583,N_7817,N_7739);
nand U8584 (N_8584,N_7090,N_7786);
and U8585 (N_8585,N_7326,N_7930);
and U8586 (N_8586,N_7510,N_7135);
nand U8587 (N_8587,N_7554,N_7916);
and U8588 (N_8588,N_7234,N_7764);
nor U8589 (N_8589,N_7306,N_7100);
nand U8590 (N_8590,N_7853,N_7937);
xor U8591 (N_8591,N_7160,N_7556);
or U8592 (N_8592,N_7356,N_7503);
and U8593 (N_8593,N_7156,N_7270);
nand U8594 (N_8594,N_7852,N_7303);
nor U8595 (N_8595,N_7266,N_7679);
or U8596 (N_8596,N_7206,N_7454);
nor U8597 (N_8597,N_7063,N_7068);
and U8598 (N_8598,N_7741,N_7217);
xnor U8599 (N_8599,N_7931,N_7619);
and U8600 (N_8600,N_7938,N_7179);
nand U8601 (N_8601,N_7188,N_7631);
or U8602 (N_8602,N_7373,N_7861);
nor U8603 (N_8603,N_7778,N_7617);
nor U8604 (N_8604,N_7145,N_7872);
nor U8605 (N_8605,N_7635,N_7661);
nor U8606 (N_8606,N_7321,N_7065);
and U8607 (N_8607,N_7757,N_7374);
nand U8608 (N_8608,N_7377,N_7897);
xor U8609 (N_8609,N_7334,N_7219);
xor U8610 (N_8610,N_7644,N_7278);
or U8611 (N_8611,N_7002,N_7866);
or U8612 (N_8612,N_7569,N_7516);
nor U8613 (N_8613,N_7450,N_7367);
xnor U8614 (N_8614,N_7708,N_7491);
nand U8615 (N_8615,N_7455,N_7944);
nand U8616 (N_8616,N_7704,N_7813);
nand U8617 (N_8617,N_7266,N_7819);
nor U8618 (N_8618,N_7911,N_7627);
and U8619 (N_8619,N_7312,N_7193);
nor U8620 (N_8620,N_7216,N_7384);
nand U8621 (N_8621,N_7791,N_7117);
xor U8622 (N_8622,N_7706,N_7406);
nor U8623 (N_8623,N_7485,N_7043);
nor U8624 (N_8624,N_7106,N_7074);
xnor U8625 (N_8625,N_7982,N_7469);
or U8626 (N_8626,N_7240,N_7339);
or U8627 (N_8627,N_7564,N_7887);
or U8628 (N_8628,N_7575,N_7447);
or U8629 (N_8629,N_7022,N_7899);
nand U8630 (N_8630,N_7740,N_7606);
or U8631 (N_8631,N_7350,N_7301);
nor U8632 (N_8632,N_7553,N_7247);
nor U8633 (N_8633,N_7168,N_7945);
and U8634 (N_8634,N_7917,N_7239);
nor U8635 (N_8635,N_7197,N_7203);
nand U8636 (N_8636,N_7954,N_7654);
nand U8637 (N_8637,N_7959,N_7559);
or U8638 (N_8638,N_7478,N_7788);
and U8639 (N_8639,N_7863,N_7528);
and U8640 (N_8640,N_7324,N_7556);
and U8641 (N_8641,N_7477,N_7719);
nor U8642 (N_8642,N_7252,N_7868);
nor U8643 (N_8643,N_7536,N_7446);
xnor U8644 (N_8644,N_7327,N_7239);
nand U8645 (N_8645,N_7327,N_7452);
and U8646 (N_8646,N_7395,N_7741);
and U8647 (N_8647,N_7880,N_7686);
or U8648 (N_8648,N_7960,N_7453);
nor U8649 (N_8649,N_7021,N_7708);
or U8650 (N_8650,N_7882,N_7988);
and U8651 (N_8651,N_7359,N_7362);
nand U8652 (N_8652,N_7515,N_7569);
or U8653 (N_8653,N_7395,N_7780);
nor U8654 (N_8654,N_7061,N_7035);
or U8655 (N_8655,N_7083,N_7285);
xnor U8656 (N_8656,N_7250,N_7299);
or U8657 (N_8657,N_7705,N_7361);
or U8658 (N_8658,N_7916,N_7967);
or U8659 (N_8659,N_7047,N_7548);
xor U8660 (N_8660,N_7811,N_7276);
and U8661 (N_8661,N_7307,N_7574);
or U8662 (N_8662,N_7969,N_7288);
or U8663 (N_8663,N_7452,N_7520);
nand U8664 (N_8664,N_7768,N_7621);
or U8665 (N_8665,N_7940,N_7441);
nand U8666 (N_8666,N_7883,N_7641);
nand U8667 (N_8667,N_7302,N_7013);
nor U8668 (N_8668,N_7601,N_7314);
nand U8669 (N_8669,N_7060,N_7110);
or U8670 (N_8670,N_7501,N_7311);
nand U8671 (N_8671,N_7756,N_7559);
nand U8672 (N_8672,N_7121,N_7368);
nor U8673 (N_8673,N_7820,N_7185);
xnor U8674 (N_8674,N_7257,N_7908);
or U8675 (N_8675,N_7768,N_7160);
nand U8676 (N_8676,N_7232,N_7498);
or U8677 (N_8677,N_7755,N_7340);
nand U8678 (N_8678,N_7271,N_7322);
nand U8679 (N_8679,N_7112,N_7057);
xnor U8680 (N_8680,N_7731,N_7240);
nand U8681 (N_8681,N_7905,N_7525);
or U8682 (N_8682,N_7352,N_7291);
or U8683 (N_8683,N_7531,N_7205);
and U8684 (N_8684,N_7582,N_7157);
nand U8685 (N_8685,N_7970,N_7624);
nand U8686 (N_8686,N_7621,N_7080);
and U8687 (N_8687,N_7461,N_7599);
nor U8688 (N_8688,N_7744,N_7406);
or U8689 (N_8689,N_7492,N_7369);
nor U8690 (N_8690,N_7366,N_7926);
or U8691 (N_8691,N_7705,N_7009);
nand U8692 (N_8692,N_7428,N_7954);
nor U8693 (N_8693,N_7733,N_7328);
or U8694 (N_8694,N_7583,N_7442);
and U8695 (N_8695,N_7824,N_7405);
and U8696 (N_8696,N_7546,N_7685);
and U8697 (N_8697,N_7483,N_7891);
nand U8698 (N_8698,N_7918,N_7275);
and U8699 (N_8699,N_7864,N_7901);
nor U8700 (N_8700,N_7056,N_7181);
nor U8701 (N_8701,N_7334,N_7793);
nand U8702 (N_8702,N_7925,N_7489);
nand U8703 (N_8703,N_7942,N_7667);
nor U8704 (N_8704,N_7476,N_7562);
nor U8705 (N_8705,N_7029,N_7341);
or U8706 (N_8706,N_7980,N_7685);
and U8707 (N_8707,N_7870,N_7824);
or U8708 (N_8708,N_7785,N_7032);
nand U8709 (N_8709,N_7368,N_7671);
nand U8710 (N_8710,N_7178,N_7798);
nand U8711 (N_8711,N_7631,N_7442);
nand U8712 (N_8712,N_7395,N_7630);
nand U8713 (N_8713,N_7432,N_7177);
nand U8714 (N_8714,N_7157,N_7423);
or U8715 (N_8715,N_7946,N_7555);
and U8716 (N_8716,N_7967,N_7177);
or U8717 (N_8717,N_7878,N_7563);
nor U8718 (N_8718,N_7492,N_7678);
and U8719 (N_8719,N_7675,N_7899);
nor U8720 (N_8720,N_7148,N_7642);
and U8721 (N_8721,N_7057,N_7337);
xor U8722 (N_8722,N_7965,N_7327);
nand U8723 (N_8723,N_7430,N_7830);
or U8724 (N_8724,N_7344,N_7199);
or U8725 (N_8725,N_7203,N_7693);
nor U8726 (N_8726,N_7691,N_7597);
or U8727 (N_8727,N_7242,N_7893);
nand U8728 (N_8728,N_7019,N_7809);
and U8729 (N_8729,N_7359,N_7298);
or U8730 (N_8730,N_7897,N_7581);
xnor U8731 (N_8731,N_7352,N_7580);
or U8732 (N_8732,N_7898,N_7304);
nor U8733 (N_8733,N_7273,N_7844);
nand U8734 (N_8734,N_7273,N_7855);
nor U8735 (N_8735,N_7074,N_7790);
nand U8736 (N_8736,N_7578,N_7865);
nor U8737 (N_8737,N_7212,N_7481);
nand U8738 (N_8738,N_7374,N_7547);
and U8739 (N_8739,N_7975,N_7035);
nand U8740 (N_8740,N_7380,N_7599);
xnor U8741 (N_8741,N_7590,N_7593);
nand U8742 (N_8742,N_7191,N_7797);
and U8743 (N_8743,N_7409,N_7172);
nand U8744 (N_8744,N_7452,N_7831);
and U8745 (N_8745,N_7849,N_7312);
and U8746 (N_8746,N_7396,N_7884);
and U8747 (N_8747,N_7361,N_7737);
or U8748 (N_8748,N_7555,N_7307);
nand U8749 (N_8749,N_7565,N_7039);
nor U8750 (N_8750,N_7932,N_7654);
nand U8751 (N_8751,N_7999,N_7642);
and U8752 (N_8752,N_7985,N_7155);
and U8753 (N_8753,N_7592,N_7507);
nor U8754 (N_8754,N_7802,N_7623);
xnor U8755 (N_8755,N_7429,N_7224);
nand U8756 (N_8756,N_7042,N_7770);
and U8757 (N_8757,N_7006,N_7130);
and U8758 (N_8758,N_7080,N_7136);
nor U8759 (N_8759,N_7040,N_7890);
xor U8760 (N_8760,N_7898,N_7053);
nor U8761 (N_8761,N_7865,N_7575);
and U8762 (N_8762,N_7166,N_7337);
and U8763 (N_8763,N_7897,N_7945);
nand U8764 (N_8764,N_7608,N_7789);
or U8765 (N_8765,N_7431,N_7901);
or U8766 (N_8766,N_7463,N_7435);
or U8767 (N_8767,N_7550,N_7800);
xor U8768 (N_8768,N_7741,N_7238);
and U8769 (N_8769,N_7712,N_7927);
nand U8770 (N_8770,N_7831,N_7614);
xor U8771 (N_8771,N_7261,N_7169);
nor U8772 (N_8772,N_7677,N_7399);
or U8773 (N_8773,N_7148,N_7266);
and U8774 (N_8774,N_7719,N_7544);
or U8775 (N_8775,N_7630,N_7066);
nand U8776 (N_8776,N_7933,N_7252);
nand U8777 (N_8777,N_7367,N_7683);
nor U8778 (N_8778,N_7156,N_7391);
or U8779 (N_8779,N_7654,N_7603);
and U8780 (N_8780,N_7395,N_7632);
nand U8781 (N_8781,N_7848,N_7428);
nand U8782 (N_8782,N_7513,N_7088);
nand U8783 (N_8783,N_7634,N_7828);
or U8784 (N_8784,N_7612,N_7951);
nand U8785 (N_8785,N_7821,N_7218);
nand U8786 (N_8786,N_7992,N_7074);
or U8787 (N_8787,N_7685,N_7882);
nand U8788 (N_8788,N_7996,N_7462);
xor U8789 (N_8789,N_7242,N_7006);
nor U8790 (N_8790,N_7177,N_7950);
xnor U8791 (N_8791,N_7855,N_7830);
xor U8792 (N_8792,N_7128,N_7984);
xnor U8793 (N_8793,N_7913,N_7401);
nand U8794 (N_8794,N_7028,N_7917);
nor U8795 (N_8795,N_7123,N_7712);
nor U8796 (N_8796,N_7771,N_7764);
or U8797 (N_8797,N_7465,N_7593);
nor U8798 (N_8798,N_7318,N_7290);
and U8799 (N_8799,N_7989,N_7888);
and U8800 (N_8800,N_7766,N_7536);
or U8801 (N_8801,N_7566,N_7289);
and U8802 (N_8802,N_7456,N_7271);
nand U8803 (N_8803,N_7262,N_7956);
xnor U8804 (N_8804,N_7725,N_7172);
xor U8805 (N_8805,N_7286,N_7642);
and U8806 (N_8806,N_7526,N_7279);
xnor U8807 (N_8807,N_7759,N_7964);
or U8808 (N_8808,N_7585,N_7126);
and U8809 (N_8809,N_7173,N_7251);
nor U8810 (N_8810,N_7950,N_7307);
nand U8811 (N_8811,N_7877,N_7929);
nor U8812 (N_8812,N_7093,N_7455);
nor U8813 (N_8813,N_7035,N_7786);
nor U8814 (N_8814,N_7409,N_7830);
xnor U8815 (N_8815,N_7882,N_7922);
and U8816 (N_8816,N_7855,N_7191);
nand U8817 (N_8817,N_7361,N_7398);
nor U8818 (N_8818,N_7438,N_7110);
nor U8819 (N_8819,N_7415,N_7013);
or U8820 (N_8820,N_7362,N_7474);
and U8821 (N_8821,N_7130,N_7598);
nor U8822 (N_8822,N_7329,N_7481);
or U8823 (N_8823,N_7489,N_7480);
and U8824 (N_8824,N_7142,N_7551);
nor U8825 (N_8825,N_7057,N_7816);
nand U8826 (N_8826,N_7439,N_7703);
nor U8827 (N_8827,N_7480,N_7855);
nand U8828 (N_8828,N_7169,N_7615);
nand U8829 (N_8829,N_7279,N_7451);
xor U8830 (N_8830,N_7318,N_7534);
and U8831 (N_8831,N_7494,N_7698);
or U8832 (N_8832,N_7595,N_7829);
nor U8833 (N_8833,N_7508,N_7965);
or U8834 (N_8834,N_7203,N_7926);
nand U8835 (N_8835,N_7418,N_7805);
nor U8836 (N_8836,N_7968,N_7604);
and U8837 (N_8837,N_7534,N_7919);
nor U8838 (N_8838,N_7356,N_7305);
or U8839 (N_8839,N_7899,N_7811);
and U8840 (N_8840,N_7491,N_7663);
or U8841 (N_8841,N_7154,N_7514);
or U8842 (N_8842,N_7556,N_7843);
nand U8843 (N_8843,N_7566,N_7772);
nand U8844 (N_8844,N_7020,N_7864);
nand U8845 (N_8845,N_7624,N_7285);
xor U8846 (N_8846,N_7346,N_7443);
or U8847 (N_8847,N_7495,N_7752);
and U8848 (N_8848,N_7389,N_7076);
and U8849 (N_8849,N_7240,N_7424);
nand U8850 (N_8850,N_7218,N_7231);
xnor U8851 (N_8851,N_7719,N_7247);
xor U8852 (N_8852,N_7828,N_7039);
or U8853 (N_8853,N_7445,N_7040);
and U8854 (N_8854,N_7523,N_7739);
and U8855 (N_8855,N_7287,N_7541);
and U8856 (N_8856,N_7804,N_7267);
or U8857 (N_8857,N_7841,N_7418);
or U8858 (N_8858,N_7978,N_7471);
and U8859 (N_8859,N_7449,N_7330);
xor U8860 (N_8860,N_7454,N_7706);
nor U8861 (N_8861,N_7784,N_7030);
nor U8862 (N_8862,N_7751,N_7718);
nor U8863 (N_8863,N_7011,N_7193);
or U8864 (N_8864,N_7087,N_7979);
or U8865 (N_8865,N_7465,N_7749);
and U8866 (N_8866,N_7482,N_7016);
or U8867 (N_8867,N_7725,N_7902);
nand U8868 (N_8868,N_7534,N_7770);
nor U8869 (N_8869,N_7236,N_7988);
nand U8870 (N_8870,N_7516,N_7211);
nor U8871 (N_8871,N_7512,N_7704);
nand U8872 (N_8872,N_7450,N_7804);
and U8873 (N_8873,N_7507,N_7364);
and U8874 (N_8874,N_7308,N_7255);
nand U8875 (N_8875,N_7493,N_7366);
nand U8876 (N_8876,N_7982,N_7196);
nor U8877 (N_8877,N_7169,N_7563);
or U8878 (N_8878,N_7881,N_7984);
nand U8879 (N_8879,N_7094,N_7890);
or U8880 (N_8880,N_7987,N_7580);
and U8881 (N_8881,N_7531,N_7368);
xor U8882 (N_8882,N_7122,N_7180);
or U8883 (N_8883,N_7521,N_7473);
nand U8884 (N_8884,N_7126,N_7460);
nor U8885 (N_8885,N_7293,N_7369);
or U8886 (N_8886,N_7107,N_7684);
and U8887 (N_8887,N_7774,N_7933);
or U8888 (N_8888,N_7223,N_7252);
xor U8889 (N_8889,N_7337,N_7523);
or U8890 (N_8890,N_7977,N_7585);
nor U8891 (N_8891,N_7143,N_7760);
nand U8892 (N_8892,N_7923,N_7436);
nand U8893 (N_8893,N_7319,N_7501);
nand U8894 (N_8894,N_7982,N_7214);
or U8895 (N_8895,N_7819,N_7615);
and U8896 (N_8896,N_7777,N_7269);
nand U8897 (N_8897,N_7459,N_7833);
nor U8898 (N_8898,N_7412,N_7505);
and U8899 (N_8899,N_7010,N_7148);
or U8900 (N_8900,N_7037,N_7524);
xor U8901 (N_8901,N_7901,N_7203);
xnor U8902 (N_8902,N_7879,N_7464);
nor U8903 (N_8903,N_7609,N_7435);
and U8904 (N_8904,N_7093,N_7867);
and U8905 (N_8905,N_7994,N_7837);
nor U8906 (N_8906,N_7164,N_7942);
or U8907 (N_8907,N_7153,N_7200);
or U8908 (N_8908,N_7597,N_7748);
nand U8909 (N_8909,N_7738,N_7140);
or U8910 (N_8910,N_7991,N_7195);
nand U8911 (N_8911,N_7525,N_7256);
or U8912 (N_8912,N_7642,N_7003);
or U8913 (N_8913,N_7813,N_7471);
and U8914 (N_8914,N_7237,N_7375);
nand U8915 (N_8915,N_7951,N_7808);
nand U8916 (N_8916,N_7294,N_7407);
nand U8917 (N_8917,N_7809,N_7783);
nand U8918 (N_8918,N_7133,N_7768);
nand U8919 (N_8919,N_7578,N_7834);
xor U8920 (N_8920,N_7747,N_7513);
and U8921 (N_8921,N_7051,N_7918);
or U8922 (N_8922,N_7949,N_7342);
xnor U8923 (N_8923,N_7744,N_7028);
or U8924 (N_8924,N_7729,N_7607);
or U8925 (N_8925,N_7139,N_7363);
or U8926 (N_8926,N_7322,N_7350);
and U8927 (N_8927,N_7559,N_7260);
nor U8928 (N_8928,N_7579,N_7509);
nor U8929 (N_8929,N_7209,N_7485);
or U8930 (N_8930,N_7852,N_7501);
nand U8931 (N_8931,N_7119,N_7968);
xor U8932 (N_8932,N_7570,N_7942);
and U8933 (N_8933,N_7841,N_7856);
nand U8934 (N_8934,N_7014,N_7010);
nand U8935 (N_8935,N_7138,N_7728);
and U8936 (N_8936,N_7876,N_7699);
nor U8937 (N_8937,N_7597,N_7457);
and U8938 (N_8938,N_7388,N_7263);
and U8939 (N_8939,N_7289,N_7219);
or U8940 (N_8940,N_7268,N_7663);
or U8941 (N_8941,N_7326,N_7783);
nand U8942 (N_8942,N_7937,N_7274);
and U8943 (N_8943,N_7407,N_7992);
nor U8944 (N_8944,N_7013,N_7853);
xnor U8945 (N_8945,N_7879,N_7688);
and U8946 (N_8946,N_7071,N_7657);
and U8947 (N_8947,N_7346,N_7130);
or U8948 (N_8948,N_7223,N_7871);
nor U8949 (N_8949,N_7968,N_7443);
and U8950 (N_8950,N_7428,N_7617);
or U8951 (N_8951,N_7407,N_7626);
or U8952 (N_8952,N_7413,N_7515);
nor U8953 (N_8953,N_7904,N_7510);
or U8954 (N_8954,N_7510,N_7809);
nor U8955 (N_8955,N_7581,N_7283);
nor U8956 (N_8956,N_7421,N_7576);
nor U8957 (N_8957,N_7190,N_7761);
or U8958 (N_8958,N_7677,N_7379);
and U8959 (N_8959,N_7910,N_7357);
nor U8960 (N_8960,N_7601,N_7939);
xor U8961 (N_8961,N_7318,N_7921);
or U8962 (N_8962,N_7046,N_7476);
and U8963 (N_8963,N_7600,N_7964);
and U8964 (N_8964,N_7905,N_7029);
nor U8965 (N_8965,N_7203,N_7768);
and U8966 (N_8966,N_7661,N_7170);
nor U8967 (N_8967,N_7944,N_7274);
and U8968 (N_8968,N_7918,N_7243);
and U8969 (N_8969,N_7886,N_7318);
and U8970 (N_8970,N_7649,N_7660);
nor U8971 (N_8971,N_7029,N_7992);
and U8972 (N_8972,N_7653,N_7028);
xnor U8973 (N_8973,N_7704,N_7667);
xor U8974 (N_8974,N_7643,N_7128);
or U8975 (N_8975,N_7174,N_7119);
nor U8976 (N_8976,N_7004,N_7729);
nand U8977 (N_8977,N_7782,N_7421);
nand U8978 (N_8978,N_7142,N_7024);
nor U8979 (N_8979,N_7322,N_7454);
nor U8980 (N_8980,N_7214,N_7691);
or U8981 (N_8981,N_7339,N_7392);
and U8982 (N_8982,N_7537,N_7121);
nand U8983 (N_8983,N_7082,N_7782);
nand U8984 (N_8984,N_7511,N_7916);
or U8985 (N_8985,N_7704,N_7218);
xor U8986 (N_8986,N_7439,N_7101);
nand U8987 (N_8987,N_7276,N_7765);
nor U8988 (N_8988,N_7823,N_7154);
nand U8989 (N_8989,N_7860,N_7395);
nor U8990 (N_8990,N_7082,N_7146);
nor U8991 (N_8991,N_7538,N_7582);
xor U8992 (N_8992,N_7865,N_7240);
or U8993 (N_8993,N_7248,N_7530);
nand U8994 (N_8994,N_7340,N_7307);
xor U8995 (N_8995,N_7803,N_7414);
and U8996 (N_8996,N_7342,N_7548);
nand U8997 (N_8997,N_7556,N_7995);
nor U8998 (N_8998,N_7989,N_7512);
nor U8999 (N_8999,N_7379,N_7428);
nand U9000 (N_9000,N_8724,N_8301);
xor U9001 (N_9001,N_8131,N_8084);
and U9002 (N_9002,N_8233,N_8272);
nand U9003 (N_9003,N_8840,N_8576);
or U9004 (N_9004,N_8254,N_8302);
nand U9005 (N_9005,N_8628,N_8988);
or U9006 (N_9006,N_8113,N_8954);
and U9007 (N_9007,N_8128,N_8098);
nor U9008 (N_9008,N_8490,N_8127);
and U9009 (N_9009,N_8832,N_8803);
xor U9010 (N_9010,N_8120,N_8141);
nor U9011 (N_9011,N_8067,N_8242);
nor U9012 (N_9012,N_8647,N_8294);
or U9013 (N_9013,N_8050,N_8462);
or U9014 (N_9014,N_8432,N_8826);
nand U9015 (N_9015,N_8425,N_8664);
or U9016 (N_9016,N_8444,N_8018);
xnor U9017 (N_9017,N_8718,N_8884);
or U9018 (N_9018,N_8489,N_8415);
nand U9019 (N_9019,N_8096,N_8101);
xor U9020 (N_9020,N_8692,N_8963);
xor U9021 (N_9021,N_8093,N_8971);
or U9022 (N_9022,N_8277,N_8321);
xor U9023 (N_9023,N_8017,N_8904);
xor U9024 (N_9024,N_8267,N_8269);
nor U9025 (N_9025,N_8465,N_8781);
and U9026 (N_9026,N_8195,N_8706);
nand U9027 (N_9027,N_8477,N_8299);
and U9028 (N_9028,N_8183,N_8232);
nand U9029 (N_9029,N_8944,N_8332);
nand U9030 (N_9030,N_8069,N_8589);
nor U9031 (N_9031,N_8333,N_8567);
nor U9032 (N_9032,N_8116,N_8328);
nand U9033 (N_9033,N_8418,N_8699);
and U9034 (N_9034,N_8820,N_8932);
nand U9035 (N_9035,N_8063,N_8870);
and U9036 (N_9036,N_8822,N_8685);
and U9037 (N_9037,N_8539,N_8819);
or U9038 (N_9038,N_8633,N_8732);
nand U9039 (N_9039,N_8914,N_8420);
or U9040 (N_9040,N_8105,N_8981);
or U9041 (N_9041,N_8719,N_8390);
and U9042 (N_9042,N_8160,N_8640);
and U9043 (N_9043,N_8615,N_8734);
nor U9044 (N_9044,N_8513,N_8920);
nand U9045 (N_9045,N_8305,N_8036);
nor U9046 (N_9046,N_8227,N_8872);
nand U9047 (N_9047,N_8869,N_8824);
nor U9048 (N_9048,N_8491,N_8799);
or U9049 (N_9049,N_8853,N_8358);
or U9050 (N_9050,N_8857,N_8748);
nand U9051 (N_9051,N_8148,N_8025);
or U9052 (N_9052,N_8038,N_8823);
and U9053 (N_9053,N_8902,N_8114);
or U9054 (N_9054,N_8049,N_8130);
and U9055 (N_9055,N_8778,N_8780);
or U9056 (N_9056,N_8617,N_8528);
and U9057 (N_9057,N_8897,N_8946);
or U9058 (N_9058,N_8596,N_8112);
nor U9059 (N_9059,N_8802,N_8094);
nor U9060 (N_9060,N_8608,N_8634);
or U9061 (N_9061,N_8953,N_8636);
or U9062 (N_9062,N_8968,N_8205);
xor U9063 (N_9063,N_8509,N_8313);
and U9064 (N_9064,N_8379,N_8385);
nor U9065 (N_9065,N_8405,N_8683);
xor U9066 (N_9066,N_8259,N_8976);
nand U9067 (N_9067,N_8249,N_8695);
and U9068 (N_9068,N_8179,N_8855);
and U9069 (N_9069,N_8330,N_8276);
nand U9070 (N_9070,N_8404,N_8532);
nor U9071 (N_9071,N_8403,N_8408);
or U9072 (N_9072,N_8849,N_8806);
nand U9073 (N_9073,N_8739,N_8854);
and U9074 (N_9074,N_8212,N_8893);
xor U9075 (N_9075,N_8681,N_8978);
nand U9076 (N_9076,N_8879,N_8607);
xor U9077 (N_9077,N_8810,N_8220);
or U9078 (N_9078,N_8392,N_8829);
and U9079 (N_9079,N_8632,N_8587);
nor U9080 (N_9080,N_8339,N_8429);
or U9081 (N_9081,N_8537,N_8980);
xor U9082 (N_9082,N_8317,N_8871);
xor U9083 (N_9083,N_8603,N_8037);
nor U9084 (N_9084,N_8574,N_8478);
nor U9085 (N_9085,N_8203,N_8624);
nand U9086 (N_9086,N_8035,N_8271);
or U9087 (N_9087,N_8888,N_8224);
or U9088 (N_9088,N_8763,N_8002);
nand U9089 (N_9089,N_8828,N_8554);
and U9090 (N_9090,N_8670,N_8848);
and U9091 (N_9091,N_8200,N_8785);
nor U9092 (N_9092,N_8700,N_8423);
nand U9093 (N_9093,N_8174,N_8264);
xor U9094 (N_9094,N_8899,N_8514);
or U9095 (N_9095,N_8629,N_8645);
and U9096 (N_9096,N_8436,N_8644);
and U9097 (N_9097,N_8553,N_8656);
xnor U9098 (N_9098,N_8565,N_8875);
and U9099 (N_9099,N_8312,N_8484);
and U9100 (N_9100,N_8266,N_8606);
or U9101 (N_9101,N_8421,N_8937);
or U9102 (N_9102,N_8246,N_8667);
xor U9103 (N_9103,N_8336,N_8865);
or U9104 (N_9104,N_8597,N_8862);
and U9105 (N_9105,N_8412,N_8908);
nor U9106 (N_9106,N_8440,N_8046);
and U9107 (N_9107,N_8091,N_8760);
nor U9108 (N_9108,N_8164,N_8235);
and U9109 (N_9109,N_8986,N_8204);
nand U9110 (N_9110,N_8997,N_8754);
nand U9111 (N_9111,N_8262,N_8238);
nor U9112 (N_9112,N_8199,N_8001);
nor U9113 (N_9113,N_8221,N_8279);
xnor U9114 (N_9114,N_8078,N_8555);
xnor U9115 (N_9115,N_8809,N_8163);
nor U9116 (N_9116,N_8165,N_8004);
and U9117 (N_9117,N_8327,N_8614);
nand U9118 (N_9118,N_8516,N_8438);
nor U9119 (N_9119,N_8864,N_8969);
nand U9120 (N_9120,N_8329,N_8326);
nor U9121 (N_9121,N_8061,N_8373);
or U9122 (N_9122,N_8985,N_8007);
nand U9123 (N_9123,N_8703,N_8924);
nor U9124 (N_9124,N_8213,N_8592);
or U9125 (N_9125,N_8005,N_8668);
or U9126 (N_9126,N_8189,N_8601);
nand U9127 (N_9127,N_8657,N_8545);
and U9128 (N_9128,N_8320,N_8602);
or U9129 (N_9129,N_8411,N_8619);
nor U9130 (N_9130,N_8129,N_8375);
nand U9131 (N_9131,N_8184,N_8051);
or U9132 (N_9132,N_8878,N_8814);
and U9133 (N_9133,N_8581,N_8182);
xnor U9134 (N_9134,N_8586,N_8720);
nand U9135 (N_9135,N_8752,N_8466);
nor U9136 (N_9136,N_8475,N_8361);
or U9137 (N_9137,N_8225,N_8143);
nor U9138 (N_9138,N_8137,N_8881);
nor U9139 (N_9139,N_8074,N_8835);
nor U9140 (N_9140,N_8052,N_8994);
and U9141 (N_9141,N_8790,N_8398);
or U9142 (N_9142,N_8169,N_8082);
xnor U9143 (N_9143,N_8936,N_8604);
or U9144 (N_9144,N_8691,N_8198);
or U9145 (N_9145,N_8787,N_8281);
nand U9146 (N_9146,N_8653,N_8698);
or U9147 (N_9147,N_8898,N_8907);
or U9148 (N_9148,N_8298,N_8244);
or U9149 (N_9149,N_8060,N_8159);
nor U9150 (N_9150,N_8181,N_8337);
and U9151 (N_9151,N_8563,N_8216);
or U9152 (N_9152,N_8210,N_8955);
nor U9153 (N_9153,N_8939,N_8346);
xor U9154 (N_9154,N_8967,N_8335);
or U9155 (N_9155,N_8791,N_8630);
or U9156 (N_9156,N_8000,N_8192);
nor U9157 (N_9157,N_8560,N_8541);
nor U9158 (N_9158,N_8638,N_8610);
nor U9159 (N_9159,N_8795,N_8414);
and U9160 (N_9160,N_8838,N_8021);
and U9161 (N_9161,N_8982,N_8753);
nor U9162 (N_9162,N_8759,N_8697);
or U9163 (N_9163,N_8649,N_8496);
nand U9164 (N_9164,N_8931,N_8505);
and U9165 (N_9165,N_8122,N_8369);
and U9166 (N_9166,N_8304,N_8132);
or U9167 (N_9167,N_8776,N_8564);
nor U9168 (N_9168,N_8529,N_8257);
xnor U9169 (N_9169,N_8048,N_8077);
or U9170 (N_9170,N_8627,N_8419);
and U9171 (N_9171,N_8209,N_8679);
and U9172 (N_9172,N_8155,N_8139);
or U9173 (N_9173,N_8399,N_8726);
nor U9174 (N_9174,N_8289,N_8639);
or U9175 (N_9175,N_8087,N_8171);
and U9176 (N_9176,N_8502,N_8524);
or U9177 (N_9177,N_8504,N_8463);
nor U9178 (N_9178,N_8578,N_8166);
and U9179 (N_9179,N_8901,N_8641);
or U9180 (N_9180,N_8834,N_8621);
nor U9181 (N_9181,N_8825,N_8501);
or U9182 (N_9182,N_8508,N_8661);
nor U9183 (N_9183,N_8972,N_8599);
xnor U9184 (N_9184,N_8910,N_8686);
and U9185 (N_9185,N_8290,N_8815);
and U9186 (N_9186,N_8702,N_8652);
nor U9187 (N_9187,N_8400,N_8743);
nand U9188 (N_9188,N_8530,N_8883);
and U9189 (N_9189,N_8518,N_8676);
nand U9190 (N_9190,N_8758,N_8396);
nand U9191 (N_9191,N_8561,N_8559);
and U9192 (N_9192,N_8957,N_8300);
or U9193 (N_9193,N_8856,N_8125);
or U9194 (N_9194,N_8352,N_8359);
or U9195 (N_9195,N_8033,N_8890);
and U9196 (N_9196,N_8427,N_8880);
or U9197 (N_9197,N_8913,N_8250);
nand U9198 (N_9198,N_8572,N_8993);
nand U9199 (N_9199,N_8933,N_8041);
or U9200 (N_9200,N_8767,N_8251);
or U9201 (N_9201,N_8506,N_8377);
xnor U9202 (N_9202,N_8750,N_8273);
nand U9203 (N_9203,N_8102,N_8071);
or U9204 (N_9204,N_8180,N_8345);
or U9205 (N_9205,N_8595,N_8618);
or U9206 (N_9206,N_8673,N_8858);
or U9207 (N_9207,N_8136,N_8308);
nor U9208 (N_9208,N_8847,N_8557);
and U9209 (N_9209,N_8356,N_8547);
nand U9210 (N_9210,N_8922,N_8472);
nor U9211 (N_9211,N_8208,N_8694);
or U9212 (N_9212,N_8158,N_8594);
and U9213 (N_9213,N_8651,N_8022);
nor U9214 (N_9214,N_8845,N_8935);
or U9215 (N_9215,N_8492,N_8381);
nand U9216 (N_9216,N_8135,N_8316);
nor U9217 (N_9217,N_8534,N_8911);
nand U9218 (N_9218,N_8470,N_8995);
nor U9219 (N_9219,N_8844,N_8248);
or U9220 (N_9220,N_8133,N_8680);
or U9221 (N_9221,N_8556,N_8773);
nand U9222 (N_9222,N_8196,N_8830);
and U9223 (N_9223,N_8357,N_8783);
and U9224 (N_9224,N_8324,N_8010);
nand U9225 (N_9225,N_8925,N_8533);
and U9226 (N_9226,N_8860,N_8256);
xnor U9227 (N_9227,N_8916,N_8153);
nand U9228 (N_9228,N_8873,N_8771);
or U9229 (N_9229,N_8646,N_8265);
and U9230 (N_9230,N_8999,N_8798);
or U9231 (N_9231,N_8306,N_8605);
or U9232 (N_9232,N_8637,N_8735);
or U9233 (N_9233,N_8388,N_8696);
and U9234 (N_9234,N_8031,N_8095);
nor U9235 (N_9235,N_8811,N_8311);
and U9236 (N_9236,N_8437,N_8054);
and U9237 (N_9237,N_8274,N_8416);
xor U9238 (N_9238,N_8620,N_8030);
nor U9239 (N_9239,N_8512,N_8056);
nor U9240 (N_9240,N_8146,N_8149);
or U9241 (N_9241,N_8283,N_8894);
nand U9242 (N_9242,N_8546,N_8837);
or U9243 (N_9243,N_8401,N_8684);
and U9244 (N_9244,N_8613,N_8582);
nor U9245 (N_9245,N_8756,N_8040);
nand U9246 (N_9246,N_8191,N_8973);
or U9247 (N_9247,N_8253,N_8207);
nor U9248 (N_9248,N_8288,N_8019);
nor U9249 (N_9249,N_8882,N_8471);
and U9250 (N_9250,N_8917,N_8808);
or U9251 (N_9251,N_8923,N_8104);
or U9252 (N_9252,N_8454,N_8325);
nand U9253 (N_9253,N_8186,N_8903);
nor U9254 (N_9254,N_8012,N_8173);
nand U9255 (N_9255,N_8059,N_8579);
nand U9256 (N_9256,N_8941,N_8736);
nand U9257 (N_9257,N_8663,N_8503);
or U9258 (N_9258,N_8138,N_8229);
nand U9259 (N_9259,N_8459,N_8349);
nor U9260 (N_9260,N_8804,N_8678);
xnor U9261 (N_9261,N_8023,N_8293);
or U9262 (N_9262,N_8740,N_8194);
xor U9263 (N_9263,N_8751,N_8410);
xor U9264 (N_9264,N_8831,N_8762);
or U9265 (N_9265,N_8447,N_8658);
and U9266 (N_9266,N_8494,N_8201);
and U9267 (N_9267,N_8996,N_8360);
nor U9268 (N_9268,N_8397,N_8921);
nor U9269 (N_9269,N_8446,N_8406);
and U9270 (N_9270,N_8234,N_8374);
nand U9271 (N_9271,N_8521,N_8677);
and U9272 (N_9272,N_8722,N_8744);
or U9273 (N_9273,N_8765,N_8666);
xnor U9274 (N_9274,N_8073,N_8243);
nand U9275 (N_9275,N_8115,N_8738);
nand U9276 (N_9276,N_8100,N_8708);
nor U9277 (N_9277,N_8121,N_8479);
and U9278 (N_9278,N_8867,N_8669);
nor U9279 (N_9279,N_8409,N_8382);
or U9280 (N_9280,N_8662,N_8949);
and U9281 (N_9281,N_8443,N_8542);
or U9282 (N_9282,N_8842,N_8961);
nand U9283 (N_9283,N_8473,N_8584);
nor U9284 (N_9284,N_8876,N_8571);
nor U9285 (N_9285,N_8086,N_8552);
nand U9286 (N_9286,N_8928,N_8066);
xnor U9287 (N_9287,N_8107,N_8544);
or U9288 (N_9288,N_8426,N_8593);
and U9289 (N_9289,N_8309,N_8467);
or U9290 (N_9290,N_8495,N_8286);
xor U9291 (N_9291,N_8850,N_8688);
or U9292 (N_9292,N_8989,N_8717);
or U9293 (N_9293,N_8206,N_8185);
nor U9294 (N_9294,N_8642,N_8020);
nand U9295 (N_9295,N_8951,N_8631);
or U9296 (N_9296,N_8764,N_8103);
and U9297 (N_9297,N_8623,N_8682);
or U9298 (N_9298,N_8245,N_8892);
or U9299 (N_9299,N_8827,N_8746);
nor U9300 (N_9300,N_8731,N_8043);
nor U9301 (N_9301,N_8487,N_8024);
nand U9302 (N_9302,N_8769,N_8430);
nand U9303 (N_9303,N_8612,N_8081);
xor U9304 (N_9304,N_8085,N_8455);
or U9305 (N_9305,N_8261,N_8039);
and U9306 (N_9306,N_8236,N_8956);
and U9307 (N_9307,N_8057,N_8974);
nand U9308 (N_9308,N_8347,N_8715);
or U9309 (N_9309,N_8940,N_8109);
or U9310 (N_9310,N_8222,N_8193);
nor U9311 (N_9311,N_8451,N_8315);
and U9312 (N_9312,N_8351,N_8042);
or U9313 (N_9313,N_8600,N_8768);
xor U9314 (N_9314,N_8029,N_8517);
nand U9315 (N_9315,N_8519,N_8918);
or U9316 (N_9316,N_8583,N_8497);
nand U9317 (N_9317,N_8741,N_8372);
nor U9318 (N_9318,N_8926,N_8364);
nand U9319 (N_9319,N_8919,N_8895);
nor U9320 (N_9320,N_8877,N_8239);
nor U9321 (N_9321,N_8142,N_8453);
nand U9322 (N_9322,N_8747,N_8394);
nand U9323 (N_9323,N_8480,N_8167);
and U9324 (N_9324,N_8874,N_8818);
xor U9325 (N_9325,N_8090,N_8197);
or U9326 (N_9326,N_8045,N_8395);
nor U9327 (N_9327,N_8150,N_8340);
nand U9328 (N_9328,N_8793,N_8280);
or U9329 (N_9329,N_8111,N_8585);
nor U9330 (N_9330,N_8202,N_8745);
nand U9331 (N_9331,N_8891,N_8522);
xor U9332 (N_9332,N_8089,N_8027);
nor U9333 (N_9333,N_8498,N_8106);
nand U9334 (N_9334,N_8728,N_8157);
nand U9335 (N_9335,N_8687,N_8434);
and U9336 (N_9336,N_8341,N_8441);
nand U9337 (N_9337,N_8998,N_8255);
nand U9338 (N_9338,N_8543,N_8866);
nand U9339 (N_9339,N_8723,N_8424);
and U9340 (N_9340,N_8439,N_8761);
or U9341 (N_9341,N_8943,N_8588);
or U9342 (N_9342,N_8172,N_8044);
nand U9343 (N_9343,N_8151,N_8580);
nand U9344 (N_9344,N_8782,N_8168);
or U9345 (N_9345,N_8386,N_8500);
nand U9346 (N_9346,N_8757,N_8383);
nand U9347 (N_9347,N_8821,N_8570);
xnor U9348 (N_9348,N_8162,N_8977);
xnor U9349 (N_9349,N_8843,N_8535);
nor U9350 (N_9350,N_8648,N_8609);
nand U9351 (N_9351,N_8577,N_8674);
and U9352 (N_9352,N_8493,N_8772);
and U9353 (N_9353,N_8334,N_8712);
nand U9354 (N_9354,N_8070,N_8863);
and U9355 (N_9355,N_8292,N_8231);
or U9356 (N_9356,N_8770,N_8015);
or U9357 (N_9357,N_8468,N_8034);
nor U9358 (N_9358,N_8464,N_8729);
or U9359 (N_9359,N_8575,N_8991);
and U9360 (N_9360,N_8675,N_8749);
nand U9361 (N_9361,N_8062,N_8714);
nor U9362 (N_9362,N_8178,N_8384);
nand U9363 (N_9363,N_8900,N_8896);
or U9364 (N_9364,N_8170,N_8422);
nor U9365 (N_9365,N_8065,N_8626);
nor U9366 (N_9366,N_8515,N_8672);
and U9367 (N_9367,N_8282,N_8889);
xor U9368 (N_9368,N_8456,N_8727);
and U9369 (N_9369,N_8704,N_8389);
nor U9370 (N_9370,N_8481,N_8984);
nor U9371 (N_9371,N_8268,N_8285);
and U9372 (N_9372,N_8801,N_8523);
xor U9373 (N_9373,N_8322,N_8659);
and U9374 (N_9374,N_8655,N_8807);
and U9375 (N_9375,N_8887,N_8915);
nor U9376 (N_9376,N_8469,N_8970);
or U9377 (N_9377,N_8217,N_8912);
and U9378 (N_9378,N_8278,N_8363);
nor U9379 (N_9379,N_8449,N_8975);
nand U9380 (N_9380,N_8428,N_8448);
nor U9381 (N_9381,N_8526,N_8527);
xnor U9382 (N_9382,N_8156,N_8958);
nor U9383 (N_9383,N_8241,N_8635);
and U9384 (N_9384,N_8003,N_8014);
or U9385 (N_9385,N_8794,N_8611);
nand U9386 (N_9386,N_8140,N_8538);
or U9387 (N_9387,N_8906,N_8474);
nand U9388 (N_9388,N_8486,N_8413);
xnor U9389 (N_9389,N_8549,N_8028);
nor U9390 (N_9390,N_8435,N_8344);
and U9391 (N_9391,N_8777,N_8188);
nor U9392 (N_9392,N_8391,N_8551);
xor U9393 (N_9393,N_8145,N_8228);
and U9394 (N_9394,N_8983,N_8319);
or U9395 (N_9395,N_8079,N_8287);
nor U9396 (N_9396,N_8710,N_8929);
nand U9397 (N_9397,N_8488,N_8690);
and U9398 (N_9398,N_8177,N_8009);
nand U9399 (N_9399,N_8370,N_8548);
or U9400 (N_9400,N_8053,N_8591);
or U9401 (N_9401,N_8147,N_8625);
nor U9402 (N_9402,N_8431,N_8643);
xor U9403 (N_9403,N_8836,N_8800);
nor U9404 (N_9404,N_8992,N_8671);
or U9405 (N_9405,N_8450,N_8550);
and U9406 (N_9406,N_8839,N_8965);
or U9407 (N_9407,N_8457,N_8755);
nand U9408 (N_9408,N_8792,N_8118);
or U9409 (N_9409,N_8616,N_8353);
and U9410 (N_9410,N_8721,N_8307);
nand U9411 (N_9411,N_8144,N_8789);
nand U9412 (N_9412,N_8707,N_8716);
nor U9413 (N_9413,N_8725,N_8310);
or U9414 (N_9414,N_8942,N_8371);
xnor U9415 (N_9415,N_8076,N_8367);
xor U9416 (N_9416,N_8187,N_8569);
xor U9417 (N_9417,N_8342,N_8713);
or U9418 (N_9418,N_8247,N_8947);
or U9419 (N_9419,N_8507,N_8088);
nand U9420 (N_9420,N_8796,N_8846);
xnor U9421 (N_9421,N_8097,N_8622);
xnor U9422 (N_9422,N_8562,N_8226);
nand U9423 (N_9423,N_8766,N_8258);
and U9424 (N_9424,N_8152,N_8338);
and U9425 (N_9425,N_8362,N_8237);
nand U9426 (N_9426,N_8841,N_8499);
and U9427 (N_9427,N_8303,N_8786);
and U9428 (N_9428,N_8934,N_8055);
nand U9429 (N_9429,N_8263,N_8598);
and U9430 (N_9430,N_8011,N_8689);
nor U9431 (N_9431,N_8987,N_8366);
nand U9432 (N_9432,N_8909,N_8990);
or U9433 (N_9433,N_8816,N_8013);
or U9434 (N_9434,N_8083,N_8047);
or U9435 (N_9435,N_8458,N_8154);
and U9436 (N_9436,N_8960,N_8833);
nand U9437 (N_9437,N_8540,N_8123);
nand U9438 (N_9438,N_8064,N_8460);
nor U9439 (N_9439,N_8938,N_8343);
xor U9440 (N_9440,N_8817,N_8797);
or U9441 (N_9441,N_8775,N_8950);
nand U9442 (N_9442,N_8573,N_8510);
and U9443 (N_9443,N_8566,N_8959);
xnor U9444 (N_9444,N_8378,N_8805);
or U9445 (N_9445,N_8525,N_8117);
nor U9446 (N_9446,N_8511,N_8092);
or U9447 (N_9447,N_8110,N_8119);
nor U9448 (N_9448,N_8323,N_8665);
nor U9449 (N_9449,N_8442,N_8590);
nand U9450 (N_9450,N_8393,N_8223);
nor U9451 (N_9451,N_8214,N_8660);
or U9452 (N_9452,N_8861,N_8240);
nor U9453 (N_9453,N_8006,N_8784);
and U9454 (N_9454,N_8068,N_8930);
or U9455 (N_9455,N_8387,N_8402);
nor U9456 (N_9456,N_8260,N_8774);
and U9457 (N_9457,N_8124,N_8742);
xnor U9458 (N_9458,N_8558,N_8075);
or U9459 (N_9459,N_8482,N_8365);
or U9460 (N_9460,N_8134,N_8788);
and U9461 (N_9461,N_8927,N_8215);
nor U9462 (N_9462,N_8230,N_8886);
or U9463 (N_9463,N_8008,N_8350);
nor U9464 (N_9464,N_8072,N_8531);
nor U9465 (N_9465,N_8654,N_8693);
nor U9466 (N_9466,N_8711,N_8452);
or U9467 (N_9467,N_8417,N_8885);
xor U9468 (N_9468,N_8852,N_8945);
nand U9469 (N_9469,N_8032,N_8190);
or U9470 (N_9470,N_8080,N_8380);
and U9471 (N_9471,N_8016,N_8851);
and U9472 (N_9472,N_8219,N_8126);
or U9473 (N_9473,N_8314,N_8318);
or U9474 (N_9474,N_8099,N_8568);
nor U9475 (N_9475,N_8520,N_8709);
or U9476 (N_9476,N_8368,N_8176);
nand U9477 (N_9477,N_8859,N_8058);
nor U9478 (N_9478,N_8812,N_8733);
xnor U9479 (N_9479,N_8218,N_8813);
nor U9480 (N_9480,N_8966,N_8355);
or U9481 (N_9481,N_8445,N_8275);
nand U9482 (N_9482,N_8868,N_8211);
and U9483 (N_9483,N_8284,N_8331);
and U9484 (N_9484,N_8108,N_8297);
nor U9485 (N_9485,N_8964,N_8952);
and U9486 (N_9486,N_8376,N_8779);
and U9487 (N_9487,N_8650,N_8905);
and U9488 (N_9488,N_8705,N_8485);
nand U9489 (N_9489,N_8737,N_8175);
nand U9490 (N_9490,N_8433,N_8354);
and U9491 (N_9491,N_8536,N_8161);
nand U9492 (N_9492,N_8948,N_8296);
nor U9493 (N_9493,N_8026,N_8295);
or U9494 (N_9494,N_8348,N_8730);
nand U9495 (N_9495,N_8461,N_8407);
xnor U9496 (N_9496,N_8979,N_8962);
xnor U9497 (N_9497,N_8701,N_8476);
nor U9498 (N_9498,N_8291,N_8270);
nor U9499 (N_9499,N_8483,N_8252);
xnor U9500 (N_9500,N_8089,N_8734);
nand U9501 (N_9501,N_8585,N_8791);
nor U9502 (N_9502,N_8828,N_8480);
and U9503 (N_9503,N_8768,N_8609);
nand U9504 (N_9504,N_8472,N_8295);
and U9505 (N_9505,N_8065,N_8376);
xnor U9506 (N_9506,N_8032,N_8247);
nor U9507 (N_9507,N_8562,N_8601);
nand U9508 (N_9508,N_8267,N_8044);
nand U9509 (N_9509,N_8247,N_8618);
nand U9510 (N_9510,N_8921,N_8362);
nand U9511 (N_9511,N_8085,N_8811);
or U9512 (N_9512,N_8088,N_8484);
or U9513 (N_9513,N_8312,N_8697);
or U9514 (N_9514,N_8227,N_8169);
and U9515 (N_9515,N_8624,N_8023);
or U9516 (N_9516,N_8853,N_8778);
and U9517 (N_9517,N_8382,N_8903);
nand U9518 (N_9518,N_8695,N_8672);
nand U9519 (N_9519,N_8045,N_8508);
xor U9520 (N_9520,N_8028,N_8017);
or U9521 (N_9521,N_8789,N_8498);
xnor U9522 (N_9522,N_8845,N_8968);
xnor U9523 (N_9523,N_8433,N_8154);
nor U9524 (N_9524,N_8726,N_8135);
nand U9525 (N_9525,N_8118,N_8492);
nor U9526 (N_9526,N_8340,N_8442);
and U9527 (N_9527,N_8694,N_8153);
and U9528 (N_9528,N_8918,N_8421);
or U9529 (N_9529,N_8802,N_8943);
and U9530 (N_9530,N_8702,N_8047);
and U9531 (N_9531,N_8532,N_8903);
or U9532 (N_9532,N_8628,N_8012);
nand U9533 (N_9533,N_8010,N_8079);
nand U9534 (N_9534,N_8270,N_8130);
nand U9535 (N_9535,N_8389,N_8198);
nand U9536 (N_9536,N_8009,N_8640);
nor U9537 (N_9537,N_8422,N_8763);
nand U9538 (N_9538,N_8559,N_8435);
xnor U9539 (N_9539,N_8807,N_8588);
nand U9540 (N_9540,N_8902,N_8761);
or U9541 (N_9541,N_8041,N_8364);
and U9542 (N_9542,N_8338,N_8982);
nand U9543 (N_9543,N_8730,N_8959);
xnor U9544 (N_9544,N_8951,N_8406);
nand U9545 (N_9545,N_8050,N_8857);
and U9546 (N_9546,N_8480,N_8651);
and U9547 (N_9547,N_8546,N_8402);
nand U9548 (N_9548,N_8754,N_8454);
or U9549 (N_9549,N_8865,N_8101);
and U9550 (N_9550,N_8786,N_8705);
and U9551 (N_9551,N_8933,N_8377);
nand U9552 (N_9552,N_8679,N_8473);
or U9553 (N_9553,N_8686,N_8058);
and U9554 (N_9554,N_8817,N_8749);
or U9555 (N_9555,N_8986,N_8408);
and U9556 (N_9556,N_8742,N_8487);
nand U9557 (N_9557,N_8427,N_8463);
nand U9558 (N_9558,N_8004,N_8161);
and U9559 (N_9559,N_8967,N_8752);
or U9560 (N_9560,N_8712,N_8344);
or U9561 (N_9561,N_8156,N_8775);
nor U9562 (N_9562,N_8071,N_8880);
or U9563 (N_9563,N_8841,N_8865);
nor U9564 (N_9564,N_8442,N_8283);
or U9565 (N_9565,N_8815,N_8985);
nor U9566 (N_9566,N_8313,N_8768);
and U9567 (N_9567,N_8440,N_8313);
nand U9568 (N_9568,N_8258,N_8767);
nor U9569 (N_9569,N_8196,N_8216);
nor U9570 (N_9570,N_8547,N_8275);
or U9571 (N_9571,N_8587,N_8080);
and U9572 (N_9572,N_8609,N_8628);
or U9573 (N_9573,N_8893,N_8713);
and U9574 (N_9574,N_8130,N_8466);
and U9575 (N_9575,N_8541,N_8261);
nand U9576 (N_9576,N_8015,N_8484);
nand U9577 (N_9577,N_8469,N_8127);
nor U9578 (N_9578,N_8825,N_8272);
xnor U9579 (N_9579,N_8875,N_8953);
or U9580 (N_9580,N_8121,N_8737);
or U9581 (N_9581,N_8068,N_8142);
nand U9582 (N_9582,N_8415,N_8547);
nand U9583 (N_9583,N_8029,N_8816);
or U9584 (N_9584,N_8569,N_8398);
and U9585 (N_9585,N_8554,N_8526);
xnor U9586 (N_9586,N_8365,N_8589);
nand U9587 (N_9587,N_8238,N_8362);
nor U9588 (N_9588,N_8894,N_8149);
nor U9589 (N_9589,N_8890,N_8950);
nand U9590 (N_9590,N_8253,N_8004);
or U9591 (N_9591,N_8271,N_8622);
xor U9592 (N_9592,N_8745,N_8208);
and U9593 (N_9593,N_8656,N_8776);
or U9594 (N_9594,N_8079,N_8730);
nand U9595 (N_9595,N_8395,N_8309);
or U9596 (N_9596,N_8040,N_8864);
or U9597 (N_9597,N_8290,N_8078);
or U9598 (N_9598,N_8881,N_8452);
or U9599 (N_9599,N_8075,N_8309);
and U9600 (N_9600,N_8029,N_8755);
or U9601 (N_9601,N_8188,N_8944);
nor U9602 (N_9602,N_8524,N_8853);
or U9603 (N_9603,N_8765,N_8572);
or U9604 (N_9604,N_8243,N_8996);
nand U9605 (N_9605,N_8990,N_8224);
nor U9606 (N_9606,N_8224,N_8940);
nand U9607 (N_9607,N_8118,N_8008);
or U9608 (N_9608,N_8822,N_8882);
nor U9609 (N_9609,N_8240,N_8110);
and U9610 (N_9610,N_8102,N_8286);
nand U9611 (N_9611,N_8656,N_8221);
nand U9612 (N_9612,N_8708,N_8984);
nor U9613 (N_9613,N_8730,N_8323);
nor U9614 (N_9614,N_8957,N_8470);
xnor U9615 (N_9615,N_8098,N_8674);
nor U9616 (N_9616,N_8280,N_8350);
nand U9617 (N_9617,N_8148,N_8423);
and U9618 (N_9618,N_8650,N_8385);
nand U9619 (N_9619,N_8785,N_8537);
nand U9620 (N_9620,N_8553,N_8609);
nor U9621 (N_9621,N_8255,N_8563);
nor U9622 (N_9622,N_8241,N_8967);
nand U9623 (N_9623,N_8296,N_8200);
nor U9624 (N_9624,N_8984,N_8563);
nor U9625 (N_9625,N_8407,N_8909);
nor U9626 (N_9626,N_8643,N_8438);
or U9627 (N_9627,N_8282,N_8556);
nor U9628 (N_9628,N_8531,N_8449);
or U9629 (N_9629,N_8165,N_8898);
or U9630 (N_9630,N_8471,N_8915);
nor U9631 (N_9631,N_8414,N_8114);
and U9632 (N_9632,N_8553,N_8798);
nor U9633 (N_9633,N_8889,N_8436);
or U9634 (N_9634,N_8683,N_8509);
or U9635 (N_9635,N_8701,N_8514);
or U9636 (N_9636,N_8635,N_8204);
or U9637 (N_9637,N_8800,N_8941);
xnor U9638 (N_9638,N_8067,N_8123);
or U9639 (N_9639,N_8622,N_8783);
and U9640 (N_9640,N_8702,N_8947);
or U9641 (N_9641,N_8027,N_8157);
nor U9642 (N_9642,N_8108,N_8081);
or U9643 (N_9643,N_8147,N_8456);
nor U9644 (N_9644,N_8599,N_8299);
and U9645 (N_9645,N_8930,N_8984);
or U9646 (N_9646,N_8851,N_8204);
nor U9647 (N_9647,N_8163,N_8341);
nor U9648 (N_9648,N_8379,N_8278);
and U9649 (N_9649,N_8777,N_8837);
nor U9650 (N_9650,N_8802,N_8961);
or U9651 (N_9651,N_8941,N_8641);
nand U9652 (N_9652,N_8995,N_8191);
nand U9653 (N_9653,N_8700,N_8235);
or U9654 (N_9654,N_8880,N_8844);
nand U9655 (N_9655,N_8216,N_8634);
or U9656 (N_9656,N_8028,N_8880);
or U9657 (N_9657,N_8083,N_8959);
and U9658 (N_9658,N_8280,N_8491);
and U9659 (N_9659,N_8761,N_8980);
nand U9660 (N_9660,N_8595,N_8761);
nor U9661 (N_9661,N_8460,N_8295);
and U9662 (N_9662,N_8750,N_8518);
nand U9663 (N_9663,N_8147,N_8095);
nand U9664 (N_9664,N_8536,N_8267);
or U9665 (N_9665,N_8270,N_8559);
xor U9666 (N_9666,N_8583,N_8038);
or U9667 (N_9667,N_8308,N_8409);
nand U9668 (N_9668,N_8303,N_8385);
and U9669 (N_9669,N_8488,N_8304);
or U9670 (N_9670,N_8760,N_8594);
or U9671 (N_9671,N_8001,N_8518);
or U9672 (N_9672,N_8093,N_8470);
or U9673 (N_9673,N_8696,N_8204);
nand U9674 (N_9674,N_8367,N_8495);
or U9675 (N_9675,N_8943,N_8934);
nand U9676 (N_9676,N_8453,N_8888);
nor U9677 (N_9677,N_8006,N_8785);
nand U9678 (N_9678,N_8856,N_8883);
nand U9679 (N_9679,N_8063,N_8122);
nand U9680 (N_9680,N_8114,N_8972);
nor U9681 (N_9681,N_8069,N_8545);
or U9682 (N_9682,N_8466,N_8346);
or U9683 (N_9683,N_8643,N_8472);
and U9684 (N_9684,N_8814,N_8836);
nor U9685 (N_9685,N_8438,N_8050);
and U9686 (N_9686,N_8971,N_8081);
nor U9687 (N_9687,N_8500,N_8720);
and U9688 (N_9688,N_8554,N_8251);
and U9689 (N_9689,N_8686,N_8676);
nor U9690 (N_9690,N_8201,N_8265);
nor U9691 (N_9691,N_8904,N_8146);
or U9692 (N_9692,N_8508,N_8582);
nand U9693 (N_9693,N_8210,N_8306);
or U9694 (N_9694,N_8111,N_8610);
nor U9695 (N_9695,N_8931,N_8783);
nor U9696 (N_9696,N_8945,N_8949);
nor U9697 (N_9697,N_8114,N_8692);
or U9698 (N_9698,N_8634,N_8904);
or U9699 (N_9699,N_8027,N_8250);
and U9700 (N_9700,N_8019,N_8008);
and U9701 (N_9701,N_8617,N_8897);
or U9702 (N_9702,N_8613,N_8320);
nand U9703 (N_9703,N_8299,N_8046);
or U9704 (N_9704,N_8666,N_8521);
or U9705 (N_9705,N_8790,N_8684);
nor U9706 (N_9706,N_8764,N_8133);
nand U9707 (N_9707,N_8787,N_8845);
nor U9708 (N_9708,N_8168,N_8433);
nor U9709 (N_9709,N_8855,N_8994);
or U9710 (N_9710,N_8610,N_8031);
nor U9711 (N_9711,N_8259,N_8768);
nor U9712 (N_9712,N_8470,N_8310);
nor U9713 (N_9713,N_8101,N_8048);
nor U9714 (N_9714,N_8148,N_8072);
or U9715 (N_9715,N_8538,N_8982);
xor U9716 (N_9716,N_8934,N_8135);
or U9717 (N_9717,N_8230,N_8410);
and U9718 (N_9718,N_8812,N_8806);
and U9719 (N_9719,N_8028,N_8844);
nor U9720 (N_9720,N_8079,N_8901);
nor U9721 (N_9721,N_8023,N_8684);
and U9722 (N_9722,N_8300,N_8018);
nand U9723 (N_9723,N_8335,N_8912);
nand U9724 (N_9724,N_8967,N_8612);
or U9725 (N_9725,N_8646,N_8500);
or U9726 (N_9726,N_8861,N_8438);
nand U9727 (N_9727,N_8957,N_8104);
nor U9728 (N_9728,N_8532,N_8932);
or U9729 (N_9729,N_8384,N_8013);
nor U9730 (N_9730,N_8959,N_8251);
nand U9731 (N_9731,N_8155,N_8909);
nor U9732 (N_9732,N_8021,N_8331);
and U9733 (N_9733,N_8158,N_8953);
xor U9734 (N_9734,N_8047,N_8777);
and U9735 (N_9735,N_8574,N_8806);
xor U9736 (N_9736,N_8241,N_8473);
xnor U9737 (N_9737,N_8524,N_8919);
and U9738 (N_9738,N_8038,N_8201);
or U9739 (N_9739,N_8744,N_8534);
or U9740 (N_9740,N_8656,N_8328);
nor U9741 (N_9741,N_8167,N_8184);
and U9742 (N_9742,N_8526,N_8180);
nand U9743 (N_9743,N_8185,N_8965);
nand U9744 (N_9744,N_8235,N_8702);
and U9745 (N_9745,N_8766,N_8309);
nand U9746 (N_9746,N_8603,N_8425);
nand U9747 (N_9747,N_8462,N_8577);
xor U9748 (N_9748,N_8389,N_8483);
and U9749 (N_9749,N_8568,N_8202);
and U9750 (N_9750,N_8115,N_8949);
and U9751 (N_9751,N_8784,N_8176);
nand U9752 (N_9752,N_8318,N_8964);
nor U9753 (N_9753,N_8070,N_8711);
and U9754 (N_9754,N_8700,N_8455);
or U9755 (N_9755,N_8436,N_8122);
or U9756 (N_9756,N_8069,N_8898);
nand U9757 (N_9757,N_8997,N_8216);
nand U9758 (N_9758,N_8485,N_8171);
nor U9759 (N_9759,N_8965,N_8402);
and U9760 (N_9760,N_8776,N_8939);
or U9761 (N_9761,N_8220,N_8429);
xor U9762 (N_9762,N_8236,N_8670);
nand U9763 (N_9763,N_8391,N_8854);
or U9764 (N_9764,N_8624,N_8667);
or U9765 (N_9765,N_8987,N_8118);
and U9766 (N_9766,N_8697,N_8349);
or U9767 (N_9767,N_8261,N_8937);
or U9768 (N_9768,N_8027,N_8692);
nand U9769 (N_9769,N_8413,N_8790);
nand U9770 (N_9770,N_8501,N_8416);
nand U9771 (N_9771,N_8303,N_8189);
nor U9772 (N_9772,N_8510,N_8350);
or U9773 (N_9773,N_8882,N_8307);
nor U9774 (N_9774,N_8198,N_8290);
or U9775 (N_9775,N_8516,N_8803);
nand U9776 (N_9776,N_8025,N_8837);
or U9777 (N_9777,N_8218,N_8567);
nor U9778 (N_9778,N_8845,N_8777);
nand U9779 (N_9779,N_8271,N_8423);
and U9780 (N_9780,N_8596,N_8452);
xnor U9781 (N_9781,N_8264,N_8179);
nor U9782 (N_9782,N_8883,N_8351);
or U9783 (N_9783,N_8410,N_8961);
nor U9784 (N_9784,N_8644,N_8473);
or U9785 (N_9785,N_8828,N_8921);
nand U9786 (N_9786,N_8865,N_8105);
nand U9787 (N_9787,N_8739,N_8468);
and U9788 (N_9788,N_8698,N_8999);
nand U9789 (N_9789,N_8316,N_8224);
and U9790 (N_9790,N_8127,N_8415);
nand U9791 (N_9791,N_8993,N_8553);
nor U9792 (N_9792,N_8097,N_8352);
nand U9793 (N_9793,N_8489,N_8603);
nand U9794 (N_9794,N_8432,N_8612);
and U9795 (N_9795,N_8767,N_8278);
nand U9796 (N_9796,N_8071,N_8823);
and U9797 (N_9797,N_8682,N_8404);
and U9798 (N_9798,N_8468,N_8301);
xnor U9799 (N_9799,N_8383,N_8582);
and U9800 (N_9800,N_8556,N_8571);
nor U9801 (N_9801,N_8996,N_8078);
nor U9802 (N_9802,N_8184,N_8206);
nor U9803 (N_9803,N_8715,N_8874);
xor U9804 (N_9804,N_8097,N_8130);
and U9805 (N_9805,N_8804,N_8636);
nand U9806 (N_9806,N_8740,N_8591);
or U9807 (N_9807,N_8288,N_8490);
nor U9808 (N_9808,N_8263,N_8011);
and U9809 (N_9809,N_8123,N_8651);
or U9810 (N_9810,N_8276,N_8098);
xnor U9811 (N_9811,N_8773,N_8800);
nor U9812 (N_9812,N_8624,N_8117);
nand U9813 (N_9813,N_8390,N_8603);
nand U9814 (N_9814,N_8534,N_8662);
or U9815 (N_9815,N_8059,N_8584);
or U9816 (N_9816,N_8838,N_8079);
nand U9817 (N_9817,N_8481,N_8564);
and U9818 (N_9818,N_8565,N_8534);
nand U9819 (N_9819,N_8481,N_8072);
nand U9820 (N_9820,N_8751,N_8548);
or U9821 (N_9821,N_8098,N_8736);
xnor U9822 (N_9822,N_8776,N_8121);
and U9823 (N_9823,N_8649,N_8051);
nor U9824 (N_9824,N_8071,N_8800);
nand U9825 (N_9825,N_8404,N_8047);
or U9826 (N_9826,N_8948,N_8619);
xor U9827 (N_9827,N_8954,N_8048);
nand U9828 (N_9828,N_8712,N_8361);
nand U9829 (N_9829,N_8831,N_8705);
or U9830 (N_9830,N_8030,N_8648);
nand U9831 (N_9831,N_8395,N_8527);
nand U9832 (N_9832,N_8847,N_8849);
or U9833 (N_9833,N_8710,N_8900);
nand U9834 (N_9834,N_8180,N_8643);
nor U9835 (N_9835,N_8570,N_8023);
or U9836 (N_9836,N_8087,N_8999);
and U9837 (N_9837,N_8488,N_8020);
and U9838 (N_9838,N_8097,N_8555);
xor U9839 (N_9839,N_8852,N_8260);
or U9840 (N_9840,N_8892,N_8548);
or U9841 (N_9841,N_8088,N_8663);
or U9842 (N_9842,N_8693,N_8865);
nand U9843 (N_9843,N_8038,N_8821);
nand U9844 (N_9844,N_8459,N_8139);
xnor U9845 (N_9845,N_8926,N_8367);
and U9846 (N_9846,N_8445,N_8949);
nor U9847 (N_9847,N_8875,N_8084);
or U9848 (N_9848,N_8247,N_8905);
xor U9849 (N_9849,N_8878,N_8980);
nor U9850 (N_9850,N_8789,N_8046);
or U9851 (N_9851,N_8235,N_8888);
nand U9852 (N_9852,N_8612,N_8963);
nand U9853 (N_9853,N_8202,N_8670);
or U9854 (N_9854,N_8350,N_8946);
nand U9855 (N_9855,N_8294,N_8516);
nand U9856 (N_9856,N_8868,N_8743);
or U9857 (N_9857,N_8125,N_8771);
nand U9858 (N_9858,N_8825,N_8727);
and U9859 (N_9859,N_8927,N_8884);
or U9860 (N_9860,N_8575,N_8401);
and U9861 (N_9861,N_8304,N_8936);
nand U9862 (N_9862,N_8997,N_8781);
xnor U9863 (N_9863,N_8985,N_8122);
and U9864 (N_9864,N_8119,N_8936);
or U9865 (N_9865,N_8781,N_8733);
nor U9866 (N_9866,N_8249,N_8104);
nor U9867 (N_9867,N_8094,N_8162);
nand U9868 (N_9868,N_8957,N_8671);
and U9869 (N_9869,N_8766,N_8162);
and U9870 (N_9870,N_8330,N_8811);
or U9871 (N_9871,N_8918,N_8500);
nor U9872 (N_9872,N_8313,N_8869);
nand U9873 (N_9873,N_8094,N_8445);
nor U9874 (N_9874,N_8297,N_8010);
and U9875 (N_9875,N_8410,N_8108);
and U9876 (N_9876,N_8572,N_8176);
or U9877 (N_9877,N_8043,N_8092);
and U9878 (N_9878,N_8175,N_8728);
nand U9879 (N_9879,N_8672,N_8703);
and U9880 (N_9880,N_8127,N_8041);
and U9881 (N_9881,N_8022,N_8516);
and U9882 (N_9882,N_8350,N_8156);
and U9883 (N_9883,N_8041,N_8302);
and U9884 (N_9884,N_8480,N_8136);
xnor U9885 (N_9885,N_8006,N_8841);
or U9886 (N_9886,N_8761,N_8159);
or U9887 (N_9887,N_8600,N_8917);
xnor U9888 (N_9888,N_8817,N_8558);
nor U9889 (N_9889,N_8642,N_8541);
or U9890 (N_9890,N_8457,N_8780);
or U9891 (N_9891,N_8596,N_8369);
or U9892 (N_9892,N_8516,N_8479);
and U9893 (N_9893,N_8835,N_8421);
or U9894 (N_9894,N_8402,N_8938);
nand U9895 (N_9895,N_8160,N_8063);
and U9896 (N_9896,N_8235,N_8690);
and U9897 (N_9897,N_8695,N_8995);
nand U9898 (N_9898,N_8758,N_8374);
or U9899 (N_9899,N_8069,N_8483);
and U9900 (N_9900,N_8565,N_8324);
and U9901 (N_9901,N_8366,N_8770);
and U9902 (N_9902,N_8449,N_8925);
nor U9903 (N_9903,N_8596,N_8758);
xor U9904 (N_9904,N_8170,N_8125);
or U9905 (N_9905,N_8479,N_8957);
nand U9906 (N_9906,N_8420,N_8739);
nand U9907 (N_9907,N_8982,N_8109);
or U9908 (N_9908,N_8307,N_8413);
and U9909 (N_9909,N_8842,N_8053);
or U9910 (N_9910,N_8191,N_8710);
nor U9911 (N_9911,N_8885,N_8383);
nand U9912 (N_9912,N_8240,N_8567);
nand U9913 (N_9913,N_8354,N_8129);
xor U9914 (N_9914,N_8268,N_8861);
nor U9915 (N_9915,N_8854,N_8149);
nor U9916 (N_9916,N_8192,N_8505);
nand U9917 (N_9917,N_8773,N_8185);
nand U9918 (N_9918,N_8168,N_8662);
and U9919 (N_9919,N_8334,N_8727);
nand U9920 (N_9920,N_8486,N_8014);
xnor U9921 (N_9921,N_8061,N_8019);
nor U9922 (N_9922,N_8181,N_8490);
and U9923 (N_9923,N_8378,N_8967);
and U9924 (N_9924,N_8215,N_8292);
or U9925 (N_9925,N_8960,N_8723);
nor U9926 (N_9926,N_8437,N_8734);
or U9927 (N_9927,N_8142,N_8896);
and U9928 (N_9928,N_8258,N_8494);
xnor U9929 (N_9929,N_8409,N_8938);
and U9930 (N_9930,N_8129,N_8760);
and U9931 (N_9931,N_8248,N_8463);
xnor U9932 (N_9932,N_8260,N_8976);
nand U9933 (N_9933,N_8136,N_8486);
or U9934 (N_9934,N_8725,N_8320);
or U9935 (N_9935,N_8378,N_8715);
and U9936 (N_9936,N_8950,N_8491);
and U9937 (N_9937,N_8160,N_8556);
nor U9938 (N_9938,N_8047,N_8212);
and U9939 (N_9939,N_8042,N_8332);
and U9940 (N_9940,N_8256,N_8756);
nand U9941 (N_9941,N_8953,N_8167);
xor U9942 (N_9942,N_8606,N_8375);
nand U9943 (N_9943,N_8637,N_8871);
nor U9944 (N_9944,N_8395,N_8798);
nor U9945 (N_9945,N_8908,N_8609);
or U9946 (N_9946,N_8027,N_8160);
and U9947 (N_9947,N_8515,N_8915);
nand U9948 (N_9948,N_8611,N_8566);
nand U9949 (N_9949,N_8732,N_8237);
or U9950 (N_9950,N_8376,N_8998);
and U9951 (N_9951,N_8921,N_8645);
or U9952 (N_9952,N_8523,N_8757);
or U9953 (N_9953,N_8404,N_8385);
and U9954 (N_9954,N_8716,N_8065);
nand U9955 (N_9955,N_8568,N_8406);
or U9956 (N_9956,N_8103,N_8674);
or U9957 (N_9957,N_8179,N_8349);
nand U9958 (N_9958,N_8318,N_8572);
nand U9959 (N_9959,N_8028,N_8617);
and U9960 (N_9960,N_8420,N_8989);
nor U9961 (N_9961,N_8592,N_8692);
or U9962 (N_9962,N_8807,N_8394);
nand U9963 (N_9963,N_8648,N_8785);
xor U9964 (N_9964,N_8214,N_8582);
nor U9965 (N_9965,N_8968,N_8260);
or U9966 (N_9966,N_8898,N_8070);
and U9967 (N_9967,N_8658,N_8371);
nand U9968 (N_9968,N_8203,N_8518);
nand U9969 (N_9969,N_8456,N_8846);
xor U9970 (N_9970,N_8560,N_8829);
xor U9971 (N_9971,N_8368,N_8148);
or U9972 (N_9972,N_8788,N_8912);
nor U9973 (N_9973,N_8190,N_8378);
nor U9974 (N_9974,N_8883,N_8027);
or U9975 (N_9975,N_8916,N_8065);
nor U9976 (N_9976,N_8225,N_8218);
or U9977 (N_9977,N_8118,N_8093);
or U9978 (N_9978,N_8958,N_8760);
xnor U9979 (N_9979,N_8818,N_8346);
xnor U9980 (N_9980,N_8755,N_8057);
and U9981 (N_9981,N_8603,N_8991);
xor U9982 (N_9982,N_8079,N_8832);
or U9983 (N_9983,N_8368,N_8768);
nor U9984 (N_9984,N_8281,N_8131);
nor U9985 (N_9985,N_8092,N_8647);
nand U9986 (N_9986,N_8781,N_8535);
and U9987 (N_9987,N_8217,N_8689);
nor U9988 (N_9988,N_8548,N_8240);
nand U9989 (N_9989,N_8419,N_8758);
or U9990 (N_9990,N_8732,N_8693);
and U9991 (N_9991,N_8202,N_8767);
and U9992 (N_9992,N_8638,N_8338);
or U9993 (N_9993,N_8097,N_8703);
nand U9994 (N_9994,N_8182,N_8135);
nor U9995 (N_9995,N_8087,N_8480);
and U9996 (N_9996,N_8522,N_8464);
xor U9997 (N_9997,N_8145,N_8233);
nor U9998 (N_9998,N_8654,N_8275);
nor U9999 (N_9999,N_8761,N_8453);
nor UO_0 (O_0,N_9275,N_9114);
and UO_1 (O_1,N_9146,N_9700);
xnor UO_2 (O_2,N_9753,N_9799);
nor UO_3 (O_3,N_9750,N_9542);
nor UO_4 (O_4,N_9718,N_9116);
nand UO_5 (O_5,N_9384,N_9537);
or UO_6 (O_6,N_9771,N_9027);
or UO_7 (O_7,N_9199,N_9941);
nand UO_8 (O_8,N_9181,N_9659);
nor UO_9 (O_9,N_9556,N_9948);
nor UO_10 (O_10,N_9924,N_9862);
and UO_11 (O_11,N_9947,N_9967);
or UO_12 (O_12,N_9066,N_9647);
and UO_13 (O_13,N_9124,N_9264);
xnor UO_14 (O_14,N_9785,N_9974);
nand UO_15 (O_15,N_9787,N_9470);
xnor UO_16 (O_16,N_9156,N_9694);
or UO_17 (O_17,N_9676,N_9227);
or UO_18 (O_18,N_9857,N_9225);
nand UO_19 (O_19,N_9747,N_9819);
nand UO_20 (O_20,N_9381,N_9080);
nor UO_21 (O_21,N_9772,N_9793);
and UO_22 (O_22,N_9092,N_9311);
nand UO_23 (O_23,N_9539,N_9257);
or UO_24 (O_24,N_9707,N_9855);
and UO_25 (O_25,N_9786,N_9474);
or UO_26 (O_26,N_9581,N_9651);
nand UO_27 (O_27,N_9251,N_9303);
or UO_28 (O_28,N_9844,N_9729);
nor UO_29 (O_29,N_9286,N_9258);
or UO_30 (O_30,N_9428,N_9397);
nand UO_31 (O_31,N_9921,N_9529);
nor UO_32 (O_32,N_9219,N_9134);
and UO_33 (O_33,N_9353,N_9062);
nor UO_34 (O_34,N_9861,N_9169);
and UO_35 (O_35,N_9567,N_9839);
xnor UO_36 (O_36,N_9763,N_9640);
nor UO_37 (O_37,N_9795,N_9490);
nor UO_38 (O_38,N_9285,N_9500);
nand UO_39 (O_39,N_9505,N_9028);
nand UO_40 (O_40,N_9807,N_9248);
nor UO_41 (O_41,N_9705,N_9421);
nor UO_42 (O_42,N_9409,N_9089);
xnor UO_43 (O_43,N_9626,N_9522);
or UO_44 (O_44,N_9082,N_9748);
or UO_45 (O_45,N_9063,N_9527);
and UO_46 (O_46,N_9991,N_9675);
and UO_47 (O_47,N_9933,N_9130);
nor UO_48 (O_48,N_9761,N_9329);
and UO_49 (O_49,N_9570,N_9448);
nor UO_50 (O_50,N_9436,N_9135);
or UO_51 (O_51,N_9593,N_9657);
nor UO_52 (O_52,N_9240,N_9084);
and UO_53 (O_53,N_9590,N_9325);
or UO_54 (O_54,N_9741,N_9427);
xnor UO_55 (O_55,N_9493,N_9633);
or UO_56 (O_56,N_9038,N_9953);
and UO_57 (O_57,N_9402,N_9830);
or UO_58 (O_58,N_9404,N_9764);
nor UO_59 (O_59,N_9091,N_9456);
nor UO_60 (O_60,N_9186,N_9698);
and UO_61 (O_61,N_9685,N_9480);
or UO_62 (O_62,N_9843,N_9681);
or UO_63 (O_63,N_9669,N_9702);
and UO_64 (O_64,N_9157,N_9895);
or UO_65 (O_65,N_9616,N_9461);
nor UO_66 (O_66,N_9762,N_9552);
or UO_67 (O_67,N_9252,N_9191);
nand UO_68 (O_68,N_9936,N_9105);
nor UO_69 (O_69,N_9532,N_9337);
or UO_70 (O_70,N_9610,N_9547);
nand UO_71 (O_71,N_9417,N_9858);
or UO_72 (O_72,N_9719,N_9208);
and UO_73 (O_73,N_9393,N_9880);
nand UO_74 (O_74,N_9333,N_9809);
or UO_75 (O_75,N_9003,N_9064);
nor UO_76 (O_76,N_9473,N_9435);
and UO_77 (O_77,N_9206,N_9929);
nor UO_78 (O_78,N_9608,N_9018);
and UO_79 (O_79,N_9366,N_9371);
xor UO_80 (O_80,N_9395,N_9587);
nand UO_81 (O_81,N_9853,N_9665);
nand UO_82 (O_82,N_9232,N_9937);
and UO_83 (O_83,N_9842,N_9036);
nand UO_84 (O_84,N_9602,N_9917);
nor UO_85 (O_85,N_9611,N_9289);
nand UO_86 (O_86,N_9033,N_9348);
nand UO_87 (O_87,N_9363,N_9376);
and UO_88 (O_88,N_9488,N_9686);
nand UO_89 (O_89,N_9399,N_9449);
nor UO_90 (O_90,N_9182,N_9851);
and UO_91 (O_91,N_9160,N_9727);
nor UO_92 (O_92,N_9714,N_9392);
nand UO_93 (O_93,N_9189,N_9101);
or UO_94 (O_94,N_9560,N_9489);
nor UO_95 (O_95,N_9165,N_9030);
or UO_96 (O_96,N_9068,N_9260);
and UO_97 (O_97,N_9850,N_9108);
xor UO_98 (O_98,N_9596,N_9554);
nor UO_99 (O_99,N_9731,N_9503);
or UO_100 (O_100,N_9241,N_9841);
nand UO_101 (O_101,N_9072,N_9013);
or UO_102 (O_102,N_9815,N_9901);
nor UO_103 (O_103,N_9242,N_9943);
nand UO_104 (O_104,N_9831,N_9653);
and UO_105 (O_105,N_9388,N_9346);
or UO_106 (O_106,N_9774,N_9722);
and UO_107 (O_107,N_9978,N_9153);
and UO_108 (O_108,N_9960,N_9804);
and UO_109 (O_109,N_9541,N_9273);
and UO_110 (O_110,N_9450,N_9012);
nor UO_111 (O_111,N_9483,N_9071);
nand UO_112 (O_112,N_9387,N_9380);
nand UO_113 (O_113,N_9999,N_9414);
xor UO_114 (O_114,N_9689,N_9284);
nor UO_115 (O_115,N_9416,N_9954);
nor UO_116 (O_116,N_9663,N_9778);
and UO_117 (O_117,N_9276,N_9755);
or UO_118 (O_118,N_9229,N_9073);
nand UO_119 (O_119,N_9057,N_9496);
or UO_120 (O_120,N_9674,N_9245);
and UO_121 (O_121,N_9837,N_9408);
nand UO_122 (O_122,N_9594,N_9897);
or UO_123 (O_123,N_9695,N_9744);
xor UO_124 (O_124,N_9400,N_9870);
xor UO_125 (O_125,N_9952,N_9998);
xnor UO_126 (O_126,N_9234,N_9144);
or UO_127 (O_127,N_9495,N_9730);
and UO_128 (O_128,N_9128,N_9099);
or UO_129 (O_129,N_9223,N_9846);
and UO_130 (O_130,N_9670,N_9106);
nor UO_131 (O_131,N_9713,N_9899);
and UO_132 (O_132,N_9055,N_9194);
or UO_133 (O_133,N_9131,N_9925);
nor UO_134 (O_134,N_9886,N_9386);
nand UO_135 (O_135,N_9765,N_9792);
nor UO_136 (O_136,N_9088,N_9865);
and UO_137 (O_137,N_9053,N_9928);
and UO_138 (O_138,N_9025,N_9354);
nor UO_139 (O_139,N_9530,N_9005);
and UO_140 (O_140,N_9783,N_9178);
or UO_141 (O_141,N_9715,N_9565);
nor UO_142 (O_142,N_9228,N_9618);
nand UO_143 (O_143,N_9817,N_9211);
xnor UO_144 (O_144,N_9017,N_9379);
nand UO_145 (O_145,N_9320,N_9918);
and UO_146 (O_146,N_9782,N_9562);
or UO_147 (O_147,N_9797,N_9652);
nor UO_148 (O_148,N_9332,N_9544);
or UO_149 (O_149,N_9634,N_9323);
nor UO_150 (O_150,N_9293,N_9508);
and UO_151 (O_151,N_9236,N_9979);
nand UO_152 (O_152,N_9210,N_9636);
nand UO_153 (O_153,N_9048,N_9989);
nand UO_154 (O_154,N_9790,N_9358);
or UO_155 (O_155,N_9056,N_9893);
xnor UO_156 (O_156,N_9294,N_9336);
nand UO_157 (O_157,N_9872,N_9423);
nor UO_158 (O_158,N_9906,N_9357);
and UO_159 (O_159,N_9022,N_9845);
and UO_160 (O_160,N_9269,N_9511);
and UO_161 (O_161,N_9331,N_9654);
nor UO_162 (O_162,N_9758,N_9350);
nand UO_163 (O_163,N_9009,N_9733);
nand UO_164 (O_164,N_9006,N_9487);
nor UO_165 (O_165,N_9356,N_9254);
or UO_166 (O_166,N_9310,N_9342);
or UO_167 (O_167,N_9283,N_9672);
xor UO_168 (O_168,N_9262,N_9919);
nand UO_169 (O_169,N_9368,N_9892);
xnor UO_170 (O_170,N_9679,N_9412);
nor UO_171 (O_171,N_9205,N_9008);
nand UO_172 (O_172,N_9308,N_9244);
nor UO_173 (O_173,N_9396,N_9445);
nor UO_174 (O_174,N_9187,N_9297);
nand UO_175 (O_175,N_9971,N_9370);
and UO_176 (O_176,N_9859,N_9724);
nand UO_177 (O_177,N_9045,N_9760);
xnor UO_178 (O_178,N_9407,N_9805);
nand UO_179 (O_179,N_9280,N_9996);
xnor UO_180 (O_180,N_9621,N_9406);
nor UO_181 (O_181,N_9338,N_9459);
nand UO_182 (O_182,N_9891,N_9172);
and UO_183 (O_183,N_9136,N_9141);
nor UO_184 (O_184,N_9198,N_9439);
and UO_185 (O_185,N_9024,N_9347);
or UO_186 (O_186,N_9641,N_9019);
nor UO_187 (O_187,N_9646,N_9316);
or UO_188 (O_188,N_9137,N_9355);
and UO_189 (O_189,N_9246,N_9163);
nand UO_190 (O_190,N_9566,N_9582);
xor UO_191 (O_191,N_9606,N_9528);
xnor UO_192 (O_192,N_9808,N_9438);
nand UO_193 (O_193,N_9442,N_9923);
and UO_194 (O_194,N_9769,N_9301);
xnor UO_195 (O_195,N_9094,N_9812);
and UO_196 (O_196,N_9341,N_9649);
or UO_197 (O_197,N_9213,N_9235);
or UO_198 (O_198,N_9279,N_9548);
or UO_199 (O_199,N_9540,N_9834);
or UO_200 (O_200,N_9613,N_9271);
or UO_201 (O_201,N_9209,N_9935);
and UO_202 (O_202,N_9796,N_9000);
or UO_203 (O_203,N_9349,N_9391);
or UO_204 (O_204,N_9723,N_9123);
nand UO_205 (O_205,N_9946,N_9875);
or UO_206 (O_206,N_9307,N_9553);
nand UO_207 (O_207,N_9510,N_9468);
nor UO_208 (O_208,N_9390,N_9903);
xor UO_209 (O_209,N_9170,N_9523);
nand UO_210 (O_210,N_9838,N_9878);
and UO_211 (O_211,N_9564,N_9453);
or UO_212 (O_212,N_9249,N_9112);
or UO_213 (O_213,N_9230,N_9981);
and UO_214 (O_214,N_9010,N_9572);
nand UO_215 (O_215,N_9430,N_9300);
nor UO_216 (O_216,N_9874,N_9043);
or UO_217 (O_217,N_9079,N_9096);
and UO_218 (O_218,N_9561,N_9711);
nor UO_219 (O_219,N_9531,N_9315);
xnor UO_220 (O_220,N_9951,N_9321);
and UO_221 (O_221,N_9635,N_9431);
xor UO_222 (O_222,N_9437,N_9344);
nor UO_223 (O_223,N_9288,N_9111);
and UO_224 (O_224,N_9688,N_9330);
and UO_225 (O_225,N_9476,N_9151);
nor UO_226 (O_226,N_9351,N_9983);
or UO_227 (O_227,N_9039,N_9167);
nand UO_228 (O_228,N_9215,N_9995);
and UO_229 (O_229,N_9848,N_9418);
nand UO_230 (O_230,N_9049,N_9619);
nor UO_231 (O_231,N_9014,N_9318);
nand UO_232 (O_232,N_9429,N_9985);
or UO_233 (O_233,N_9377,N_9040);
and UO_234 (O_234,N_9988,N_9963);
and UO_235 (O_235,N_9585,N_9142);
nor UO_236 (O_236,N_9526,N_9823);
xor UO_237 (O_237,N_9682,N_9067);
nand UO_238 (O_238,N_9352,N_9756);
or UO_239 (O_239,N_9692,N_9592);
xnor UO_240 (O_240,N_9847,N_9680);
and UO_241 (O_241,N_9287,N_9910);
nor UO_242 (O_242,N_9509,N_9104);
or UO_243 (O_243,N_9023,N_9638);
or UO_244 (O_244,N_9882,N_9890);
or UO_245 (O_245,N_9441,N_9274);
and UO_246 (O_246,N_9803,N_9888);
and UO_247 (O_247,N_9224,N_9029);
or UO_248 (O_248,N_9779,N_9949);
and UO_249 (O_249,N_9202,N_9990);
or UO_250 (O_250,N_9422,N_9662);
nand UO_251 (O_251,N_9885,N_9502);
nand UO_252 (O_252,N_9455,N_9993);
nor UO_253 (O_253,N_9827,N_9766);
and UO_254 (O_254,N_9643,N_9607);
or UO_255 (O_255,N_9873,N_9220);
and UO_256 (O_256,N_9908,N_9717);
nand UO_257 (O_257,N_9664,N_9265);
or UO_258 (O_258,N_9405,N_9375);
nand UO_259 (O_259,N_9726,N_9369);
or UO_260 (O_260,N_9575,N_9693);
nand UO_261 (O_261,N_9343,N_9942);
or UO_262 (O_262,N_9233,N_9047);
or UO_263 (O_263,N_9469,N_9026);
and UO_264 (O_264,N_9075,N_9295);
nand UO_265 (O_265,N_9155,N_9628);
or UO_266 (O_266,N_9869,N_9577);
and UO_267 (O_267,N_9021,N_9322);
and UO_268 (O_268,N_9583,N_9648);
or UO_269 (O_269,N_9403,N_9655);
nand UO_270 (O_270,N_9317,N_9780);
and UO_271 (O_271,N_9401,N_9624);
nor UO_272 (O_272,N_9207,N_9866);
or UO_273 (O_273,N_9849,N_9970);
or UO_274 (O_274,N_9630,N_9856);
or UO_275 (O_275,N_9078,N_9661);
and UO_276 (O_276,N_9464,N_9296);
or UO_277 (O_277,N_9477,N_9513);
nor UO_278 (O_278,N_9113,N_9835);
or UO_279 (O_279,N_9125,N_9568);
nand UO_280 (O_280,N_9833,N_9639);
or UO_281 (O_281,N_9121,N_9745);
nand UO_282 (O_282,N_9451,N_9465);
xnor UO_283 (O_283,N_9515,N_9867);
nand UO_284 (O_284,N_9927,N_9081);
or UO_285 (O_285,N_9304,N_9701);
nand UO_286 (O_286,N_9256,N_9054);
nand UO_287 (O_287,N_9133,N_9810);
and UO_288 (O_288,N_9696,N_9822);
xnor UO_289 (O_289,N_9050,N_9253);
or UO_290 (O_290,N_9749,N_9573);
xor UO_291 (O_291,N_9632,N_9904);
or UO_292 (O_292,N_9190,N_9148);
and UO_293 (O_293,N_9980,N_9902);
and UO_294 (O_294,N_9595,N_9140);
and UO_295 (O_295,N_9298,N_9982);
xor UO_296 (O_296,N_9267,N_9800);
and UO_297 (O_297,N_9992,N_9217);
nand UO_298 (O_298,N_9197,N_9314);
nand UO_299 (O_299,N_9864,N_9166);
nor UO_300 (O_300,N_9521,N_9704);
nand UO_301 (O_301,N_9597,N_9860);
and UO_302 (O_302,N_9759,N_9277);
or UO_303 (O_303,N_9374,N_9997);
nor UO_304 (O_304,N_9291,N_9746);
or UO_305 (O_305,N_9328,N_9306);
nor UO_306 (O_306,N_9788,N_9305);
and UO_307 (O_307,N_9533,N_9884);
and UO_308 (O_308,N_9150,N_9961);
nor UO_309 (O_309,N_9203,N_9896);
and UO_310 (O_310,N_9212,N_9912);
or UO_311 (O_311,N_9339,N_9754);
and UO_312 (O_312,N_9334,N_9907);
nor UO_313 (O_313,N_9446,N_9986);
nor UO_314 (O_314,N_9117,N_9032);
nand UO_315 (O_315,N_9491,N_9770);
and UO_316 (O_316,N_9725,N_9102);
nor UO_317 (O_317,N_9829,N_9964);
nor UO_318 (O_318,N_9889,N_9041);
and UO_319 (O_319,N_9176,N_9828);
nor UO_320 (O_320,N_9868,N_9097);
or UO_321 (O_321,N_9580,N_9721);
and UO_322 (O_322,N_9781,N_9854);
xor UO_323 (O_323,N_9668,N_9922);
and UO_324 (O_324,N_9378,N_9667);
and UO_325 (O_325,N_9627,N_9697);
nor UO_326 (O_326,N_9767,N_9196);
nand UO_327 (O_327,N_9525,N_9460);
and UO_328 (O_328,N_9266,N_9327);
nand UO_329 (O_329,N_9625,N_9179);
nor UO_330 (O_330,N_9973,N_9058);
nor UO_331 (O_331,N_9752,N_9103);
nor UO_332 (O_332,N_9716,N_9604);
or UO_333 (O_333,N_9440,N_9571);
or UO_334 (O_334,N_9020,N_9751);
xor UO_335 (O_335,N_9263,N_9802);
xor UO_336 (O_336,N_9703,N_9950);
or UO_337 (O_337,N_9814,N_9433);
nor UO_338 (O_338,N_9085,N_9945);
and UO_339 (O_339,N_9193,N_9454);
xnor UO_340 (O_340,N_9699,N_9852);
nor UO_341 (O_341,N_9494,N_9143);
nor UO_342 (O_342,N_9312,N_9535);
xor UO_343 (O_343,N_9507,N_9076);
nand UO_344 (O_344,N_9472,N_9385);
and UO_345 (O_345,N_9367,N_9550);
or UO_346 (O_346,N_9876,N_9966);
and UO_347 (O_347,N_9574,N_9938);
or UO_348 (O_348,N_9518,N_9415);
or UO_349 (O_349,N_9313,N_9840);
xor UO_350 (O_350,N_9962,N_9660);
nand UO_351 (O_351,N_9877,N_9900);
nand UO_352 (O_352,N_9557,N_9359);
or UO_353 (O_353,N_9683,N_9420);
nand UO_354 (O_354,N_9994,N_9777);
and UO_355 (O_355,N_9984,N_9383);
or UO_356 (O_356,N_9620,N_9958);
or UO_357 (O_357,N_9965,N_9836);
or UO_358 (O_358,N_9093,N_9784);
and UO_359 (O_359,N_9791,N_9268);
or UO_360 (O_360,N_9498,N_9881);
nand UO_361 (O_361,N_9955,N_9920);
and UO_362 (O_362,N_9195,N_9204);
or UO_363 (O_363,N_9832,N_9158);
or UO_364 (O_364,N_9132,N_9740);
xnor UO_365 (O_365,N_9086,N_9536);
and UO_366 (O_366,N_9545,N_9444);
and UO_367 (O_367,N_9011,N_9364);
xor UO_368 (O_368,N_9601,N_9161);
or UO_369 (O_369,N_9598,N_9466);
and UO_370 (O_370,N_9292,N_9658);
nand UO_371 (O_371,N_9909,N_9326);
nand UO_372 (O_372,N_9044,N_9650);
or UO_373 (O_373,N_9237,N_9255);
and UO_374 (O_374,N_9410,N_9389);
nand UO_375 (O_375,N_9743,N_9637);
or UO_376 (O_376,N_9738,N_9478);
nor UO_377 (O_377,N_9180,N_9871);
or UO_378 (O_378,N_9734,N_9120);
xor UO_379 (O_379,N_9690,N_9914);
or UO_380 (O_380,N_9776,N_9046);
nor UO_381 (O_381,N_9411,N_9934);
nand UO_382 (O_382,N_9159,N_9558);
nand UO_383 (O_383,N_9492,N_9584);
nand UO_384 (O_384,N_9247,N_9671);
nor UO_385 (O_385,N_9119,N_9164);
or UO_386 (O_386,N_9090,N_9479);
or UO_387 (O_387,N_9145,N_9972);
nand UO_388 (O_388,N_9149,N_9152);
nor UO_389 (O_389,N_9462,N_9007);
or UO_390 (O_390,N_9789,N_9324);
nor UO_391 (O_391,N_9037,N_9485);
nor UO_392 (O_392,N_9617,N_9259);
nor UO_393 (O_393,N_9818,N_9015);
nand UO_394 (O_394,N_9801,N_9569);
nor UO_395 (O_395,N_9184,N_9911);
nand UO_396 (O_396,N_9070,N_9188);
nor UO_397 (O_397,N_9278,N_9516);
nand UO_398 (O_398,N_9302,N_9673);
nand UO_399 (O_399,N_9642,N_9239);
or UO_400 (O_400,N_9394,N_9742);
and UO_401 (O_401,N_9578,N_9192);
or UO_402 (O_402,N_9452,N_9319);
or UO_403 (O_403,N_9052,N_9340);
nor UO_404 (O_404,N_9957,N_9272);
and UO_405 (O_405,N_9563,N_9576);
nor UO_406 (O_406,N_9811,N_9138);
and UO_407 (O_407,N_9824,N_9361);
nand UO_408 (O_408,N_9069,N_9042);
nand UO_409 (O_409,N_9736,N_9739);
nor UO_410 (O_410,N_9218,N_9579);
nor UO_411 (O_411,N_9107,N_9684);
nand UO_412 (O_412,N_9915,N_9559);
nand UO_413 (O_413,N_9001,N_9710);
nand UO_414 (O_414,N_9335,N_9471);
or UO_415 (O_415,N_9926,N_9939);
xor UO_416 (O_416,N_9126,N_9820);
and UO_417 (O_417,N_9631,N_9720);
nor UO_418 (O_418,N_9129,N_9887);
nand UO_419 (O_419,N_9250,N_9174);
or UO_420 (O_420,N_9645,N_9309);
nor UO_421 (O_421,N_9426,N_9365);
or UO_422 (O_422,N_9497,N_9709);
or UO_423 (O_423,N_9629,N_9463);
xnor UO_424 (O_424,N_9735,N_9588);
nor UO_425 (O_425,N_9447,N_9775);
nand UO_426 (O_426,N_9110,N_9768);
or UO_427 (O_427,N_9603,N_9969);
and UO_428 (O_428,N_9894,N_9061);
nand UO_429 (O_429,N_9586,N_9034);
and UO_430 (O_430,N_9931,N_9728);
nand UO_431 (O_431,N_9656,N_9794);
xnor UO_432 (O_432,N_9214,N_9913);
or UO_433 (O_433,N_9419,N_9712);
and UO_434 (O_434,N_9481,N_9517);
nand UO_435 (O_435,N_9200,N_9976);
nand UO_436 (O_436,N_9898,N_9299);
nand UO_437 (O_437,N_9002,N_9183);
and UO_438 (O_438,N_9373,N_9524);
nor UO_439 (O_439,N_9757,N_9231);
and UO_440 (O_440,N_9074,N_9031);
and UO_441 (O_441,N_9372,N_9175);
nand UO_442 (O_442,N_9501,N_9457);
nand UO_443 (O_443,N_9879,N_9773);
and UO_444 (O_444,N_9806,N_9065);
nor UO_445 (O_445,N_9863,N_9968);
or UO_446 (O_446,N_9139,N_9519);
nor UO_447 (O_447,N_9977,N_9600);
or UO_448 (O_448,N_9813,N_9261);
and UO_449 (O_449,N_9591,N_9987);
and UO_450 (O_450,N_9514,N_9098);
nand UO_451 (O_451,N_9243,N_9398);
and UO_452 (O_452,N_9060,N_9916);
nor UO_453 (O_453,N_9605,N_9171);
or UO_454 (O_454,N_9825,N_9467);
nor UO_455 (O_455,N_9538,N_9425);
and UO_456 (O_456,N_9382,N_9185);
and UO_457 (O_457,N_9609,N_9162);
nor UO_458 (O_458,N_9475,N_9216);
or UO_459 (O_459,N_9100,N_9932);
nand UO_460 (O_460,N_9222,N_9115);
nor UO_461 (O_461,N_9512,N_9706);
or UO_462 (O_462,N_9546,N_9482);
xor UO_463 (O_463,N_9551,N_9816);
and UO_464 (O_464,N_9798,N_9083);
nand UO_465 (O_465,N_9118,N_9432);
nor UO_466 (O_466,N_9959,N_9226);
or UO_467 (O_467,N_9173,N_9543);
and UO_468 (O_468,N_9424,N_9221);
or UO_469 (O_469,N_9944,N_9678);
or UO_470 (O_470,N_9095,N_9122);
nand UO_471 (O_471,N_9077,N_9270);
and UO_472 (O_472,N_9282,N_9484);
or UO_473 (O_473,N_9687,N_9599);
nor UO_474 (O_474,N_9016,N_9177);
xor UO_475 (O_475,N_9930,N_9486);
nand UO_476 (O_476,N_9737,N_9168);
and UO_477 (O_477,N_9534,N_9732);
or UO_478 (O_478,N_9499,N_9154);
or UO_479 (O_479,N_9147,N_9677);
nand UO_480 (O_480,N_9290,N_9623);
nor UO_481 (O_481,N_9434,N_9826);
and UO_482 (O_482,N_9458,N_9506);
nor UO_483 (O_483,N_9666,N_9956);
nor UO_484 (O_484,N_9362,N_9644);
xor UO_485 (O_485,N_9035,N_9975);
nand UO_486 (O_486,N_9051,N_9549);
nand UO_487 (O_487,N_9555,N_9622);
nand UO_488 (O_488,N_9201,N_9443);
xnor UO_489 (O_489,N_9504,N_9087);
nor UO_490 (O_490,N_9004,N_9905);
and UO_491 (O_491,N_9360,N_9708);
and UO_492 (O_492,N_9413,N_9614);
nor UO_493 (O_493,N_9109,N_9940);
and UO_494 (O_494,N_9691,N_9127);
nand UO_495 (O_495,N_9520,N_9615);
nor UO_496 (O_496,N_9345,N_9281);
nand UO_497 (O_497,N_9821,N_9612);
nand UO_498 (O_498,N_9059,N_9238);
and UO_499 (O_499,N_9589,N_9883);
xnor UO_500 (O_500,N_9049,N_9602);
and UO_501 (O_501,N_9050,N_9893);
nor UO_502 (O_502,N_9925,N_9073);
nand UO_503 (O_503,N_9080,N_9067);
and UO_504 (O_504,N_9353,N_9192);
and UO_505 (O_505,N_9193,N_9176);
nor UO_506 (O_506,N_9608,N_9775);
nand UO_507 (O_507,N_9838,N_9566);
nor UO_508 (O_508,N_9559,N_9135);
nand UO_509 (O_509,N_9144,N_9111);
or UO_510 (O_510,N_9724,N_9094);
nor UO_511 (O_511,N_9283,N_9006);
nor UO_512 (O_512,N_9493,N_9073);
nor UO_513 (O_513,N_9712,N_9290);
or UO_514 (O_514,N_9784,N_9702);
xor UO_515 (O_515,N_9825,N_9445);
nand UO_516 (O_516,N_9907,N_9048);
or UO_517 (O_517,N_9173,N_9163);
nor UO_518 (O_518,N_9302,N_9287);
nor UO_519 (O_519,N_9053,N_9300);
nor UO_520 (O_520,N_9522,N_9635);
or UO_521 (O_521,N_9380,N_9343);
or UO_522 (O_522,N_9892,N_9192);
and UO_523 (O_523,N_9619,N_9191);
or UO_524 (O_524,N_9850,N_9274);
nor UO_525 (O_525,N_9450,N_9504);
and UO_526 (O_526,N_9427,N_9823);
xor UO_527 (O_527,N_9512,N_9578);
or UO_528 (O_528,N_9475,N_9132);
nor UO_529 (O_529,N_9893,N_9116);
nand UO_530 (O_530,N_9698,N_9667);
nand UO_531 (O_531,N_9566,N_9118);
and UO_532 (O_532,N_9085,N_9301);
nor UO_533 (O_533,N_9458,N_9448);
nand UO_534 (O_534,N_9746,N_9429);
nand UO_535 (O_535,N_9293,N_9709);
or UO_536 (O_536,N_9233,N_9859);
and UO_537 (O_537,N_9925,N_9712);
nand UO_538 (O_538,N_9828,N_9250);
and UO_539 (O_539,N_9647,N_9329);
or UO_540 (O_540,N_9635,N_9508);
xor UO_541 (O_541,N_9181,N_9329);
xnor UO_542 (O_542,N_9114,N_9060);
and UO_543 (O_543,N_9784,N_9667);
or UO_544 (O_544,N_9140,N_9290);
or UO_545 (O_545,N_9205,N_9127);
xor UO_546 (O_546,N_9787,N_9548);
and UO_547 (O_547,N_9625,N_9095);
nand UO_548 (O_548,N_9348,N_9771);
or UO_549 (O_549,N_9015,N_9981);
and UO_550 (O_550,N_9363,N_9875);
xnor UO_551 (O_551,N_9777,N_9438);
xor UO_552 (O_552,N_9675,N_9337);
nand UO_553 (O_553,N_9565,N_9819);
or UO_554 (O_554,N_9949,N_9064);
xnor UO_555 (O_555,N_9120,N_9331);
nand UO_556 (O_556,N_9045,N_9360);
nor UO_557 (O_557,N_9515,N_9772);
nor UO_558 (O_558,N_9086,N_9429);
and UO_559 (O_559,N_9314,N_9118);
nor UO_560 (O_560,N_9904,N_9347);
nand UO_561 (O_561,N_9065,N_9138);
xnor UO_562 (O_562,N_9530,N_9207);
nand UO_563 (O_563,N_9732,N_9784);
or UO_564 (O_564,N_9005,N_9004);
or UO_565 (O_565,N_9180,N_9649);
nand UO_566 (O_566,N_9326,N_9217);
nor UO_567 (O_567,N_9708,N_9119);
xor UO_568 (O_568,N_9470,N_9333);
nand UO_569 (O_569,N_9196,N_9887);
nor UO_570 (O_570,N_9543,N_9675);
and UO_571 (O_571,N_9751,N_9022);
nand UO_572 (O_572,N_9574,N_9857);
nor UO_573 (O_573,N_9135,N_9883);
nand UO_574 (O_574,N_9722,N_9106);
or UO_575 (O_575,N_9848,N_9500);
nand UO_576 (O_576,N_9349,N_9303);
nor UO_577 (O_577,N_9543,N_9210);
or UO_578 (O_578,N_9549,N_9218);
xnor UO_579 (O_579,N_9735,N_9430);
nand UO_580 (O_580,N_9324,N_9057);
nand UO_581 (O_581,N_9655,N_9718);
nor UO_582 (O_582,N_9079,N_9185);
nand UO_583 (O_583,N_9288,N_9227);
and UO_584 (O_584,N_9278,N_9422);
or UO_585 (O_585,N_9616,N_9186);
nor UO_586 (O_586,N_9559,N_9292);
nand UO_587 (O_587,N_9760,N_9146);
nor UO_588 (O_588,N_9336,N_9136);
nor UO_589 (O_589,N_9761,N_9701);
and UO_590 (O_590,N_9833,N_9568);
nand UO_591 (O_591,N_9309,N_9887);
or UO_592 (O_592,N_9904,N_9593);
nand UO_593 (O_593,N_9541,N_9529);
or UO_594 (O_594,N_9573,N_9568);
and UO_595 (O_595,N_9358,N_9351);
nor UO_596 (O_596,N_9140,N_9680);
and UO_597 (O_597,N_9293,N_9261);
and UO_598 (O_598,N_9557,N_9351);
xor UO_599 (O_599,N_9170,N_9175);
xor UO_600 (O_600,N_9508,N_9562);
nor UO_601 (O_601,N_9133,N_9874);
nand UO_602 (O_602,N_9113,N_9100);
or UO_603 (O_603,N_9296,N_9655);
and UO_604 (O_604,N_9328,N_9905);
or UO_605 (O_605,N_9502,N_9452);
xnor UO_606 (O_606,N_9009,N_9791);
and UO_607 (O_607,N_9699,N_9831);
and UO_608 (O_608,N_9886,N_9944);
nor UO_609 (O_609,N_9592,N_9205);
nor UO_610 (O_610,N_9118,N_9986);
nand UO_611 (O_611,N_9464,N_9583);
xnor UO_612 (O_612,N_9476,N_9641);
and UO_613 (O_613,N_9285,N_9527);
nor UO_614 (O_614,N_9590,N_9251);
or UO_615 (O_615,N_9167,N_9126);
nand UO_616 (O_616,N_9142,N_9765);
or UO_617 (O_617,N_9066,N_9733);
nand UO_618 (O_618,N_9059,N_9845);
or UO_619 (O_619,N_9290,N_9728);
nand UO_620 (O_620,N_9889,N_9873);
and UO_621 (O_621,N_9353,N_9938);
or UO_622 (O_622,N_9166,N_9029);
or UO_623 (O_623,N_9681,N_9696);
and UO_624 (O_624,N_9737,N_9162);
nor UO_625 (O_625,N_9107,N_9518);
nand UO_626 (O_626,N_9401,N_9847);
or UO_627 (O_627,N_9806,N_9742);
xnor UO_628 (O_628,N_9979,N_9416);
and UO_629 (O_629,N_9431,N_9301);
or UO_630 (O_630,N_9693,N_9378);
and UO_631 (O_631,N_9659,N_9890);
and UO_632 (O_632,N_9701,N_9269);
nor UO_633 (O_633,N_9003,N_9359);
nor UO_634 (O_634,N_9333,N_9307);
nand UO_635 (O_635,N_9148,N_9304);
and UO_636 (O_636,N_9156,N_9584);
nor UO_637 (O_637,N_9299,N_9469);
or UO_638 (O_638,N_9069,N_9419);
nand UO_639 (O_639,N_9031,N_9868);
or UO_640 (O_640,N_9694,N_9438);
nand UO_641 (O_641,N_9583,N_9861);
and UO_642 (O_642,N_9330,N_9286);
xor UO_643 (O_643,N_9287,N_9165);
or UO_644 (O_644,N_9980,N_9675);
nand UO_645 (O_645,N_9526,N_9980);
nor UO_646 (O_646,N_9863,N_9941);
or UO_647 (O_647,N_9588,N_9904);
nor UO_648 (O_648,N_9708,N_9518);
nor UO_649 (O_649,N_9081,N_9050);
nand UO_650 (O_650,N_9979,N_9413);
nor UO_651 (O_651,N_9057,N_9263);
nor UO_652 (O_652,N_9190,N_9478);
nor UO_653 (O_653,N_9210,N_9658);
or UO_654 (O_654,N_9126,N_9761);
and UO_655 (O_655,N_9168,N_9005);
nand UO_656 (O_656,N_9768,N_9453);
nand UO_657 (O_657,N_9939,N_9500);
or UO_658 (O_658,N_9836,N_9394);
nand UO_659 (O_659,N_9599,N_9851);
or UO_660 (O_660,N_9584,N_9506);
and UO_661 (O_661,N_9168,N_9500);
nand UO_662 (O_662,N_9522,N_9614);
xnor UO_663 (O_663,N_9427,N_9955);
or UO_664 (O_664,N_9025,N_9825);
nand UO_665 (O_665,N_9962,N_9246);
nor UO_666 (O_666,N_9636,N_9922);
and UO_667 (O_667,N_9242,N_9037);
nand UO_668 (O_668,N_9433,N_9096);
xnor UO_669 (O_669,N_9996,N_9671);
nor UO_670 (O_670,N_9585,N_9260);
nand UO_671 (O_671,N_9397,N_9406);
and UO_672 (O_672,N_9738,N_9669);
and UO_673 (O_673,N_9338,N_9232);
nand UO_674 (O_674,N_9234,N_9985);
nand UO_675 (O_675,N_9992,N_9958);
nor UO_676 (O_676,N_9255,N_9290);
nand UO_677 (O_677,N_9527,N_9382);
nor UO_678 (O_678,N_9953,N_9103);
nor UO_679 (O_679,N_9484,N_9160);
and UO_680 (O_680,N_9743,N_9589);
nand UO_681 (O_681,N_9888,N_9030);
nor UO_682 (O_682,N_9002,N_9949);
nand UO_683 (O_683,N_9009,N_9113);
xnor UO_684 (O_684,N_9510,N_9148);
and UO_685 (O_685,N_9967,N_9366);
nor UO_686 (O_686,N_9550,N_9571);
and UO_687 (O_687,N_9842,N_9856);
nor UO_688 (O_688,N_9735,N_9276);
nor UO_689 (O_689,N_9634,N_9373);
nor UO_690 (O_690,N_9524,N_9813);
or UO_691 (O_691,N_9785,N_9534);
and UO_692 (O_692,N_9453,N_9030);
or UO_693 (O_693,N_9001,N_9277);
or UO_694 (O_694,N_9344,N_9559);
nor UO_695 (O_695,N_9399,N_9223);
or UO_696 (O_696,N_9776,N_9938);
or UO_697 (O_697,N_9277,N_9980);
or UO_698 (O_698,N_9486,N_9820);
or UO_699 (O_699,N_9047,N_9636);
and UO_700 (O_700,N_9802,N_9206);
nor UO_701 (O_701,N_9227,N_9911);
or UO_702 (O_702,N_9211,N_9851);
xor UO_703 (O_703,N_9900,N_9696);
nand UO_704 (O_704,N_9784,N_9379);
nor UO_705 (O_705,N_9424,N_9422);
xor UO_706 (O_706,N_9996,N_9577);
or UO_707 (O_707,N_9438,N_9742);
nand UO_708 (O_708,N_9511,N_9086);
and UO_709 (O_709,N_9163,N_9423);
and UO_710 (O_710,N_9514,N_9950);
and UO_711 (O_711,N_9778,N_9777);
nand UO_712 (O_712,N_9056,N_9016);
and UO_713 (O_713,N_9286,N_9871);
and UO_714 (O_714,N_9757,N_9074);
and UO_715 (O_715,N_9789,N_9004);
or UO_716 (O_716,N_9665,N_9520);
and UO_717 (O_717,N_9585,N_9261);
nand UO_718 (O_718,N_9045,N_9654);
nor UO_719 (O_719,N_9197,N_9726);
nand UO_720 (O_720,N_9920,N_9635);
nand UO_721 (O_721,N_9028,N_9899);
or UO_722 (O_722,N_9103,N_9936);
xnor UO_723 (O_723,N_9603,N_9260);
nand UO_724 (O_724,N_9685,N_9651);
or UO_725 (O_725,N_9694,N_9402);
and UO_726 (O_726,N_9595,N_9337);
nand UO_727 (O_727,N_9236,N_9815);
nand UO_728 (O_728,N_9157,N_9386);
and UO_729 (O_729,N_9379,N_9402);
or UO_730 (O_730,N_9901,N_9148);
or UO_731 (O_731,N_9664,N_9078);
and UO_732 (O_732,N_9327,N_9322);
nor UO_733 (O_733,N_9359,N_9772);
or UO_734 (O_734,N_9257,N_9644);
nand UO_735 (O_735,N_9179,N_9334);
nand UO_736 (O_736,N_9392,N_9375);
nor UO_737 (O_737,N_9923,N_9383);
and UO_738 (O_738,N_9034,N_9573);
nand UO_739 (O_739,N_9055,N_9519);
and UO_740 (O_740,N_9529,N_9120);
nor UO_741 (O_741,N_9708,N_9638);
nand UO_742 (O_742,N_9833,N_9009);
xor UO_743 (O_743,N_9458,N_9492);
nor UO_744 (O_744,N_9273,N_9852);
and UO_745 (O_745,N_9826,N_9899);
nor UO_746 (O_746,N_9199,N_9814);
and UO_747 (O_747,N_9026,N_9783);
nand UO_748 (O_748,N_9301,N_9427);
nand UO_749 (O_749,N_9891,N_9282);
nor UO_750 (O_750,N_9508,N_9148);
or UO_751 (O_751,N_9600,N_9800);
or UO_752 (O_752,N_9351,N_9491);
nor UO_753 (O_753,N_9701,N_9848);
xor UO_754 (O_754,N_9881,N_9312);
xor UO_755 (O_755,N_9220,N_9596);
nand UO_756 (O_756,N_9877,N_9752);
and UO_757 (O_757,N_9006,N_9882);
and UO_758 (O_758,N_9391,N_9039);
and UO_759 (O_759,N_9404,N_9008);
or UO_760 (O_760,N_9863,N_9507);
xor UO_761 (O_761,N_9011,N_9398);
nand UO_762 (O_762,N_9841,N_9875);
nor UO_763 (O_763,N_9993,N_9707);
nand UO_764 (O_764,N_9429,N_9504);
nor UO_765 (O_765,N_9823,N_9024);
or UO_766 (O_766,N_9357,N_9143);
nand UO_767 (O_767,N_9442,N_9523);
nand UO_768 (O_768,N_9081,N_9248);
or UO_769 (O_769,N_9251,N_9697);
and UO_770 (O_770,N_9986,N_9586);
nand UO_771 (O_771,N_9943,N_9226);
nand UO_772 (O_772,N_9663,N_9246);
or UO_773 (O_773,N_9109,N_9366);
or UO_774 (O_774,N_9232,N_9968);
or UO_775 (O_775,N_9119,N_9299);
or UO_776 (O_776,N_9134,N_9444);
and UO_777 (O_777,N_9237,N_9220);
nor UO_778 (O_778,N_9511,N_9793);
nor UO_779 (O_779,N_9607,N_9902);
or UO_780 (O_780,N_9735,N_9768);
nand UO_781 (O_781,N_9452,N_9619);
nor UO_782 (O_782,N_9969,N_9891);
nand UO_783 (O_783,N_9603,N_9508);
and UO_784 (O_784,N_9439,N_9082);
and UO_785 (O_785,N_9794,N_9690);
nand UO_786 (O_786,N_9341,N_9047);
or UO_787 (O_787,N_9252,N_9976);
nor UO_788 (O_788,N_9744,N_9705);
and UO_789 (O_789,N_9023,N_9455);
and UO_790 (O_790,N_9060,N_9184);
nor UO_791 (O_791,N_9684,N_9532);
and UO_792 (O_792,N_9929,N_9710);
nand UO_793 (O_793,N_9161,N_9512);
or UO_794 (O_794,N_9609,N_9668);
and UO_795 (O_795,N_9972,N_9018);
and UO_796 (O_796,N_9899,N_9153);
or UO_797 (O_797,N_9572,N_9378);
and UO_798 (O_798,N_9611,N_9980);
nor UO_799 (O_799,N_9309,N_9420);
nand UO_800 (O_800,N_9394,N_9013);
and UO_801 (O_801,N_9426,N_9795);
nand UO_802 (O_802,N_9250,N_9784);
nand UO_803 (O_803,N_9815,N_9750);
nor UO_804 (O_804,N_9563,N_9325);
and UO_805 (O_805,N_9345,N_9672);
nor UO_806 (O_806,N_9609,N_9905);
nand UO_807 (O_807,N_9252,N_9966);
nand UO_808 (O_808,N_9478,N_9937);
and UO_809 (O_809,N_9981,N_9997);
and UO_810 (O_810,N_9924,N_9690);
or UO_811 (O_811,N_9685,N_9432);
xor UO_812 (O_812,N_9332,N_9476);
and UO_813 (O_813,N_9366,N_9757);
and UO_814 (O_814,N_9033,N_9387);
or UO_815 (O_815,N_9179,N_9546);
or UO_816 (O_816,N_9272,N_9563);
nand UO_817 (O_817,N_9161,N_9533);
and UO_818 (O_818,N_9378,N_9487);
and UO_819 (O_819,N_9877,N_9284);
and UO_820 (O_820,N_9430,N_9886);
or UO_821 (O_821,N_9576,N_9969);
nor UO_822 (O_822,N_9589,N_9073);
nor UO_823 (O_823,N_9035,N_9839);
nand UO_824 (O_824,N_9180,N_9706);
nand UO_825 (O_825,N_9728,N_9085);
nor UO_826 (O_826,N_9128,N_9323);
xor UO_827 (O_827,N_9674,N_9962);
nand UO_828 (O_828,N_9370,N_9376);
nand UO_829 (O_829,N_9612,N_9987);
nor UO_830 (O_830,N_9578,N_9342);
and UO_831 (O_831,N_9372,N_9023);
and UO_832 (O_832,N_9373,N_9792);
nand UO_833 (O_833,N_9858,N_9678);
nor UO_834 (O_834,N_9808,N_9773);
nor UO_835 (O_835,N_9139,N_9548);
or UO_836 (O_836,N_9191,N_9480);
nand UO_837 (O_837,N_9787,N_9486);
and UO_838 (O_838,N_9674,N_9394);
nor UO_839 (O_839,N_9522,N_9394);
and UO_840 (O_840,N_9334,N_9069);
nand UO_841 (O_841,N_9328,N_9453);
or UO_842 (O_842,N_9517,N_9459);
nor UO_843 (O_843,N_9912,N_9057);
and UO_844 (O_844,N_9927,N_9966);
nor UO_845 (O_845,N_9959,N_9218);
nand UO_846 (O_846,N_9708,N_9542);
nor UO_847 (O_847,N_9747,N_9392);
nor UO_848 (O_848,N_9392,N_9531);
or UO_849 (O_849,N_9000,N_9163);
or UO_850 (O_850,N_9492,N_9572);
xor UO_851 (O_851,N_9259,N_9253);
xnor UO_852 (O_852,N_9885,N_9612);
and UO_853 (O_853,N_9654,N_9288);
nand UO_854 (O_854,N_9252,N_9540);
nand UO_855 (O_855,N_9935,N_9887);
xor UO_856 (O_856,N_9221,N_9439);
or UO_857 (O_857,N_9362,N_9540);
nor UO_858 (O_858,N_9852,N_9221);
nor UO_859 (O_859,N_9652,N_9706);
and UO_860 (O_860,N_9819,N_9469);
and UO_861 (O_861,N_9959,N_9221);
nand UO_862 (O_862,N_9046,N_9009);
and UO_863 (O_863,N_9506,N_9888);
and UO_864 (O_864,N_9799,N_9810);
or UO_865 (O_865,N_9622,N_9652);
nand UO_866 (O_866,N_9487,N_9889);
or UO_867 (O_867,N_9760,N_9145);
nor UO_868 (O_868,N_9612,N_9735);
nand UO_869 (O_869,N_9448,N_9697);
and UO_870 (O_870,N_9255,N_9666);
or UO_871 (O_871,N_9373,N_9281);
and UO_872 (O_872,N_9892,N_9035);
nor UO_873 (O_873,N_9584,N_9789);
xor UO_874 (O_874,N_9779,N_9330);
xor UO_875 (O_875,N_9539,N_9984);
or UO_876 (O_876,N_9566,N_9290);
xnor UO_877 (O_877,N_9270,N_9297);
and UO_878 (O_878,N_9899,N_9646);
xnor UO_879 (O_879,N_9087,N_9056);
or UO_880 (O_880,N_9192,N_9649);
nand UO_881 (O_881,N_9404,N_9583);
and UO_882 (O_882,N_9248,N_9496);
and UO_883 (O_883,N_9163,N_9309);
or UO_884 (O_884,N_9737,N_9633);
nor UO_885 (O_885,N_9618,N_9564);
nor UO_886 (O_886,N_9075,N_9910);
or UO_887 (O_887,N_9024,N_9726);
nand UO_888 (O_888,N_9329,N_9578);
or UO_889 (O_889,N_9225,N_9181);
or UO_890 (O_890,N_9054,N_9948);
or UO_891 (O_891,N_9520,N_9476);
or UO_892 (O_892,N_9442,N_9827);
or UO_893 (O_893,N_9563,N_9136);
xnor UO_894 (O_894,N_9842,N_9199);
nand UO_895 (O_895,N_9388,N_9878);
nor UO_896 (O_896,N_9948,N_9578);
or UO_897 (O_897,N_9974,N_9319);
or UO_898 (O_898,N_9084,N_9281);
xnor UO_899 (O_899,N_9539,N_9607);
nand UO_900 (O_900,N_9711,N_9762);
nand UO_901 (O_901,N_9206,N_9898);
nand UO_902 (O_902,N_9246,N_9044);
nand UO_903 (O_903,N_9307,N_9384);
or UO_904 (O_904,N_9008,N_9260);
and UO_905 (O_905,N_9581,N_9352);
and UO_906 (O_906,N_9896,N_9382);
nand UO_907 (O_907,N_9935,N_9625);
or UO_908 (O_908,N_9165,N_9926);
nor UO_909 (O_909,N_9055,N_9115);
nand UO_910 (O_910,N_9326,N_9775);
and UO_911 (O_911,N_9601,N_9583);
nand UO_912 (O_912,N_9218,N_9102);
xnor UO_913 (O_913,N_9422,N_9992);
and UO_914 (O_914,N_9812,N_9806);
nand UO_915 (O_915,N_9732,N_9350);
or UO_916 (O_916,N_9982,N_9798);
nand UO_917 (O_917,N_9486,N_9575);
and UO_918 (O_918,N_9102,N_9547);
nor UO_919 (O_919,N_9367,N_9150);
nor UO_920 (O_920,N_9097,N_9268);
nand UO_921 (O_921,N_9012,N_9954);
and UO_922 (O_922,N_9259,N_9826);
nor UO_923 (O_923,N_9278,N_9537);
or UO_924 (O_924,N_9164,N_9906);
and UO_925 (O_925,N_9934,N_9184);
xor UO_926 (O_926,N_9038,N_9042);
nand UO_927 (O_927,N_9208,N_9352);
xor UO_928 (O_928,N_9799,N_9456);
xor UO_929 (O_929,N_9902,N_9094);
nand UO_930 (O_930,N_9014,N_9185);
and UO_931 (O_931,N_9565,N_9292);
or UO_932 (O_932,N_9776,N_9694);
or UO_933 (O_933,N_9862,N_9177);
nand UO_934 (O_934,N_9911,N_9292);
and UO_935 (O_935,N_9644,N_9553);
and UO_936 (O_936,N_9703,N_9672);
nor UO_937 (O_937,N_9676,N_9555);
nand UO_938 (O_938,N_9395,N_9953);
nor UO_939 (O_939,N_9278,N_9126);
or UO_940 (O_940,N_9729,N_9349);
nand UO_941 (O_941,N_9619,N_9846);
nor UO_942 (O_942,N_9907,N_9388);
and UO_943 (O_943,N_9893,N_9565);
or UO_944 (O_944,N_9292,N_9261);
and UO_945 (O_945,N_9304,N_9126);
and UO_946 (O_946,N_9792,N_9236);
xnor UO_947 (O_947,N_9144,N_9517);
nor UO_948 (O_948,N_9943,N_9638);
nor UO_949 (O_949,N_9980,N_9873);
nand UO_950 (O_950,N_9989,N_9146);
nand UO_951 (O_951,N_9917,N_9143);
nand UO_952 (O_952,N_9860,N_9771);
or UO_953 (O_953,N_9065,N_9826);
or UO_954 (O_954,N_9869,N_9082);
and UO_955 (O_955,N_9623,N_9302);
or UO_956 (O_956,N_9447,N_9938);
nand UO_957 (O_957,N_9951,N_9679);
and UO_958 (O_958,N_9448,N_9565);
and UO_959 (O_959,N_9424,N_9302);
nand UO_960 (O_960,N_9727,N_9641);
or UO_961 (O_961,N_9679,N_9305);
and UO_962 (O_962,N_9567,N_9372);
nand UO_963 (O_963,N_9677,N_9668);
xnor UO_964 (O_964,N_9532,N_9390);
or UO_965 (O_965,N_9972,N_9614);
and UO_966 (O_966,N_9902,N_9887);
and UO_967 (O_967,N_9521,N_9825);
nor UO_968 (O_968,N_9137,N_9642);
and UO_969 (O_969,N_9659,N_9738);
xnor UO_970 (O_970,N_9982,N_9570);
xnor UO_971 (O_971,N_9754,N_9256);
or UO_972 (O_972,N_9978,N_9958);
nor UO_973 (O_973,N_9135,N_9197);
or UO_974 (O_974,N_9094,N_9512);
and UO_975 (O_975,N_9455,N_9203);
and UO_976 (O_976,N_9563,N_9574);
or UO_977 (O_977,N_9434,N_9645);
or UO_978 (O_978,N_9875,N_9093);
or UO_979 (O_979,N_9765,N_9170);
and UO_980 (O_980,N_9071,N_9418);
or UO_981 (O_981,N_9686,N_9815);
xnor UO_982 (O_982,N_9773,N_9509);
or UO_983 (O_983,N_9132,N_9110);
xor UO_984 (O_984,N_9020,N_9134);
and UO_985 (O_985,N_9890,N_9196);
nor UO_986 (O_986,N_9805,N_9880);
nor UO_987 (O_987,N_9308,N_9529);
nand UO_988 (O_988,N_9884,N_9857);
nand UO_989 (O_989,N_9919,N_9496);
nor UO_990 (O_990,N_9704,N_9324);
nor UO_991 (O_991,N_9382,N_9470);
and UO_992 (O_992,N_9862,N_9252);
or UO_993 (O_993,N_9008,N_9095);
xor UO_994 (O_994,N_9664,N_9198);
and UO_995 (O_995,N_9997,N_9279);
nor UO_996 (O_996,N_9869,N_9026);
nor UO_997 (O_997,N_9318,N_9877);
xor UO_998 (O_998,N_9038,N_9842);
or UO_999 (O_999,N_9999,N_9517);
or UO_1000 (O_1000,N_9260,N_9932);
xnor UO_1001 (O_1001,N_9521,N_9797);
or UO_1002 (O_1002,N_9690,N_9689);
nor UO_1003 (O_1003,N_9155,N_9938);
xor UO_1004 (O_1004,N_9267,N_9794);
nor UO_1005 (O_1005,N_9915,N_9623);
nand UO_1006 (O_1006,N_9610,N_9320);
nand UO_1007 (O_1007,N_9503,N_9928);
or UO_1008 (O_1008,N_9411,N_9860);
and UO_1009 (O_1009,N_9942,N_9509);
and UO_1010 (O_1010,N_9483,N_9211);
or UO_1011 (O_1011,N_9455,N_9185);
xnor UO_1012 (O_1012,N_9440,N_9102);
and UO_1013 (O_1013,N_9821,N_9841);
nand UO_1014 (O_1014,N_9237,N_9355);
nor UO_1015 (O_1015,N_9611,N_9165);
and UO_1016 (O_1016,N_9956,N_9733);
nand UO_1017 (O_1017,N_9036,N_9209);
and UO_1018 (O_1018,N_9517,N_9249);
nand UO_1019 (O_1019,N_9492,N_9929);
nand UO_1020 (O_1020,N_9018,N_9733);
and UO_1021 (O_1021,N_9492,N_9589);
and UO_1022 (O_1022,N_9250,N_9984);
nor UO_1023 (O_1023,N_9636,N_9987);
nand UO_1024 (O_1024,N_9282,N_9621);
nor UO_1025 (O_1025,N_9201,N_9504);
or UO_1026 (O_1026,N_9090,N_9612);
or UO_1027 (O_1027,N_9657,N_9930);
and UO_1028 (O_1028,N_9646,N_9572);
or UO_1029 (O_1029,N_9504,N_9884);
or UO_1030 (O_1030,N_9077,N_9122);
nand UO_1031 (O_1031,N_9951,N_9760);
or UO_1032 (O_1032,N_9596,N_9738);
or UO_1033 (O_1033,N_9520,N_9139);
nand UO_1034 (O_1034,N_9890,N_9727);
nand UO_1035 (O_1035,N_9868,N_9972);
nor UO_1036 (O_1036,N_9404,N_9300);
or UO_1037 (O_1037,N_9635,N_9095);
and UO_1038 (O_1038,N_9996,N_9118);
and UO_1039 (O_1039,N_9818,N_9373);
and UO_1040 (O_1040,N_9375,N_9035);
or UO_1041 (O_1041,N_9158,N_9035);
nor UO_1042 (O_1042,N_9625,N_9052);
xnor UO_1043 (O_1043,N_9773,N_9361);
and UO_1044 (O_1044,N_9682,N_9423);
nand UO_1045 (O_1045,N_9861,N_9962);
and UO_1046 (O_1046,N_9895,N_9425);
and UO_1047 (O_1047,N_9840,N_9344);
or UO_1048 (O_1048,N_9192,N_9618);
and UO_1049 (O_1049,N_9125,N_9885);
xor UO_1050 (O_1050,N_9216,N_9400);
nor UO_1051 (O_1051,N_9884,N_9653);
nor UO_1052 (O_1052,N_9928,N_9262);
nor UO_1053 (O_1053,N_9803,N_9238);
xnor UO_1054 (O_1054,N_9701,N_9854);
and UO_1055 (O_1055,N_9583,N_9944);
or UO_1056 (O_1056,N_9163,N_9077);
nor UO_1057 (O_1057,N_9622,N_9502);
or UO_1058 (O_1058,N_9912,N_9182);
or UO_1059 (O_1059,N_9444,N_9886);
nor UO_1060 (O_1060,N_9980,N_9189);
nor UO_1061 (O_1061,N_9173,N_9116);
or UO_1062 (O_1062,N_9222,N_9618);
nor UO_1063 (O_1063,N_9560,N_9643);
or UO_1064 (O_1064,N_9693,N_9737);
xor UO_1065 (O_1065,N_9643,N_9658);
nor UO_1066 (O_1066,N_9952,N_9119);
nand UO_1067 (O_1067,N_9550,N_9651);
or UO_1068 (O_1068,N_9254,N_9793);
or UO_1069 (O_1069,N_9588,N_9835);
nor UO_1070 (O_1070,N_9498,N_9913);
or UO_1071 (O_1071,N_9438,N_9155);
nor UO_1072 (O_1072,N_9825,N_9814);
and UO_1073 (O_1073,N_9724,N_9126);
nor UO_1074 (O_1074,N_9926,N_9861);
or UO_1075 (O_1075,N_9018,N_9056);
or UO_1076 (O_1076,N_9127,N_9904);
nand UO_1077 (O_1077,N_9679,N_9359);
and UO_1078 (O_1078,N_9165,N_9177);
or UO_1079 (O_1079,N_9004,N_9328);
and UO_1080 (O_1080,N_9970,N_9193);
or UO_1081 (O_1081,N_9150,N_9227);
nand UO_1082 (O_1082,N_9688,N_9244);
nor UO_1083 (O_1083,N_9911,N_9434);
nand UO_1084 (O_1084,N_9876,N_9273);
nor UO_1085 (O_1085,N_9206,N_9251);
or UO_1086 (O_1086,N_9657,N_9323);
or UO_1087 (O_1087,N_9508,N_9374);
nor UO_1088 (O_1088,N_9185,N_9478);
nor UO_1089 (O_1089,N_9696,N_9212);
nor UO_1090 (O_1090,N_9420,N_9424);
nor UO_1091 (O_1091,N_9916,N_9865);
and UO_1092 (O_1092,N_9722,N_9094);
nand UO_1093 (O_1093,N_9310,N_9783);
and UO_1094 (O_1094,N_9465,N_9495);
and UO_1095 (O_1095,N_9251,N_9964);
nor UO_1096 (O_1096,N_9132,N_9470);
and UO_1097 (O_1097,N_9621,N_9847);
nand UO_1098 (O_1098,N_9483,N_9112);
or UO_1099 (O_1099,N_9691,N_9436);
and UO_1100 (O_1100,N_9747,N_9173);
nor UO_1101 (O_1101,N_9618,N_9253);
and UO_1102 (O_1102,N_9663,N_9571);
nor UO_1103 (O_1103,N_9455,N_9747);
nor UO_1104 (O_1104,N_9342,N_9817);
and UO_1105 (O_1105,N_9455,N_9221);
nand UO_1106 (O_1106,N_9934,N_9083);
nand UO_1107 (O_1107,N_9104,N_9630);
or UO_1108 (O_1108,N_9885,N_9256);
and UO_1109 (O_1109,N_9182,N_9389);
nand UO_1110 (O_1110,N_9546,N_9142);
nand UO_1111 (O_1111,N_9373,N_9870);
or UO_1112 (O_1112,N_9557,N_9518);
and UO_1113 (O_1113,N_9833,N_9645);
nor UO_1114 (O_1114,N_9300,N_9117);
nor UO_1115 (O_1115,N_9630,N_9249);
or UO_1116 (O_1116,N_9749,N_9057);
or UO_1117 (O_1117,N_9038,N_9887);
and UO_1118 (O_1118,N_9135,N_9368);
nand UO_1119 (O_1119,N_9905,N_9626);
nand UO_1120 (O_1120,N_9948,N_9759);
or UO_1121 (O_1121,N_9619,N_9089);
or UO_1122 (O_1122,N_9240,N_9783);
nand UO_1123 (O_1123,N_9668,N_9997);
nand UO_1124 (O_1124,N_9486,N_9552);
nand UO_1125 (O_1125,N_9735,N_9762);
nand UO_1126 (O_1126,N_9656,N_9795);
or UO_1127 (O_1127,N_9745,N_9592);
nand UO_1128 (O_1128,N_9935,N_9501);
xnor UO_1129 (O_1129,N_9431,N_9310);
and UO_1130 (O_1130,N_9307,N_9550);
nor UO_1131 (O_1131,N_9435,N_9167);
nor UO_1132 (O_1132,N_9515,N_9289);
and UO_1133 (O_1133,N_9306,N_9451);
nor UO_1134 (O_1134,N_9921,N_9987);
or UO_1135 (O_1135,N_9645,N_9429);
nand UO_1136 (O_1136,N_9782,N_9165);
nor UO_1137 (O_1137,N_9813,N_9830);
or UO_1138 (O_1138,N_9564,N_9738);
and UO_1139 (O_1139,N_9019,N_9132);
nand UO_1140 (O_1140,N_9430,N_9825);
nand UO_1141 (O_1141,N_9361,N_9789);
and UO_1142 (O_1142,N_9099,N_9934);
or UO_1143 (O_1143,N_9155,N_9337);
and UO_1144 (O_1144,N_9698,N_9543);
nor UO_1145 (O_1145,N_9704,N_9154);
or UO_1146 (O_1146,N_9840,N_9642);
or UO_1147 (O_1147,N_9350,N_9110);
nand UO_1148 (O_1148,N_9526,N_9631);
nand UO_1149 (O_1149,N_9382,N_9243);
and UO_1150 (O_1150,N_9521,N_9502);
nor UO_1151 (O_1151,N_9229,N_9696);
nand UO_1152 (O_1152,N_9892,N_9842);
nand UO_1153 (O_1153,N_9671,N_9500);
and UO_1154 (O_1154,N_9681,N_9987);
nand UO_1155 (O_1155,N_9765,N_9705);
and UO_1156 (O_1156,N_9477,N_9654);
and UO_1157 (O_1157,N_9913,N_9531);
xor UO_1158 (O_1158,N_9580,N_9702);
and UO_1159 (O_1159,N_9243,N_9412);
or UO_1160 (O_1160,N_9713,N_9884);
or UO_1161 (O_1161,N_9591,N_9198);
nor UO_1162 (O_1162,N_9958,N_9670);
nor UO_1163 (O_1163,N_9046,N_9052);
nor UO_1164 (O_1164,N_9554,N_9644);
nor UO_1165 (O_1165,N_9178,N_9978);
nand UO_1166 (O_1166,N_9415,N_9971);
or UO_1167 (O_1167,N_9103,N_9675);
or UO_1168 (O_1168,N_9775,N_9367);
xor UO_1169 (O_1169,N_9467,N_9204);
nand UO_1170 (O_1170,N_9854,N_9722);
nand UO_1171 (O_1171,N_9816,N_9569);
nand UO_1172 (O_1172,N_9239,N_9753);
xor UO_1173 (O_1173,N_9379,N_9638);
and UO_1174 (O_1174,N_9632,N_9628);
nor UO_1175 (O_1175,N_9921,N_9966);
and UO_1176 (O_1176,N_9086,N_9603);
or UO_1177 (O_1177,N_9253,N_9708);
nor UO_1178 (O_1178,N_9009,N_9765);
and UO_1179 (O_1179,N_9206,N_9827);
nor UO_1180 (O_1180,N_9000,N_9389);
nand UO_1181 (O_1181,N_9964,N_9018);
or UO_1182 (O_1182,N_9781,N_9501);
nor UO_1183 (O_1183,N_9310,N_9694);
xnor UO_1184 (O_1184,N_9042,N_9255);
and UO_1185 (O_1185,N_9272,N_9600);
or UO_1186 (O_1186,N_9328,N_9540);
and UO_1187 (O_1187,N_9575,N_9891);
nand UO_1188 (O_1188,N_9728,N_9098);
nor UO_1189 (O_1189,N_9048,N_9634);
or UO_1190 (O_1190,N_9998,N_9289);
and UO_1191 (O_1191,N_9465,N_9219);
or UO_1192 (O_1192,N_9103,N_9025);
nand UO_1193 (O_1193,N_9068,N_9417);
nand UO_1194 (O_1194,N_9713,N_9005);
xor UO_1195 (O_1195,N_9358,N_9266);
nor UO_1196 (O_1196,N_9161,N_9732);
and UO_1197 (O_1197,N_9468,N_9933);
or UO_1198 (O_1198,N_9494,N_9222);
nor UO_1199 (O_1199,N_9345,N_9018);
and UO_1200 (O_1200,N_9062,N_9555);
and UO_1201 (O_1201,N_9486,N_9554);
nand UO_1202 (O_1202,N_9223,N_9445);
or UO_1203 (O_1203,N_9319,N_9050);
xnor UO_1204 (O_1204,N_9047,N_9048);
or UO_1205 (O_1205,N_9144,N_9622);
or UO_1206 (O_1206,N_9362,N_9048);
nand UO_1207 (O_1207,N_9409,N_9767);
or UO_1208 (O_1208,N_9137,N_9332);
or UO_1209 (O_1209,N_9017,N_9714);
nor UO_1210 (O_1210,N_9928,N_9376);
nand UO_1211 (O_1211,N_9154,N_9647);
or UO_1212 (O_1212,N_9226,N_9106);
or UO_1213 (O_1213,N_9358,N_9262);
nand UO_1214 (O_1214,N_9868,N_9142);
and UO_1215 (O_1215,N_9538,N_9111);
nand UO_1216 (O_1216,N_9191,N_9721);
and UO_1217 (O_1217,N_9025,N_9990);
or UO_1218 (O_1218,N_9782,N_9347);
xnor UO_1219 (O_1219,N_9193,N_9683);
nand UO_1220 (O_1220,N_9993,N_9921);
nor UO_1221 (O_1221,N_9397,N_9374);
or UO_1222 (O_1222,N_9158,N_9615);
and UO_1223 (O_1223,N_9182,N_9003);
nand UO_1224 (O_1224,N_9636,N_9868);
or UO_1225 (O_1225,N_9926,N_9089);
or UO_1226 (O_1226,N_9491,N_9071);
nand UO_1227 (O_1227,N_9228,N_9704);
nor UO_1228 (O_1228,N_9460,N_9342);
xor UO_1229 (O_1229,N_9755,N_9873);
and UO_1230 (O_1230,N_9197,N_9953);
nor UO_1231 (O_1231,N_9602,N_9052);
or UO_1232 (O_1232,N_9804,N_9516);
or UO_1233 (O_1233,N_9628,N_9000);
and UO_1234 (O_1234,N_9334,N_9636);
xnor UO_1235 (O_1235,N_9085,N_9259);
nor UO_1236 (O_1236,N_9102,N_9036);
and UO_1237 (O_1237,N_9799,N_9071);
and UO_1238 (O_1238,N_9838,N_9003);
and UO_1239 (O_1239,N_9648,N_9234);
nor UO_1240 (O_1240,N_9802,N_9323);
and UO_1241 (O_1241,N_9475,N_9771);
xor UO_1242 (O_1242,N_9742,N_9905);
or UO_1243 (O_1243,N_9766,N_9572);
nand UO_1244 (O_1244,N_9186,N_9916);
or UO_1245 (O_1245,N_9863,N_9784);
or UO_1246 (O_1246,N_9974,N_9914);
and UO_1247 (O_1247,N_9821,N_9596);
and UO_1248 (O_1248,N_9631,N_9811);
or UO_1249 (O_1249,N_9082,N_9435);
or UO_1250 (O_1250,N_9382,N_9922);
or UO_1251 (O_1251,N_9828,N_9139);
nor UO_1252 (O_1252,N_9040,N_9050);
nor UO_1253 (O_1253,N_9626,N_9270);
nor UO_1254 (O_1254,N_9605,N_9184);
nand UO_1255 (O_1255,N_9688,N_9485);
nor UO_1256 (O_1256,N_9752,N_9560);
and UO_1257 (O_1257,N_9947,N_9172);
or UO_1258 (O_1258,N_9212,N_9289);
or UO_1259 (O_1259,N_9571,N_9762);
xor UO_1260 (O_1260,N_9690,N_9956);
nor UO_1261 (O_1261,N_9232,N_9667);
nand UO_1262 (O_1262,N_9654,N_9246);
nand UO_1263 (O_1263,N_9055,N_9359);
nand UO_1264 (O_1264,N_9177,N_9478);
or UO_1265 (O_1265,N_9576,N_9116);
xnor UO_1266 (O_1266,N_9411,N_9327);
nand UO_1267 (O_1267,N_9972,N_9246);
and UO_1268 (O_1268,N_9656,N_9124);
and UO_1269 (O_1269,N_9834,N_9005);
or UO_1270 (O_1270,N_9144,N_9521);
and UO_1271 (O_1271,N_9886,N_9038);
nor UO_1272 (O_1272,N_9205,N_9100);
nor UO_1273 (O_1273,N_9842,N_9719);
or UO_1274 (O_1274,N_9266,N_9817);
nor UO_1275 (O_1275,N_9088,N_9826);
nor UO_1276 (O_1276,N_9870,N_9248);
or UO_1277 (O_1277,N_9854,N_9582);
xnor UO_1278 (O_1278,N_9033,N_9671);
nor UO_1279 (O_1279,N_9210,N_9467);
nor UO_1280 (O_1280,N_9689,N_9839);
and UO_1281 (O_1281,N_9920,N_9423);
and UO_1282 (O_1282,N_9922,N_9642);
or UO_1283 (O_1283,N_9223,N_9597);
nor UO_1284 (O_1284,N_9174,N_9100);
nand UO_1285 (O_1285,N_9247,N_9085);
and UO_1286 (O_1286,N_9234,N_9399);
or UO_1287 (O_1287,N_9250,N_9979);
and UO_1288 (O_1288,N_9816,N_9560);
nor UO_1289 (O_1289,N_9393,N_9341);
xnor UO_1290 (O_1290,N_9265,N_9964);
or UO_1291 (O_1291,N_9639,N_9758);
xor UO_1292 (O_1292,N_9290,N_9358);
and UO_1293 (O_1293,N_9857,N_9414);
nor UO_1294 (O_1294,N_9714,N_9110);
and UO_1295 (O_1295,N_9362,N_9025);
and UO_1296 (O_1296,N_9298,N_9944);
xnor UO_1297 (O_1297,N_9044,N_9412);
and UO_1298 (O_1298,N_9620,N_9703);
or UO_1299 (O_1299,N_9959,N_9176);
nor UO_1300 (O_1300,N_9112,N_9896);
xnor UO_1301 (O_1301,N_9221,N_9194);
nor UO_1302 (O_1302,N_9304,N_9567);
nor UO_1303 (O_1303,N_9100,N_9494);
nor UO_1304 (O_1304,N_9850,N_9380);
nor UO_1305 (O_1305,N_9477,N_9563);
nand UO_1306 (O_1306,N_9072,N_9185);
nand UO_1307 (O_1307,N_9158,N_9784);
and UO_1308 (O_1308,N_9824,N_9007);
and UO_1309 (O_1309,N_9668,N_9302);
or UO_1310 (O_1310,N_9534,N_9592);
and UO_1311 (O_1311,N_9322,N_9739);
nor UO_1312 (O_1312,N_9767,N_9205);
or UO_1313 (O_1313,N_9385,N_9818);
nor UO_1314 (O_1314,N_9332,N_9470);
nand UO_1315 (O_1315,N_9788,N_9519);
nor UO_1316 (O_1316,N_9728,N_9507);
nand UO_1317 (O_1317,N_9936,N_9564);
nor UO_1318 (O_1318,N_9223,N_9912);
or UO_1319 (O_1319,N_9427,N_9428);
nand UO_1320 (O_1320,N_9919,N_9989);
nand UO_1321 (O_1321,N_9407,N_9449);
and UO_1322 (O_1322,N_9974,N_9766);
nand UO_1323 (O_1323,N_9760,N_9772);
nand UO_1324 (O_1324,N_9362,N_9509);
nand UO_1325 (O_1325,N_9027,N_9497);
nand UO_1326 (O_1326,N_9458,N_9284);
and UO_1327 (O_1327,N_9786,N_9876);
or UO_1328 (O_1328,N_9241,N_9194);
and UO_1329 (O_1329,N_9489,N_9749);
or UO_1330 (O_1330,N_9221,N_9349);
xnor UO_1331 (O_1331,N_9406,N_9905);
nand UO_1332 (O_1332,N_9661,N_9347);
nand UO_1333 (O_1333,N_9396,N_9183);
or UO_1334 (O_1334,N_9374,N_9263);
and UO_1335 (O_1335,N_9445,N_9496);
nor UO_1336 (O_1336,N_9389,N_9122);
nor UO_1337 (O_1337,N_9458,N_9872);
and UO_1338 (O_1338,N_9370,N_9849);
nor UO_1339 (O_1339,N_9507,N_9780);
or UO_1340 (O_1340,N_9219,N_9917);
or UO_1341 (O_1341,N_9068,N_9182);
xnor UO_1342 (O_1342,N_9670,N_9539);
and UO_1343 (O_1343,N_9102,N_9731);
nand UO_1344 (O_1344,N_9031,N_9663);
nand UO_1345 (O_1345,N_9272,N_9323);
and UO_1346 (O_1346,N_9365,N_9766);
or UO_1347 (O_1347,N_9711,N_9430);
or UO_1348 (O_1348,N_9676,N_9596);
or UO_1349 (O_1349,N_9740,N_9356);
nand UO_1350 (O_1350,N_9763,N_9327);
and UO_1351 (O_1351,N_9781,N_9776);
nand UO_1352 (O_1352,N_9901,N_9838);
and UO_1353 (O_1353,N_9467,N_9033);
and UO_1354 (O_1354,N_9734,N_9532);
nor UO_1355 (O_1355,N_9844,N_9275);
nor UO_1356 (O_1356,N_9421,N_9930);
nand UO_1357 (O_1357,N_9374,N_9839);
nor UO_1358 (O_1358,N_9060,N_9705);
nor UO_1359 (O_1359,N_9951,N_9568);
nand UO_1360 (O_1360,N_9085,N_9895);
nand UO_1361 (O_1361,N_9672,N_9022);
and UO_1362 (O_1362,N_9604,N_9655);
nand UO_1363 (O_1363,N_9241,N_9855);
and UO_1364 (O_1364,N_9420,N_9711);
nor UO_1365 (O_1365,N_9315,N_9897);
and UO_1366 (O_1366,N_9023,N_9694);
xnor UO_1367 (O_1367,N_9874,N_9598);
or UO_1368 (O_1368,N_9889,N_9416);
nor UO_1369 (O_1369,N_9953,N_9700);
and UO_1370 (O_1370,N_9793,N_9825);
xor UO_1371 (O_1371,N_9949,N_9136);
nand UO_1372 (O_1372,N_9427,N_9594);
nand UO_1373 (O_1373,N_9061,N_9064);
nor UO_1374 (O_1374,N_9692,N_9301);
nor UO_1375 (O_1375,N_9970,N_9198);
and UO_1376 (O_1376,N_9976,N_9984);
xor UO_1377 (O_1377,N_9513,N_9882);
nand UO_1378 (O_1378,N_9011,N_9554);
nor UO_1379 (O_1379,N_9716,N_9317);
and UO_1380 (O_1380,N_9398,N_9663);
or UO_1381 (O_1381,N_9269,N_9929);
and UO_1382 (O_1382,N_9684,N_9111);
xor UO_1383 (O_1383,N_9186,N_9554);
or UO_1384 (O_1384,N_9735,N_9253);
nand UO_1385 (O_1385,N_9861,N_9819);
or UO_1386 (O_1386,N_9328,N_9245);
and UO_1387 (O_1387,N_9994,N_9503);
xnor UO_1388 (O_1388,N_9305,N_9367);
and UO_1389 (O_1389,N_9408,N_9931);
nor UO_1390 (O_1390,N_9309,N_9508);
and UO_1391 (O_1391,N_9781,N_9127);
nand UO_1392 (O_1392,N_9632,N_9930);
or UO_1393 (O_1393,N_9130,N_9592);
or UO_1394 (O_1394,N_9615,N_9023);
and UO_1395 (O_1395,N_9961,N_9441);
and UO_1396 (O_1396,N_9986,N_9994);
and UO_1397 (O_1397,N_9417,N_9689);
or UO_1398 (O_1398,N_9793,N_9638);
nor UO_1399 (O_1399,N_9468,N_9451);
and UO_1400 (O_1400,N_9949,N_9848);
and UO_1401 (O_1401,N_9896,N_9949);
and UO_1402 (O_1402,N_9155,N_9585);
nor UO_1403 (O_1403,N_9865,N_9164);
and UO_1404 (O_1404,N_9375,N_9002);
and UO_1405 (O_1405,N_9595,N_9044);
and UO_1406 (O_1406,N_9015,N_9068);
or UO_1407 (O_1407,N_9936,N_9455);
and UO_1408 (O_1408,N_9860,N_9020);
and UO_1409 (O_1409,N_9789,N_9041);
nor UO_1410 (O_1410,N_9695,N_9256);
nor UO_1411 (O_1411,N_9920,N_9684);
nor UO_1412 (O_1412,N_9285,N_9553);
xor UO_1413 (O_1413,N_9476,N_9338);
nor UO_1414 (O_1414,N_9322,N_9915);
nor UO_1415 (O_1415,N_9551,N_9141);
xor UO_1416 (O_1416,N_9659,N_9279);
or UO_1417 (O_1417,N_9082,N_9104);
and UO_1418 (O_1418,N_9479,N_9102);
or UO_1419 (O_1419,N_9124,N_9512);
nor UO_1420 (O_1420,N_9642,N_9940);
xnor UO_1421 (O_1421,N_9429,N_9628);
and UO_1422 (O_1422,N_9093,N_9593);
nor UO_1423 (O_1423,N_9335,N_9049);
and UO_1424 (O_1424,N_9276,N_9533);
xnor UO_1425 (O_1425,N_9987,N_9162);
and UO_1426 (O_1426,N_9916,N_9619);
nor UO_1427 (O_1427,N_9713,N_9199);
and UO_1428 (O_1428,N_9466,N_9571);
nor UO_1429 (O_1429,N_9954,N_9378);
or UO_1430 (O_1430,N_9340,N_9653);
nand UO_1431 (O_1431,N_9219,N_9367);
nor UO_1432 (O_1432,N_9116,N_9024);
xnor UO_1433 (O_1433,N_9940,N_9266);
nand UO_1434 (O_1434,N_9992,N_9841);
and UO_1435 (O_1435,N_9351,N_9680);
xnor UO_1436 (O_1436,N_9187,N_9664);
and UO_1437 (O_1437,N_9255,N_9074);
nor UO_1438 (O_1438,N_9281,N_9250);
and UO_1439 (O_1439,N_9879,N_9259);
xor UO_1440 (O_1440,N_9754,N_9508);
or UO_1441 (O_1441,N_9302,N_9496);
nor UO_1442 (O_1442,N_9737,N_9754);
xnor UO_1443 (O_1443,N_9184,N_9722);
and UO_1444 (O_1444,N_9075,N_9355);
nor UO_1445 (O_1445,N_9431,N_9253);
and UO_1446 (O_1446,N_9065,N_9829);
nand UO_1447 (O_1447,N_9513,N_9694);
xnor UO_1448 (O_1448,N_9526,N_9650);
nor UO_1449 (O_1449,N_9481,N_9628);
nand UO_1450 (O_1450,N_9001,N_9977);
and UO_1451 (O_1451,N_9618,N_9693);
nor UO_1452 (O_1452,N_9064,N_9151);
and UO_1453 (O_1453,N_9867,N_9762);
nor UO_1454 (O_1454,N_9407,N_9967);
and UO_1455 (O_1455,N_9999,N_9900);
or UO_1456 (O_1456,N_9469,N_9911);
or UO_1457 (O_1457,N_9316,N_9903);
xnor UO_1458 (O_1458,N_9841,N_9768);
nor UO_1459 (O_1459,N_9958,N_9872);
or UO_1460 (O_1460,N_9246,N_9417);
and UO_1461 (O_1461,N_9324,N_9098);
or UO_1462 (O_1462,N_9836,N_9954);
nor UO_1463 (O_1463,N_9095,N_9874);
or UO_1464 (O_1464,N_9903,N_9386);
nor UO_1465 (O_1465,N_9125,N_9545);
nand UO_1466 (O_1466,N_9279,N_9890);
or UO_1467 (O_1467,N_9882,N_9428);
nor UO_1468 (O_1468,N_9890,N_9840);
xor UO_1469 (O_1469,N_9667,N_9758);
xor UO_1470 (O_1470,N_9941,N_9768);
nand UO_1471 (O_1471,N_9223,N_9669);
and UO_1472 (O_1472,N_9498,N_9370);
nand UO_1473 (O_1473,N_9503,N_9655);
or UO_1474 (O_1474,N_9482,N_9429);
nand UO_1475 (O_1475,N_9075,N_9123);
nor UO_1476 (O_1476,N_9138,N_9759);
or UO_1477 (O_1477,N_9297,N_9962);
nand UO_1478 (O_1478,N_9423,N_9146);
nor UO_1479 (O_1479,N_9284,N_9631);
and UO_1480 (O_1480,N_9098,N_9731);
and UO_1481 (O_1481,N_9903,N_9430);
nor UO_1482 (O_1482,N_9782,N_9781);
nand UO_1483 (O_1483,N_9990,N_9141);
or UO_1484 (O_1484,N_9593,N_9798);
or UO_1485 (O_1485,N_9265,N_9127);
nand UO_1486 (O_1486,N_9961,N_9904);
nor UO_1487 (O_1487,N_9429,N_9045);
nand UO_1488 (O_1488,N_9428,N_9259);
nand UO_1489 (O_1489,N_9110,N_9117);
or UO_1490 (O_1490,N_9836,N_9790);
nand UO_1491 (O_1491,N_9764,N_9631);
and UO_1492 (O_1492,N_9843,N_9746);
or UO_1493 (O_1493,N_9981,N_9716);
xnor UO_1494 (O_1494,N_9348,N_9342);
nand UO_1495 (O_1495,N_9651,N_9472);
and UO_1496 (O_1496,N_9017,N_9079);
and UO_1497 (O_1497,N_9418,N_9430);
and UO_1498 (O_1498,N_9364,N_9162);
and UO_1499 (O_1499,N_9658,N_9286);
endmodule