module basic_750_5000_1000_50_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_232,In_93);
nor U1 (N_1,In_581,In_181);
nor U2 (N_2,In_452,In_360);
nor U3 (N_3,In_578,In_545);
or U4 (N_4,In_561,In_251);
or U5 (N_5,In_107,In_285);
xor U6 (N_6,In_229,In_341);
and U7 (N_7,In_27,In_701);
xnor U8 (N_8,In_128,In_358);
and U9 (N_9,In_306,In_391);
nand U10 (N_10,In_161,In_156);
and U11 (N_11,In_670,In_470);
and U12 (N_12,In_237,In_318);
nor U13 (N_13,In_130,In_323);
and U14 (N_14,In_515,In_523);
nor U15 (N_15,In_176,In_448);
nor U16 (N_16,In_586,In_335);
nand U17 (N_17,In_2,In_34);
and U18 (N_18,In_673,In_635);
nor U19 (N_19,In_148,In_377);
and U20 (N_20,In_589,In_608);
nor U21 (N_21,In_493,In_423);
nor U22 (N_22,In_276,In_469);
nand U23 (N_23,In_268,In_711);
and U24 (N_24,In_173,In_398);
nor U25 (N_25,In_567,In_612);
xor U26 (N_26,In_476,In_544);
nand U27 (N_27,In_10,In_81);
and U28 (N_28,In_265,In_228);
xnor U29 (N_29,In_208,In_63);
nand U30 (N_30,In_668,In_112);
or U31 (N_31,In_693,In_409);
nand U32 (N_32,In_244,In_273);
xnor U33 (N_33,In_82,In_392);
or U34 (N_34,In_147,In_304);
and U35 (N_35,In_433,In_205);
and U36 (N_36,In_464,In_362);
and U37 (N_37,In_291,In_256);
nor U38 (N_38,In_631,In_399);
nor U39 (N_39,In_337,In_346);
xor U40 (N_40,In_692,In_85);
nor U41 (N_41,In_332,In_472);
nand U42 (N_42,In_384,In_97);
and U43 (N_43,In_35,In_51);
and U44 (N_44,In_704,In_21);
or U45 (N_45,In_108,In_569);
and U46 (N_46,In_109,In_465);
xnor U47 (N_47,In_488,In_595);
nand U48 (N_48,In_184,In_553);
nand U49 (N_49,In_623,In_720);
and U50 (N_50,In_618,In_422);
nor U51 (N_51,In_301,In_633);
xor U52 (N_52,In_94,In_497);
and U53 (N_53,In_83,In_560);
nand U54 (N_54,In_46,In_695);
or U55 (N_55,In_606,In_400);
nand U56 (N_56,In_307,In_709);
nor U57 (N_57,In_52,In_290);
xnor U58 (N_58,In_235,In_659);
nand U59 (N_59,In_505,In_15);
nand U60 (N_60,In_619,In_137);
xnor U61 (N_61,In_30,In_463);
or U62 (N_62,In_520,In_461);
nor U63 (N_63,In_195,In_177);
and U64 (N_64,In_654,In_738);
nor U65 (N_65,In_729,In_639);
xnor U66 (N_66,In_115,In_458);
nand U67 (N_67,In_253,In_707);
nand U68 (N_68,In_664,In_548);
nor U69 (N_69,In_343,In_604);
or U70 (N_70,In_79,In_165);
and U71 (N_71,In_313,In_363);
or U72 (N_72,In_694,In_153);
and U73 (N_73,In_54,In_474);
or U74 (N_74,In_473,In_716);
nand U75 (N_75,In_4,In_5);
nor U76 (N_76,In_224,In_684);
or U77 (N_77,In_727,In_271);
nor U78 (N_78,In_340,In_640);
or U79 (N_79,In_401,In_376);
xnor U80 (N_80,In_518,In_70);
nand U81 (N_81,In_60,In_282);
xor U82 (N_82,In_522,In_577);
nand U83 (N_83,In_23,In_55);
nand U84 (N_84,In_28,In_598);
or U85 (N_85,In_555,In_566);
or U86 (N_86,In_141,In_725);
nand U87 (N_87,In_215,In_713);
or U88 (N_88,In_95,In_140);
nor U89 (N_89,In_226,In_286);
xnor U90 (N_90,In_733,In_585);
or U91 (N_91,In_104,In_26);
xnor U92 (N_92,In_33,In_502);
nand U93 (N_93,In_499,In_267);
or U94 (N_94,In_76,In_186);
xnor U95 (N_95,In_272,In_39);
or U96 (N_96,In_219,In_180);
xor U97 (N_97,In_411,In_702);
and U98 (N_98,In_397,In_258);
or U99 (N_99,In_353,In_266);
or U100 (N_100,In_428,In_621);
nor U101 (N_101,N_12,In_672);
or U102 (N_102,In_432,In_526);
nand U103 (N_103,In_248,In_718);
or U104 (N_104,In_152,In_201);
nor U105 (N_105,In_274,In_333);
nand U106 (N_106,In_536,In_216);
and U107 (N_107,In_281,In_622);
and U108 (N_108,N_74,In_642);
nand U109 (N_109,In_559,In_390);
nand U110 (N_110,In_414,N_69);
nand U111 (N_111,In_434,In_185);
nor U112 (N_112,In_749,In_261);
and U113 (N_113,In_513,In_349);
nand U114 (N_114,In_20,In_435);
nand U115 (N_115,In_416,In_468);
xor U116 (N_116,In_731,In_671);
xor U117 (N_117,In_457,In_375);
nor U118 (N_118,In_573,In_591);
and U119 (N_119,N_2,In_431);
and U120 (N_120,N_33,N_10);
and U121 (N_121,In_171,N_55);
and U122 (N_122,In_239,In_86);
xor U123 (N_123,In_596,N_3);
nor U124 (N_124,In_269,In_351);
and U125 (N_125,In_212,In_601);
nor U126 (N_126,In_501,In_649);
and U127 (N_127,N_67,In_31);
and U128 (N_128,In_644,In_84);
nor U129 (N_129,N_52,In_734);
or U130 (N_130,N_29,In_225);
or U131 (N_131,In_78,In_627);
nand U132 (N_132,N_41,In_344);
xnor U133 (N_133,In_645,In_188);
nor U134 (N_134,In_710,In_582);
xor U135 (N_135,In_588,In_125);
and U136 (N_136,In_41,N_25);
nand U137 (N_137,In_223,In_724);
and U138 (N_138,In_617,In_355);
nand U139 (N_139,N_47,In_489);
nand U140 (N_140,In_207,In_529);
or U141 (N_141,In_443,In_38);
xnor U142 (N_142,In_445,In_697);
nor U143 (N_143,In_218,In_227);
nand U144 (N_144,In_365,In_118);
or U145 (N_145,In_175,In_172);
nor U146 (N_146,In_72,In_426);
or U147 (N_147,In_316,N_82);
or U148 (N_148,In_625,In_283);
xor U149 (N_149,In_342,In_43);
nor U150 (N_150,In_562,In_66);
or U151 (N_151,N_86,In_348);
nand U152 (N_152,In_372,In_96);
xnor U153 (N_153,In_471,N_50);
xnor U154 (N_154,In_679,In_278);
or U155 (N_155,In_62,In_387);
or U156 (N_156,In_453,N_64);
or U157 (N_157,In_677,In_53);
nor U158 (N_158,N_81,In_303);
and U159 (N_159,In_490,In_441);
nand U160 (N_160,In_685,In_18);
nand U161 (N_161,In_231,In_299);
xor U162 (N_162,In_57,In_530);
or U163 (N_163,In_728,In_209);
nor U164 (N_164,In_320,In_217);
and U165 (N_165,In_568,In_420);
xor U166 (N_166,In_356,In_389);
xor U167 (N_167,In_47,In_65);
xor U168 (N_168,In_748,N_53);
xor U169 (N_169,N_7,In_289);
and U170 (N_170,In_630,In_494);
and U171 (N_171,In_556,In_134);
or U172 (N_172,In_626,In_747);
and U173 (N_173,In_178,In_92);
or U174 (N_174,In_179,In_482);
nor U175 (N_175,In_517,In_1);
xnor U176 (N_176,In_17,In_549);
nor U177 (N_177,In_59,In_419);
or U178 (N_178,In_326,In_480);
nand U179 (N_179,In_0,N_56);
xor U180 (N_180,In_402,In_519);
xnor U181 (N_181,In_280,In_16);
or U182 (N_182,In_146,N_98);
nor U183 (N_183,In_683,In_603);
nor U184 (N_184,N_21,In_48);
and U185 (N_185,N_49,In_123);
xor U186 (N_186,N_8,In_540);
nand U187 (N_187,In_132,In_680);
and U188 (N_188,In_150,In_506);
or U189 (N_189,In_42,N_91);
or U190 (N_190,In_240,In_297);
xor U191 (N_191,In_330,In_145);
or U192 (N_192,In_12,In_607);
and U193 (N_193,In_352,In_194);
xnor U194 (N_194,In_552,In_587);
nand U195 (N_195,In_327,In_541);
xor U196 (N_196,In_264,In_558);
xnor U197 (N_197,In_485,In_9);
nor U198 (N_198,In_287,In_381);
xnor U199 (N_199,In_706,In_315);
xnor U200 (N_200,N_30,In_538);
or U201 (N_201,In_496,N_51);
and U202 (N_202,In_388,In_164);
xor U203 (N_203,In_120,In_277);
xor U204 (N_204,N_143,N_77);
and U205 (N_205,N_185,In_405);
nand U206 (N_206,In_539,N_0);
or U207 (N_207,In_350,In_745);
and U208 (N_208,N_182,In_334);
or U209 (N_209,In_44,In_296);
and U210 (N_210,In_666,In_570);
nor U211 (N_211,In_396,N_160);
xnor U212 (N_212,N_16,In_620);
or U213 (N_213,In_158,N_93);
nand U214 (N_214,In_259,N_152);
nor U215 (N_215,In_646,In_317);
xor U216 (N_216,In_440,In_149);
nor U217 (N_217,In_602,In_191);
or U218 (N_218,N_73,In_32);
nor U219 (N_219,In_708,N_183);
nand U220 (N_220,In_667,In_19);
nor U221 (N_221,N_63,N_37);
xnor U222 (N_222,In_691,In_647);
or U223 (N_223,In_742,In_521);
nor U224 (N_224,In_305,N_48);
and U225 (N_225,In_64,In_124);
nand U226 (N_226,In_324,N_155);
xnor U227 (N_227,In_222,N_193);
xor U228 (N_228,In_255,N_38);
and U229 (N_229,N_71,In_592);
xor U230 (N_230,In_359,In_615);
xor U231 (N_231,In_740,In_467);
xor U232 (N_232,In_739,In_447);
nand U233 (N_233,N_80,In_183);
xor U234 (N_234,N_156,In_437);
xnor U235 (N_235,N_138,In_236);
xor U236 (N_236,In_257,In_584);
and U237 (N_237,In_503,In_122);
and U238 (N_238,In_288,In_628);
or U239 (N_239,N_11,N_169);
nand U240 (N_240,In_746,In_557);
xor U241 (N_241,In_254,In_221);
and U242 (N_242,In_127,In_138);
xor U243 (N_243,In_418,N_120);
nand U244 (N_244,In_114,In_22);
nand U245 (N_245,N_174,N_104);
or U246 (N_246,N_85,In_504);
and U247 (N_247,In_661,N_149);
xor U248 (N_248,N_162,N_58);
nand U249 (N_249,N_107,In_477);
and U250 (N_250,In_721,In_382);
or U251 (N_251,In_71,In_211);
nand U252 (N_252,In_486,In_113);
nor U253 (N_253,In_69,In_260);
or U254 (N_254,In_325,In_571);
or U255 (N_255,N_110,In_714);
nor U256 (N_256,In_583,N_137);
nand U257 (N_257,In_624,In_590);
or U258 (N_258,In_110,N_118);
or U259 (N_259,In_241,In_688);
nor U260 (N_260,In_406,In_368);
nand U261 (N_261,N_45,In_427);
xor U262 (N_262,N_168,N_95);
and U263 (N_263,In_336,In_528);
nand U264 (N_264,N_173,In_357);
or U265 (N_265,In_743,In_698);
and U266 (N_266,N_194,In_651);
or U267 (N_267,In_117,In_614);
xnor U268 (N_268,In_386,In_163);
xnor U269 (N_269,In_14,N_5);
nand U270 (N_270,N_34,In_36);
or U271 (N_271,In_610,In_563);
xnor U272 (N_272,In_413,In_302);
nand U273 (N_273,In_8,N_175);
nand U274 (N_274,In_653,In_424);
nand U275 (N_275,In_364,N_197);
xor U276 (N_276,N_167,In_723);
xnor U277 (N_277,In_616,In_246);
or U278 (N_278,N_170,In_88);
nand U279 (N_279,In_155,In_157);
nor U280 (N_280,In_715,In_532);
xor U281 (N_281,In_367,N_59);
xor U282 (N_282,N_78,In_726);
nor U283 (N_283,In_245,In_25);
or U284 (N_284,N_106,In_430);
or U285 (N_285,In_682,N_140);
nand U286 (N_286,In_546,N_159);
nand U287 (N_287,N_139,In_295);
and U288 (N_288,N_131,N_75);
nand U289 (N_289,In_100,N_70);
xor U290 (N_290,In_144,N_109);
xor U291 (N_291,In_162,In_67);
or U292 (N_292,In_293,In_193);
or U293 (N_293,In_331,In_579);
and U294 (N_294,N_66,N_115);
or U295 (N_295,In_198,In_170);
or U296 (N_296,N_192,In_354);
or U297 (N_297,N_166,N_26);
nand U298 (N_298,In_404,In_735);
or U299 (N_299,In_74,In_547);
nand U300 (N_300,In_703,N_102);
or U301 (N_301,N_178,In_294);
or U302 (N_302,In_407,In_370);
xnor U303 (N_303,N_299,N_288);
xnor U304 (N_304,N_17,In_449);
and U305 (N_305,In_509,In_102);
xor U306 (N_306,In_234,N_205);
and U307 (N_307,In_143,In_637);
nor U308 (N_308,In_322,In_643);
or U309 (N_309,N_289,In_466);
or U310 (N_310,In_37,N_28);
or U311 (N_311,N_132,In_136);
nand U312 (N_312,In_663,N_292);
xnor U313 (N_313,N_271,N_43);
nand U314 (N_314,In_674,N_150);
nor U315 (N_315,In_712,N_281);
and U316 (N_316,N_191,In_498);
xnor U317 (N_317,In_483,In_220);
nand U318 (N_318,In_732,N_261);
xor U319 (N_319,N_39,N_124);
nand U320 (N_320,N_268,N_231);
nor U321 (N_321,In_524,N_285);
xnor U322 (N_322,In_263,N_293);
or U323 (N_323,N_97,N_245);
and U324 (N_324,N_144,In_99);
nor U325 (N_325,N_133,N_136);
nand U326 (N_326,In_516,In_133);
xnor U327 (N_327,In_13,In_508);
and U328 (N_328,In_314,N_36);
xnor U329 (N_329,N_198,N_273);
and U330 (N_330,In_374,In_270);
nor U331 (N_331,N_135,N_188);
and U332 (N_332,In_233,In_262);
xnor U333 (N_333,N_207,In_380);
or U334 (N_334,In_373,In_491);
nor U335 (N_335,In_298,N_225);
and U336 (N_336,In_705,N_123);
nor U337 (N_337,In_594,In_613);
xnor U338 (N_338,In_169,In_210);
nor U339 (N_339,In_527,N_187);
xor U340 (N_340,In_238,In_50);
and U341 (N_341,N_158,N_221);
nand U342 (N_342,In_510,In_393);
and U343 (N_343,N_265,N_112);
and U344 (N_344,In_730,N_54);
or U345 (N_345,N_254,In_279);
and U346 (N_346,In_687,N_249);
and U347 (N_347,In_174,In_403);
xor U348 (N_348,In_699,N_296);
xor U349 (N_349,N_237,In_657);
xnor U350 (N_350,N_266,In_425);
nor U351 (N_351,In_89,N_20);
nand U352 (N_352,In_690,N_105);
xor U353 (N_353,N_190,N_228);
nand U354 (N_354,N_206,N_125);
or U355 (N_355,In_68,N_79);
or U356 (N_356,In_40,In_554);
and U357 (N_357,N_244,In_329);
nand U358 (N_358,N_210,In_656);
and U359 (N_359,In_154,N_240);
xnor U360 (N_360,N_236,N_269);
and U361 (N_361,N_157,N_108);
xnor U362 (N_362,In_311,N_72);
or U363 (N_363,N_264,In_537);
nand U364 (N_364,N_246,In_61);
nor U365 (N_365,N_215,N_61);
xor U366 (N_366,In_717,N_278);
nor U367 (N_367,N_57,In_543);
or U368 (N_368,N_248,In_611);
and U369 (N_369,N_280,N_119);
and U370 (N_370,In_487,In_131);
and U371 (N_371,In_204,In_339);
or U372 (N_372,N_35,N_253);
nand U373 (N_373,N_274,N_89);
xnor U374 (N_374,N_176,In_605);
xor U375 (N_375,N_226,In_460);
or U376 (N_376,N_241,In_87);
or U377 (N_377,In_681,N_272);
nand U378 (N_378,In_45,In_676);
or U379 (N_379,In_347,In_455);
or U380 (N_380,In_593,N_277);
xor U381 (N_381,In_686,In_514);
nand U382 (N_382,N_113,N_76);
nor U383 (N_383,In_456,N_100);
xnor U384 (N_384,N_154,In_91);
and U385 (N_385,In_658,N_227);
xnor U386 (N_386,In_213,N_147);
and U387 (N_387,In_292,In_249);
or U388 (N_388,In_580,In_121);
nand U389 (N_389,N_220,In_160);
and U390 (N_390,In_534,In_182);
or U391 (N_391,In_310,N_263);
or U392 (N_392,N_229,In_192);
and U393 (N_393,In_383,In_655);
or U394 (N_394,In_300,In_203);
nor U395 (N_395,N_242,In_214);
and U396 (N_396,N_212,In_75);
nand U397 (N_397,In_500,N_291);
nand U398 (N_398,In_459,In_190);
and U399 (N_399,N_101,N_282);
or U400 (N_400,N_103,N_243);
or U401 (N_401,In_662,N_161);
nand U402 (N_402,In_116,N_294);
and U403 (N_403,N_366,N_252);
nand U404 (N_404,N_216,N_351);
nand U405 (N_405,In_565,N_337);
nand U406 (N_406,In_429,N_365);
nand U407 (N_407,In_77,In_436);
xnor U408 (N_408,N_303,N_329);
nand U409 (N_409,In_319,N_307);
nand U410 (N_410,In_652,In_101);
and U411 (N_411,N_374,N_22);
and U412 (N_412,In_328,N_18);
and U413 (N_413,In_111,N_84);
xor U414 (N_414,N_311,In_139);
xor U415 (N_415,N_340,N_325);
nand U416 (N_416,In_199,N_301);
nor U417 (N_417,In_533,N_94);
or U418 (N_418,N_341,N_364);
and U419 (N_419,N_370,N_347);
nor U420 (N_420,In_696,N_355);
or U421 (N_421,In_438,N_358);
nand U422 (N_422,In_525,N_65);
xnor U423 (N_423,N_394,N_369);
or U424 (N_424,N_232,N_270);
nor U425 (N_425,N_40,N_284);
nor U426 (N_426,N_313,In_159);
or U427 (N_427,N_163,N_260);
or U428 (N_428,N_362,In_369);
xnor U429 (N_429,In_638,N_129);
nor U430 (N_430,In_56,N_19);
and U431 (N_431,In_98,N_195);
xor U432 (N_432,In_250,In_242);
nand U433 (N_433,N_333,In_200);
xor U434 (N_434,In_609,In_722);
or U435 (N_435,N_4,In_206);
nand U436 (N_436,N_111,N_153);
xor U437 (N_437,In_572,In_7);
and U438 (N_438,N_381,N_262);
and U439 (N_439,In_252,N_310);
or U440 (N_440,N_46,N_372);
nand U441 (N_441,In_550,N_367);
nor U442 (N_442,N_257,N_377);
xnor U443 (N_443,In_371,N_13);
or U444 (N_444,In_535,N_234);
or U445 (N_445,In_312,N_300);
xnor U446 (N_446,N_315,In_542);
nand U447 (N_447,N_83,In_492);
or U448 (N_448,In_511,In_478);
xnor U449 (N_449,In_417,N_378);
nor U450 (N_450,N_208,In_135);
and U451 (N_451,In_167,In_166);
xnor U452 (N_452,N_302,In_379);
and U453 (N_453,N_368,N_304);
nand U454 (N_454,N_177,In_196);
xnor U455 (N_455,In_669,N_224);
nor U456 (N_456,In_126,In_415);
and U457 (N_457,In_564,In_189);
nor U458 (N_458,In_103,N_165);
xnor U459 (N_459,N_322,N_360);
nand U460 (N_460,In_648,N_114);
xor U461 (N_461,In_385,In_507);
or U462 (N_462,In_475,N_346);
nor U463 (N_463,In_338,N_297);
and U464 (N_464,N_312,In_495);
or U465 (N_465,N_92,N_335);
or U466 (N_466,N_222,In_197);
and U467 (N_467,N_117,N_376);
xor U468 (N_468,N_230,N_343);
nand U469 (N_469,N_202,N_395);
nor U470 (N_470,In_412,N_141);
nand U471 (N_471,N_99,N_218);
nand U472 (N_472,N_27,N_87);
or U473 (N_473,N_116,In_275);
nor U474 (N_474,N_90,N_24);
nor U475 (N_475,N_88,N_353);
xor U476 (N_476,N_276,In_678);
or U477 (N_477,N_238,N_9);
or U478 (N_478,In_168,In_361);
nor U479 (N_479,In_650,N_134);
and U480 (N_480,In_284,N_342);
nand U481 (N_481,N_375,In_309);
nor U482 (N_482,In_454,N_275);
or U483 (N_483,In_636,N_214);
xor U484 (N_484,In_11,N_199);
xnor U485 (N_485,In_187,N_171);
xnor U486 (N_486,N_345,N_391);
or U487 (N_487,N_217,N_60);
or U488 (N_488,N_356,N_203);
or U489 (N_489,In_247,N_349);
xor U490 (N_490,N_363,In_129);
nor U491 (N_491,N_15,N_339);
and U492 (N_492,N_145,In_481);
nor U493 (N_493,In_345,In_24);
nor U494 (N_494,N_373,N_327);
or U495 (N_495,N_219,N_6);
and U496 (N_496,N_1,N_328);
nor U497 (N_497,N_14,In_142);
and U498 (N_498,In_80,N_279);
and U499 (N_499,N_298,In_641);
nand U500 (N_500,N_352,N_464);
xor U501 (N_501,N_477,N_196);
or U502 (N_502,N_148,In_675);
xnor U503 (N_503,N_429,N_400);
nand U504 (N_504,N_209,N_305);
xor U505 (N_505,N_320,In_243);
and U506 (N_506,N_223,N_250);
nor U507 (N_507,N_444,N_485);
xnor U508 (N_508,In_321,In_736);
or U509 (N_509,N_399,N_130);
nand U510 (N_510,In_665,N_424);
nor U511 (N_511,N_412,N_330);
xor U512 (N_512,N_392,N_433);
nand U513 (N_513,N_487,N_380);
xor U514 (N_514,N_468,N_350);
nor U515 (N_515,In_90,N_318);
and U516 (N_516,N_459,N_344);
xor U517 (N_517,N_383,In_629);
nor U518 (N_518,N_122,N_482);
nor U519 (N_519,In_202,N_450);
nor U520 (N_520,N_290,N_31);
nand U521 (N_521,In_446,N_172);
or U522 (N_522,N_452,N_473);
xor U523 (N_523,N_357,In_700);
nand U524 (N_524,N_239,N_68);
xnor U525 (N_525,N_251,N_494);
nor U526 (N_526,N_470,In_29);
nand U527 (N_527,N_427,N_428);
nand U528 (N_528,In_744,N_179);
nor U529 (N_529,N_306,N_471);
nor U530 (N_530,N_393,In_58);
nand U531 (N_531,N_443,In_462);
xor U532 (N_532,N_186,N_425);
nor U533 (N_533,N_461,N_434);
nand U534 (N_534,N_44,N_235);
or U535 (N_535,In_442,N_321);
or U536 (N_536,N_414,In_576);
nor U537 (N_537,In_574,In_105);
or U538 (N_538,In_719,N_490);
nand U539 (N_539,N_426,N_354);
nor U540 (N_540,In_73,In_450);
xnor U541 (N_541,N_326,N_404);
nand U542 (N_542,N_483,N_436);
and U543 (N_543,N_415,N_432);
nor U544 (N_544,N_258,N_406);
xnor U545 (N_545,In_512,N_201);
and U546 (N_546,N_338,N_480);
and U547 (N_547,In_394,N_204);
nor U548 (N_548,In_106,N_498);
xor U549 (N_549,N_440,N_180);
nand U550 (N_550,N_420,N_397);
and U551 (N_551,N_466,N_474);
or U552 (N_552,N_421,In_741);
nor U553 (N_553,N_361,N_255);
and U554 (N_554,N_371,N_359);
nor U555 (N_555,N_462,N_385);
nor U556 (N_556,In_395,N_126);
xor U557 (N_557,N_491,N_435);
xnor U558 (N_558,N_295,N_486);
xor U559 (N_559,N_151,N_437);
nor U560 (N_560,N_316,N_441);
or U561 (N_561,N_396,N_402);
nor U562 (N_562,N_331,N_431);
nand U563 (N_563,N_419,N_488);
xor U564 (N_564,N_472,N_489);
xnor U565 (N_565,N_442,N_475);
nor U566 (N_566,In_444,N_454);
or U567 (N_567,N_416,In_230);
xnor U568 (N_568,N_411,N_121);
nand U569 (N_569,In_366,N_409);
and U570 (N_570,N_332,N_42);
xnor U571 (N_571,In_551,N_267);
or U572 (N_572,N_446,N_460);
nand U573 (N_573,N_319,N_164);
and U574 (N_574,In_408,In_632);
xor U575 (N_575,N_492,N_413);
and U576 (N_576,N_499,In_597);
nand U577 (N_577,N_181,N_32);
nor U578 (N_578,N_481,N_324);
or U579 (N_579,N_96,N_407);
and U580 (N_580,In_439,N_334);
nand U581 (N_581,In_6,In_410);
xnor U582 (N_582,N_465,N_62);
or U583 (N_583,N_247,N_495);
nor U584 (N_584,N_213,In_634);
or U585 (N_585,In_378,N_388);
and U586 (N_586,N_410,N_463);
nor U587 (N_587,N_314,N_348);
nor U588 (N_588,In_3,N_467);
or U589 (N_589,N_478,N_317);
or U590 (N_590,N_387,N_458);
or U591 (N_591,N_389,N_497);
xnor U592 (N_592,N_453,N_142);
nand U593 (N_593,N_233,N_476);
nor U594 (N_594,In_599,N_417);
or U595 (N_595,N_423,N_479);
and U596 (N_596,N_455,In_737);
xnor U597 (N_597,N_493,N_403);
nor U598 (N_598,N_256,N_496);
or U599 (N_599,N_200,N_323);
nand U600 (N_600,N_573,N_519);
nor U601 (N_601,N_524,N_551);
and U602 (N_602,N_559,N_599);
or U603 (N_603,N_558,N_510);
xor U604 (N_604,N_513,N_530);
nor U605 (N_605,N_596,N_501);
or U606 (N_606,N_500,N_544);
or U607 (N_607,N_469,N_422);
nor U608 (N_608,N_146,N_523);
or U609 (N_609,N_517,N_336);
or U610 (N_610,N_520,N_507);
nand U611 (N_611,In_575,N_591);
nand U612 (N_612,In_421,N_566);
or U613 (N_613,N_555,N_259);
and U614 (N_614,N_590,N_438);
or U615 (N_615,In_308,N_580);
nand U616 (N_616,N_592,N_386);
and U617 (N_617,N_521,N_308);
or U618 (N_618,N_451,N_408);
nand U619 (N_619,In_451,N_570);
xor U620 (N_620,N_540,N_529);
nor U621 (N_621,N_595,N_502);
nand U622 (N_622,N_430,N_563);
xor U623 (N_623,N_588,N_553);
xor U624 (N_624,N_594,N_542);
and U625 (N_625,N_379,In_119);
and U626 (N_626,N_550,N_543);
or U627 (N_627,N_578,N_565);
nor U628 (N_628,N_538,N_516);
and U629 (N_629,N_184,N_448);
nor U630 (N_630,N_398,In_484);
nor U631 (N_631,N_598,N_574);
and U632 (N_632,In_531,N_526);
nor U633 (N_633,N_569,In_479);
and U634 (N_634,N_552,N_548);
and U635 (N_635,N_575,N_589);
xor U636 (N_636,N_560,N_128);
nand U637 (N_637,N_528,N_418);
nand U638 (N_638,N_518,N_283);
xnor U639 (N_639,N_506,N_579);
xnor U640 (N_640,N_583,N_522);
and U641 (N_641,N_525,N_449);
and U642 (N_642,N_445,N_401);
xor U643 (N_643,N_504,N_557);
or U644 (N_644,N_584,In_151);
nor U645 (N_645,N_549,N_508);
nand U646 (N_646,N_554,N_382);
nand U647 (N_647,N_515,N_534);
nand U648 (N_648,N_384,N_484);
or U649 (N_649,N_577,N_287);
nand U650 (N_650,N_582,N_457);
or U651 (N_651,N_539,N_390);
or U652 (N_652,N_531,N_571);
nor U653 (N_653,N_536,N_572);
xnor U654 (N_654,N_503,N_439);
nor U655 (N_655,N_509,N_535);
and U656 (N_656,In_689,N_541);
nor U657 (N_657,N_556,N_532);
nand U658 (N_658,N_585,N_567);
nor U659 (N_659,N_447,N_546);
xnor U660 (N_660,N_405,N_576);
xnor U661 (N_661,N_505,N_514);
and U662 (N_662,N_511,N_547);
xnor U663 (N_663,In_660,N_456);
xor U664 (N_664,N_581,N_587);
nand U665 (N_665,In_49,N_533);
nor U666 (N_666,N_593,N_286);
and U667 (N_667,N_564,N_309);
or U668 (N_668,N_23,In_600);
and U669 (N_669,N_127,N_597);
nand U670 (N_670,N_537,N_189);
nor U671 (N_671,N_586,N_561);
nor U672 (N_672,N_211,N_512);
or U673 (N_673,N_568,N_562);
and U674 (N_674,N_527,N_545);
xor U675 (N_675,N_528,N_545);
or U676 (N_676,N_577,N_398);
and U677 (N_677,N_127,N_540);
and U678 (N_678,N_534,N_544);
xor U679 (N_679,N_504,N_398);
and U680 (N_680,N_510,N_514);
and U681 (N_681,In_484,N_545);
or U682 (N_682,N_379,N_513);
and U683 (N_683,N_526,In_660);
and U684 (N_684,N_555,N_405);
xnor U685 (N_685,N_558,N_514);
or U686 (N_686,N_561,N_581);
xnor U687 (N_687,N_578,N_405);
xnor U688 (N_688,In_119,N_554);
nand U689 (N_689,N_510,N_515);
xnor U690 (N_690,N_566,N_558);
or U691 (N_691,N_538,N_577);
xnor U692 (N_692,N_582,N_596);
nor U693 (N_693,N_570,N_564);
nand U694 (N_694,N_531,N_576);
nand U695 (N_695,N_584,N_535);
nor U696 (N_696,N_556,N_570);
nand U697 (N_697,N_568,N_286);
and U698 (N_698,N_590,N_541);
nor U699 (N_699,N_588,N_544);
nor U700 (N_700,N_662,N_697);
nor U701 (N_701,N_619,N_666);
or U702 (N_702,N_674,N_601);
or U703 (N_703,N_681,N_667);
or U704 (N_704,N_695,N_675);
and U705 (N_705,N_627,N_685);
xnor U706 (N_706,N_636,N_610);
xor U707 (N_707,N_677,N_658);
and U708 (N_708,N_648,N_679);
nor U709 (N_709,N_631,N_646);
nand U710 (N_710,N_657,N_614);
nand U711 (N_711,N_686,N_664);
or U712 (N_712,N_692,N_617);
or U713 (N_713,N_641,N_615);
or U714 (N_714,N_604,N_687);
and U715 (N_715,N_654,N_690);
xor U716 (N_716,N_651,N_645);
xnor U717 (N_717,N_694,N_699);
nand U718 (N_718,N_649,N_612);
nor U719 (N_719,N_611,N_688);
nor U720 (N_720,N_609,N_671);
and U721 (N_721,N_602,N_606);
and U722 (N_722,N_616,N_625);
xor U723 (N_723,N_644,N_633);
nor U724 (N_724,N_659,N_632);
and U725 (N_725,N_656,N_621);
nor U726 (N_726,N_676,N_672);
and U727 (N_727,N_682,N_652);
xnor U728 (N_728,N_643,N_607);
nor U729 (N_729,N_655,N_670);
or U730 (N_730,N_663,N_661);
or U731 (N_731,N_623,N_634);
xnor U732 (N_732,N_629,N_650);
nor U733 (N_733,N_638,N_603);
nor U734 (N_734,N_628,N_680);
nor U735 (N_735,N_693,N_626);
xor U736 (N_736,N_691,N_600);
nand U737 (N_737,N_653,N_639);
nor U738 (N_738,N_668,N_678);
nand U739 (N_739,N_635,N_665);
or U740 (N_740,N_630,N_660);
or U741 (N_741,N_689,N_618);
nand U742 (N_742,N_620,N_683);
xnor U743 (N_743,N_696,N_622);
and U744 (N_744,N_669,N_640);
xor U745 (N_745,N_624,N_605);
nand U746 (N_746,N_608,N_673);
and U747 (N_747,N_698,N_613);
nand U748 (N_748,N_684,N_642);
nor U749 (N_749,N_637,N_647);
nand U750 (N_750,N_662,N_626);
and U751 (N_751,N_679,N_651);
nor U752 (N_752,N_616,N_682);
nand U753 (N_753,N_691,N_646);
nand U754 (N_754,N_664,N_670);
nand U755 (N_755,N_628,N_674);
and U756 (N_756,N_633,N_637);
and U757 (N_757,N_655,N_667);
nand U758 (N_758,N_615,N_669);
xor U759 (N_759,N_602,N_696);
and U760 (N_760,N_646,N_656);
nor U761 (N_761,N_628,N_613);
or U762 (N_762,N_651,N_634);
nor U763 (N_763,N_663,N_628);
and U764 (N_764,N_643,N_649);
and U765 (N_765,N_671,N_603);
nand U766 (N_766,N_642,N_647);
nor U767 (N_767,N_692,N_635);
nand U768 (N_768,N_612,N_650);
xor U769 (N_769,N_621,N_683);
and U770 (N_770,N_627,N_610);
nand U771 (N_771,N_681,N_661);
nor U772 (N_772,N_664,N_684);
nand U773 (N_773,N_610,N_687);
or U774 (N_774,N_630,N_622);
or U775 (N_775,N_620,N_670);
xnor U776 (N_776,N_614,N_688);
nand U777 (N_777,N_698,N_661);
nor U778 (N_778,N_688,N_668);
and U779 (N_779,N_605,N_691);
and U780 (N_780,N_679,N_690);
xnor U781 (N_781,N_668,N_616);
nand U782 (N_782,N_600,N_630);
and U783 (N_783,N_661,N_603);
nor U784 (N_784,N_655,N_613);
xor U785 (N_785,N_693,N_620);
nor U786 (N_786,N_687,N_638);
or U787 (N_787,N_697,N_623);
or U788 (N_788,N_656,N_678);
nor U789 (N_789,N_616,N_624);
nand U790 (N_790,N_612,N_656);
and U791 (N_791,N_692,N_624);
nor U792 (N_792,N_663,N_677);
nor U793 (N_793,N_684,N_635);
nor U794 (N_794,N_609,N_605);
and U795 (N_795,N_679,N_650);
or U796 (N_796,N_629,N_631);
or U797 (N_797,N_689,N_681);
or U798 (N_798,N_602,N_685);
nand U799 (N_799,N_617,N_669);
nor U800 (N_800,N_788,N_729);
xor U801 (N_801,N_784,N_707);
and U802 (N_802,N_737,N_705);
nand U803 (N_803,N_766,N_711);
and U804 (N_804,N_786,N_767);
and U805 (N_805,N_762,N_779);
or U806 (N_806,N_768,N_718);
and U807 (N_807,N_743,N_772);
or U808 (N_808,N_719,N_787);
or U809 (N_809,N_763,N_709);
nand U810 (N_810,N_791,N_769);
nand U811 (N_811,N_778,N_795);
nand U812 (N_812,N_783,N_712);
nor U813 (N_813,N_716,N_715);
xnor U814 (N_814,N_714,N_710);
xnor U815 (N_815,N_706,N_757);
xor U816 (N_816,N_750,N_722);
and U817 (N_817,N_792,N_745);
and U818 (N_818,N_731,N_702);
and U819 (N_819,N_739,N_798);
xor U820 (N_820,N_785,N_744);
nand U821 (N_821,N_751,N_794);
and U822 (N_822,N_720,N_701);
and U823 (N_823,N_759,N_700);
xor U824 (N_824,N_746,N_755);
xor U825 (N_825,N_777,N_749);
nor U826 (N_826,N_734,N_758);
xnor U827 (N_827,N_782,N_727);
nor U828 (N_828,N_799,N_754);
nor U829 (N_829,N_741,N_781);
nand U830 (N_830,N_704,N_797);
or U831 (N_831,N_728,N_753);
or U832 (N_832,N_733,N_713);
nor U833 (N_833,N_738,N_723);
and U834 (N_834,N_790,N_776);
or U835 (N_835,N_735,N_748);
or U836 (N_836,N_771,N_730);
and U837 (N_837,N_793,N_747);
and U838 (N_838,N_789,N_761);
nand U839 (N_839,N_764,N_732);
nand U840 (N_840,N_740,N_708);
nand U841 (N_841,N_780,N_770);
or U842 (N_842,N_736,N_726);
xnor U843 (N_843,N_752,N_742);
or U844 (N_844,N_756,N_765);
or U845 (N_845,N_703,N_717);
and U846 (N_846,N_724,N_773);
nor U847 (N_847,N_796,N_774);
nand U848 (N_848,N_725,N_721);
and U849 (N_849,N_775,N_760);
or U850 (N_850,N_735,N_739);
nor U851 (N_851,N_712,N_770);
xor U852 (N_852,N_776,N_711);
or U853 (N_853,N_763,N_701);
or U854 (N_854,N_747,N_774);
nor U855 (N_855,N_767,N_761);
xor U856 (N_856,N_776,N_734);
nor U857 (N_857,N_735,N_737);
and U858 (N_858,N_799,N_743);
nand U859 (N_859,N_752,N_739);
and U860 (N_860,N_784,N_775);
or U861 (N_861,N_716,N_783);
or U862 (N_862,N_709,N_706);
nand U863 (N_863,N_734,N_783);
and U864 (N_864,N_766,N_786);
or U865 (N_865,N_746,N_784);
and U866 (N_866,N_719,N_783);
or U867 (N_867,N_700,N_736);
xnor U868 (N_868,N_722,N_727);
xnor U869 (N_869,N_728,N_707);
and U870 (N_870,N_760,N_793);
xnor U871 (N_871,N_720,N_748);
and U872 (N_872,N_713,N_787);
or U873 (N_873,N_715,N_772);
and U874 (N_874,N_722,N_790);
or U875 (N_875,N_760,N_717);
or U876 (N_876,N_736,N_735);
or U877 (N_877,N_736,N_704);
and U878 (N_878,N_761,N_716);
nand U879 (N_879,N_756,N_730);
nor U880 (N_880,N_706,N_786);
nand U881 (N_881,N_718,N_712);
or U882 (N_882,N_761,N_776);
and U883 (N_883,N_779,N_789);
nor U884 (N_884,N_709,N_741);
or U885 (N_885,N_724,N_753);
nor U886 (N_886,N_729,N_778);
xor U887 (N_887,N_701,N_722);
and U888 (N_888,N_799,N_723);
nor U889 (N_889,N_723,N_715);
nor U890 (N_890,N_752,N_753);
nand U891 (N_891,N_727,N_787);
xnor U892 (N_892,N_705,N_769);
nand U893 (N_893,N_790,N_785);
or U894 (N_894,N_779,N_784);
or U895 (N_895,N_739,N_724);
nor U896 (N_896,N_780,N_742);
or U897 (N_897,N_700,N_737);
or U898 (N_898,N_740,N_757);
and U899 (N_899,N_793,N_770);
nand U900 (N_900,N_868,N_880);
nand U901 (N_901,N_863,N_856);
nor U902 (N_902,N_876,N_815);
xor U903 (N_903,N_823,N_811);
and U904 (N_904,N_829,N_869);
nand U905 (N_905,N_899,N_883);
nor U906 (N_906,N_886,N_820);
and U907 (N_907,N_841,N_865);
or U908 (N_908,N_813,N_877);
nor U909 (N_909,N_844,N_803);
nand U910 (N_910,N_804,N_832);
nor U911 (N_911,N_852,N_871);
and U912 (N_912,N_818,N_882);
xnor U913 (N_913,N_870,N_896);
and U914 (N_914,N_836,N_894);
xor U915 (N_915,N_866,N_833);
and U916 (N_916,N_861,N_858);
and U917 (N_917,N_830,N_897);
nor U918 (N_918,N_890,N_879);
or U919 (N_919,N_859,N_801);
or U920 (N_920,N_831,N_898);
or U921 (N_921,N_862,N_812);
nor U922 (N_922,N_878,N_885);
xor U923 (N_923,N_827,N_806);
nor U924 (N_924,N_849,N_808);
nor U925 (N_925,N_846,N_809);
xnor U926 (N_926,N_891,N_875);
and U927 (N_927,N_893,N_855);
nor U928 (N_928,N_842,N_881);
or U929 (N_929,N_860,N_810);
xor U930 (N_930,N_843,N_888);
nor U931 (N_931,N_828,N_864);
nand U932 (N_932,N_807,N_802);
nor U933 (N_933,N_826,N_837);
and U934 (N_934,N_851,N_848);
and U935 (N_935,N_853,N_805);
nor U936 (N_936,N_819,N_892);
xnor U937 (N_937,N_835,N_884);
nor U938 (N_938,N_867,N_887);
xor U939 (N_939,N_838,N_834);
nor U940 (N_940,N_845,N_800);
or U941 (N_941,N_814,N_857);
nand U942 (N_942,N_872,N_824);
xor U943 (N_943,N_821,N_847);
and U944 (N_944,N_840,N_822);
nand U945 (N_945,N_850,N_825);
or U946 (N_946,N_873,N_874);
nand U947 (N_947,N_889,N_895);
nor U948 (N_948,N_817,N_816);
nand U949 (N_949,N_839,N_854);
xor U950 (N_950,N_843,N_817);
nand U951 (N_951,N_839,N_879);
nand U952 (N_952,N_838,N_809);
nor U953 (N_953,N_838,N_824);
xnor U954 (N_954,N_883,N_821);
nor U955 (N_955,N_806,N_860);
xor U956 (N_956,N_805,N_839);
and U957 (N_957,N_806,N_844);
and U958 (N_958,N_856,N_841);
nor U959 (N_959,N_863,N_821);
xnor U960 (N_960,N_815,N_875);
and U961 (N_961,N_846,N_832);
or U962 (N_962,N_866,N_882);
and U963 (N_963,N_848,N_856);
xnor U964 (N_964,N_836,N_855);
or U965 (N_965,N_878,N_893);
or U966 (N_966,N_848,N_859);
and U967 (N_967,N_847,N_872);
and U968 (N_968,N_802,N_837);
and U969 (N_969,N_837,N_868);
and U970 (N_970,N_804,N_877);
nor U971 (N_971,N_887,N_837);
xor U972 (N_972,N_888,N_853);
and U973 (N_973,N_886,N_811);
nand U974 (N_974,N_868,N_873);
and U975 (N_975,N_816,N_855);
xnor U976 (N_976,N_860,N_887);
xnor U977 (N_977,N_859,N_816);
nand U978 (N_978,N_879,N_896);
and U979 (N_979,N_837,N_811);
nor U980 (N_980,N_870,N_885);
nor U981 (N_981,N_836,N_873);
xor U982 (N_982,N_804,N_887);
or U983 (N_983,N_816,N_891);
and U984 (N_984,N_899,N_884);
and U985 (N_985,N_880,N_801);
xor U986 (N_986,N_868,N_851);
nand U987 (N_987,N_892,N_855);
xor U988 (N_988,N_835,N_848);
and U989 (N_989,N_899,N_806);
and U990 (N_990,N_857,N_877);
nor U991 (N_991,N_859,N_851);
nand U992 (N_992,N_885,N_884);
and U993 (N_993,N_856,N_844);
or U994 (N_994,N_895,N_809);
and U995 (N_995,N_810,N_881);
nor U996 (N_996,N_868,N_898);
and U997 (N_997,N_886,N_814);
or U998 (N_998,N_830,N_829);
and U999 (N_999,N_804,N_879);
and U1000 (N_1000,N_957,N_950);
and U1001 (N_1001,N_900,N_975);
nand U1002 (N_1002,N_960,N_968);
and U1003 (N_1003,N_971,N_910);
xor U1004 (N_1004,N_941,N_951);
xnor U1005 (N_1005,N_988,N_936);
or U1006 (N_1006,N_917,N_912);
or U1007 (N_1007,N_987,N_955);
xnor U1008 (N_1008,N_923,N_914);
or U1009 (N_1009,N_908,N_978);
nand U1010 (N_1010,N_925,N_964);
nand U1011 (N_1011,N_932,N_940);
or U1012 (N_1012,N_903,N_970);
nor U1013 (N_1013,N_956,N_926);
or U1014 (N_1014,N_973,N_924);
or U1015 (N_1015,N_992,N_974);
or U1016 (N_1016,N_958,N_909);
and U1017 (N_1017,N_930,N_927);
nand U1018 (N_1018,N_999,N_942);
or U1019 (N_1019,N_922,N_986);
nand U1020 (N_1020,N_943,N_939);
xnor U1021 (N_1021,N_946,N_994);
and U1022 (N_1022,N_996,N_916);
and U1023 (N_1023,N_915,N_920);
xnor U1024 (N_1024,N_913,N_949);
or U1025 (N_1025,N_931,N_921);
xor U1026 (N_1026,N_982,N_907);
xor U1027 (N_1027,N_995,N_981);
or U1028 (N_1028,N_904,N_911);
nand U1029 (N_1029,N_977,N_954);
and U1030 (N_1030,N_947,N_985);
xnor U1031 (N_1031,N_962,N_929);
and U1032 (N_1032,N_905,N_961);
nand U1033 (N_1033,N_934,N_967);
and U1034 (N_1034,N_984,N_980);
and U1035 (N_1035,N_933,N_966);
xor U1036 (N_1036,N_902,N_919);
nand U1037 (N_1037,N_976,N_965);
or U1038 (N_1038,N_969,N_918);
and U1039 (N_1039,N_998,N_948);
or U1040 (N_1040,N_963,N_953);
xnor U1041 (N_1041,N_991,N_945);
nor U1042 (N_1042,N_997,N_901);
xnor U1043 (N_1043,N_959,N_938);
or U1044 (N_1044,N_906,N_937);
or U1045 (N_1045,N_952,N_983);
and U1046 (N_1046,N_928,N_989);
or U1047 (N_1047,N_944,N_979);
nand U1048 (N_1048,N_935,N_990);
nor U1049 (N_1049,N_993,N_972);
xor U1050 (N_1050,N_901,N_975);
or U1051 (N_1051,N_976,N_921);
nor U1052 (N_1052,N_919,N_969);
nor U1053 (N_1053,N_970,N_957);
or U1054 (N_1054,N_954,N_942);
nand U1055 (N_1055,N_920,N_980);
and U1056 (N_1056,N_959,N_914);
nand U1057 (N_1057,N_946,N_958);
xnor U1058 (N_1058,N_940,N_928);
or U1059 (N_1059,N_987,N_945);
and U1060 (N_1060,N_937,N_985);
nor U1061 (N_1061,N_971,N_958);
xnor U1062 (N_1062,N_953,N_946);
or U1063 (N_1063,N_961,N_959);
and U1064 (N_1064,N_918,N_945);
nand U1065 (N_1065,N_953,N_973);
xor U1066 (N_1066,N_951,N_947);
xnor U1067 (N_1067,N_912,N_934);
nor U1068 (N_1068,N_965,N_986);
and U1069 (N_1069,N_994,N_963);
and U1070 (N_1070,N_978,N_946);
nor U1071 (N_1071,N_906,N_956);
or U1072 (N_1072,N_931,N_974);
xor U1073 (N_1073,N_918,N_908);
nor U1074 (N_1074,N_974,N_917);
nor U1075 (N_1075,N_992,N_986);
or U1076 (N_1076,N_900,N_949);
xnor U1077 (N_1077,N_945,N_917);
and U1078 (N_1078,N_900,N_905);
nand U1079 (N_1079,N_981,N_978);
nand U1080 (N_1080,N_920,N_945);
and U1081 (N_1081,N_949,N_933);
xor U1082 (N_1082,N_941,N_938);
nand U1083 (N_1083,N_932,N_972);
and U1084 (N_1084,N_913,N_937);
and U1085 (N_1085,N_971,N_989);
or U1086 (N_1086,N_988,N_920);
nor U1087 (N_1087,N_965,N_991);
nand U1088 (N_1088,N_965,N_921);
or U1089 (N_1089,N_970,N_930);
or U1090 (N_1090,N_910,N_983);
nor U1091 (N_1091,N_986,N_960);
nor U1092 (N_1092,N_977,N_932);
xor U1093 (N_1093,N_980,N_911);
or U1094 (N_1094,N_936,N_999);
nand U1095 (N_1095,N_999,N_958);
xnor U1096 (N_1096,N_982,N_929);
nand U1097 (N_1097,N_995,N_947);
nand U1098 (N_1098,N_946,N_961);
or U1099 (N_1099,N_902,N_956);
or U1100 (N_1100,N_1000,N_1093);
or U1101 (N_1101,N_1018,N_1050);
or U1102 (N_1102,N_1080,N_1077);
xnor U1103 (N_1103,N_1078,N_1043);
nor U1104 (N_1104,N_1066,N_1003);
nor U1105 (N_1105,N_1019,N_1024);
xnor U1106 (N_1106,N_1021,N_1008);
nand U1107 (N_1107,N_1068,N_1035);
xor U1108 (N_1108,N_1056,N_1065);
and U1109 (N_1109,N_1099,N_1087);
or U1110 (N_1110,N_1013,N_1067);
xnor U1111 (N_1111,N_1096,N_1063);
xor U1112 (N_1112,N_1086,N_1098);
or U1113 (N_1113,N_1082,N_1057);
or U1114 (N_1114,N_1059,N_1025);
nor U1115 (N_1115,N_1010,N_1036);
nor U1116 (N_1116,N_1088,N_1034);
nand U1117 (N_1117,N_1031,N_1092);
or U1118 (N_1118,N_1070,N_1004);
and U1119 (N_1119,N_1069,N_1083);
nand U1120 (N_1120,N_1015,N_1047);
xnor U1121 (N_1121,N_1045,N_1064);
nand U1122 (N_1122,N_1055,N_1030);
and U1123 (N_1123,N_1085,N_1052);
and U1124 (N_1124,N_1075,N_1072);
nand U1125 (N_1125,N_1079,N_1091);
nor U1126 (N_1126,N_1033,N_1090);
or U1127 (N_1127,N_1007,N_1095);
nand U1128 (N_1128,N_1014,N_1023);
and U1129 (N_1129,N_1060,N_1022);
nor U1130 (N_1130,N_1006,N_1001);
and U1131 (N_1131,N_1073,N_1038);
or U1132 (N_1132,N_1053,N_1011);
xor U1133 (N_1133,N_1012,N_1042);
nor U1134 (N_1134,N_1029,N_1048);
and U1135 (N_1135,N_1032,N_1009);
nand U1136 (N_1136,N_1039,N_1020);
xor U1137 (N_1137,N_1040,N_1076);
nor U1138 (N_1138,N_1074,N_1002);
and U1139 (N_1139,N_1071,N_1028);
nand U1140 (N_1140,N_1097,N_1044);
or U1141 (N_1141,N_1046,N_1054);
xnor U1142 (N_1142,N_1005,N_1041);
nor U1143 (N_1143,N_1027,N_1084);
and U1144 (N_1144,N_1058,N_1051);
nor U1145 (N_1145,N_1037,N_1089);
and U1146 (N_1146,N_1094,N_1062);
and U1147 (N_1147,N_1061,N_1081);
and U1148 (N_1148,N_1049,N_1016);
or U1149 (N_1149,N_1026,N_1017);
xor U1150 (N_1150,N_1057,N_1036);
xnor U1151 (N_1151,N_1001,N_1053);
xor U1152 (N_1152,N_1013,N_1005);
or U1153 (N_1153,N_1009,N_1001);
xnor U1154 (N_1154,N_1007,N_1005);
nand U1155 (N_1155,N_1044,N_1085);
and U1156 (N_1156,N_1012,N_1082);
nor U1157 (N_1157,N_1012,N_1004);
nand U1158 (N_1158,N_1063,N_1020);
nor U1159 (N_1159,N_1046,N_1068);
xor U1160 (N_1160,N_1090,N_1048);
nor U1161 (N_1161,N_1027,N_1077);
nand U1162 (N_1162,N_1054,N_1043);
and U1163 (N_1163,N_1016,N_1025);
and U1164 (N_1164,N_1009,N_1031);
nor U1165 (N_1165,N_1039,N_1030);
nor U1166 (N_1166,N_1088,N_1029);
or U1167 (N_1167,N_1035,N_1027);
nand U1168 (N_1168,N_1080,N_1002);
nand U1169 (N_1169,N_1083,N_1061);
nor U1170 (N_1170,N_1061,N_1088);
nand U1171 (N_1171,N_1089,N_1006);
or U1172 (N_1172,N_1080,N_1075);
nand U1173 (N_1173,N_1076,N_1084);
nand U1174 (N_1174,N_1045,N_1032);
or U1175 (N_1175,N_1097,N_1026);
or U1176 (N_1176,N_1050,N_1068);
xnor U1177 (N_1177,N_1072,N_1021);
or U1178 (N_1178,N_1063,N_1003);
or U1179 (N_1179,N_1012,N_1057);
xor U1180 (N_1180,N_1095,N_1008);
or U1181 (N_1181,N_1094,N_1002);
nor U1182 (N_1182,N_1054,N_1061);
nor U1183 (N_1183,N_1002,N_1057);
xor U1184 (N_1184,N_1092,N_1022);
xnor U1185 (N_1185,N_1075,N_1013);
nand U1186 (N_1186,N_1063,N_1091);
xor U1187 (N_1187,N_1098,N_1030);
or U1188 (N_1188,N_1057,N_1080);
xnor U1189 (N_1189,N_1020,N_1003);
and U1190 (N_1190,N_1022,N_1098);
and U1191 (N_1191,N_1033,N_1086);
or U1192 (N_1192,N_1091,N_1087);
and U1193 (N_1193,N_1070,N_1080);
xor U1194 (N_1194,N_1039,N_1084);
or U1195 (N_1195,N_1087,N_1009);
or U1196 (N_1196,N_1072,N_1044);
or U1197 (N_1197,N_1049,N_1067);
and U1198 (N_1198,N_1015,N_1095);
and U1199 (N_1199,N_1033,N_1060);
or U1200 (N_1200,N_1191,N_1124);
and U1201 (N_1201,N_1127,N_1139);
and U1202 (N_1202,N_1197,N_1153);
and U1203 (N_1203,N_1141,N_1163);
xor U1204 (N_1204,N_1115,N_1159);
or U1205 (N_1205,N_1107,N_1129);
nand U1206 (N_1206,N_1177,N_1170);
and U1207 (N_1207,N_1189,N_1101);
and U1208 (N_1208,N_1116,N_1181);
or U1209 (N_1209,N_1118,N_1111);
nand U1210 (N_1210,N_1112,N_1121);
or U1211 (N_1211,N_1157,N_1152);
and U1212 (N_1212,N_1109,N_1167);
nand U1213 (N_1213,N_1193,N_1176);
xor U1214 (N_1214,N_1156,N_1195);
xnor U1215 (N_1215,N_1155,N_1135);
or U1216 (N_1216,N_1150,N_1113);
or U1217 (N_1217,N_1145,N_1126);
nor U1218 (N_1218,N_1132,N_1138);
nor U1219 (N_1219,N_1168,N_1100);
nor U1220 (N_1220,N_1144,N_1137);
and U1221 (N_1221,N_1174,N_1134);
or U1222 (N_1222,N_1154,N_1180);
xor U1223 (N_1223,N_1192,N_1199);
and U1224 (N_1224,N_1196,N_1165);
and U1225 (N_1225,N_1158,N_1166);
xor U1226 (N_1226,N_1125,N_1160);
xor U1227 (N_1227,N_1147,N_1120);
and U1228 (N_1228,N_1103,N_1187);
nand U1229 (N_1229,N_1148,N_1198);
nand U1230 (N_1230,N_1114,N_1133);
or U1231 (N_1231,N_1105,N_1104);
and U1232 (N_1232,N_1179,N_1117);
or U1233 (N_1233,N_1178,N_1183);
xnor U1234 (N_1234,N_1142,N_1164);
nand U1235 (N_1235,N_1173,N_1184);
or U1236 (N_1236,N_1169,N_1190);
xor U1237 (N_1237,N_1131,N_1130);
nand U1238 (N_1238,N_1119,N_1106);
nor U1239 (N_1239,N_1143,N_1161);
xor U1240 (N_1240,N_1162,N_1186);
nand U1241 (N_1241,N_1110,N_1182);
and U1242 (N_1242,N_1194,N_1185);
nand U1243 (N_1243,N_1140,N_1188);
xnor U1244 (N_1244,N_1172,N_1149);
xnor U1245 (N_1245,N_1128,N_1122);
and U1246 (N_1246,N_1102,N_1123);
or U1247 (N_1247,N_1136,N_1108);
or U1248 (N_1248,N_1151,N_1175);
xor U1249 (N_1249,N_1146,N_1171);
nor U1250 (N_1250,N_1174,N_1154);
and U1251 (N_1251,N_1189,N_1176);
nand U1252 (N_1252,N_1146,N_1144);
or U1253 (N_1253,N_1113,N_1191);
and U1254 (N_1254,N_1189,N_1159);
nand U1255 (N_1255,N_1171,N_1139);
xnor U1256 (N_1256,N_1168,N_1142);
nor U1257 (N_1257,N_1189,N_1196);
xnor U1258 (N_1258,N_1162,N_1165);
xnor U1259 (N_1259,N_1179,N_1143);
nor U1260 (N_1260,N_1109,N_1173);
xnor U1261 (N_1261,N_1154,N_1184);
nor U1262 (N_1262,N_1195,N_1107);
and U1263 (N_1263,N_1186,N_1196);
nor U1264 (N_1264,N_1182,N_1150);
and U1265 (N_1265,N_1160,N_1105);
nor U1266 (N_1266,N_1194,N_1158);
or U1267 (N_1267,N_1157,N_1131);
nor U1268 (N_1268,N_1173,N_1170);
xor U1269 (N_1269,N_1197,N_1176);
and U1270 (N_1270,N_1171,N_1138);
nand U1271 (N_1271,N_1162,N_1172);
or U1272 (N_1272,N_1118,N_1105);
or U1273 (N_1273,N_1151,N_1136);
nand U1274 (N_1274,N_1178,N_1145);
nor U1275 (N_1275,N_1112,N_1152);
xnor U1276 (N_1276,N_1108,N_1156);
xnor U1277 (N_1277,N_1113,N_1185);
xnor U1278 (N_1278,N_1162,N_1189);
nand U1279 (N_1279,N_1191,N_1132);
and U1280 (N_1280,N_1157,N_1100);
xnor U1281 (N_1281,N_1127,N_1186);
nand U1282 (N_1282,N_1198,N_1145);
xor U1283 (N_1283,N_1157,N_1166);
xor U1284 (N_1284,N_1149,N_1126);
xor U1285 (N_1285,N_1168,N_1153);
nor U1286 (N_1286,N_1194,N_1136);
nor U1287 (N_1287,N_1178,N_1168);
xor U1288 (N_1288,N_1184,N_1141);
xor U1289 (N_1289,N_1150,N_1195);
nor U1290 (N_1290,N_1102,N_1162);
nor U1291 (N_1291,N_1113,N_1183);
nand U1292 (N_1292,N_1130,N_1106);
nor U1293 (N_1293,N_1148,N_1180);
or U1294 (N_1294,N_1128,N_1180);
nor U1295 (N_1295,N_1147,N_1197);
or U1296 (N_1296,N_1139,N_1193);
nand U1297 (N_1297,N_1100,N_1156);
nor U1298 (N_1298,N_1132,N_1185);
or U1299 (N_1299,N_1101,N_1130);
xnor U1300 (N_1300,N_1223,N_1291);
or U1301 (N_1301,N_1274,N_1234);
and U1302 (N_1302,N_1278,N_1253);
or U1303 (N_1303,N_1293,N_1258);
nor U1304 (N_1304,N_1213,N_1222);
nand U1305 (N_1305,N_1245,N_1231);
nand U1306 (N_1306,N_1212,N_1268);
nor U1307 (N_1307,N_1255,N_1276);
and U1308 (N_1308,N_1282,N_1228);
nand U1309 (N_1309,N_1266,N_1264);
or U1310 (N_1310,N_1239,N_1273);
nand U1311 (N_1311,N_1247,N_1299);
or U1312 (N_1312,N_1243,N_1220);
nand U1313 (N_1313,N_1275,N_1205);
and U1314 (N_1314,N_1246,N_1229);
nand U1315 (N_1315,N_1203,N_1209);
nand U1316 (N_1316,N_1269,N_1221);
or U1317 (N_1317,N_1207,N_1232);
or U1318 (N_1318,N_1200,N_1280);
xnor U1319 (N_1319,N_1206,N_1236);
nand U1320 (N_1320,N_1286,N_1249);
nand U1321 (N_1321,N_1272,N_1225);
nand U1322 (N_1322,N_1281,N_1267);
and U1323 (N_1323,N_1208,N_1287);
nand U1324 (N_1324,N_1204,N_1298);
xor U1325 (N_1325,N_1260,N_1297);
nor U1326 (N_1326,N_1241,N_1202);
xor U1327 (N_1327,N_1215,N_1288);
nor U1328 (N_1328,N_1262,N_1252);
and U1329 (N_1329,N_1271,N_1235);
or U1330 (N_1330,N_1261,N_1289);
or U1331 (N_1331,N_1211,N_1295);
xnor U1332 (N_1332,N_1226,N_1214);
and U1333 (N_1333,N_1284,N_1224);
or U1334 (N_1334,N_1216,N_1217);
xnor U1335 (N_1335,N_1263,N_1277);
xnor U1336 (N_1336,N_1283,N_1201);
nor U1337 (N_1337,N_1237,N_1285);
or U1338 (N_1338,N_1251,N_1244);
or U1339 (N_1339,N_1257,N_1227);
xnor U1340 (N_1340,N_1238,N_1279);
nand U1341 (N_1341,N_1230,N_1250);
nor U1342 (N_1342,N_1256,N_1292);
xnor U1343 (N_1343,N_1240,N_1210);
nand U1344 (N_1344,N_1248,N_1296);
nand U1345 (N_1345,N_1242,N_1265);
nand U1346 (N_1346,N_1219,N_1259);
or U1347 (N_1347,N_1270,N_1294);
and U1348 (N_1348,N_1218,N_1233);
and U1349 (N_1349,N_1254,N_1290);
nand U1350 (N_1350,N_1291,N_1220);
and U1351 (N_1351,N_1275,N_1267);
nand U1352 (N_1352,N_1219,N_1264);
and U1353 (N_1353,N_1239,N_1256);
nor U1354 (N_1354,N_1213,N_1291);
xnor U1355 (N_1355,N_1281,N_1269);
xor U1356 (N_1356,N_1295,N_1245);
xnor U1357 (N_1357,N_1251,N_1282);
nor U1358 (N_1358,N_1257,N_1212);
and U1359 (N_1359,N_1259,N_1208);
or U1360 (N_1360,N_1260,N_1201);
or U1361 (N_1361,N_1203,N_1226);
nand U1362 (N_1362,N_1239,N_1277);
nor U1363 (N_1363,N_1240,N_1244);
and U1364 (N_1364,N_1247,N_1255);
nand U1365 (N_1365,N_1217,N_1227);
or U1366 (N_1366,N_1275,N_1278);
nand U1367 (N_1367,N_1218,N_1225);
nor U1368 (N_1368,N_1275,N_1219);
and U1369 (N_1369,N_1291,N_1261);
nand U1370 (N_1370,N_1288,N_1278);
and U1371 (N_1371,N_1296,N_1221);
xor U1372 (N_1372,N_1266,N_1291);
nor U1373 (N_1373,N_1278,N_1213);
nand U1374 (N_1374,N_1248,N_1267);
and U1375 (N_1375,N_1276,N_1200);
nor U1376 (N_1376,N_1249,N_1273);
and U1377 (N_1377,N_1274,N_1208);
nor U1378 (N_1378,N_1285,N_1296);
nor U1379 (N_1379,N_1258,N_1253);
and U1380 (N_1380,N_1259,N_1277);
nor U1381 (N_1381,N_1260,N_1209);
xor U1382 (N_1382,N_1282,N_1216);
xor U1383 (N_1383,N_1240,N_1277);
and U1384 (N_1384,N_1275,N_1207);
nand U1385 (N_1385,N_1278,N_1258);
xor U1386 (N_1386,N_1212,N_1271);
nand U1387 (N_1387,N_1205,N_1286);
or U1388 (N_1388,N_1280,N_1211);
nor U1389 (N_1389,N_1272,N_1248);
nor U1390 (N_1390,N_1201,N_1214);
or U1391 (N_1391,N_1265,N_1252);
or U1392 (N_1392,N_1258,N_1234);
and U1393 (N_1393,N_1220,N_1236);
nor U1394 (N_1394,N_1240,N_1253);
xnor U1395 (N_1395,N_1242,N_1260);
and U1396 (N_1396,N_1236,N_1259);
nor U1397 (N_1397,N_1255,N_1275);
nand U1398 (N_1398,N_1224,N_1295);
xor U1399 (N_1399,N_1234,N_1232);
nor U1400 (N_1400,N_1374,N_1343);
and U1401 (N_1401,N_1312,N_1383);
nand U1402 (N_1402,N_1340,N_1380);
xor U1403 (N_1403,N_1315,N_1332);
nor U1404 (N_1404,N_1386,N_1308);
xnor U1405 (N_1405,N_1327,N_1365);
and U1406 (N_1406,N_1321,N_1398);
or U1407 (N_1407,N_1302,N_1376);
nor U1408 (N_1408,N_1310,N_1364);
nand U1409 (N_1409,N_1344,N_1358);
xor U1410 (N_1410,N_1330,N_1309);
nand U1411 (N_1411,N_1377,N_1322);
or U1412 (N_1412,N_1381,N_1318);
nor U1413 (N_1413,N_1379,N_1351);
or U1414 (N_1414,N_1385,N_1326);
xnor U1415 (N_1415,N_1362,N_1363);
or U1416 (N_1416,N_1389,N_1366);
nand U1417 (N_1417,N_1367,N_1353);
or U1418 (N_1418,N_1320,N_1369);
or U1419 (N_1419,N_1390,N_1341);
nand U1420 (N_1420,N_1307,N_1333);
xor U1421 (N_1421,N_1347,N_1303);
nand U1422 (N_1422,N_1348,N_1304);
xnor U1423 (N_1423,N_1350,N_1388);
and U1424 (N_1424,N_1338,N_1395);
nor U1425 (N_1425,N_1317,N_1334);
or U1426 (N_1426,N_1301,N_1399);
or U1427 (N_1427,N_1393,N_1375);
and U1428 (N_1428,N_1361,N_1382);
and U1429 (N_1429,N_1342,N_1356);
or U1430 (N_1430,N_1359,N_1325);
or U1431 (N_1431,N_1370,N_1372);
xor U1432 (N_1432,N_1314,N_1345);
and U1433 (N_1433,N_1371,N_1336);
nand U1434 (N_1434,N_1337,N_1329);
or U1435 (N_1435,N_1397,N_1355);
xor U1436 (N_1436,N_1360,N_1300);
or U1437 (N_1437,N_1313,N_1378);
nand U1438 (N_1438,N_1305,N_1331);
nand U1439 (N_1439,N_1387,N_1396);
xor U1440 (N_1440,N_1357,N_1324);
or U1441 (N_1441,N_1311,N_1384);
nor U1442 (N_1442,N_1339,N_1346);
nor U1443 (N_1443,N_1319,N_1354);
nand U1444 (N_1444,N_1323,N_1349);
nor U1445 (N_1445,N_1335,N_1391);
xor U1446 (N_1446,N_1352,N_1394);
xor U1447 (N_1447,N_1328,N_1306);
nor U1448 (N_1448,N_1316,N_1373);
nor U1449 (N_1449,N_1368,N_1392);
nor U1450 (N_1450,N_1335,N_1313);
and U1451 (N_1451,N_1339,N_1387);
and U1452 (N_1452,N_1322,N_1343);
nand U1453 (N_1453,N_1336,N_1386);
and U1454 (N_1454,N_1398,N_1326);
nor U1455 (N_1455,N_1334,N_1302);
and U1456 (N_1456,N_1342,N_1351);
nand U1457 (N_1457,N_1372,N_1308);
xor U1458 (N_1458,N_1318,N_1328);
xnor U1459 (N_1459,N_1387,N_1315);
nor U1460 (N_1460,N_1303,N_1336);
xor U1461 (N_1461,N_1360,N_1333);
or U1462 (N_1462,N_1319,N_1371);
or U1463 (N_1463,N_1311,N_1345);
xnor U1464 (N_1464,N_1313,N_1337);
or U1465 (N_1465,N_1381,N_1315);
or U1466 (N_1466,N_1398,N_1342);
xor U1467 (N_1467,N_1349,N_1377);
nor U1468 (N_1468,N_1323,N_1362);
nand U1469 (N_1469,N_1357,N_1350);
nor U1470 (N_1470,N_1339,N_1328);
nor U1471 (N_1471,N_1391,N_1376);
nor U1472 (N_1472,N_1350,N_1361);
xnor U1473 (N_1473,N_1309,N_1380);
nor U1474 (N_1474,N_1314,N_1302);
xor U1475 (N_1475,N_1376,N_1371);
nand U1476 (N_1476,N_1354,N_1391);
or U1477 (N_1477,N_1321,N_1338);
xnor U1478 (N_1478,N_1394,N_1377);
nand U1479 (N_1479,N_1378,N_1396);
nand U1480 (N_1480,N_1356,N_1345);
xnor U1481 (N_1481,N_1359,N_1336);
or U1482 (N_1482,N_1315,N_1305);
xor U1483 (N_1483,N_1322,N_1335);
nor U1484 (N_1484,N_1353,N_1374);
or U1485 (N_1485,N_1308,N_1398);
nand U1486 (N_1486,N_1308,N_1309);
or U1487 (N_1487,N_1314,N_1370);
nor U1488 (N_1488,N_1334,N_1375);
nand U1489 (N_1489,N_1374,N_1317);
xnor U1490 (N_1490,N_1381,N_1365);
or U1491 (N_1491,N_1309,N_1315);
or U1492 (N_1492,N_1395,N_1362);
or U1493 (N_1493,N_1325,N_1323);
nand U1494 (N_1494,N_1386,N_1379);
or U1495 (N_1495,N_1310,N_1367);
xor U1496 (N_1496,N_1304,N_1305);
or U1497 (N_1497,N_1399,N_1371);
or U1498 (N_1498,N_1306,N_1355);
xnor U1499 (N_1499,N_1369,N_1395);
nor U1500 (N_1500,N_1499,N_1475);
or U1501 (N_1501,N_1413,N_1400);
xnor U1502 (N_1502,N_1422,N_1496);
xor U1503 (N_1503,N_1441,N_1402);
xnor U1504 (N_1504,N_1486,N_1464);
xnor U1505 (N_1505,N_1424,N_1494);
nor U1506 (N_1506,N_1453,N_1489);
xor U1507 (N_1507,N_1470,N_1412);
xnor U1508 (N_1508,N_1479,N_1420);
or U1509 (N_1509,N_1403,N_1417);
xnor U1510 (N_1510,N_1481,N_1446);
or U1511 (N_1511,N_1466,N_1469);
and U1512 (N_1512,N_1425,N_1460);
nand U1513 (N_1513,N_1411,N_1450);
nor U1514 (N_1514,N_1451,N_1493);
nor U1515 (N_1515,N_1431,N_1444);
and U1516 (N_1516,N_1435,N_1448);
nor U1517 (N_1517,N_1455,N_1476);
nor U1518 (N_1518,N_1438,N_1401);
and U1519 (N_1519,N_1443,N_1445);
nand U1520 (N_1520,N_1432,N_1409);
and U1521 (N_1521,N_1419,N_1447);
or U1522 (N_1522,N_1405,N_1463);
nand U1523 (N_1523,N_1492,N_1415);
or U1524 (N_1524,N_1461,N_1468);
and U1525 (N_1525,N_1423,N_1483);
xnor U1526 (N_1526,N_1428,N_1497);
nand U1527 (N_1527,N_1440,N_1457);
xnor U1528 (N_1528,N_1472,N_1485);
nand U1529 (N_1529,N_1452,N_1449);
nor U1530 (N_1530,N_1487,N_1430);
nand U1531 (N_1531,N_1416,N_1491);
xor U1532 (N_1532,N_1442,N_1459);
or U1533 (N_1533,N_1458,N_1488);
nor U1534 (N_1534,N_1477,N_1404);
and U1535 (N_1535,N_1426,N_1410);
and U1536 (N_1536,N_1406,N_1495);
xor U1537 (N_1537,N_1434,N_1427);
nand U1538 (N_1538,N_1471,N_1484);
nand U1539 (N_1539,N_1407,N_1421);
nor U1540 (N_1540,N_1436,N_1478);
or U1541 (N_1541,N_1498,N_1473);
nor U1542 (N_1542,N_1437,N_1433);
nand U1543 (N_1543,N_1418,N_1480);
nor U1544 (N_1544,N_1462,N_1414);
and U1545 (N_1545,N_1490,N_1439);
and U1546 (N_1546,N_1454,N_1482);
nor U1547 (N_1547,N_1429,N_1408);
nor U1548 (N_1548,N_1456,N_1474);
nor U1549 (N_1549,N_1465,N_1467);
or U1550 (N_1550,N_1454,N_1484);
or U1551 (N_1551,N_1461,N_1481);
nor U1552 (N_1552,N_1423,N_1430);
xnor U1553 (N_1553,N_1442,N_1416);
or U1554 (N_1554,N_1409,N_1418);
and U1555 (N_1555,N_1425,N_1426);
xor U1556 (N_1556,N_1481,N_1459);
or U1557 (N_1557,N_1448,N_1468);
or U1558 (N_1558,N_1403,N_1433);
or U1559 (N_1559,N_1433,N_1444);
xor U1560 (N_1560,N_1460,N_1480);
nor U1561 (N_1561,N_1428,N_1482);
and U1562 (N_1562,N_1421,N_1416);
nand U1563 (N_1563,N_1415,N_1487);
nand U1564 (N_1564,N_1490,N_1495);
xor U1565 (N_1565,N_1416,N_1497);
and U1566 (N_1566,N_1495,N_1415);
nor U1567 (N_1567,N_1419,N_1496);
nand U1568 (N_1568,N_1411,N_1400);
xnor U1569 (N_1569,N_1413,N_1447);
nor U1570 (N_1570,N_1477,N_1491);
xnor U1571 (N_1571,N_1442,N_1438);
and U1572 (N_1572,N_1488,N_1417);
xor U1573 (N_1573,N_1442,N_1425);
and U1574 (N_1574,N_1441,N_1420);
or U1575 (N_1575,N_1400,N_1488);
nand U1576 (N_1576,N_1454,N_1481);
xor U1577 (N_1577,N_1474,N_1438);
xnor U1578 (N_1578,N_1422,N_1444);
and U1579 (N_1579,N_1462,N_1404);
nor U1580 (N_1580,N_1402,N_1428);
nor U1581 (N_1581,N_1459,N_1453);
or U1582 (N_1582,N_1443,N_1485);
or U1583 (N_1583,N_1461,N_1455);
and U1584 (N_1584,N_1462,N_1486);
nand U1585 (N_1585,N_1491,N_1420);
and U1586 (N_1586,N_1499,N_1483);
or U1587 (N_1587,N_1472,N_1439);
and U1588 (N_1588,N_1459,N_1411);
xnor U1589 (N_1589,N_1475,N_1465);
nor U1590 (N_1590,N_1495,N_1418);
nand U1591 (N_1591,N_1443,N_1429);
and U1592 (N_1592,N_1481,N_1477);
or U1593 (N_1593,N_1434,N_1480);
or U1594 (N_1594,N_1421,N_1404);
and U1595 (N_1595,N_1472,N_1429);
or U1596 (N_1596,N_1449,N_1455);
nor U1597 (N_1597,N_1462,N_1469);
nor U1598 (N_1598,N_1452,N_1444);
xor U1599 (N_1599,N_1459,N_1418);
nor U1600 (N_1600,N_1548,N_1510);
and U1601 (N_1601,N_1566,N_1522);
or U1602 (N_1602,N_1539,N_1511);
nor U1603 (N_1603,N_1572,N_1533);
or U1604 (N_1604,N_1581,N_1593);
nand U1605 (N_1605,N_1559,N_1546);
nand U1606 (N_1606,N_1505,N_1565);
and U1607 (N_1607,N_1528,N_1506);
and U1608 (N_1608,N_1540,N_1590);
or U1609 (N_1609,N_1538,N_1534);
xnor U1610 (N_1610,N_1532,N_1587);
nand U1611 (N_1611,N_1518,N_1579);
xor U1612 (N_1612,N_1563,N_1586);
or U1613 (N_1613,N_1567,N_1545);
and U1614 (N_1614,N_1524,N_1585);
and U1615 (N_1615,N_1573,N_1584);
and U1616 (N_1616,N_1551,N_1508);
and U1617 (N_1617,N_1568,N_1509);
xor U1618 (N_1618,N_1594,N_1507);
nand U1619 (N_1619,N_1575,N_1578);
nand U1620 (N_1620,N_1597,N_1526);
nor U1621 (N_1621,N_1516,N_1500);
nor U1622 (N_1622,N_1504,N_1595);
xor U1623 (N_1623,N_1515,N_1582);
xor U1624 (N_1624,N_1547,N_1530);
or U1625 (N_1625,N_1574,N_1550);
and U1626 (N_1626,N_1544,N_1580);
nand U1627 (N_1627,N_1561,N_1521);
nor U1628 (N_1628,N_1549,N_1513);
nor U1629 (N_1629,N_1557,N_1553);
xnor U1630 (N_1630,N_1537,N_1589);
nor U1631 (N_1631,N_1583,N_1570);
xor U1632 (N_1632,N_1599,N_1552);
nor U1633 (N_1633,N_1517,N_1596);
xor U1634 (N_1634,N_1571,N_1525);
and U1635 (N_1635,N_1556,N_1554);
nor U1636 (N_1636,N_1558,N_1592);
and U1637 (N_1637,N_1512,N_1523);
or U1638 (N_1638,N_1501,N_1543);
nand U1639 (N_1639,N_1536,N_1555);
or U1640 (N_1640,N_1535,N_1564);
nor U1641 (N_1641,N_1541,N_1529);
nand U1642 (N_1642,N_1562,N_1514);
and U1643 (N_1643,N_1531,N_1569);
nand U1644 (N_1644,N_1503,N_1542);
and U1645 (N_1645,N_1502,N_1588);
xor U1646 (N_1646,N_1591,N_1598);
xnor U1647 (N_1647,N_1527,N_1520);
nor U1648 (N_1648,N_1560,N_1519);
nand U1649 (N_1649,N_1577,N_1576);
nor U1650 (N_1650,N_1594,N_1574);
xor U1651 (N_1651,N_1584,N_1568);
or U1652 (N_1652,N_1588,N_1505);
and U1653 (N_1653,N_1515,N_1545);
or U1654 (N_1654,N_1572,N_1503);
nor U1655 (N_1655,N_1567,N_1530);
and U1656 (N_1656,N_1506,N_1547);
and U1657 (N_1657,N_1544,N_1545);
xor U1658 (N_1658,N_1518,N_1566);
and U1659 (N_1659,N_1576,N_1552);
nor U1660 (N_1660,N_1576,N_1583);
and U1661 (N_1661,N_1508,N_1574);
and U1662 (N_1662,N_1527,N_1562);
nand U1663 (N_1663,N_1551,N_1583);
or U1664 (N_1664,N_1526,N_1518);
and U1665 (N_1665,N_1557,N_1578);
nand U1666 (N_1666,N_1567,N_1548);
or U1667 (N_1667,N_1568,N_1519);
xnor U1668 (N_1668,N_1588,N_1586);
xor U1669 (N_1669,N_1543,N_1506);
xnor U1670 (N_1670,N_1575,N_1545);
nor U1671 (N_1671,N_1575,N_1555);
and U1672 (N_1672,N_1531,N_1520);
or U1673 (N_1673,N_1537,N_1543);
nand U1674 (N_1674,N_1557,N_1562);
nand U1675 (N_1675,N_1566,N_1557);
nand U1676 (N_1676,N_1522,N_1528);
xnor U1677 (N_1677,N_1576,N_1572);
and U1678 (N_1678,N_1565,N_1562);
and U1679 (N_1679,N_1599,N_1579);
xnor U1680 (N_1680,N_1523,N_1571);
and U1681 (N_1681,N_1518,N_1568);
xor U1682 (N_1682,N_1583,N_1514);
or U1683 (N_1683,N_1568,N_1502);
or U1684 (N_1684,N_1564,N_1510);
nand U1685 (N_1685,N_1594,N_1566);
or U1686 (N_1686,N_1581,N_1583);
nor U1687 (N_1687,N_1517,N_1536);
nor U1688 (N_1688,N_1550,N_1510);
nand U1689 (N_1689,N_1511,N_1596);
xnor U1690 (N_1690,N_1555,N_1529);
and U1691 (N_1691,N_1557,N_1585);
xnor U1692 (N_1692,N_1593,N_1549);
nor U1693 (N_1693,N_1576,N_1579);
or U1694 (N_1694,N_1518,N_1511);
and U1695 (N_1695,N_1585,N_1523);
or U1696 (N_1696,N_1501,N_1509);
or U1697 (N_1697,N_1587,N_1514);
nor U1698 (N_1698,N_1540,N_1529);
nor U1699 (N_1699,N_1508,N_1558);
nor U1700 (N_1700,N_1627,N_1645);
nand U1701 (N_1701,N_1675,N_1606);
or U1702 (N_1702,N_1680,N_1671);
or U1703 (N_1703,N_1649,N_1623);
or U1704 (N_1704,N_1653,N_1676);
nor U1705 (N_1705,N_1691,N_1658);
nor U1706 (N_1706,N_1613,N_1622);
nor U1707 (N_1707,N_1641,N_1637);
nor U1708 (N_1708,N_1634,N_1624);
nand U1709 (N_1709,N_1607,N_1630);
nand U1710 (N_1710,N_1603,N_1657);
and U1711 (N_1711,N_1644,N_1611);
or U1712 (N_1712,N_1619,N_1602);
nor U1713 (N_1713,N_1609,N_1681);
or U1714 (N_1714,N_1628,N_1678);
xnor U1715 (N_1715,N_1632,N_1654);
nor U1716 (N_1716,N_1694,N_1686);
nor U1717 (N_1717,N_1672,N_1618);
xnor U1718 (N_1718,N_1659,N_1650);
or U1719 (N_1719,N_1677,N_1605);
xor U1720 (N_1720,N_1652,N_1636);
xnor U1721 (N_1721,N_1640,N_1696);
nor U1722 (N_1722,N_1638,N_1679);
and U1723 (N_1723,N_1662,N_1635);
or U1724 (N_1724,N_1682,N_1669);
nor U1725 (N_1725,N_1651,N_1688);
nand U1726 (N_1726,N_1621,N_1664);
or U1727 (N_1727,N_1626,N_1648);
nand U1728 (N_1728,N_1667,N_1692);
or U1729 (N_1729,N_1684,N_1625);
and U1730 (N_1730,N_1666,N_1604);
nor U1731 (N_1731,N_1698,N_1612);
xnor U1732 (N_1732,N_1693,N_1663);
nor U1733 (N_1733,N_1642,N_1668);
and U1734 (N_1734,N_1661,N_1674);
and U1735 (N_1735,N_1695,N_1673);
nand U1736 (N_1736,N_1646,N_1615);
and U1737 (N_1737,N_1633,N_1690);
xor U1738 (N_1738,N_1614,N_1670);
or U1739 (N_1739,N_1683,N_1665);
xnor U1740 (N_1740,N_1600,N_1656);
nor U1741 (N_1741,N_1617,N_1689);
nor U1742 (N_1742,N_1660,N_1616);
nor U1743 (N_1743,N_1647,N_1608);
nand U1744 (N_1744,N_1697,N_1601);
nand U1745 (N_1745,N_1610,N_1643);
xor U1746 (N_1746,N_1699,N_1685);
or U1747 (N_1747,N_1655,N_1629);
nand U1748 (N_1748,N_1687,N_1620);
nor U1749 (N_1749,N_1631,N_1639);
nor U1750 (N_1750,N_1696,N_1638);
and U1751 (N_1751,N_1679,N_1660);
xnor U1752 (N_1752,N_1689,N_1684);
or U1753 (N_1753,N_1652,N_1626);
xor U1754 (N_1754,N_1683,N_1694);
or U1755 (N_1755,N_1655,N_1660);
nor U1756 (N_1756,N_1611,N_1698);
and U1757 (N_1757,N_1697,N_1687);
nor U1758 (N_1758,N_1683,N_1676);
nor U1759 (N_1759,N_1653,N_1665);
nand U1760 (N_1760,N_1620,N_1615);
xnor U1761 (N_1761,N_1697,N_1608);
and U1762 (N_1762,N_1664,N_1612);
and U1763 (N_1763,N_1602,N_1640);
nand U1764 (N_1764,N_1692,N_1621);
and U1765 (N_1765,N_1668,N_1681);
or U1766 (N_1766,N_1621,N_1683);
xnor U1767 (N_1767,N_1688,N_1680);
nand U1768 (N_1768,N_1643,N_1676);
and U1769 (N_1769,N_1642,N_1614);
nor U1770 (N_1770,N_1635,N_1647);
nor U1771 (N_1771,N_1646,N_1608);
or U1772 (N_1772,N_1652,N_1696);
xor U1773 (N_1773,N_1612,N_1671);
xor U1774 (N_1774,N_1678,N_1636);
nand U1775 (N_1775,N_1663,N_1617);
nand U1776 (N_1776,N_1698,N_1663);
xor U1777 (N_1777,N_1661,N_1672);
or U1778 (N_1778,N_1652,N_1603);
nor U1779 (N_1779,N_1639,N_1626);
nand U1780 (N_1780,N_1667,N_1649);
xnor U1781 (N_1781,N_1613,N_1628);
and U1782 (N_1782,N_1635,N_1640);
or U1783 (N_1783,N_1647,N_1680);
xor U1784 (N_1784,N_1629,N_1671);
and U1785 (N_1785,N_1681,N_1683);
nor U1786 (N_1786,N_1691,N_1675);
or U1787 (N_1787,N_1686,N_1632);
and U1788 (N_1788,N_1600,N_1668);
nand U1789 (N_1789,N_1640,N_1657);
nor U1790 (N_1790,N_1616,N_1664);
and U1791 (N_1791,N_1612,N_1647);
nand U1792 (N_1792,N_1625,N_1683);
xnor U1793 (N_1793,N_1686,N_1678);
nor U1794 (N_1794,N_1674,N_1673);
nand U1795 (N_1795,N_1640,N_1665);
xor U1796 (N_1796,N_1699,N_1674);
xnor U1797 (N_1797,N_1684,N_1658);
or U1798 (N_1798,N_1648,N_1666);
nand U1799 (N_1799,N_1600,N_1678);
xnor U1800 (N_1800,N_1709,N_1796);
and U1801 (N_1801,N_1799,N_1728);
xnor U1802 (N_1802,N_1716,N_1730);
or U1803 (N_1803,N_1776,N_1762);
and U1804 (N_1804,N_1767,N_1778);
xnor U1805 (N_1805,N_1739,N_1727);
or U1806 (N_1806,N_1759,N_1764);
nor U1807 (N_1807,N_1777,N_1718);
xnor U1808 (N_1808,N_1789,N_1783);
nand U1809 (N_1809,N_1754,N_1701);
or U1810 (N_1810,N_1786,N_1790);
nand U1811 (N_1811,N_1711,N_1703);
xnor U1812 (N_1812,N_1717,N_1774);
nand U1813 (N_1813,N_1760,N_1704);
or U1814 (N_1814,N_1795,N_1723);
xor U1815 (N_1815,N_1794,N_1769);
nor U1816 (N_1816,N_1710,N_1782);
or U1817 (N_1817,N_1787,N_1744);
nand U1818 (N_1818,N_1745,N_1705);
and U1819 (N_1819,N_1756,N_1788);
xor U1820 (N_1820,N_1731,N_1752);
nand U1821 (N_1821,N_1766,N_1765);
and U1822 (N_1822,N_1798,N_1751);
nand U1823 (N_1823,N_1746,N_1749);
xnor U1824 (N_1824,N_1772,N_1753);
and U1825 (N_1825,N_1715,N_1714);
and U1826 (N_1826,N_1708,N_1758);
nand U1827 (N_1827,N_1742,N_1768);
xor U1828 (N_1828,N_1779,N_1713);
or U1829 (N_1829,N_1702,N_1738);
and U1830 (N_1830,N_1733,N_1712);
or U1831 (N_1831,N_1721,N_1793);
nand U1832 (N_1832,N_1792,N_1720);
or U1833 (N_1833,N_1791,N_1732);
xnor U1834 (N_1834,N_1763,N_1722);
nand U1835 (N_1835,N_1770,N_1748);
and U1836 (N_1836,N_1736,N_1757);
nor U1837 (N_1837,N_1737,N_1780);
and U1838 (N_1838,N_1734,N_1750);
nor U1839 (N_1839,N_1781,N_1700);
xor U1840 (N_1840,N_1729,N_1797);
nor U1841 (N_1841,N_1785,N_1725);
and U1842 (N_1842,N_1747,N_1740);
xnor U1843 (N_1843,N_1761,N_1741);
and U1844 (N_1844,N_1706,N_1775);
nand U1845 (N_1845,N_1719,N_1773);
and U1846 (N_1846,N_1735,N_1726);
nand U1847 (N_1847,N_1724,N_1743);
or U1848 (N_1848,N_1707,N_1771);
or U1849 (N_1849,N_1784,N_1755);
nand U1850 (N_1850,N_1717,N_1712);
nor U1851 (N_1851,N_1799,N_1790);
and U1852 (N_1852,N_1717,N_1728);
or U1853 (N_1853,N_1747,N_1767);
nor U1854 (N_1854,N_1797,N_1783);
xnor U1855 (N_1855,N_1733,N_1708);
nand U1856 (N_1856,N_1745,N_1784);
nand U1857 (N_1857,N_1725,N_1737);
nor U1858 (N_1858,N_1796,N_1741);
or U1859 (N_1859,N_1722,N_1730);
nand U1860 (N_1860,N_1770,N_1783);
and U1861 (N_1861,N_1741,N_1793);
or U1862 (N_1862,N_1723,N_1736);
or U1863 (N_1863,N_1722,N_1726);
nor U1864 (N_1864,N_1760,N_1750);
xor U1865 (N_1865,N_1786,N_1730);
nand U1866 (N_1866,N_1769,N_1746);
or U1867 (N_1867,N_1746,N_1725);
or U1868 (N_1868,N_1703,N_1775);
or U1869 (N_1869,N_1722,N_1759);
nand U1870 (N_1870,N_1742,N_1795);
and U1871 (N_1871,N_1796,N_1745);
and U1872 (N_1872,N_1730,N_1787);
or U1873 (N_1873,N_1718,N_1782);
xnor U1874 (N_1874,N_1724,N_1796);
nand U1875 (N_1875,N_1717,N_1740);
nor U1876 (N_1876,N_1774,N_1748);
nand U1877 (N_1877,N_1787,N_1738);
nor U1878 (N_1878,N_1710,N_1762);
and U1879 (N_1879,N_1768,N_1749);
or U1880 (N_1880,N_1791,N_1798);
nor U1881 (N_1881,N_1778,N_1782);
xor U1882 (N_1882,N_1708,N_1731);
or U1883 (N_1883,N_1704,N_1733);
nor U1884 (N_1884,N_1731,N_1782);
and U1885 (N_1885,N_1713,N_1764);
or U1886 (N_1886,N_1709,N_1718);
nor U1887 (N_1887,N_1767,N_1763);
nor U1888 (N_1888,N_1758,N_1722);
nand U1889 (N_1889,N_1724,N_1774);
xor U1890 (N_1890,N_1793,N_1711);
and U1891 (N_1891,N_1721,N_1715);
and U1892 (N_1892,N_1759,N_1713);
nor U1893 (N_1893,N_1795,N_1786);
or U1894 (N_1894,N_1726,N_1778);
nor U1895 (N_1895,N_1785,N_1738);
and U1896 (N_1896,N_1768,N_1738);
xor U1897 (N_1897,N_1738,N_1764);
nor U1898 (N_1898,N_1740,N_1784);
or U1899 (N_1899,N_1770,N_1766);
or U1900 (N_1900,N_1859,N_1894);
or U1901 (N_1901,N_1818,N_1893);
nor U1902 (N_1902,N_1887,N_1883);
xor U1903 (N_1903,N_1849,N_1898);
nand U1904 (N_1904,N_1868,N_1837);
xnor U1905 (N_1905,N_1848,N_1891);
xnor U1906 (N_1906,N_1852,N_1889);
or U1907 (N_1907,N_1884,N_1864);
xor U1908 (N_1908,N_1890,N_1882);
xnor U1909 (N_1909,N_1832,N_1812);
and U1910 (N_1910,N_1850,N_1878);
nor U1911 (N_1911,N_1829,N_1853);
and U1912 (N_1912,N_1819,N_1825);
and U1913 (N_1913,N_1841,N_1831);
nor U1914 (N_1914,N_1870,N_1875);
nor U1915 (N_1915,N_1845,N_1846);
xor U1916 (N_1916,N_1855,N_1851);
xor U1917 (N_1917,N_1897,N_1857);
or U1918 (N_1918,N_1821,N_1862);
xnor U1919 (N_1919,N_1858,N_1807);
nand U1920 (N_1920,N_1880,N_1802);
nor U1921 (N_1921,N_1861,N_1844);
or U1922 (N_1922,N_1895,N_1804);
nand U1923 (N_1923,N_1816,N_1881);
nor U1924 (N_1924,N_1847,N_1869);
nand U1925 (N_1925,N_1840,N_1834);
and U1926 (N_1926,N_1874,N_1836);
or U1927 (N_1927,N_1813,N_1800);
and U1928 (N_1928,N_1805,N_1801);
and U1929 (N_1929,N_1810,N_1839);
or U1930 (N_1930,N_1817,N_1888);
nand U1931 (N_1931,N_1899,N_1896);
and U1932 (N_1932,N_1823,N_1860);
and U1933 (N_1933,N_1885,N_1843);
xor U1934 (N_1934,N_1866,N_1872);
nand U1935 (N_1935,N_1809,N_1856);
nor U1936 (N_1936,N_1828,N_1876);
and U1937 (N_1937,N_1822,N_1871);
xnor U1938 (N_1938,N_1803,N_1833);
nand U1939 (N_1939,N_1892,N_1842);
or U1940 (N_1940,N_1811,N_1838);
and U1941 (N_1941,N_1808,N_1830);
nand U1942 (N_1942,N_1826,N_1854);
nand U1943 (N_1943,N_1815,N_1877);
nor U1944 (N_1944,N_1865,N_1863);
or U1945 (N_1945,N_1806,N_1820);
and U1946 (N_1946,N_1827,N_1867);
nor U1947 (N_1947,N_1879,N_1835);
or U1948 (N_1948,N_1814,N_1873);
or U1949 (N_1949,N_1824,N_1886);
and U1950 (N_1950,N_1848,N_1816);
or U1951 (N_1951,N_1832,N_1828);
or U1952 (N_1952,N_1897,N_1839);
nor U1953 (N_1953,N_1860,N_1896);
nor U1954 (N_1954,N_1853,N_1826);
nand U1955 (N_1955,N_1896,N_1833);
and U1956 (N_1956,N_1844,N_1837);
nand U1957 (N_1957,N_1890,N_1866);
nor U1958 (N_1958,N_1896,N_1827);
nand U1959 (N_1959,N_1811,N_1814);
nor U1960 (N_1960,N_1875,N_1866);
and U1961 (N_1961,N_1840,N_1896);
and U1962 (N_1962,N_1899,N_1863);
nand U1963 (N_1963,N_1845,N_1838);
nand U1964 (N_1964,N_1854,N_1808);
xnor U1965 (N_1965,N_1864,N_1818);
xor U1966 (N_1966,N_1805,N_1840);
nor U1967 (N_1967,N_1889,N_1894);
nand U1968 (N_1968,N_1801,N_1892);
nand U1969 (N_1969,N_1877,N_1873);
and U1970 (N_1970,N_1827,N_1882);
or U1971 (N_1971,N_1826,N_1887);
xnor U1972 (N_1972,N_1845,N_1837);
or U1973 (N_1973,N_1888,N_1877);
nor U1974 (N_1974,N_1834,N_1860);
or U1975 (N_1975,N_1850,N_1897);
or U1976 (N_1976,N_1859,N_1892);
nand U1977 (N_1977,N_1849,N_1809);
xnor U1978 (N_1978,N_1821,N_1877);
and U1979 (N_1979,N_1818,N_1861);
or U1980 (N_1980,N_1884,N_1885);
xor U1981 (N_1981,N_1878,N_1863);
or U1982 (N_1982,N_1811,N_1831);
and U1983 (N_1983,N_1852,N_1855);
xor U1984 (N_1984,N_1826,N_1866);
nand U1985 (N_1985,N_1830,N_1883);
or U1986 (N_1986,N_1876,N_1851);
or U1987 (N_1987,N_1898,N_1859);
or U1988 (N_1988,N_1830,N_1876);
xnor U1989 (N_1989,N_1854,N_1816);
nand U1990 (N_1990,N_1884,N_1813);
nand U1991 (N_1991,N_1869,N_1809);
nor U1992 (N_1992,N_1817,N_1839);
nand U1993 (N_1993,N_1806,N_1860);
or U1994 (N_1994,N_1891,N_1865);
nand U1995 (N_1995,N_1873,N_1826);
nor U1996 (N_1996,N_1817,N_1862);
or U1997 (N_1997,N_1801,N_1876);
and U1998 (N_1998,N_1833,N_1883);
or U1999 (N_1999,N_1873,N_1839);
xor U2000 (N_2000,N_1938,N_1949);
xnor U2001 (N_2001,N_1982,N_1941);
nor U2002 (N_2002,N_1911,N_1970);
xnor U2003 (N_2003,N_1904,N_1947);
nor U2004 (N_2004,N_1936,N_1914);
xor U2005 (N_2005,N_1932,N_1998);
and U2006 (N_2006,N_1925,N_1928);
nand U2007 (N_2007,N_1964,N_1996);
or U2008 (N_2008,N_1975,N_1930);
and U2009 (N_2009,N_1905,N_1994);
nor U2010 (N_2010,N_1983,N_1943);
nand U2011 (N_2011,N_1997,N_1992);
and U2012 (N_2012,N_1954,N_1957);
or U2013 (N_2013,N_1934,N_1903);
nand U2014 (N_2014,N_1965,N_1961);
nand U2015 (N_2015,N_1956,N_1946);
nand U2016 (N_2016,N_1929,N_1969);
nor U2017 (N_2017,N_1953,N_1967);
xnor U2018 (N_2018,N_1902,N_1910);
nor U2019 (N_2019,N_1966,N_1976);
or U2020 (N_2020,N_1962,N_1990);
or U2021 (N_2021,N_1974,N_1924);
or U2022 (N_2022,N_1906,N_1959);
xor U2023 (N_2023,N_1919,N_1991);
xnor U2024 (N_2024,N_1917,N_1944);
nor U2025 (N_2025,N_1955,N_1916);
nor U2026 (N_2026,N_1989,N_1951);
and U2027 (N_2027,N_1958,N_1981);
xor U2028 (N_2028,N_1926,N_1921);
nand U2029 (N_2029,N_1937,N_1979);
and U2030 (N_2030,N_1971,N_1909);
and U2031 (N_2031,N_1920,N_1933);
nor U2032 (N_2032,N_1985,N_1980);
xor U2033 (N_2033,N_1995,N_1923);
nor U2034 (N_2034,N_1935,N_1950);
and U2035 (N_2035,N_1927,N_1922);
and U2036 (N_2036,N_1908,N_1912);
xnor U2037 (N_2037,N_1977,N_1940);
and U2038 (N_2038,N_1915,N_1945);
nor U2039 (N_2039,N_1942,N_1952);
nor U2040 (N_2040,N_1999,N_1960);
and U2041 (N_2041,N_1973,N_1972);
nor U2042 (N_2042,N_1978,N_1993);
or U2043 (N_2043,N_1913,N_1968);
nand U2044 (N_2044,N_1907,N_1901);
nor U2045 (N_2045,N_1963,N_1988);
xor U2046 (N_2046,N_1948,N_1931);
and U2047 (N_2047,N_1918,N_1939);
nand U2048 (N_2048,N_1987,N_1984);
or U2049 (N_2049,N_1900,N_1986);
or U2050 (N_2050,N_1935,N_1901);
and U2051 (N_2051,N_1917,N_1973);
and U2052 (N_2052,N_1922,N_1910);
nor U2053 (N_2053,N_1900,N_1970);
or U2054 (N_2054,N_1910,N_1965);
xor U2055 (N_2055,N_1930,N_1992);
or U2056 (N_2056,N_1913,N_1946);
nor U2057 (N_2057,N_1948,N_1907);
xnor U2058 (N_2058,N_1942,N_1925);
xnor U2059 (N_2059,N_1942,N_1916);
or U2060 (N_2060,N_1937,N_1900);
xnor U2061 (N_2061,N_1999,N_1992);
or U2062 (N_2062,N_1938,N_1966);
or U2063 (N_2063,N_1905,N_1940);
or U2064 (N_2064,N_1938,N_1908);
or U2065 (N_2065,N_1902,N_1960);
nor U2066 (N_2066,N_1998,N_1906);
nand U2067 (N_2067,N_1969,N_1922);
or U2068 (N_2068,N_1909,N_1936);
nand U2069 (N_2069,N_1906,N_1938);
and U2070 (N_2070,N_1971,N_1948);
and U2071 (N_2071,N_1987,N_1933);
xnor U2072 (N_2072,N_1946,N_1938);
and U2073 (N_2073,N_1951,N_1980);
and U2074 (N_2074,N_1931,N_1986);
or U2075 (N_2075,N_1900,N_1932);
and U2076 (N_2076,N_1984,N_1916);
nor U2077 (N_2077,N_1913,N_1931);
or U2078 (N_2078,N_1956,N_1966);
and U2079 (N_2079,N_1992,N_1923);
or U2080 (N_2080,N_1901,N_1984);
nor U2081 (N_2081,N_1979,N_1964);
and U2082 (N_2082,N_1991,N_1913);
xor U2083 (N_2083,N_1982,N_1981);
nor U2084 (N_2084,N_1986,N_1946);
and U2085 (N_2085,N_1964,N_1955);
or U2086 (N_2086,N_1976,N_1939);
nand U2087 (N_2087,N_1938,N_1931);
and U2088 (N_2088,N_1917,N_1907);
xnor U2089 (N_2089,N_1940,N_1932);
nor U2090 (N_2090,N_1922,N_1937);
and U2091 (N_2091,N_1996,N_1966);
nand U2092 (N_2092,N_1908,N_1997);
xnor U2093 (N_2093,N_1941,N_1949);
nor U2094 (N_2094,N_1907,N_1979);
or U2095 (N_2095,N_1922,N_1960);
or U2096 (N_2096,N_1976,N_1978);
nor U2097 (N_2097,N_1933,N_1901);
xnor U2098 (N_2098,N_1935,N_1915);
and U2099 (N_2099,N_1936,N_1919);
or U2100 (N_2100,N_2032,N_2068);
nand U2101 (N_2101,N_2086,N_2079);
nand U2102 (N_2102,N_2061,N_2051);
nor U2103 (N_2103,N_2035,N_2097);
xor U2104 (N_2104,N_2058,N_2074);
nor U2105 (N_2105,N_2089,N_2018);
or U2106 (N_2106,N_2038,N_2084);
and U2107 (N_2107,N_2025,N_2012);
and U2108 (N_2108,N_2065,N_2013);
or U2109 (N_2109,N_2057,N_2010);
xnor U2110 (N_2110,N_2098,N_2029);
nand U2111 (N_2111,N_2030,N_2066);
or U2112 (N_2112,N_2088,N_2076);
nor U2113 (N_2113,N_2042,N_2083);
and U2114 (N_2114,N_2019,N_2027);
nand U2115 (N_2115,N_2022,N_2008);
or U2116 (N_2116,N_2092,N_2085);
or U2117 (N_2117,N_2007,N_2005);
xor U2118 (N_2118,N_2052,N_2003);
xnor U2119 (N_2119,N_2039,N_2072);
xnor U2120 (N_2120,N_2044,N_2073);
nor U2121 (N_2121,N_2071,N_2095);
nor U2122 (N_2122,N_2048,N_2040);
and U2123 (N_2123,N_2014,N_2099);
or U2124 (N_2124,N_2036,N_2002);
nor U2125 (N_2125,N_2028,N_2006);
nor U2126 (N_2126,N_2011,N_2041);
xnor U2127 (N_2127,N_2023,N_2015);
or U2128 (N_2128,N_2090,N_2047);
and U2129 (N_2129,N_2069,N_2016);
or U2130 (N_2130,N_2055,N_2063);
and U2131 (N_2131,N_2024,N_2062);
nand U2132 (N_2132,N_2054,N_2080);
and U2133 (N_2133,N_2056,N_2009);
nor U2134 (N_2134,N_2001,N_2096);
xor U2135 (N_2135,N_2037,N_2045);
xor U2136 (N_2136,N_2075,N_2026);
or U2137 (N_2137,N_2059,N_2091);
nor U2138 (N_2138,N_2082,N_2060);
or U2139 (N_2139,N_2087,N_2034);
and U2140 (N_2140,N_2050,N_2078);
or U2141 (N_2141,N_2020,N_2093);
and U2142 (N_2142,N_2049,N_2081);
and U2143 (N_2143,N_2053,N_2031);
nor U2144 (N_2144,N_2000,N_2046);
or U2145 (N_2145,N_2021,N_2094);
and U2146 (N_2146,N_2043,N_2077);
nand U2147 (N_2147,N_2064,N_2004);
nand U2148 (N_2148,N_2017,N_2033);
or U2149 (N_2149,N_2067,N_2070);
or U2150 (N_2150,N_2024,N_2066);
or U2151 (N_2151,N_2036,N_2099);
and U2152 (N_2152,N_2081,N_2068);
nand U2153 (N_2153,N_2003,N_2049);
nand U2154 (N_2154,N_2029,N_2095);
or U2155 (N_2155,N_2013,N_2068);
xor U2156 (N_2156,N_2089,N_2098);
and U2157 (N_2157,N_2016,N_2020);
or U2158 (N_2158,N_2067,N_2026);
nand U2159 (N_2159,N_2019,N_2041);
or U2160 (N_2160,N_2059,N_2024);
nand U2161 (N_2161,N_2077,N_2058);
nor U2162 (N_2162,N_2067,N_2078);
nand U2163 (N_2163,N_2034,N_2043);
and U2164 (N_2164,N_2034,N_2072);
xnor U2165 (N_2165,N_2074,N_2022);
xor U2166 (N_2166,N_2065,N_2014);
and U2167 (N_2167,N_2010,N_2079);
xor U2168 (N_2168,N_2081,N_2048);
nor U2169 (N_2169,N_2068,N_2088);
nor U2170 (N_2170,N_2061,N_2024);
xnor U2171 (N_2171,N_2085,N_2023);
or U2172 (N_2172,N_2088,N_2071);
xnor U2173 (N_2173,N_2030,N_2083);
and U2174 (N_2174,N_2022,N_2058);
nand U2175 (N_2175,N_2019,N_2032);
or U2176 (N_2176,N_2018,N_2047);
nor U2177 (N_2177,N_2044,N_2023);
nand U2178 (N_2178,N_2004,N_2045);
or U2179 (N_2179,N_2048,N_2094);
nand U2180 (N_2180,N_2015,N_2052);
or U2181 (N_2181,N_2096,N_2033);
nand U2182 (N_2182,N_2093,N_2019);
xor U2183 (N_2183,N_2016,N_2034);
nand U2184 (N_2184,N_2099,N_2013);
nor U2185 (N_2185,N_2048,N_2047);
nor U2186 (N_2186,N_2003,N_2076);
nor U2187 (N_2187,N_2094,N_2028);
xnor U2188 (N_2188,N_2010,N_2038);
or U2189 (N_2189,N_2071,N_2067);
or U2190 (N_2190,N_2091,N_2015);
or U2191 (N_2191,N_2019,N_2026);
nand U2192 (N_2192,N_2023,N_2068);
nor U2193 (N_2193,N_2082,N_2093);
nand U2194 (N_2194,N_2024,N_2029);
nor U2195 (N_2195,N_2006,N_2002);
or U2196 (N_2196,N_2043,N_2010);
xnor U2197 (N_2197,N_2071,N_2096);
xor U2198 (N_2198,N_2061,N_2071);
or U2199 (N_2199,N_2067,N_2079);
or U2200 (N_2200,N_2150,N_2135);
or U2201 (N_2201,N_2152,N_2140);
nor U2202 (N_2202,N_2170,N_2117);
nand U2203 (N_2203,N_2185,N_2193);
xor U2204 (N_2204,N_2154,N_2141);
nor U2205 (N_2205,N_2123,N_2105);
xor U2206 (N_2206,N_2155,N_2132);
nand U2207 (N_2207,N_2113,N_2166);
or U2208 (N_2208,N_2176,N_2108);
and U2209 (N_2209,N_2180,N_2129);
and U2210 (N_2210,N_2133,N_2102);
nor U2211 (N_2211,N_2192,N_2196);
or U2212 (N_2212,N_2134,N_2171);
nand U2213 (N_2213,N_2158,N_2194);
or U2214 (N_2214,N_2191,N_2173);
and U2215 (N_2215,N_2122,N_2167);
or U2216 (N_2216,N_2157,N_2137);
and U2217 (N_2217,N_2115,N_2151);
nand U2218 (N_2218,N_2146,N_2127);
and U2219 (N_2219,N_2164,N_2109);
xnor U2220 (N_2220,N_2149,N_2195);
xor U2221 (N_2221,N_2183,N_2100);
and U2222 (N_2222,N_2186,N_2116);
and U2223 (N_2223,N_2131,N_2199);
and U2224 (N_2224,N_2107,N_2101);
and U2225 (N_2225,N_2188,N_2153);
or U2226 (N_2226,N_2120,N_2178);
nor U2227 (N_2227,N_2174,N_2175);
or U2228 (N_2228,N_2197,N_2104);
xor U2229 (N_2229,N_2163,N_2125);
or U2230 (N_2230,N_2142,N_2148);
and U2231 (N_2231,N_2126,N_2103);
xor U2232 (N_2232,N_2144,N_2130);
xor U2233 (N_2233,N_2172,N_2160);
xnor U2234 (N_2234,N_2143,N_2114);
and U2235 (N_2235,N_2187,N_2184);
nand U2236 (N_2236,N_2121,N_2159);
and U2237 (N_2237,N_2111,N_2179);
and U2238 (N_2238,N_2145,N_2147);
nand U2239 (N_2239,N_2169,N_2128);
or U2240 (N_2240,N_2106,N_2165);
nor U2241 (N_2241,N_2181,N_2118);
xor U2242 (N_2242,N_2189,N_2177);
nor U2243 (N_2243,N_2124,N_2110);
nor U2244 (N_2244,N_2190,N_2182);
nor U2245 (N_2245,N_2119,N_2156);
nand U2246 (N_2246,N_2138,N_2198);
nor U2247 (N_2247,N_2139,N_2168);
or U2248 (N_2248,N_2162,N_2112);
nand U2249 (N_2249,N_2136,N_2161);
nor U2250 (N_2250,N_2190,N_2169);
and U2251 (N_2251,N_2137,N_2134);
or U2252 (N_2252,N_2157,N_2160);
or U2253 (N_2253,N_2102,N_2117);
nand U2254 (N_2254,N_2196,N_2133);
nor U2255 (N_2255,N_2153,N_2191);
nand U2256 (N_2256,N_2190,N_2143);
or U2257 (N_2257,N_2164,N_2197);
nand U2258 (N_2258,N_2143,N_2196);
nand U2259 (N_2259,N_2118,N_2153);
nor U2260 (N_2260,N_2196,N_2141);
nor U2261 (N_2261,N_2149,N_2179);
nand U2262 (N_2262,N_2112,N_2120);
xnor U2263 (N_2263,N_2101,N_2189);
and U2264 (N_2264,N_2174,N_2116);
nand U2265 (N_2265,N_2187,N_2119);
xnor U2266 (N_2266,N_2178,N_2143);
or U2267 (N_2267,N_2124,N_2166);
nand U2268 (N_2268,N_2169,N_2124);
or U2269 (N_2269,N_2114,N_2187);
or U2270 (N_2270,N_2140,N_2155);
xnor U2271 (N_2271,N_2130,N_2183);
nand U2272 (N_2272,N_2195,N_2140);
nand U2273 (N_2273,N_2180,N_2175);
xnor U2274 (N_2274,N_2145,N_2127);
or U2275 (N_2275,N_2170,N_2198);
nor U2276 (N_2276,N_2182,N_2144);
or U2277 (N_2277,N_2148,N_2156);
and U2278 (N_2278,N_2173,N_2116);
nor U2279 (N_2279,N_2103,N_2162);
nor U2280 (N_2280,N_2192,N_2136);
nor U2281 (N_2281,N_2108,N_2162);
nand U2282 (N_2282,N_2108,N_2166);
and U2283 (N_2283,N_2146,N_2106);
nor U2284 (N_2284,N_2119,N_2162);
nand U2285 (N_2285,N_2105,N_2148);
or U2286 (N_2286,N_2101,N_2177);
nor U2287 (N_2287,N_2105,N_2122);
and U2288 (N_2288,N_2192,N_2190);
nor U2289 (N_2289,N_2136,N_2189);
and U2290 (N_2290,N_2173,N_2130);
or U2291 (N_2291,N_2171,N_2173);
nor U2292 (N_2292,N_2115,N_2193);
and U2293 (N_2293,N_2127,N_2153);
nand U2294 (N_2294,N_2175,N_2171);
nand U2295 (N_2295,N_2101,N_2190);
nand U2296 (N_2296,N_2102,N_2105);
xnor U2297 (N_2297,N_2109,N_2104);
and U2298 (N_2298,N_2109,N_2138);
xor U2299 (N_2299,N_2190,N_2174);
xor U2300 (N_2300,N_2200,N_2260);
xnor U2301 (N_2301,N_2250,N_2238);
and U2302 (N_2302,N_2229,N_2299);
xor U2303 (N_2303,N_2234,N_2265);
nor U2304 (N_2304,N_2277,N_2243);
xnor U2305 (N_2305,N_2251,N_2271);
xor U2306 (N_2306,N_2298,N_2264);
nor U2307 (N_2307,N_2285,N_2228);
and U2308 (N_2308,N_2256,N_2205);
xor U2309 (N_2309,N_2246,N_2221);
nand U2310 (N_2310,N_2293,N_2248);
or U2311 (N_2311,N_2276,N_2270);
nand U2312 (N_2312,N_2279,N_2295);
and U2313 (N_2313,N_2219,N_2239);
nand U2314 (N_2314,N_2252,N_2213);
nand U2315 (N_2315,N_2263,N_2261);
nor U2316 (N_2316,N_2280,N_2236);
nand U2317 (N_2317,N_2286,N_2284);
nand U2318 (N_2318,N_2258,N_2201);
nand U2319 (N_2319,N_2220,N_2267);
nor U2320 (N_2320,N_2259,N_2273);
or U2321 (N_2321,N_2296,N_2240);
nand U2322 (N_2322,N_2289,N_2241);
nand U2323 (N_2323,N_2202,N_2245);
and U2324 (N_2324,N_2257,N_2247);
xnor U2325 (N_2325,N_2216,N_2275);
xor U2326 (N_2326,N_2214,N_2203);
nor U2327 (N_2327,N_2288,N_2231);
nand U2328 (N_2328,N_2209,N_2215);
nand U2329 (N_2329,N_2269,N_2292);
nor U2330 (N_2330,N_2232,N_2274);
xor U2331 (N_2331,N_2272,N_2233);
and U2332 (N_2332,N_2254,N_2268);
xnor U2333 (N_2333,N_2222,N_2283);
nand U2334 (N_2334,N_2224,N_2297);
nand U2335 (N_2335,N_2208,N_2225);
and U2336 (N_2336,N_2218,N_2235);
nor U2337 (N_2337,N_2206,N_2282);
nand U2338 (N_2338,N_2237,N_2207);
and U2339 (N_2339,N_2290,N_2217);
xnor U2340 (N_2340,N_2262,N_2212);
xnor U2341 (N_2341,N_2242,N_2244);
and U2342 (N_2342,N_2249,N_2287);
xor U2343 (N_2343,N_2223,N_2291);
xnor U2344 (N_2344,N_2281,N_2227);
or U2345 (N_2345,N_2255,N_2211);
and U2346 (N_2346,N_2253,N_2210);
or U2347 (N_2347,N_2278,N_2266);
xnor U2348 (N_2348,N_2294,N_2204);
nor U2349 (N_2349,N_2230,N_2226);
or U2350 (N_2350,N_2252,N_2241);
xnor U2351 (N_2351,N_2204,N_2289);
nor U2352 (N_2352,N_2209,N_2224);
and U2353 (N_2353,N_2283,N_2299);
and U2354 (N_2354,N_2202,N_2211);
or U2355 (N_2355,N_2285,N_2206);
or U2356 (N_2356,N_2248,N_2227);
and U2357 (N_2357,N_2263,N_2206);
or U2358 (N_2358,N_2293,N_2245);
and U2359 (N_2359,N_2278,N_2227);
nand U2360 (N_2360,N_2226,N_2218);
or U2361 (N_2361,N_2256,N_2245);
xor U2362 (N_2362,N_2262,N_2217);
xor U2363 (N_2363,N_2282,N_2271);
or U2364 (N_2364,N_2263,N_2230);
and U2365 (N_2365,N_2260,N_2275);
xor U2366 (N_2366,N_2299,N_2227);
xnor U2367 (N_2367,N_2288,N_2218);
xnor U2368 (N_2368,N_2246,N_2216);
or U2369 (N_2369,N_2244,N_2232);
or U2370 (N_2370,N_2273,N_2205);
xor U2371 (N_2371,N_2234,N_2288);
nand U2372 (N_2372,N_2231,N_2296);
nand U2373 (N_2373,N_2227,N_2252);
nor U2374 (N_2374,N_2281,N_2201);
and U2375 (N_2375,N_2239,N_2207);
and U2376 (N_2376,N_2250,N_2284);
and U2377 (N_2377,N_2230,N_2210);
or U2378 (N_2378,N_2250,N_2267);
and U2379 (N_2379,N_2293,N_2220);
and U2380 (N_2380,N_2235,N_2230);
xnor U2381 (N_2381,N_2200,N_2296);
nand U2382 (N_2382,N_2266,N_2214);
and U2383 (N_2383,N_2205,N_2253);
or U2384 (N_2384,N_2298,N_2249);
nand U2385 (N_2385,N_2208,N_2280);
and U2386 (N_2386,N_2296,N_2261);
nor U2387 (N_2387,N_2274,N_2264);
nor U2388 (N_2388,N_2286,N_2285);
xor U2389 (N_2389,N_2266,N_2232);
nor U2390 (N_2390,N_2209,N_2251);
or U2391 (N_2391,N_2292,N_2257);
and U2392 (N_2392,N_2219,N_2216);
and U2393 (N_2393,N_2225,N_2240);
nor U2394 (N_2394,N_2259,N_2200);
xnor U2395 (N_2395,N_2257,N_2222);
nand U2396 (N_2396,N_2216,N_2241);
xnor U2397 (N_2397,N_2213,N_2216);
xor U2398 (N_2398,N_2258,N_2227);
or U2399 (N_2399,N_2297,N_2228);
nand U2400 (N_2400,N_2359,N_2369);
nand U2401 (N_2401,N_2306,N_2371);
or U2402 (N_2402,N_2325,N_2364);
nand U2403 (N_2403,N_2391,N_2356);
xnor U2404 (N_2404,N_2311,N_2337);
or U2405 (N_2405,N_2326,N_2310);
nand U2406 (N_2406,N_2386,N_2397);
nor U2407 (N_2407,N_2342,N_2333);
xnor U2408 (N_2408,N_2318,N_2366);
nand U2409 (N_2409,N_2316,N_2381);
or U2410 (N_2410,N_2330,N_2301);
xor U2411 (N_2411,N_2377,N_2376);
and U2412 (N_2412,N_2322,N_2302);
or U2413 (N_2413,N_2320,N_2334);
and U2414 (N_2414,N_2388,N_2354);
nand U2415 (N_2415,N_2383,N_2358);
nand U2416 (N_2416,N_2379,N_2343);
nand U2417 (N_2417,N_2355,N_2387);
or U2418 (N_2418,N_2378,N_2393);
nand U2419 (N_2419,N_2347,N_2372);
nand U2420 (N_2420,N_2396,N_2319);
xnor U2421 (N_2421,N_2307,N_2394);
nor U2422 (N_2422,N_2340,N_2346);
nor U2423 (N_2423,N_2367,N_2314);
xnor U2424 (N_2424,N_2350,N_2308);
and U2425 (N_2425,N_2336,N_2363);
and U2426 (N_2426,N_2321,N_2352);
nand U2427 (N_2427,N_2360,N_2373);
nand U2428 (N_2428,N_2380,N_2365);
or U2429 (N_2429,N_2390,N_2362);
nand U2430 (N_2430,N_2312,N_2324);
or U2431 (N_2431,N_2385,N_2348);
xnor U2432 (N_2432,N_2305,N_2370);
nand U2433 (N_2433,N_2399,N_2328);
and U2434 (N_2434,N_2304,N_2395);
nor U2435 (N_2435,N_2392,N_2353);
or U2436 (N_2436,N_2398,N_2357);
xor U2437 (N_2437,N_2374,N_2315);
nand U2438 (N_2438,N_2313,N_2317);
xnor U2439 (N_2439,N_2331,N_2382);
nand U2440 (N_2440,N_2309,N_2345);
xnor U2441 (N_2441,N_2338,N_2384);
xor U2442 (N_2442,N_2323,N_2341);
nand U2443 (N_2443,N_2389,N_2335);
xor U2444 (N_2444,N_2329,N_2303);
xnor U2445 (N_2445,N_2349,N_2361);
and U2446 (N_2446,N_2339,N_2368);
nor U2447 (N_2447,N_2327,N_2332);
or U2448 (N_2448,N_2351,N_2344);
nand U2449 (N_2449,N_2375,N_2300);
nand U2450 (N_2450,N_2348,N_2375);
nand U2451 (N_2451,N_2350,N_2368);
and U2452 (N_2452,N_2393,N_2321);
xnor U2453 (N_2453,N_2350,N_2355);
nor U2454 (N_2454,N_2324,N_2311);
nand U2455 (N_2455,N_2396,N_2370);
and U2456 (N_2456,N_2382,N_2363);
or U2457 (N_2457,N_2379,N_2399);
xnor U2458 (N_2458,N_2391,N_2347);
nor U2459 (N_2459,N_2358,N_2363);
nand U2460 (N_2460,N_2370,N_2335);
nand U2461 (N_2461,N_2353,N_2312);
nor U2462 (N_2462,N_2396,N_2374);
xnor U2463 (N_2463,N_2367,N_2363);
and U2464 (N_2464,N_2332,N_2318);
or U2465 (N_2465,N_2347,N_2332);
or U2466 (N_2466,N_2371,N_2309);
and U2467 (N_2467,N_2312,N_2304);
or U2468 (N_2468,N_2351,N_2361);
nor U2469 (N_2469,N_2337,N_2320);
nor U2470 (N_2470,N_2307,N_2324);
and U2471 (N_2471,N_2300,N_2383);
xor U2472 (N_2472,N_2370,N_2345);
nor U2473 (N_2473,N_2321,N_2344);
nand U2474 (N_2474,N_2329,N_2353);
or U2475 (N_2475,N_2348,N_2387);
or U2476 (N_2476,N_2337,N_2358);
and U2477 (N_2477,N_2321,N_2315);
nand U2478 (N_2478,N_2319,N_2355);
or U2479 (N_2479,N_2301,N_2358);
or U2480 (N_2480,N_2347,N_2338);
nor U2481 (N_2481,N_2363,N_2312);
nor U2482 (N_2482,N_2393,N_2358);
and U2483 (N_2483,N_2347,N_2364);
xnor U2484 (N_2484,N_2336,N_2393);
nand U2485 (N_2485,N_2380,N_2314);
and U2486 (N_2486,N_2373,N_2312);
and U2487 (N_2487,N_2330,N_2352);
and U2488 (N_2488,N_2380,N_2304);
nor U2489 (N_2489,N_2333,N_2322);
nand U2490 (N_2490,N_2337,N_2398);
or U2491 (N_2491,N_2330,N_2326);
nand U2492 (N_2492,N_2379,N_2323);
and U2493 (N_2493,N_2305,N_2350);
and U2494 (N_2494,N_2375,N_2311);
nor U2495 (N_2495,N_2330,N_2373);
nand U2496 (N_2496,N_2373,N_2340);
and U2497 (N_2497,N_2316,N_2324);
nand U2498 (N_2498,N_2315,N_2313);
or U2499 (N_2499,N_2325,N_2330);
or U2500 (N_2500,N_2487,N_2414);
nand U2501 (N_2501,N_2402,N_2475);
or U2502 (N_2502,N_2412,N_2477);
nand U2503 (N_2503,N_2406,N_2443);
nor U2504 (N_2504,N_2459,N_2405);
xnor U2505 (N_2505,N_2411,N_2426);
and U2506 (N_2506,N_2438,N_2403);
nand U2507 (N_2507,N_2499,N_2495);
or U2508 (N_2508,N_2498,N_2481);
nor U2509 (N_2509,N_2488,N_2408);
nor U2510 (N_2510,N_2482,N_2424);
and U2511 (N_2511,N_2450,N_2478);
xor U2512 (N_2512,N_2452,N_2439);
xor U2513 (N_2513,N_2430,N_2471);
nand U2514 (N_2514,N_2431,N_2422);
nand U2515 (N_2515,N_2456,N_2444);
or U2516 (N_2516,N_2446,N_2483);
nand U2517 (N_2517,N_2416,N_2453);
and U2518 (N_2518,N_2428,N_2476);
and U2519 (N_2519,N_2436,N_2404);
nand U2520 (N_2520,N_2473,N_2465);
xor U2521 (N_2521,N_2448,N_2493);
and U2522 (N_2522,N_2485,N_2437);
or U2523 (N_2523,N_2409,N_2401);
and U2524 (N_2524,N_2464,N_2466);
or U2525 (N_2525,N_2479,N_2441);
xor U2526 (N_2526,N_2474,N_2492);
nor U2527 (N_2527,N_2467,N_2463);
nand U2528 (N_2528,N_2429,N_2421);
xnor U2529 (N_2529,N_2497,N_2461);
nor U2530 (N_2530,N_2420,N_2472);
and U2531 (N_2531,N_2410,N_2491);
or U2532 (N_2532,N_2417,N_2451);
nand U2533 (N_2533,N_2457,N_2469);
nand U2534 (N_2534,N_2486,N_2413);
nand U2535 (N_2535,N_2449,N_2445);
nand U2536 (N_2536,N_2480,N_2468);
or U2537 (N_2537,N_2489,N_2496);
and U2538 (N_2538,N_2460,N_2415);
xnor U2539 (N_2539,N_2454,N_2407);
nand U2540 (N_2540,N_2470,N_2484);
nor U2541 (N_2541,N_2435,N_2494);
nor U2542 (N_2542,N_2458,N_2432);
xnor U2543 (N_2543,N_2462,N_2418);
xnor U2544 (N_2544,N_2447,N_2442);
and U2545 (N_2545,N_2419,N_2423);
and U2546 (N_2546,N_2434,N_2425);
or U2547 (N_2547,N_2400,N_2433);
or U2548 (N_2548,N_2427,N_2490);
or U2549 (N_2549,N_2455,N_2440);
nor U2550 (N_2550,N_2494,N_2436);
or U2551 (N_2551,N_2460,N_2422);
xor U2552 (N_2552,N_2442,N_2479);
nand U2553 (N_2553,N_2436,N_2442);
nand U2554 (N_2554,N_2466,N_2446);
nand U2555 (N_2555,N_2471,N_2468);
or U2556 (N_2556,N_2426,N_2475);
nor U2557 (N_2557,N_2417,N_2459);
and U2558 (N_2558,N_2465,N_2405);
nand U2559 (N_2559,N_2418,N_2447);
nand U2560 (N_2560,N_2471,N_2490);
or U2561 (N_2561,N_2471,N_2480);
nor U2562 (N_2562,N_2419,N_2438);
xor U2563 (N_2563,N_2408,N_2468);
and U2564 (N_2564,N_2435,N_2414);
xor U2565 (N_2565,N_2438,N_2456);
or U2566 (N_2566,N_2424,N_2452);
nor U2567 (N_2567,N_2472,N_2441);
nand U2568 (N_2568,N_2463,N_2471);
xnor U2569 (N_2569,N_2400,N_2423);
nand U2570 (N_2570,N_2457,N_2499);
nor U2571 (N_2571,N_2418,N_2415);
nand U2572 (N_2572,N_2467,N_2446);
nand U2573 (N_2573,N_2495,N_2482);
and U2574 (N_2574,N_2441,N_2424);
nor U2575 (N_2575,N_2464,N_2472);
nor U2576 (N_2576,N_2451,N_2497);
and U2577 (N_2577,N_2440,N_2461);
or U2578 (N_2578,N_2466,N_2404);
nor U2579 (N_2579,N_2465,N_2438);
and U2580 (N_2580,N_2497,N_2431);
nor U2581 (N_2581,N_2473,N_2411);
nand U2582 (N_2582,N_2402,N_2449);
and U2583 (N_2583,N_2411,N_2498);
and U2584 (N_2584,N_2479,N_2498);
nor U2585 (N_2585,N_2436,N_2435);
xor U2586 (N_2586,N_2412,N_2426);
or U2587 (N_2587,N_2496,N_2499);
and U2588 (N_2588,N_2472,N_2474);
nor U2589 (N_2589,N_2421,N_2410);
or U2590 (N_2590,N_2435,N_2419);
nand U2591 (N_2591,N_2467,N_2414);
xor U2592 (N_2592,N_2465,N_2490);
nand U2593 (N_2593,N_2444,N_2415);
nor U2594 (N_2594,N_2427,N_2435);
or U2595 (N_2595,N_2443,N_2442);
or U2596 (N_2596,N_2460,N_2429);
or U2597 (N_2597,N_2446,N_2470);
nand U2598 (N_2598,N_2431,N_2454);
nand U2599 (N_2599,N_2483,N_2469);
or U2600 (N_2600,N_2599,N_2501);
or U2601 (N_2601,N_2576,N_2530);
xor U2602 (N_2602,N_2564,N_2557);
xor U2603 (N_2603,N_2529,N_2512);
xnor U2604 (N_2604,N_2594,N_2536);
nand U2605 (N_2605,N_2510,N_2524);
or U2606 (N_2606,N_2582,N_2586);
nand U2607 (N_2607,N_2548,N_2554);
nand U2608 (N_2608,N_2535,N_2587);
nor U2609 (N_2609,N_2571,N_2552);
nand U2610 (N_2610,N_2577,N_2598);
xnor U2611 (N_2611,N_2514,N_2511);
xor U2612 (N_2612,N_2589,N_2537);
nor U2613 (N_2613,N_2540,N_2561);
nor U2614 (N_2614,N_2555,N_2583);
and U2615 (N_2615,N_2585,N_2549);
xor U2616 (N_2616,N_2500,N_2580);
or U2617 (N_2617,N_2528,N_2525);
xor U2618 (N_2618,N_2559,N_2574);
and U2619 (N_2619,N_2568,N_2505);
and U2620 (N_2620,N_2547,N_2516);
nor U2621 (N_2621,N_2513,N_2575);
or U2622 (N_2622,N_2518,N_2523);
xor U2623 (N_2623,N_2543,N_2502);
nor U2624 (N_2624,N_2565,N_2531);
nor U2625 (N_2625,N_2515,N_2546);
and U2626 (N_2626,N_2504,N_2556);
xnor U2627 (N_2627,N_2590,N_2591);
or U2628 (N_2628,N_2592,N_2522);
nand U2629 (N_2629,N_2596,N_2541);
xor U2630 (N_2630,N_2527,N_2584);
or U2631 (N_2631,N_2508,N_2520);
xnor U2632 (N_2632,N_2534,N_2597);
or U2633 (N_2633,N_2569,N_2509);
or U2634 (N_2634,N_2566,N_2573);
nor U2635 (N_2635,N_2578,N_2538);
nor U2636 (N_2636,N_2570,N_2521);
xnor U2637 (N_2637,N_2506,N_2539);
and U2638 (N_2638,N_2579,N_2545);
nand U2639 (N_2639,N_2507,N_2595);
xnor U2640 (N_2640,N_2526,N_2567);
or U2641 (N_2641,N_2558,N_2542);
or U2642 (N_2642,N_2588,N_2581);
and U2643 (N_2643,N_2550,N_2533);
xor U2644 (N_2644,N_2560,N_2544);
xor U2645 (N_2645,N_2503,N_2572);
and U2646 (N_2646,N_2562,N_2593);
or U2647 (N_2647,N_2563,N_2553);
nand U2648 (N_2648,N_2532,N_2519);
nand U2649 (N_2649,N_2551,N_2517);
or U2650 (N_2650,N_2599,N_2593);
nand U2651 (N_2651,N_2512,N_2554);
nor U2652 (N_2652,N_2586,N_2552);
nand U2653 (N_2653,N_2526,N_2530);
nor U2654 (N_2654,N_2598,N_2535);
or U2655 (N_2655,N_2525,N_2562);
nor U2656 (N_2656,N_2580,N_2522);
or U2657 (N_2657,N_2521,N_2548);
nand U2658 (N_2658,N_2574,N_2543);
xnor U2659 (N_2659,N_2556,N_2527);
nand U2660 (N_2660,N_2551,N_2571);
xnor U2661 (N_2661,N_2539,N_2547);
and U2662 (N_2662,N_2546,N_2569);
nor U2663 (N_2663,N_2562,N_2581);
or U2664 (N_2664,N_2520,N_2533);
and U2665 (N_2665,N_2512,N_2578);
and U2666 (N_2666,N_2540,N_2578);
or U2667 (N_2667,N_2573,N_2506);
xnor U2668 (N_2668,N_2502,N_2535);
and U2669 (N_2669,N_2585,N_2519);
nand U2670 (N_2670,N_2544,N_2513);
nand U2671 (N_2671,N_2576,N_2511);
and U2672 (N_2672,N_2585,N_2507);
nor U2673 (N_2673,N_2518,N_2571);
xnor U2674 (N_2674,N_2558,N_2508);
nand U2675 (N_2675,N_2507,N_2584);
or U2676 (N_2676,N_2575,N_2591);
nor U2677 (N_2677,N_2549,N_2563);
and U2678 (N_2678,N_2530,N_2575);
nand U2679 (N_2679,N_2554,N_2577);
xor U2680 (N_2680,N_2528,N_2548);
nand U2681 (N_2681,N_2579,N_2529);
and U2682 (N_2682,N_2500,N_2565);
xor U2683 (N_2683,N_2515,N_2525);
and U2684 (N_2684,N_2571,N_2559);
nor U2685 (N_2685,N_2530,N_2522);
or U2686 (N_2686,N_2553,N_2545);
nand U2687 (N_2687,N_2521,N_2580);
nor U2688 (N_2688,N_2508,N_2501);
xor U2689 (N_2689,N_2516,N_2505);
xnor U2690 (N_2690,N_2598,N_2518);
nand U2691 (N_2691,N_2544,N_2583);
nand U2692 (N_2692,N_2556,N_2528);
and U2693 (N_2693,N_2581,N_2535);
xnor U2694 (N_2694,N_2510,N_2581);
xnor U2695 (N_2695,N_2597,N_2572);
and U2696 (N_2696,N_2509,N_2572);
or U2697 (N_2697,N_2550,N_2575);
or U2698 (N_2698,N_2586,N_2556);
xor U2699 (N_2699,N_2543,N_2558);
and U2700 (N_2700,N_2627,N_2661);
nand U2701 (N_2701,N_2656,N_2606);
and U2702 (N_2702,N_2605,N_2643);
or U2703 (N_2703,N_2624,N_2630);
and U2704 (N_2704,N_2611,N_2694);
nor U2705 (N_2705,N_2665,N_2684);
and U2706 (N_2706,N_2646,N_2629);
and U2707 (N_2707,N_2613,N_2600);
nand U2708 (N_2708,N_2692,N_2638);
nor U2709 (N_2709,N_2622,N_2648);
xor U2710 (N_2710,N_2663,N_2687);
nand U2711 (N_2711,N_2670,N_2659);
or U2712 (N_2712,N_2641,N_2653);
and U2713 (N_2713,N_2603,N_2657);
nor U2714 (N_2714,N_2676,N_2637);
nand U2715 (N_2715,N_2677,N_2655);
xor U2716 (N_2716,N_2602,N_2680);
and U2717 (N_2717,N_2635,N_2652);
or U2718 (N_2718,N_2612,N_2668);
xnor U2719 (N_2719,N_2673,N_2632);
xor U2720 (N_2720,N_2640,N_2697);
nor U2721 (N_2721,N_2626,N_2689);
xnor U2722 (N_2722,N_2617,N_2662);
nor U2723 (N_2723,N_2685,N_2628);
nand U2724 (N_2724,N_2696,N_2667);
nand U2725 (N_2725,N_2682,N_2647);
xor U2726 (N_2726,N_2679,N_2672);
xor U2727 (N_2727,N_2642,N_2671);
and U2728 (N_2728,N_2639,N_2690);
nand U2729 (N_2729,N_2660,N_2645);
nand U2730 (N_2730,N_2688,N_2601);
and U2731 (N_2731,N_2604,N_2619);
or U2732 (N_2732,N_2698,N_2669);
and U2733 (N_2733,N_2654,N_2631);
nor U2734 (N_2734,N_2650,N_2664);
nand U2735 (N_2735,N_2691,N_2681);
xnor U2736 (N_2736,N_2609,N_2699);
nand U2737 (N_2737,N_2678,N_2633);
or U2738 (N_2738,N_2651,N_2634);
and U2739 (N_2739,N_2674,N_2675);
nand U2740 (N_2740,N_2683,N_2658);
nand U2741 (N_2741,N_2644,N_2618);
nor U2742 (N_2742,N_2608,N_2666);
or U2743 (N_2743,N_2625,N_2623);
or U2744 (N_2744,N_2620,N_2610);
xnor U2745 (N_2745,N_2621,N_2615);
nand U2746 (N_2746,N_2616,N_2649);
xor U2747 (N_2747,N_2686,N_2636);
or U2748 (N_2748,N_2614,N_2607);
and U2749 (N_2749,N_2693,N_2695);
xnor U2750 (N_2750,N_2660,N_2623);
nor U2751 (N_2751,N_2661,N_2688);
or U2752 (N_2752,N_2637,N_2610);
nand U2753 (N_2753,N_2677,N_2603);
or U2754 (N_2754,N_2665,N_2643);
or U2755 (N_2755,N_2659,N_2678);
and U2756 (N_2756,N_2643,N_2677);
nor U2757 (N_2757,N_2608,N_2628);
and U2758 (N_2758,N_2687,N_2698);
and U2759 (N_2759,N_2658,N_2619);
or U2760 (N_2760,N_2674,N_2654);
or U2761 (N_2761,N_2646,N_2612);
nor U2762 (N_2762,N_2661,N_2640);
xnor U2763 (N_2763,N_2659,N_2615);
or U2764 (N_2764,N_2645,N_2661);
and U2765 (N_2765,N_2695,N_2617);
nor U2766 (N_2766,N_2637,N_2687);
and U2767 (N_2767,N_2630,N_2610);
nor U2768 (N_2768,N_2659,N_2652);
and U2769 (N_2769,N_2653,N_2608);
or U2770 (N_2770,N_2651,N_2696);
and U2771 (N_2771,N_2619,N_2663);
nand U2772 (N_2772,N_2661,N_2637);
nand U2773 (N_2773,N_2631,N_2649);
nor U2774 (N_2774,N_2677,N_2630);
nand U2775 (N_2775,N_2654,N_2623);
and U2776 (N_2776,N_2609,N_2634);
nand U2777 (N_2777,N_2609,N_2650);
and U2778 (N_2778,N_2668,N_2662);
or U2779 (N_2779,N_2688,N_2694);
nor U2780 (N_2780,N_2691,N_2649);
and U2781 (N_2781,N_2680,N_2630);
xor U2782 (N_2782,N_2607,N_2652);
and U2783 (N_2783,N_2631,N_2612);
and U2784 (N_2784,N_2647,N_2631);
nand U2785 (N_2785,N_2694,N_2666);
xor U2786 (N_2786,N_2662,N_2676);
nor U2787 (N_2787,N_2693,N_2680);
and U2788 (N_2788,N_2651,N_2695);
or U2789 (N_2789,N_2621,N_2680);
xor U2790 (N_2790,N_2668,N_2672);
nand U2791 (N_2791,N_2641,N_2690);
xnor U2792 (N_2792,N_2647,N_2628);
or U2793 (N_2793,N_2668,N_2673);
and U2794 (N_2794,N_2673,N_2636);
or U2795 (N_2795,N_2661,N_2606);
xor U2796 (N_2796,N_2604,N_2679);
and U2797 (N_2797,N_2632,N_2661);
and U2798 (N_2798,N_2637,N_2670);
xnor U2799 (N_2799,N_2666,N_2652);
nor U2800 (N_2800,N_2793,N_2775);
nand U2801 (N_2801,N_2791,N_2722);
and U2802 (N_2802,N_2726,N_2706);
and U2803 (N_2803,N_2748,N_2730);
nand U2804 (N_2804,N_2777,N_2733);
nand U2805 (N_2805,N_2717,N_2729);
nand U2806 (N_2806,N_2792,N_2786);
and U2807 (N_2807,N_2737,N_2742);
nand U2808 (N_2808,N_2788,N_2721);
nand U2809 (N_2809,N_2732,N_2746);
or U2810 (N_2810,N_2728,N_2707);
nand U2811 (N_2811,N_2709,N_2738);
nand U2812 (N_2812,N_2781,N_2795);
and U2813 (N_2813,N_2711,N_2714);
or U2814 (N_2814,N_2704,N_2794);
or U2815 (N_2815,N_2718,N_2713);
nand U2816 (N_2816,N_2778,N_2789);
nand U2817 (N_2817,N_2770,N_2710);
nor U2818 (N_2818,N_2797,N_2725);
nor U2819 (N_2819,N_2752,N_2767);
xor U2820 (N_2820,N_2749,N_2796);
nor U2821 (N_2821,N_2739,N_2702);
xnor U2822 (N_2822,N_2774,N_2762);
and U2823 (N_2823,N_2727,N_2772);
nand U2824 (N_2824,N_2741,N_2724);
and U2825 (N_2825,N_2712,N_2745);
or U2826 (N_2826,N_2785,N_2740);
and U2827 (N_2827,N_2780,N_2716);
xor U2828 (N_2828,N_2769,N_2759);
nand U2829 (N_2829,N_2735,N_2719);
or U2830 (N_2830,N_2768,N_2743);
nor U2831 (N_2831,N_2723,N_2708);
nand U2832 (N_2832,N_2771,N_2753);
and U2833 (N_2833,N_2734,N_2715);
xor U2834 (N_2834,N_2701,N_2736);
xor U2835 (N_2835,N_2757,N_2790);
xor U2836 (N_2836,N_2744,N_2798);
nand U2837 (N_2837,N_2705,N_2765);
or U2838 (N_2838,N_2766,N_2750);
nor U2839 (N_2839,N_2756,N_2760);
or U2840 (N_2840,N_2700,N_2754);
or U2841 (N_2841,N_2720,N_2773);
and U2842 (N_2842,N_2761,N_2783);
nor U2843 (N_2843,N_2755,N_2776);
nand U2844 (N_2844,N_2764,N_2763);
xnor U2845 (N_2845,N_2703,N_2751);
xnor U2846 (N_2846,N_2799,N_2782);
xor U2847 (N_2847,N_2731,N_2787);
or U2848 (N_2848,N_2779,N_2784);
nand U2849 (N_2849,N_2747,N_2758);
nand U2850 (N_2850,N_2799,N_2722);
and U2851 (N_2851,N_2765,N_2775);
or U2852 (N_2852,N_2763,N_2731);
and U2853 (N_2853,N_2763,N_2769);
and U2854 (N_2854,N_2799,N_2703);
nand U2855 (N_2855,N_2753,N_2782);
xor U2856 (N_2856,N_2706,N_2750);
and U2857 (N_2857,N_2733,N_2740);
nand U2858 (N_2858,N_2731,N_2798);
nor U2859 (N_2859,N_2700,N_2783);
or U2860 (N_2860,N_2789,N_2795);
nand U2861 (N_2861,N_2794,N_2754);
and U2862 (N_2862,N_2744,N_2758);
nor U2863 (N_2863,N_2750,N_2707);
nand U2864 (N_2864,N_2756,N_2700);
nor U2865 (N_2865,N_2739,N_2767);
nor U2866 (N_2866,N_2765,N_2744);
and U2867 (N_2867,N_2783,N_2725);
and U2868 (N_2868,N_2790,N_2780);
nand U2869 (N_2869,N_2702,N_2772);
nand U2870 (N_2870,N_2782,N_2739);
or U2871 (N_2871,N_2798,N_2758);
and U2872 (N_2872,N_2755,N_2739);
nand U2873 (N_2873,N_2700,N_2722);
nor U2874 (N_2874,N_2754,N_2779);
and U2875 (N_2875,N_2745,N_2748);
or U2876 (N_2876,N_2770,N_2781);
nor U2877 (N_2877,N_2736,N_2722);
nor U2878 (N_2878,N_2768,N_2795);
or U2879 (N_2879,N_2783,N_2740);
or U2880 (N_2880,N_2783,N_2798);
and U2881 (N_2881,N_2741,N_2737);
or U2882 (N_2882,N_2720,N_2778);
nand U2883 (N_2883,N_2761,N_2702);
and U2884 (N_2884,N_2731,N_2702);
or U2885 (N_2885,N_2725,N_2722);
or U2886 (N_2886,N_2705,N_2779);
xor U2887 (N_2887,N_2778,N_2770);
or U2888 (N_2888,N_2798,N_2716);
nand U2889 (N_2889,N_2772,N_2793);
nor U2890 (N_2890,N_2721,N_2767);
and U2891 (N_2891,N_2764,N_2760);
nor U2892 (N_2892,N_2739,N_2789);
xnor U2893 (N_2893,N_2704,N_2740);
xnor U2894 (N_2894,N_2753,N_2731);
xnor U2895 (N_2895,N_2749,N_2751);
xor U2896 (N_2896,N_2786,N_2740);
nand U2897 (N_2897,N_2775,N_2784);
or U2898 (N_2898,N_2747,N_2704);
nor U2899 (N_2899,N_2720,N_2743);
and U2900 (N_2900,N_2830,N_2805);
or U2901 (N_2901,N_2823,N_2887);
and U2902 (N_2902,N_2814,N_2860);
and U2903 (N_2903,N_2884,N_2897);
and U2904 (N_2904,N_2820,N_2877);
or U2905 (N_2905,N_2876,N_2826);
nand U2906 (N_2906,N_2899,N_2852);
and U2907 (N_2907,N_2881,N_2813);
xor U2908 (N_2908,N_2893,N_2828);
and U2909 (N_2909,N_2803,N_2840);
nor U2910 (N_2910,N_2888,N_2800);
xor U2911 (N_2911,N_2812,N_2836);
xnor U2912 (N_2912,N_2817,N_2844);
or U2913 (N_2913,N_2848,N_2802);
nor U2914 (N_2914,N_2846,N_2853);
nor U2915 (N_2915,N_2895,N_2808);
nor U2916 (N_2916,N_2815,N_2850);
xnor U2917 (N_2917,N_2870,N_2890);
or U2918 (N_2918,N_2874,N_2818);
or U2919 (N_2919,N_2863,N_2861);
or U2920 (N_2920,N_2891,N_2898);
xor U2921 (N_2921,N_2824,N_2885);
xor U2922 (N_2922,N_2892,N_2859);
xnor U2923 (N_2923,N_2886,N_2810);
xnor U2924 (N_2924,N_2883,N_2829);
xnor U2925 (N_2925,N_2879,N_2894);
xor U2926 (N_2926,N_2831,N_2875);
nor U2927 (N_2927,N_2871,N_2867);
nor U2928 (N_2928,N_2849,N_2842);
or U2929 (N_2929,N_2845,N_2839);
and U2930 (N_2930,N_2841,N_2851);
nor U2931 (N_2931,N_2809,N_2832);
nor U2932 (N_2932,N_2827,N_2864);
and U2933 (N_2933,N_2835,N_2837);
xor U2934 (N_2934,N_2866,N_2825);
or U2935 (N_2935,N_2843,N_2855);
nor U2936 (N_2936,N_2807,N_2847);
xnor U2937 (N_2937,N_2857,N_2821);
nand U2938 (N_2938,N_2896,N_2872);
xor U2939 (N_2939,N_2819,N_2889);
or U2940 (N_2940,N_2873,N_2834);
nand U2941 (N_2941,N_2865,N_2854);
and U2942 (N_2942,N_2811,N_2868);
or U2943 (N_2943,N_2858,N_2862);
nand U2944 (N_2944,N_2838,N_2822);
nand U2945 (N_2945,N_2816,N_2804);
nor U2946 (N_2946,N_2880,N_2856);
and U2947 (N_2947,N_2869,N_2878);
nor U2948 (N_2948,N_2806,N_2833);
nand U2949 (N_2949,N_2801,N_2882);
nor U2950 (N_2950,N_2820,N_2895);
xnor U2951 (N_2951,N_2850,N_2863);
xor U2952 (N_2952,N_2816,N_2836);
xor U2953 (N_2953,N_2856,N_2841);
nor U2954 (N_2954,N_2861,N_2834);
xnor U2955 (N_2955,N_2847,N_2831);
xor U2956 (N_2956,N_2853,N_2830);
xnor U2957 (N_2957,N_2870,N_2810);
and U2958 (N_2958,N_2815,N_2878);
nor U2959 (N_2959,N_2816,N_2834);
nand U2960 (N_2960,N_2851,N_2890);
or U2961 (N_2961,N_2822,N_2899);
nor U2962 (N_2962,N_2883,N_2881);
nor U2963 (N_2963,N_2862,N_2861);
and U2964 (N_2964,N_2890,N_2858);
and U2965 (N_2965,N_2896,N_2866);
nor U2966 (N_2966,N_2802,N_2865);
nor U2967 (N_2967,N_2875,N_2852);
nor U2968 (N_2968,N_2839,N_2854);
nor U2969 (N_2969,N_2835,N_2832);
and U2970 (N_2970,N_2855,N_2881);
and U2971 (N_2971,N_2833,N_2857);
and U2972 (N_2972,N_2888,N_2805);
nor U2973 (N_2973,N_2839,N_2851);
and U2974 (N_2974,N_2892,N_2823);
xnor U2975 (N_2975,N_2800,N_2866);
or U2976 (N_2976,N_2849,N_2882);
xor U2977 (N_2977,N_2821,N_2853);
and U2978 (N_2978,N_2868,N_2858);
nor U2979 (N_2979,N_2818,N_2856);
and U2980 (N_2980,N_2807,N_2819);
nor U2981 (N_2981,N_2842,N_2839);
nor U2982 (N_2982,N_2818,N_2862);
or U2983 (N_2983,N_2816,N_2841);
nor U2984 (N_2984,N_2888,N_2822);
or U2985 (N_2985,N_2820,N_2804);
nor U2986 (N_2986,N_2889,N_2837);
and U2987 (N_2987,N_2888,N_2899);
or U2988 (N_2988,N_2886,N_2877);
and U2989 (N_2989,N_2867,N_2801);
nor U2990 (N_2990,N_2886,N_2887);
and U2991 (N_2991,N_2871,N_2834);
xor U2992 (N_2992,N_2800,N_2869);
xor U2993 (N_2993,N_2849,N_2846);
xnor U2994 (N_2994,N_2850,N_2875);
and U2995 (N_2995,N_2864,N_2863);
or U2996 (N_2996,N_2894,N_2874);
or U2997 (N_2997,N_2884,N_2886);
and U2998 (N_2998,N_2839,N_2807);
nand U2999 (N_2999,N_2827,N_2808);
nor U3000 (N_3000,N_2923,N_2968);
or U3001 (N_3001,N_2951,N_2907);
and U3002 (N_3002,N_2902,N_2988);
nor U3003 (N_3003,N_2904,N_2986);
or U3004 (N_3004,N_2917,N_2950);
or U3005 (N_3005,N_2937,N_2928);
xor U3006 (N_3006,N_2945,N_2962);
xor U3007 (N_3007,N_2956,N_2933);
nand U3008 (N_3008,N_2948,N_2903);
xor U3009 (N_3009,N_2957,N_2967);
or U3010 (N_3010,N_2906,N_2999);
or U3011 (N_3011,N_2946,N_2905);
nor U3012 (N_3012,N_2949,N_2911);
nand U3013 (N_3013,N_2970,N_2974);
nor U3014 (N_3014,N_2920,N_2958);
and U3015 (N_3015,N_2916,N_2922);
nor U3016 (N_3016,N_2924,N_2984);
xnor U3017 (N_3017,N_2982,N_2979);
xor U3018 (N_3018,N_2925,N_2981);
xor U3019 (N_3019,N_2991,N_2936);
or U3020 (N_3020,N_2919,N_2989);
xor U3021 (N_3021,N_2966,N_2901);
nor U3022 (N_3022,N_2963,N_2934);
or U3023 (N_3023,N_2929,N_2975);
and U3024 (N_3024,N_2995,N_2947);
nand U3025 (N_3025,N_2927,N_2913);
or U3026 (N_3026,N_2943,N_2940);
nor U3027 (N_3027,N_2985,N_2910);
xor U3028 (N_3028,N_2930,N_2980);
and U3029 (N_3029,N_2977,N_2973);
xor U3030 (N_3030,N_2965,N_2909);
or U3031 (N_3031,N_2972,N_2976);
xor U3032 (N_3032,N_2944,N_2953);
nor U3033 (N_3033,N_2938,N_2939);
nor U3034 (N_3034,N_2996,N_2954);
or U3035 (N_3035,N_2918,N_2915);
nand U3036 (N_3036,N_2969,N_2900);
and U3037 (N_3037,N_2912,N_2990);
and U3038 (N_3038,N_2932,N_2960);
xor U3039 (N_3039,N_2971,N_2942);
and U3040 (N_3040,N_2993,N_2955);
or U3041 (N_3041,N_2992,N_2983);
or U3042 (N_3042,N_2921,N_2959);
nor U3043 (N_3043,N_2978,N_2926);
nor U3044 (N_3044,N_2935,N_2941);
nand U3045 (N_3045,N_2961,N_2908);
or U3046 (N_3046,N_2914,N_2994);
nor U3047 (N_3047,N_2997,N_2998);
and U3048 (N_3048,N_2964,N_2987);
or U3049 (N_3049,N_2931,N_2952);
xor U3050 (N_3050,N_2981,N_2998);
and U3051 (N_3051,N_2929,N_2944);
xor U3052 (N_3052,N_2945,N_2994);
nand U3053 (N_3053,N_2978,N_2921);
and U3054 (N_3054,N_2983,N_2947);
nor U3055 (N_3055,N_2911,N_2992);
or U3056 (N_3056,N_2967,N_2934);
nor U3057 (N_3057,N_2962,N_2912);
nand U3058 (N_3058,N_2932,N_2951);
and U3059 (N_3059,N_2913,N_2949);
nor U3060 (N_3060,N_2953,N_2905);
or U3061 (N_3061,N_2928,N_2976);
and U3062 (N_3062,N_2963,N_2980);
xnor U3063 (N_3063,N_2974,N_2961);
or U3064 (N_3064,N_2942,N_2951);
nor U3065 (N_3065,N_2950,N_2954);
or U3066 (N_3066,N_2944,N_2974);
or U3067 (N_3067,N_2919,N_2914);
xor U3068 (N_3068,N_2922,N_2947);
or U3069 (N_3069,N_2980,N_2961);
nand U3070 (N_3070,N_2990,N_2954);
nand U3071 (N_3071,N_2997,N_2957);
or U3072 (N_3072,N_2980,N_2967);
nand U3073 (N_3073,N_2963,N_2935);
or U3074 (N_3074,N_2915,N_2938);
xor U3075 (N_3075,N_2986,N_2925);
nand U3076 (N_3076,N_2914,N_2988);
xor U3077 (N_3077,N_2938,N_2943);
xnor U3078 (N_3078,N_2903,N_2969);
or U3079 (N_3079,N_2914,N_2923);
nand U3080 (N_3080,N_2953,N_2951);
and U3081 (N_3081,N_2900,N_2967);
nand U3082 (N_3082,N_2912,N_2953);
xnor U3083 (N_3083,N_2980,N_2925);
xnor U3084 (N_3084,N_2909,N_2945);
nand U3085 (N_3085,N_2931,N_2961);
nor U3086 (N_3086,N_2904,N_2994);
nand U3087 (N_3087,N_2944,N_2981);
or U3088 (N_3088,N_2988,N_2958);
xor U3089 (N_3089,N_2933,N_2963);
or U3090 (N_3090,N_2906,N_2965);
nor U3091 (N_3091,N_2936,N_2924);
nand U3092 (N_3092,N_2932,N_2905);
nor U3093 (N_3093,N_2975,N_2987);
nand U3094 (N_3094,N_2956,N_2988);
nand U3095 (N_3095,N_2907,N_2977);
or U3096 (N_3096,N_2943,N_2906);
nand U3097 (N_3097,N_2932,N_2926);
and U3098 (N_3098,N_2998,N_2974);
nand U3099 (N_3099,N_2912,N_2917);
nor U3100 (N_3100,N_3065,N_3082);
nand U3101 (N_3101,N_3009,N_3042);
nand U3102 (N_3102,N_3030,N_3001);
nand U3103 (N_3103,N_3018,N_3043);
nand U3104 (N_3104,N_3036,N_3053);
and U3105 (N_3105,N_3067,N_3070);
nor U3106 (N_3106,N_3072,N_3081);
or U3107 (N_3107,N_3025,N_3013);
xor U3108 (N_3108,N_3061,N_3089);
nand U3109 (N_3109,N_3074,N_3052);
and U3110 (N_3110,N_3088,N_3083);
xnor U3111 (N_3111,N_3022,N_3050);
and U3112 (N_3112,N_3044,N_3020);
nand U3113 (N_3113,N_3079,N_3077);
nand U3114 (N_3114,N_3029,N_3031);
nand U3115 (N_3115,N_3023,N_3017);
nor U3116 (N_3116,N_3008,N_3028);
or U3117 (N_3117,N_3026,N_3024);
nand U3118 (N_3118,N_3096,N_3002);
xnor U3119 (N_3119,N_3095,N_3071);
xor U3120 (N_3120,N_3099,N_3038);
nand U3121 (N_3121,N_3098,N_3048);
nand U3122 (N_3122,N_3045,N_3078);
nor U3123 (N_3123,N_3085,N_3004);
or U3124 (N_3124,N_3019,N_3016);
nor U3125 (N_3125,N_3039,N_3040);
and U3126 (N_3126,N_3094,N_3051);
and U3127 (N_3127,N_3059,N_3092);
and U3128 (N_3128,N_3033,N_3027);
nand U3129 (N_3129,N_3069,N_3010);
xor U3130 (N_3130,N_3047,N_3063);
and U3131 (N_3131,N_3003,N_3037);
xnor U3132 (N_3132,N_3005,N_3090);
nor U3133 (N_3133,N_3014,N_3056);
xor U3134 (N_3134,N_3073,N_3093);
or U3135 (N_3135,N_3011,N_3087);
nor U3136 (N_3136,N_3076,N_3064);
or U3137 (N_3137,N_3097,N_3068);
nor U3138 (N_3138,N_3021,N_3006);
or U3139 (N_3139,N_3049,N_3046);
nand U3140 (N_3140,N_3086,N_3000);
nor U3141 (N_3141,N_3057,N_3041);
nor U3142 (N_3142,N_3012,N_3015);
xnor U3143 (N_3143,N_3055,N_3054);
or U3144 (N_3144,N_3066,N_3007);
xnor U3145 (N_3145,N_3062,N_3080);
nor U3146 (N_3146,N_3091,N_3084);
and U3147 (N_3147,N_3075,N_3058);
and U3148 (N_3148,N_3035,N_3060);
or U3149 (N_3149,N_3034,N_3032);
or U3150 (N_3150,N_3021,N_3061);
nand U3151 (N_3151,N_3045,N_3093);
nand U3152 (N_3152,N_3086,N_3095);
xor U3153 (N_3153,N_3087,N_3010);
xnor U3154 (N_3154,N_3025,N_3004);
nand U3155 (N_3155,N_3027,N_3073);
and U3156 (N_3156,N_3070,N_3022);
nor U3157 (N_3157,N_3051,N_3075);
xnor U3158 (N_3158,N_3003,N_3023);
or U3159 (N_3159,N_3050,N_3096);
nand U3160 (N_3160,N_3087,N_3013);
nand U3161 (N_3161,N_3059,N_3027);
and U3162 (N_3162,N_3095,N_3064);
xnor U3163 (N_3163,N_3058,N_3022);
or U3164 (N_3164,N_3084,N_3019);
xor U3165 (N_3165,N_3001,N_3062);
xnor U3166 (N_3166,N_3067,N_3082);
nor U3167 (N_3167,N_3073,N_3020);
nand U3168 (N_3168,N_3001,N_3012);
and U3169 (N_3169,N_3088,N_3036);
nor U3170 (N_3170,N_3016,N_3000);
xor U3171 (N_3171,N_3038,N_3031);
xor U3172 (N_3172,N_3054,N_3022);
and U3173 (N_3173,N_3000,N_3040);
xor U3174 (N_3174,N_3029,N_3003);
nand U3175 (N_3175,N_3018,N_3090);
or U3176 (N_3176,N_3001,N_3041);
or U3177 (N_3177,N_3060,N_3081);
xor U3178 (N_3178,N_3004,N_3068);
xnor U3179 (N_3179,N_3082,N_3010);
nor U3180 (N_3180,N_3015,N_3075);
nor U3181 (N_3181,N_3076,N_3060);
xnor U3182 (N_3182,N_3046,N_3050);
nand U3183 (N_3183,N_3082,N_3050);
xor U3184 (N_3184,N_3052,N_3043);
nand U3185 (N_3185,N_3039,N_3002);
and U3186 (N_3186,N_3061,N_3001);
and U3187 (N_3187,N_3089,N_3001);
and U3188 (N_3188,N_3050,N_3064);
and U3189 (N_3189,N_3064,N_3019);
and U3190 (N_3190,N_3043,N_3086);
or U3191 (N_3191,N_3060,N_3017);
or U3192 (N_3192,N_3060,N_3091);
nor U3193 (N_3193,N_3001,N_3085);
and U3194 (N_3194,N_3038,N_3026);
nor U3195 (N_3195,N_3078,N_3096);
and U3196 (N_3196,N_3068,N_3053);
xnor U3197 (N_3197,N_3035,N_3075);
and U3198 (N_3198,N_3029,N_3097);
nor U3199 (N_3199,N_3092,N_3001);
nand U3200 (N_3200,N_3137,N_3197);
or U3201 (N_3201,N_3149,N_3143);
and U3202 (N_3202,N_3180,N_3103);
or U3203 (N_3203,N_3161,N_3100);
nand U3204 (N_3204,N_3151,N_3112);
or U3205 (N_3205,N_3158,N_3111);
nor U3206 (N_3206,N_3101,N_3173);
xor U3207 (N_3207,N_3171,N_3157);
and U3208 (N_3208,N_3136,N_3133);
or U3209 (N_3209,N_3167,N_3123);
nor U3210 (N_3210,N_3169,N_3144);
xnor U3211 (N_3211,N_3147,N_3138);
xor U3212 (N_3212,N_3119,N_3162);
nor U3213 (N_3213,N_3128,N_3126);
nand U3214 (N_3214,N_3193,N_3125);
or U3215 (N_3215,N_3145,N_3155);
or U3216 (N_3216,N_3189,N_3175);
nand U3217 (N_3217,N_3131,N_3122);
nand U3218 (N_3218,N_3134,N_3176);
xnor U3219 (N_3219,N_3168,N_3114);
nor U3220 (N_3220,N_3130,N_3104);
xnor U3221 (N_3221,N_3115,N_3184);
nand U3222 (N_3222,N_3153,N_3170);
or U3223 (N_3223,N_3198,N_3113);
nand U3224 (N_3224,N_3199,N_3163);
and U3225 (N_3225,N_3183,N_3118);
nor U3226 (N_3226,N_3117,N_3186);
xnor U3227 (N_3227,N_3106,N_3146);
nor U3228 (N_3228,N_3172,N_3124);
and U3229 (N_3229,N_3188,N_3174);
and U3230 (N_3230,N_3105,N_3152);
and U3231 (N_3231,N_3121,N_3177);
and U3232 (N_3232,N_3142,N_3107);
xnor U3233 (N_3233,N_3194,N_3102);
or U3234 (N_3234,N_3190,N_3110);
and U3235 (N_3235,N_3148,N_3196);
or U3236 (N_3236,N_3140,N_3109);
xor U3237 (N_3237,N_3178,N_3141);
nor U3238 (N_3238,N_3120,N_3129);
and U3239 (N_3239,N_3185,N_3154);
or U3240 (N_3240,N_3159,N_3187);
nand U3241 (N_3241,N_3192,N_3164);
xor U3242 (N_3242,N_3127,N_3182);
xnor U3243 (N_3243,N_3139,N_3132);
or U3244 (N_3244,N_3160,N_3165);
and U3245 (N_3245,N_3156,N_3166);
xor U3246 (N_3246,N_3181,N_3191);
xor U3247 (N_3247,N_3150,N_3195);
xor U3248 (N_3248,N_3108,N_3116);
and U3249 (N_3249,N_3135,N_3179);
or U3250 (N_3250,N_3164,N_3101);
nor U3251 (N_3251,N_3188,N_3190);
xor U3252 (N_3252,N_3141,N_3121);
nand U3253 (N_3253,N_3199,N_3162);
or U3254 (N_3254,N_3165,N_3116);
or U3255 (N_3255,N_3164,N_3107);
and U3256 (N_3256,N_3157,N_3116);
and U3257 (N_3257,N_3138,N_3134);
xnor U3258 (N_3258,N_3158,N_3183);
xnor U3259 (N_3259,N_3184,N_3125);
or U3260 (N_3260,N_3110,N_3148);
nor U3261 (N_3261,N_3174,N_3164);
nand U3262 (N_3262,N_3117,N_3197);
or U3263 (N_3263,N_3185,N_3131);
or U3264 (N_3264,N_3196,N_3185);
and U3265 (N_3265,N_3184,N_3119);
or U3266 (N_3266,N_3154,N_3101);
xor U3267 (N_3267,N_3146,N_3126);
xnor U3268 (N_3268,N_3130,N_3176);
xnor U3269 (N_3269,N_3175,N_3124);
xor U3270 (N_3270,N_3114,N_3175);
and U3271 (N_3271,N_3183,N_3132);
or U3272 (N_3272,N_3178,N_3155);
xnor U3273 (N_3273,N_3190,N_3102);
nand U3274 (N_3274,N_3117,N_3122);
xor U3275 (N_3275,N_3150,N_3173);
and U3276 (N_3276,N_3142,N_3119);
or U3277 (N_3277,N_3194,N_3177);
nor U3278 (N_3278,N_3163,N_3172);
nor U3279 (N_3279,N_3185,N_3109);
and U3280 (N_3280,N_3138,N_3124);
nand U3281 (N_3281,N_3166,N_3147);
nor U3282 (N_3282,N_3104,N_3174);
xnor U3283 (N_3283,N_3144,N_3153);
xor U3284 (N_3284,N_3119,N_3156);
nand U3285 (N_3285,N_3131,N_3105);
and U3286 (N_3286,N_3109,N_3102);
nand U3287 (N_3287,N_3195,N_3172);
or U3288 (N_3288,N_3147,N_3111);
nor U3289 (N_3289,N_3134,N_3104);
nand U3290 (N_3290,N_3196,N_3125);
or U3291 (N_3291,N_3183,N_3126);
nand U3292 (N_3292,N_3149,N_3158);
and U3293 (N_3293,N_3155,N_3180);
xor U3294 (N_3294,N_3152,N_3137);
xnor U3295 (N_3295,N_3137,N_3130);
or U3296 (N_3296,N_3107,N_3118);
nand U3297 (N_3297,N_3169,N_3142);
nor U3298 (N_3298,N_3159,N_3100);
xor U3299 (N_3299,N_3133,N_3159);
nand U3300 (N_3300,N_3230,N_3298);
nand U3301 (N_3301,N_3225,N_3299);
nand U3302 (N_3302,N_3264,N_3255);
xnor U3303 (N_3303,N_3290,N_3281);
or U3304 (N_3304,N_3291,N_3235);
nand U3305 (N_3305,N_3215,N_3260);
and U3306 (N_3306,N_3295,N_3293);
xor U3307 (N_3307,N_3214,N_3251);
nand U3308 (N_3308,N_3268,N_3237);
and U3309 (N_3309,N_3284,N_3252);
nand U3310 (N_3310,N_3204,N_3242);
xnor U3311 (N_3311,N_3211,N_3283);
or U3312 (N_3312,N_3285,N_3223);
nor U3313 (N_3313,N_3269,N_3253);
or U3314 (N_3314,N_3238,N_3256);
and U3315 (N_3315,N_3288,N_3226);
xnor U3316 (N_3316,N_3279,N_3239);
or U3317 (N_3317,N_3267,N_3259);
nand U3318 (N_3318,N_3263,N_3286);
nor U3319 (N_3319,N_3202,N_3292);
and U3320 (N_3320,N_3207,N_3247);
or U3321 (N_3321,N_3212,N_3206);
and U3322 (N_3322,N_3219,N_3200);
and U3323 (N_3323,N_3233,N_3278);
nor U3324 (N_3324,N_3276,N_3289);
nor U3325 (N_3325,N_3217,N_3201);
nand U3326 (N_3326,N_3209,N_3266);
and U3327 (N_3327,N_3272,N_3287);
nor U3328 (N_3328,N_3224,N_3216);
nand U3329 (N_3329,N_3218,N_3265);
nand U3330 (N_3330,N_3250,N_3243);
nand U3331 (N_3331,N_3221,N_3249);
nor U3332 (N_3332,N_3274,N_3270);
or U3333 (N_3333,N_3220,N_3245);
xor U3334 (N_3334,N_3228,N_3222);
nand U3335 (N_3335,N_3257,N_3261);
nor U3336 (N_3336,N_3203,N_3277);
nor U3337 (N_3337,N_3232,N_3254);
nand U3338 (N_3338,N_3244,N_3297);
and U3339 (N_3339,N_3296,N_3231);
and U3340 (N_3340,N_3246,N_3210);
or U3341 (N_3341,N_3258,N_3227);
nor U3342 (N_3342,N_3241,N_3248);
nand U3343 (N_3343,N_3229,N_3273);
nor U3344 (N_3344,N_3282,N_3271);
nand U3345 (N_3345,N_3294,N_3213);
xnor U3346 (N_3346,N_3275,N_3262);
or U3347 (N_3347,N_3240,N_3205);
and U3348 (N_3348,N_3236,N_3234);
or U3349 (N_3349,N_3208,N_3280);
or U3350 (N_3350,N_3213,N_3203);
nand U3351 (N_3351,N_3227,N_3213);
and U3352 (N_3352,N_3266,N_3263);
or U3353 (N_3353,N_3216,N_3282);
nand U3354 (N_3354,N_3227,N_3295);
xor U3355 (N_3355,N_3269,N_3240);
nor U3356 (N_3356,N_3247,N_3291);
and U3357 (N_3357,N_3243,N_3223);
nand U3358 (N_3358,N_3286,N_3236);
xnor U3359 (N_3359,N_3218,N_3270);
xnor U3360 (N_3360,N_3209,N_3225);
and U3361 (N_3361,N_3293,N_3234);
and U3362 (N_3362,N_3234,N_3226);
nor U3363 (N_3363,N_3255,N_3299);
and U3364 (N_3364,N_3267,N_3262);
xnor U3365 (N_3365,N_3208,N_3298);
or U3366 (N_3366,N_3206,N_3294);
xnor U3367 (N_3367,N_3205,N_3291);
xor U3368 (N_3368,N_3295,N_3253);
xor U3369 (N_3369,N_3237,N_3272);
nand U3370 (N_3370,N_3216,N_3271);
or U3371 (N_3371,N_3287,N_3286);
nor U3372 (N_3372,N_3232,N_3217);
and U3373 (N_3373,N_3203,N_3274);
nand U3374 (N_3374,N_3209,N_3220);
and U3375 (N_3375,N_3206,N_3284);
xnor U3376 (N_3376,N_3212,N_3290);
or U3377 (N_3377,N_3277,N_3245);
nor U3378 (N_3378,N_3292,N_3279);
nand U3379 (N_3379,N_3288,N_3204);
and U3380 (N_3380,N_3205,N_3208);
nand U3381 (N_3381,N_3201,N_3206);
nor U3382 (N_3382,N_3287,N_3274);
nor U3383 (N_3383,N_3200,N_3233);
or U3384 (N_3384,N_3204,N_3211);
xor U3385 (N_3385,N_3224,N_3211);
or U3386 (N_3386,N_3213,N_3289);
and U3387 (N_3387,N_3260,N_3220);
nor U3388 (N_3388,N_3296,N_3230);
nor U3389 (N_3389,N_3228,N_3296);
nand U3390 (N_3390,N_3200,N_3282);
nand U3391 (N_3391,N_3242,N_3286);
xor U3392 (N_3392,N_3251,N_3289);
nand U3393 (N_3393,N_3237,N_3215);
xnor U3394 (N_3394,N_3225,N_3269);
nor U3395 (N_3395,N_3208,N_3236);
or U3396 (N_3396,N_3242,N_3292);
and U3397 (N_3397,N_3295,N_3215);
nor U3398 (N_3398,N_3299,N_3221);
and U3399 (N_3399,N_3214,N_3241);
nand U3400 (N_3400,N_3330,N_3386);
and U3401 (N_3401,N_3334,N_3357);
nor U3402 (N_3402,N_3333,N_3303);
and U3403 (N_3403,N_3396,N_3364);
nand U3404 (N_3404,N_3382,N_3374);
nor U3405 (N_3405,N_3392,N_3324);
and U3406 (N_3406,N_3359,N_3341);
xor U3407 (N_3407,N_3320,N_3337);
xnor U3408 (N_3408,N_3376,N_3358);
xnor U3409 (N_3409,N_3328,N_3375);
nand U3410 (N_3410,N_3347,N_3371);
or U3411 (N_3411,N_3389,N_3356);
or U3412 (N_3412,N_3352,N_3323);
or U3413 (N_3413,N_3302,N_3349);
nor U3414 (N_3414,N_3312,N_3350);
nor U3415 (N_3415,N_3351,N_3390);
xnor U3416 (N_3416,N_3327,N_3354);
or U3417 (N_3417,N_3316,N_3339);
nand U3418 (N_3418,N_3306,N_3398);
nor U3419 (N_3419,N_3366,N_3345);
nand U3420 (N_3420,N_3311,N_3301);
xor U3421 (N_3421,N_3326,N_3372);
and U3422 (N_3422,N_3377,N_3304);
nor U3423 (N_3423,N_3365,N_3336);
xnor U3424 (N_3424,N_3368,N_3380);
xnor U3425 (N_3425,N_3305,N_3370);
and U3426 (N_3426,N_3342,N_3313);
or U3427 (N_3427,N_3344,N_3310);
xor U3428 (N_3428,N_3321,N_3322);
nand U3429 (N_3429,N_3395,N_3329);
nor U3430 (N_3430,N_3369,N_3373);
or U3431 (N_3431,N_3314,N_3397);
nand U3432 (N_3432,N_3361,N_3387);
nand U3433 (N_3433,N_3391,N_3383);
xor U3434 (N_3434,N_3363,N_3378);
nor U3435 (N_3435,N_3381,N_3394);
and U3436 (N_3436,N_3319,N_3353);
nand U3437 (N_3437,N_3399,N_3393);
nor U3438 (N_3438,N_3332,N_3308);
xor U3439 (N_3439,N_3385,N_3360);
nor U3440 (N_3440,N_3340,N_3346);
nand U3441 (N_3441,N_3300,N_3309);
or U3442 (N_3442,N_3317,N_3331);
xor U3443 (N_3443,N_3343,N_3325);
nor U3444 (N_3444,N_3355,N_3307);
xnor U3445 (N_3445,N_3379,N_3362);
or U3446 (N_3446,N_3388,N_3348);
or U3447 (N_3447,N_3367,N_3318);
and U3448 (N_3448,N_3384,N_3335);
nor U3449 (N_3449,N_3315,N_3338);
nand U3450 (N_3450,N_3342,N_3316);
xnor U3451 (N_3451,N_3362,N_3325);
or U3452 (N_3452,N_3317,N_3332);
xor U3453 (N_3453,N_3365,N_3398);
nand U3454 (N_3454,N_3309,N_3331);
or U3455 (N_3455,N_3327,N_3385);
xnor U3456 (N_3456,N_3343,N_3387);
nor U3457 (N_3457,N_3388,N_3310);
or U3458 (N_3458,N_3325,N_3373);
and U3459 (N_3459,N_3388,N_3342);
or U3460 (N_3460,N_3361,N_3317);
nand U3461 (N_3461,N_3385,N_3356);
and U3462 (N_3462,N_3344,N_3341);
or U3463 (N_3463,N_3308,N_3334);
and U3464 (N_3464,N_3323,N_3333);
or U3465 (N_3465,N_3343,N_3327);
or U3466 (N_3466,N_3325,N_3317);
or U3467 (N_3467,N_3394,N_3325);
xnor U3468 (N_3468,N_3333,N_3345);
or U3469 (N_3469,N_3318,N_3380);
nand U3470 (N_3470,N_3375,N_3303);
xnor U3471 (N_3471,N_3311,N_3331);
and U3472 (N_3472,N_3306,N_3367);
nand U3473 (N_3473,N_3347,N_3325);
or U3474 (N_3474,N_3347,N_3329);
or U3475 (N_3475,N_3318,N_3362);
nand U3476 (N_3476,N_3350,N_3341);
nor U3477 (N_3477,N_3380,N_3335);
nor U3478 (N_3478,N_3354,N_3332);
nor U3479 (N_3479,N_3373,N_3389);
xnor U3480 (N_3480,N_3396,N_3302);
and U3481 (N_3481,N_3355,N_3328);
nor U3482 (N_3482,N_3350,N_3337);
or U3483 (N_3483,N_3334,N_3375);
nand U3484 (N_3484,N_3300,N_3369);
nor U3485 (N_3485,N_3391,N_3354);
or U3486 (N_3486,N_3346,N_3399);
and U3487 (N_3487,N_3359,N_3363);
nand U3488 (N_3488,N_3393,N_3334);
or U3489 (N_3489,N_3357,N_3315);
nand U3490 (N_3490,N_3317,N_3375);
xnor U3491 (N_3491,N_3301,N_3318);
nor U3492 (N_3492,N_3367,N_3356);
nand U3493 (N_3493,N_3304,N_3352);
and U3494 (N_3494,N_3361,N_3357);
and U3495 (N_3495,N_3379,N_3380);
or U3496 (N_3496,N_3324,N_3318);
or U3497 (N_3497,N_3333,N_3327);
or U3498 (N_3498,N_3324,N_3379);
nand U3499 (N_3499,N_3328,N_3357);
xor U3500 (N_3500,N_3429,N_3451);
xnor U3501 (N_3501,N_3498,N_3484);
xor U3502 (N_3502,N_3448,N_3415);
or U3503 (N_3503,N_3432,N_3417);
nor U3504 (N_3504,N_3406,N_3475);
nand U3505 (N_3505,N_3485,N_3420);
xor U3506 (N_3506,N_3492,N_3468);
and U3507 (N_3507,N_3489,N_3499);
or U3508 (N_3508,N_3445,N_3443);
nor U3509 (N_3509,N_3472,N_3491);
nor U3510 (N_3510,N_3488,N_3423);
nor U3511 (N_3511,N_3438,N_3437);
xor U3512 (N_3512,N_3404,N_3441);
nor U3513 (N_3513,N_3407,N_3431);
xor U3514 (N_3514,N_3455,N_3410);
and U3515 (N_3515,N_3464,N_3467);
nor U3516 (N_3516,N_3466,N_3402);
nor U3517 (N_3517,N_3456,N_3458);
or U3518 (N_3518,N_3401,N_3444);
or U3519 (N_3519,N_3494,N_3446);
and U3520 (N_3520,N_3453,N_3465);
nor U3521 (N_3521,N_3421,N_3478);
and U3522 (N_3522,N_3418,N_3436);
or U3523 (N_3523,N_3425,N_3426);
nor U3524 (N_3524,N_3493,N_3408);
and U3525 (N_3525,N_3440,N_3481);
xor U3526 (N_3526,N_3403,N_3479);
xnor U3527 (N_3527,N_3434,N_3480);
nor U3528 (N_3528,N_3477,N_3461);
or U3529 (N_3529,N_3433,N_3496);
and U3530 (N_3530,N_3497,N_3439);
xor U3531 (N_3531,N_3411,N_3473);
nor U3532 (N_3532,N_3405,N_3449);
or U3533 (N_3533,N_3428,N_3412);
nor U3534 (N_3534,N_3462,N_3424);
and U3535 (N_3535,N_3454,N_3495);
xnor U3536 (N_3536,N_3416,N_3486);
xnor U3537 (N_3537,N_3450,N_3419);
nor U3538 (N_3538,N_3470,N_3471);
or U3539 (N_3539,N_3447,N_3427);
or U3540 (N_3540,N_3435,N_3460);
nand U3541 (N_3541,N_3463,N_3414);
nand U3542 (N_3542,N_3409,N_3487);
and U3543 (N_3543,N_3483,N_3442);
and U3544 (N_3544,N_3422,N_3482);
nand U3545 (N_3545,N_3490,N_3413);
and U3546 (N_3546,N_3430,N_3452);
xor U3547 (N_3547,N_3400,N_3474);
xnor U3548 (N_3548,N_3469,N_3459);
xor U3549 (N_3549,N_3457,N_3476);
and U3550 (N_3550,N_3405,N_3438);
or U3551 (N_3551,N_3435,N_3452);
xor U3552 (N_3552,N_3476,N_3499);
nand U3553 (N_3553,N_3469,N_3412);
or U3554 (N_3554,N_3434,N_3497);
and U3555 (N_3555,N_3443,N_3408);
nor U3556 (N_3556,N_3431,N_3495);
and U3557 (N_3557,N_3436,N_3476);
xor U3558 (N_3558,N_3440,N_3435);
or U3559 (N_3559,N_3447,N_3441);
nor U3560 (N_3560,N_3465,N_3489);
and U3561 (N_3561,N_3479,N_3415);
and U3562 (N_3562,N_3475,N_3405);
xor U3563 (N_3563,N_3401,N_3416);
or U3564 (N_3564,N_3479,N_3429);
nor U3565 (N_3565,N_3441,N_3476);
and U3566 (N_3566,N_3436,N_3428);
nor U3567 (N_3567,N_3431,N_3468);
xor U3568 (N_3568,N_3448,N_3437);
nand U3569 (N_3569,N_3421,N_3487);
nand U3570 (N_3570,N_3423,N_3412);
and U3571 (N_3571,N_3461,N_3407);
nand U3572 (N_3572,N_3494,N_3435);
nor U3573 (N_3573,N_3450,N_3402);
xnor U3574 (N_3574,N_3444,N_3464);
or U3575 (N_3575,N_3424,N_3415);
xor U3576 (N_3576,N_3427,N_3438);
xor U3577 (N_3577,N_3457,N_3462);
nand U3578 (N_3578,N_3463,N_3420);
nor U3579 (N_3579,N_3426,N_3401);
or U3580 (N_3580,N_3441,N_3471);
xor U3581 (N_3581,N_3459,N_3433);
or U3582 (N_3582,N_3455,N_3467);
xor U3583 (N_3583,N_3473,N_3433);
xor U3584 (N_3584,N_3488,N_3469);
nand U3585 (N_3585,N_3431,N_3442);
or U3586 (N_3586,N_3401,N_3480);
or U3587 (N_3587,N_3425,N_3450);
xnor U3588 (N_3588,N_3422,N_3492);
or U3589 (N_3589,N_3437,N_3427);
nand U3590 (N_3590,N_3469,N_3466);
or U3591 (N_3591,N_3443,N_3436);
nor U3592 (N_3592,N_3422,N_3426);
nand U3593 (N_3593,N_3414,N_3430);
nor U3594 (N_3594,N_3427,N_3485);
nand U3595 (N_3595,N_3490,N_3477);
nand U3596 (N_3596,N_3446,N_3402);
or U3597 (N_3597,N_3490,N_3495);
nand U3598 (N_3598,N_3452,N_3413);
nor U3599 (N_3599,N_3427,N_3461);
nand U3600 (N_3600,N_3528,N_3565);
or U3601 (N_3601,N_3552,N_3531);
or U3602 (N_3602,N_3569,N_3574);
nor U3603 (N_3603,N_3564,N_3516);
xnor U3604 (N_3604,N_3581,N_3521);
nor U3605 (N_3605,N_3535,N_3591);
or U3606 (N_3606,N_3539,N_3553);
xnor U3607 (N_3607,N_3536,N_3573);
and U3608 (N_3608,N_3505,N_3504);
nand U3609 (N_3609,N_3517,N_3586);
nand U3610 (N_3610,N_3550,N_3538);
or U3611 (N_3611,N_3596,N_3582);
nor U3612 (N_3612,N_3597,N_3551);
nor U3613 (N_3613,N_3558,N_3583);
nand U3614 (N_3614,N_3560,N_3509);
and U3615 (N_3615,N_3562,N_3549);
nor U3616 (N_3616,N_3594,N_3587);
and U3617 (N_3617,N_3554,N_3593);
and U3618 (N_3618,N_3592,N_3527);
nand U3619 (N_3619,N_3559,N_3530);
nor U3620 (N_3620,N_3557,N_3501);
or U3621 (N_3621,N_3544,N_3567);
or U3622 (N_3622,N_3580,N_3506);
nor U3623 (N_3623,N_3570,N_3510);
xor U3624 (N_3624,N_3598,N_3540);
and U3625 (N_3625,N_3519,N_3532);
nand U3626 (N_3626,N_3500,N_3534);
nor U3627 (N_3627,N_3575,N_3595);
nand U3628 (N_3628,N_3590,N_3503);
nor U3629 (N_3629,N_3518,N_3561);
and U3630 (N_3630,N_3589,N_3576);
xnor U3631 (N_3631,N_3599,N_3547);
nor U3632 (N_3632,N_3556,N_3523);
nand U3633 (N_3633,N_3502,N_3515);
xor U3634 (N_3634,N_3513,N_3514);
nor U3635 (N_3635,N_3545,N_3568);
xor U3636 (N_3636,N_3542,N_3511);
nand U3637 (N_3637,N_3585,N_3522);
nand U3638 (N_3638,N_3512,N_3537);
or U3639 (N_3639,N_3543,N_3584);
nand U3640 (N_3640,N_3529,N_3525);
nor U3641 (N_3641,N_3526,N_3578);
or U3642 (N_3642,N_3579,N_3588);
xnor U3643 (N_3643,N_3563,N_3508);
xor U3644 (N_3644,N_3533,N_3524);
or U3645 (N_3645,N_3520,N_3507);
and U3646 (N_3646,N_3541,N_3546);
or U3647 (N_3647,N_3572,N_3548);
nor U3648 (N_3648,N_3577,N_3571);
or U3649 (N_3649,N_3566,N_3555);
and U3650 (N_3650,N_3554,N_3589);
or U3651 (N_3651,N_3540,N_3559);
or U3652 (N_3652,N_3560,N_3541);
nand U3653 (N_3653,N_3528,N_3503);
or U3654 (N_3654,N_3567,N_3506);
nand U3655 (N_3655,N_3510,N_3525);
nand U3656 (N_3656,N_3578,N_3544);
nand U3657 (N_3657,N_3597,N_3510);
or U3658 (N_3658,N_3540,N_3546);
nor U3659 (N_3659,N_3580,N_3579);
or U3660 (N_3660,N_3558,N_3550);
nor U3661 (N_3661,N_3526,N_3558);
nand U3662 (N_3662,N_3516,N_3560);
or U3663 (N_3663,N_3546,N_3538);
and U3664 (N_3664,N_3581,N_3554);
xor U3665 (N_3665,N_3550,N_3525);
nor U3666 (N_3666,N_3568,N_3567);
nand U3667 (N_3667,N_3572,N_3589);
and U3668 (N_3668,N_3532,N_3583);
and U3669 (N_3669,N_3513,N_3527);
nand U3670 (N_3670,N_3547,N_3511);
and U3671 (N_3671,N_3513,N_3502);
and U3672 (N_3672,N_3590,N_3538);
and U3673 (N_3673,N_3562,N_3524);
xor U3674 (N_3674,N_3575,N_3596);
xor U3675 (N_3675,N_3575,N_3592);
xnor U3676 (N_3676,N_3523,N_3572);
and U3677 (N_3677,N_3558,N_3591);
nand U3678 (N_3678,N_3575,N_3507);
or U3679 (N_3679,N_3501,N_3526);
nor U3680 (N_3680,N_3536,N_3583);
nand U3681 (N_3681,N_3529,N_3574);
and U3682 (N_3682,N_3596,N_3564);
nand U3683 (N_3683,N_3519,N_3521);
and U3684 (N_3684,N_3514,N_3560);
xor U3685 (N_3685,N_3521,N_3536);
and U3686 (N_3686,N_3542,N_3504);
nor U3687 (N_3687,N_3565,N_3550);
nor U3688 (N_3688,N_3516,N_3517);
nand U3689 (N_3689,N_3545,N_3509);
nand U3690 (N_3690,N_3532,N_3561);
nand U3691 (N_3691,N_3557,N_3515);
nand U3692 (N_3692,N_3515,N_3517);
xor U3693 (N_3693,N_3569,N_3544);
nor U3694 (N_3694,N_3510,N_3500);
nor U3695 (N_3695,N_3596,N_3595);
or U3696 (N_3696,N_3559,N_3511);
xor U3697 (N_3697,N_3516,N_3545);
or U3698 (N_3698,N_3532,N_3511);
nand U3699 (N_3699,N_3518,N_3568);
xnor U3700 (N_3700,N_3608,N_3627);
xnor U3701 (N_3701,N_3683,N_3606);
xnor U3702 (N_3702,N_3670,N_3685);
xor U3703 (N_3703,N_3651,N_3605);
or U3704 (N_3704,N_3629,N_3632);
nor U3705 (N_3705,N_3604,N_3690);
xnor U3706 (N_3706,N_3652,N_3655);
nor U3707 (N_3707,N_3675,N_3637);
or U3708 (N_3708,N_3650,N_3626);
and U3709 (N_3709,N_3669,N_3676);
nand U3710 (N_3710,N_3648,N_3672);
or U3711 (N_3711,N_3684,N_3644);
nor U3712 (N_3712,N_3601,N_3628);
or U3713 (N_3713,N_3633,N_3622);
or U3714 (N_3714,N_3697,N_3642);
xor U3715 (N_3715,N_3658,N_3619);
nor U3716 (N_3716,N_3656,N_3673);
nand U3717 (N_3717,N_3649,N_3682);
and U3718 (N_3718,N_3691,N_3692);
or U3719 (N_3719,N_3698,N_3688);
xnor U3720 (N_3720,N_3695,N_3674);
or U3721 (N_3721,N_3624,N_3666);
xor U3722 (N_3722,N_3640,N_3699);
or U3723 (N_3723,N_3641,N_3636);
and U3724 (N_3724,N_3661,N_3689);
and U3725 (N_3725,N_3610,N_3639);
and U3726 (N_3726,N_3653,N_3603);
or U3727 (N_3727,N_3694,N_3662);
or U3728 (N_3728,N_3686,N_3679);
nand U3729 (N_3729,N_3635,N_3677);
xor U3730 (N_3730,N_3617,N_3668);
nand U3731 (N_3731,N_3638,N_3611);
nor U3732 (N_3732,N_3693,N_3600);
or U3733 (N_3733,N_3621,N_3687);
nand U3734 (N_3734,N_3634,N_3671);
nor U3735 (N_3735,N_3657,N_3607);
xor U3736 (N_3736,N_3609,N_3667);
xor U3737 (N_3737,N_3659,N_3623);
and U3738 (N_3738,N_3620,N_3696);
and U3739 (N_3739,N_3643,N_3660);
nor U3740 (N_3740,N_3647,N_3663);
or U3741 (N_3741,N_3680,N_3616);
or U3742 (N_3742,N_3645,N_3630);
nand U3743 (N_3743,N_3614,N_3665);
nand U3744 (N_3744,N_3613,N_3625);
nand U3745 (N_3745,N_3631,N_3602);
nand U3746 (N_3746,N_3615,N_3654);
nand U3747 (N_3747,N_3681,N_3678);
nor U3748 (N_3748,N_3646,N_3612);
nand U3749 (N_3749,N_3618,N_3664);
and U3750 (N_3750,N_3602,N_3660);
xor U3751 (N_3751,N_3625,N_3614);
or U3752 (N_3752,N_3680,N_3686);
nor U3753 (N_3753,N_3618,N_3627);
nand U3754 (N_3754,N_3655,N_3657);
or U3755 (N_3755,N_3659,N_3693);
nor U3756 (N_3756,N_3640,N_3610);
or U3757 (N_3757,N_3636,N_3639);
xor U3758 (N_3758,N_3635,N_3687);
nand U3759 (N_3759,N_3654,N_3674);
nand U3760 (N_3760,N_3691,N_3633);
xnor U3761 (N_3761,N_3629,N_3655);
nand U3762 (N_3762,N_3651,N_3635);
nand U3763 (N_3763,N_3621,N_3620);
and U3764 (N_3764,N_3694,N_3626);
and U3765 (N_3765,N_3606,N_3684);
xnor U3766 (N_3766,N_3688,N_3600);
and U3767 (N_3767,N_3668,N_3657);
nor U3768 (N_3768,N_3612,N_3614);
and U3769 (N_3769,N_3629,N_3662);
xnor U3770 (N_3770,N_3669,N_3681);
or U3771 (N_3771,N_3623,N_3666);
and U3772 (N_3772,N_3618,N_3657);
nand U3773 (N_3773,N_3629,N_3650);
and U3774 (N_3774,N_3635,N_3605);
nor U3775 (N_3775,N_3688,N_3604);
or U3776 (N_3776,N_3604,N_3682);
nand U3777 (N_3777,N_3622,N_3656);
nand U3778 (N_3778,N_3664,N_3683);
xnor U3779 (N_3779,N_3627,N_3649);
nand U3780 (N_3780,N_3601,N_3697);
or U3781 (N_3781,N_3652,N_3641);
or U3782 (N_3782,N_3685,N_3668);
xor U3783 (N_3783,N_3687,N_3645);
and U3784 (N_3784,N_3682,N_3644);
xor U3785 (N_3785,N_3656,N_3613);
or U3786 (N_3786,N_3644,N_3641);
and U3787 (N_3787,N_3686,N_3671);
xor U3788 (N_3788,N_3642,N_3690);
and U3789 (N_3789,N_3623,N_3633);
nor U3790 (N_3790,N_3656,N_3675);
xor U3791 (N_3791,N_3656,N_3615);
and U3792 (N_3792,N_3637,N_3634);
nand U3793 (N_3793,N_3697,N_3668);
xor U3794 (N_3794,N_3634,N_3600);
xor U3795 (N_3795,N_3680,N_3671);
xnor U3796 (N_3796,N_3631,N_3680);
xnor U3797 (N_3797,N_3629,N_3694);
nand U3798 (N_3798,N_3604,N_3696);
xnor U3799 (N_3799,N_3658,N_3692);
xnor U3800 (N_3800,N_3786,N_3706);
xnor U3801 (N_3801,N_3721,N_3785);
xnor U3802 (N_3802,N_3799,N_3766);
and U3803 (N_3803,N_3711,N_3737);
or U3804 (N_3804,N_3704,N_3740);
or U3805 (N_3805,N_3769,N_3746);
xnor U3806 (N_3806,N_3713,N_3738);
or U3807 (N_3807,N_3797,N_3759);
nand U3808 (N_3808,N_3747,N_3709);
xnor U3809 (N_3809,N_3772,N_3753);
xor U3810 (N_3810,N_3700,N_3761);
nor U3811 (N_3811,N_3791,N_3798);
or U3812 (N_3812,N_3776,N_3731);
and U3813 (N_3813,N_3767,N_3758);
nand U3814 (N_3814,N_3773,N_3796);
and U3815 (N_3815,N_3775,N_3716);
or U3816 (N_3816,N_3779,N_3730);
and U3817 (N_3817,N_3778,N_3725);
or U3818 (N_3818,N_3715,N_3762);
nand U3819 (N_3819,N_3754,N_3735);
xor U3820 (N_3820,N_3750,N_3752);
or U3821 (N_3821,N_3749,N_3717);
xor U3822 (N_3822,N_3719,N_3783);
and U3823 (N_3823,N_3736,N_3720);
or U3824 (N_3824,N_3793,N_3792);
nand U3825 (N_3825,N_3718,N_3770);
and U3826 (N_3826,N_3787,N_3765);
xnor U3827 (N_3827,N_3794,N_3756);
and U3828 (N_3828,N_3777,N_3714);
and U3829 (N_3829,N_3760,N_3705);
and U3830 (N_3830,N_3724,N_3733);
nor U3831 (N_3831,N_3745,N_3729);
and U3832 (N_3832,N_3708,N_3795);
nand U3833 (N_3833,N_3774,N_3751);
nor U3834 (N_3834,N_3781,N_3790);
or U3835 (N_3835,N_3743,N_3739);
and U3836 (N_3836,N_3771,N_3726);
xnor U3837 (N_3837,N_3757,N_3722);
or U3838 (N_3838,N_3780,N_3734);
nor U3839 (N_3839,N_3784,N_3727);
or U3840 (N_3840,N_3732,N_3728);
nor U3841 (N_3841,N_3764,N_3744);
nand U3842 (N_3842,N_3782,N_3763);
nand U3843 (N_3843,N_3748,N_3789);
and U3844 (N_3844,N_3707,N_3742);
or U3845 (N_3845,N_3768,N_3788);
xnor U3846 (N_3846,N_3741,N_3701);
xor U3847 (N_3847,N_3703,N_3710);
xor U3848 (N_3848,N_3712,N_3723);
xnor U3849 (N_3849,N_3702,N_3755);
xor U3850 (N_3850,N_3778,N_3769);
nand U3851 (N_3851,N_3742,N_3798);
or U3852 (N_3852,N_3764,N_3785);
nand U3853 (N_3853,N_3702,N_3799);
xor U3854 (N_3854,N_3767,N_3784);
and U3855 (N_3855,N_3747,N_3789);
xnor U3856 (N_3856,N_3725,N_3712);
or U3857 (N_3857,N_3755,N_3745);
and U3858 (N_3858,N_3739,N_3791);
xor U3859 (N_3859,N_3765,N_3726);
xor U3860 (N_3860,N_3764,N_3704);
nor U3861 (N_3861,N_3745,N_3790);
nand U3862 (N_3862,N_3778,N_3753);
nand U3863 (N_3863,N_3761,N_3727);
and U3864 (N_3864,N_3755,N_3727);
nor U3865 (N_3865,N_3741,N_3747);
xor U3866 (N_3866,N_3737,N_3796);
xor U3867 (N_3867,N_3758,N_3794);
or U3868 (N_3868,N_3722,N_3734);
xor U3869 (N_3869,N_3748,N_3702);
xnor U3870 (N_3870,N_3732,N_3747);
xnor U3871 (N_3871,N_3734,N_3796);
xnor U3872 (N_3872,N_3745,N_3789);
nand U3873 (N_3873,N_3724,N_3775);
nor U3874 (N_3874,N_3747,N_3752);
xor U3875 (N_3875,N_3715,N_3707);
xnor U3876 (N_3876,N_3763,N_3770);
nand U3877 (N_3877,N_3779,N_3747);
or U3878 (N_3878,N_3723,N_3732);
xnor U3879 (N_3879,N_3749,N_3757);
nor U3880 (N_3880,N_3799,N_3747);
nand U3881 (N_3881,N_3762,N_3744);
xor U3882 (N_3882,N_3788,N_3756);
nor U3883 (N_3883,N_3789,N_3792);
and U3884 (N_3884,N_3738,N_3715);
and U3885 (N_3885,N_3731,N_3797);
xnor U3886 (N_3886,N_3785,N_3775);
xnor U3887 (N_3887,N_3732,N_3770);
and U3888 (N_3888,N_3753,N_3752);
and U3889 (N_3889,N_3725,N_3752);
nand U3890 (N_3890,N_3758,N_3777);
or U3891 (N_3891,N_3760,N_3710);
xor U3892 (N_3892,N_3728,N_3798);
or U3893 (N_3893,N_3719,N_3739);
nand U3894 (N_3894,N_3719,N_3713);
nand U3895 (N_3895,N_3743,N_3763);
xor U3896 (N_3896,N_3788,N_3763);
nand U3897 (N_3897,N_3752,N_3797);
and U3898 (N_3898,N_3738,N_3722);
nor U3899 (N_3899,N_3721,N_3725);
nor U3900 (N_3900,N_3857,N_3841);
nand U3901 (N_3901,N_3885,N_3886);
nor U3902 (N_3902,N_3828,N_3853);
nand U3903 (N_3903,N_3868,N_3844);
and U3904 (N_3904,N_3862,N_3845);
xnor U3905 (N_3905,N_3892,N_3811);
xnor U3906 (N_3906,N_3891,N_3840);
or U3907 (N_3907,N_3877,N_3842);
nor U3908 (N_3908,N_3898,N_3863);
or U3909 (N_3909,N_3876,N_3855);
and U3910 (N_3910,N_3875,N_3814);
nor U3911 (N_3911,N_3893,N_3881);
or U3912 (N_3912,N_3895,N_3807);
and U3913 (N_3913,N_3899,N_3829);
nand U3914 (N_3914,N_3874,N_3860);
nor U3915 (N_3915,N_3831,N_3882);
nor U3916 (N_3916,N_3819,N_3833);
and U3917 (N_3917,N_3854,N_3843);
and U3918 (N_3918,N_3835,N_3884);
nor U3919 (N_3919,N_3834,N_3866);
xnor U3920 (N_3920,N_3847,N_3896);
or U3921 (N_3921,N_3888,N_3825);
xor U3922 (N_3922,N_3890,N_3837);
and U3923 (N_3923,N_3872,N_3894);
or U3924 (N_3924,N_3817,N_3826);
xnor U3925 (N_3925,N_3809,N_3830);
and U3926 (N_3926,N_3887,N_3801);
xor U3927 (N_3927,N_3832,N_3827);
or U3928 (N_3928,N_3858,N_3864);
and U3929 (N_3929,N_3824,N_3851);
and U3930 (N_3930,N_3823,N_3813);
nor U3931 (N_3931,N_3856,N_3804);
or U3932 (N_3932,N_3808,N_3879);
nand U3933 (N_3933,N_3848,N_3861);
and U3934 (N_3934,N_3846,N_3805);
nor U3935 (N_3935,N_3850,N_3897);
and U3936 (N_3936,N_3815,N_3810);
xnor U3937 (N_3937,N_3883,N_3852);
xnor U3938 (N_3938,N_3873,N_3820);
or U3939 (N_3939,N_3859,N_3803);
xor U3940 (N_3940,N_3816,N_3821);
and U3941 (N_3941,N_3802,N_3812);
xor U3942 (N_3942,N_3870,N_3878);
nor U3943 (N_3943,N_3865,N_3839);
or U3944 (N_3944,N_3869,N_3836);
xor U3945 (N_3945,N_3806,N_3822);
or U3946 (N_3946,N_3867,N_3838);
and U3947 (N_3947,N_3871,N_3800);
xor U3948 (N_3948,N_3849,N_3880);
nor U3949 (N_3949,N_3818,N_3889);
or U3950 (N_3950,N_3846,N_3817);
or U3951 (N_3951,N_3855,N_3821);
nand U3952 (N_3952,N_3845,N_3855);
nor U3953 (N_3953,N_3886,N_3858);
and U3954 (N_3954,N_3889,N_3820);
nor U3955 (N_3955,N_3814,N_3862);
nor U3956 (N_3956,N_3800,N_3876);
nor U3957 (N_3957,N_3844,N_3895);
nor U3958 (N_3958,N_3851,N_3808);
or U3959 (N_3959,N_3802,N_3870);
xor U3960 (N_3960,N_3842,N_3819);
or U3961 (N_3961,N_3851,N_3864);
and U3962 (N_3962,N_3831,N_3878);
nor U3963 (N_3963,N_3877,N_3846);
nor U3964 (N_3964,N_3865,N_3828);
nand U3965 (N_3965,N_3810,N_3856);
nor U3966 (N_3966,N_3805,N_3810);
and U3967 (N_3967,N_3890,N_3868);
nand U3968 (N_3968,N_3807,N_3880);
xnor U3969 (N_3969,N_3849,N_3822);
and U3970 (N_3970,N_3893,N_3863);
nor U3971 (N_3971,N_3808,N_3842);
xor U3972 (N_3972,N_3890,N_3818);
xor U3973 (N_3973,N_3867,N_3825);
and U3974 (N_3974,N_3874,N_3872);
or U3975 (N_3975,N_3837,N_3884);
or U3976 (N_3976,N_3801,N_3836);
or U3977 (N_3977,N_3804,N_3867);
nand U3978 (N_3978,N_3845,N_3829);
nor U3979 (N_3979,N_3847,N_3856);
and U3980 (N_3980,N_3824,N_3803);
or U3981 (N_3981,N_3881,N_3814);
or U3982 (N_3982,N_3801,N_3843);
nor U3983 (N_3983,N_3819,N_3860);
and U3984 (N_3984,N_3850,N_3872);
nand U3985 (N_3985,N_3860,N_3871);
nor U3986 (N_3986,N_3898,N_3893);
nor U3987 (N_3987,N_3822,N_3827);
and U3988 (N_3988,N_3836,N_3845);
nor U3989 (N_3989,N_3828,N_3834);
xnor U3990 (N_3990,N_3817,N_3854);
and U3991 (N_3991,N_3805,N_3842);
or U3992 (N_3992,N_3852,N_3819);
nor U3993 (N_3993,N_3834,N_3856);
and U3994 (N_3994,N_3897,N_3841);
and U3995 (N_3995,N_3888,N_3899);
nand U3996 (N_3996,N_3878,N_3858);
or U3997 (N_3997,N_3873,N_3834);
nand U3998 (N_3998,N_3891,N_3885);
or U3999 (N_3999,N_3835,N_3832);
xnor U4000 (N_4000,N_3988,N_3917);
and U4001 (N_4001,N_3954,N_3991);
nor U4002 (N_4002,N_3985,N_3999);
xnor U4003 (N_4003,N_3942,N_3918);
xor U4004 (N_4004,N_3997,N_3919);
or U4005 (N_4005,N_3978,N_3902);
nor U4006 (N_4006,N_3996,N_3940);
or U4007 (N_4007,N_3965,N_3903);
nand U4008 (N_4008,N_3957,N_3921);
nor U4009 (N_4009,N_3964,N_3935);
nor U4010 (N_4010,N_3911,N_3923);
nor U4011 (N_4011,N_3951,N_3992);
or U4012 (N_4012,N_3907,N_3941);
nand U4013 (N_4013,N_3948,N_3974);
nor U4014 (N_4014,N_3938,N_3995);
or U4015 (N_4015,N_3910,N_3937);
nor U4016 (N_4016,N_3947,N_3972);
and U4017 (N_4017,N_3900,N_3932);
nand U4018 (N_4018,N_3959,N_3977);
nor U4019 (N_4019,N_3933,N_3967);
nand U4020 (N_4020,N_3924,N_3987);
xor U4021 (N_4021,N_3962,N_3909);
and U4022 (N_4022,N_3906,N_3958);
nor U4023 (N_4023,N_3931,N_3908);
or U4024 (N_4024,N_3980,N_3914);
nand U4025 (N_4025,N_3949,N_3922);
xor U4026 (N_4026,N_3927,N_3901);
xor U4027 (N_4027,N_3950,N_3973);
and U4028 (N_4028,N_3970,N_3971);
nand U4029 (N_4029,N_3952,N_3989);
and U4030 (N_4030,N_3946,N_3955);
and U4031 (N_4031,N_3915,N_3963);
xor U4032 (N_4032,N_3979,N_3934);
nand U4033 (N_4033,N_3945,N_3913);
and U4034 (N_4034,N_3939,N_3925);
nand U4035 (N_4035,N_3904,N_3916);
and U4036 (N_4036,N_3998,N_3994);
nor U4037 (N_4037,N_3936,N_3968);
xor U4038 (N_4038,N_3983,N_3976);
nand U4039 (N_4039,N_3928,N_3912);
or U4040 (N_4040,N_3981,N_3926);
xnor U4041 (N_4041,N_3929,N_3993);
xor U4042 (N_4042,N_3920,N_3966);
nor U4043 (N_4043,N_3956,N_3943);
nand U4044 (N_4044,N_3986,N_3969);
nor U4045 (N_4045,N_3990,N_3905);
and U4046 (N_4046,N_3975,N_3960);
or U4047 (N_4047,N_3930,N_3984);
and U4048 (N_4048,N_3961,N_3982);
and U4049 (N_4049,N_3953,N_3944);
nand U4050 (N_4050,N_3912,N_3933);
and U4051 (N_4051,N_3954,N_3980);
nor U4052 (N_4052,N_3954,N_3940);
and U4053 (N_4053,N_3908,N_3943);
and U4054 (N_4054,N_3988,N_3977);
and U4055 (N_4055,N_3911,N_3960);
nand U4056 (N_4056,N_3950,N_3952);
xnor U4057 (N_4057,N_3960,N_3933);
and U4058 (N_4058,N_3971,N_3927);
xor U4059 (N_4059,N_3943,N_3921);
and U4060 (N_4060,N_3979,N_3916);
or U4061 (N_4061,N_3977,N_3928);
and U4062 (N_4062,N_3935,N_3902);
xor U4063 (N_4063,N_3957,N_3969);
nor U4064 (N_4064,N_3931,N_3976);
nand U4065 (N_4065,N_3965,N_3974);
nand U4066 (N_4066,N_3966,N_3934);
or U4067 (N_4067,N_3961,N_3927);
nand U4068 (N_4068,N_3957,N_3932);
nor U4069 (N_4069,N_3916,N_3962);
and U4070 (N_4070,N_3937,N_3939);
nand U4071 (N_4071,N_3913,N_3994);
nor U4072 (N_4072,N_3931,N_3901);
or U4073 (N_4073,N_3945,N_3944);
and U4074 (N_4074,N_3979,N_3987);
and U4075 (N_4075,N_3926,N_3986);
nor U4076 (N_4076,N_3987,N_3958);
xnor U4077 (N_4077,N_3978,N_3931);
xor U4078 (N_4078,N_3906,N_3992);
and U4079 (N_4079,N_3959,N_3998);
nor U4080 (N_4080,N_3938,N_3967);
xnor U4081 (N_4081,N_3982,N_3958);
nand U4082 (N_4082,N_3983,N_3945);
xor U4083 (N_4083,N_3915,N_3911);
or U4084 (N_4084,N_3922,N_3948);
nand U4085 (N_4085,N_3914,N_3911);
and U4086 (N_4086,N_3996,N_3963);
nand U4087 (N_4087,N_3914,N_3996);
nand U4088 (N_4088,N_3925,N_3912);
nand U4089 (N_4089,N_3968,N_3949);
nand U4090 (N_4090,N_3976,N_3908);
and U4091 (N_4091,N_3901,N_3935);
and U4092 (N_4092,N_3925,N_3936);
xnor U4093 (N_4093,N_3960,N_3952);
and U4094 (N_4094,N_3912,N_3962);
nor U4095 (N_4095,N_3934,N_3973);
xor U4096 (N_4096,N_3960,N_3966);
or U4097 (N_4097,N_3902,N_3973);
or U4098 (N_4098,N_3907,N_3965);
or U4099 (N_4099,N_3977,N_3915);
and U4100 (N_4100,N_4025,N_4002);
and U4101 (N_4101,N_4055,N_4067);
nor U4102 (N_4102,N_4045,N_4044);
nor U4103 (N_4103,N_4027,N_4083);
xor U4104 (N_4104,N_4033,N_4094);
and U4105 (N_4105,N_4056,N_4069);
and U4106 (N_4106,N_4029,N_4014);
or U4107 (N_4107,N_4035,N_4031);
or U4108 (N_4108,N_4077,N_4079);
nand U4109 (N_4109,N_4087,N_4024);
or U4110 (N_4110,N_4096,N_4038);
nor U4111 (N_4111,N_4074,N_4032);
xor U4112 (N_4112,N_4048,N_4093);
xor U4113 (N_4113,N_4088,N_4005);
nand U4114 (N_4114,N_4058,N_4054);
xor U4115 (N_4115,N_4061,N_4057);
xnor U4116 (N_4116,N_4066,N_4063);
and U4117 (N_4117,N_4016,N_4018);
nor U4118 (N_4118,N_4017,N_4049);
nand U4119 (N_4119,N_4006,N_4007);
xnor U4120 (N_4120,N_4026,N_4047);
nand U4121 (N_4121,N_4028,N_4073);
nor U4122 (N_4122,N_4062,N_4080);
nor U4123 (N_4123,N_4059,N_4082);
or U4124 (N_4124,N_4003,N_4011);
and U4125 (N_4125,N_4004,N_4076);
and U4126 (N_4126,N_4099,N_4065);
and U4127 (N_4127,N_4075,N_4060);
nand U4128 (N_4128,N_4034,N_4064);
nand U4129 (N_4129,N_4012,N_4091);
nand U4130 (N_4130,N_4019,N_4037);
nor U4131 (N_4131,N_4015,N_4086);
xor U4132 (N_4132,N_4081,N_4040);
nand U4133 (N_4133,N_4092,N_4097);
nor U4134 (N_4134,N_4013,N_4041);
nand U4135 (N_4135,N_4046,N_4009);
or U4136 (N_4136,N_4023,N_4039);
nor U4137 (N_4137,N_4053,N_4000);
nand U4138 (N_4138,N_4050,N_4078);
and U4139 (N_4139,N_4051,N_4021);
nand U4140 (N_4140,N_4043,N_4095);
xnor U4141 (N_4141,N_4084,N_4001);
xnor U4142 (N_4142,N_4070,N_4036);
or U4143 (N_4143,N_4072,N_4098);
or U4144 (N_4144,N_4008,N_4020);
xor U4145 (N_4145,N_4071,N_4068);
and U4146 (N_4146,N_4090,N_4052);
or U4147 (N_4147,N_4089,N_4042);
xnor U4148 (N_4148,N_4010,N_4030);
nor U4149 (N_4149,N_4085,N_4022);
xnor U4150 (N_4150,N_4002,N_4096);
xnor U4151 (N_4151,N_4018,N_4081);
nor U4152 (N_4152,N_4017,N_4073);
xor U4153 (N_4153,N_4041,N_4087);
or U4154 (N_4154,N_4069,N_4000);
nand U4155 (N_4155,N_4055,N_4096);
and U4156 (N_4156,N_4098,N_4020);
nand U4157 (N_4157,N_4022,N_4038);
and U4158 (N_4158,N_4037,N_4032);
nand U4159 (N_4159,N_4016,N_4083);
or U4160 (N_4160,N_4080,N_4021);
nand U4161 (N_4161,N_4015,N_4029);
nor U4162 (N_4162,N_4081,N_4091);
nand U4163 (N_4163,N_4044,N_4066);
nand U4164 (N_4164,N_4060,N_4026);
nand U4165 (N_4165,N_4004,N_4020);
nand U4166 (N_4166,N_4085,N_4096);
nor U4167 (N_4167,N_4066,N_4073);
nor U4168 (N_4168,N_4099,N_4031);
nor U4169 (N_4169,N_4092,N_4038);
nor U4170 (N_4170,N_4003,N_4080);
or U4171 (N_4171,N_4021,N_4022);
xnor U4172 (N_4172,N_4057,N_4085);
and U4173 (N_4173,N_4084,N_4085);
nor U4174 (N_4174,N_4043,N_4007);
and U4175 (N_4175,N_4020,N_4092);
or U4176 (N_4176,N_4028,N_4034);
nand U4177 (N_4177,N_4038,N_4089);
nor U4178 (N_4178,N_4056,N_4098);
or U4179 (N_4179,N_4054,N_4078);
nand U4180 (N_4180,N_4022,N_4065);
and U4181 (N_4181,N_4098,N_4099);
and U4182 (N_4182,N_4043,N_4010);
and U4183 (N_4183,N_4065,N_4089);
nand U4184 (N_4184,N_4098,N_4044);
xnor U4185 (N_4185,N_4052,N_4022);
xor U4186 (N_4186,N_4019,N_4035);
xnor U4187 (N_4187,N_4017,N_4048);
xor U4188 (N_4188,N_4044,N_4051);
nor U4189 (N_4189,N_4091,N_4053);
nor U4190 (N_4190,N_4002,N_4061);
nor U4191 (N_4191,N_4020,N_4056);
nand U4192 (N_4192,N_4091,N_4049);
or U4193 (N_4193,N_4014,N_4001);
nand U4194 (N_4194,N_4088,N_4022);
nor U4195 (N_4195,N_4015,N_4043);
xor U4196 (N_4196,N_4093,N_4062);
nand U4197 (N_4197,N_4089,N_4096);
nor U4198 (N_4198,N_4091,N_4046);
xor U4199 (N_4199,N_4059,N_4056);
and U4200 (N_4200,N_4134,N_4199);
or U4201 (N_4201,N_4153,N_4128);
nor U4202 (N_4202,N_4183,N_4152);
nor U4203 (N_4203,N_4157,N_4130);
nor U4204 (N_4204,N_4162,N_4169);
xnor U4205 (N_4205,N_4181,N_4186);
and U4206 (N_4206,N_4146,N_4116);
or U4207 (N_4207,N_4138,N_4120);
or U4208 (N_4208,N_4192,N_4165);
xnor U4209 (N_4209,N_4109,N_4127);
nor U4210 (N_4210,N_4139,N_4182);
xor U4211 (N_4211,N_4119,N_4133);
nand U4212 (N_4212,N_4121,N_4194);
and U4213 (N_4213,N_4137,N_4103);
nand U4214 (N_4214,N_4164,N_4177);
nand U4215 (N_4215,N_4112,N_4148);
nor U4216 (N_4216,N_4102,N_4197);
nor U4217 (N_4217,N_4175,N_4110);
nand U4218 (N_4218,N_4161,N_4123);
nand U4219 (N_4219,N_4117,N_4129);
xnor U4220 (N_4220,N_4154,N_4172);
nand U4221 (N_4221,N_4118,N_4189);
xnor U4222 (N_4222,N_4104,N_4114);
nor U4223 (N_4223,N_4179,N_4173);
nor U4224 (N_4224,N_4168,N_4125);
nor U4225 (N_4225,N_4131,N_4174);
nand U4226 (N_4226,N_4107,N_4171);
nor U4227 (N_4227,N_4188,N_4176);
nor U4228 (N_4228,N_4149,N_4106);
and U4229 (N_4229,N_4170,N_4126);
and U4230 (N_4230,N_4196,N_4105);
nor U4231 (N_4231,N_4108,N_4140);
and U4232 (N_4232,N_4191,N_4135);
xor U4233 (N_4233,N_4184,N_4145);
nor U4234 (N_4234,N_4156,N_4163);
nor U4235 (N_4235,N_4100,N_4187);
xor U4236 (N_4236,N_4185,N_4122);
and U4237 (N_4237,N_4155,N_4180);
and U4238 (N_4238,N_4151,N_4178);
or U4239 (N_4239,N_4132,N_4124);
nor U4240 (N_4240,N_4159,N_4141);
or U4241 (N_4241,N_4190,N_4193);
xnor U4242 (N_4242,N_4111,N_4158);
or U4243 (N_4243,N_4115,N_4198);
nor U4244 (N_4244,N_4195,N_4150);
or U4245 (N_4245,N_4101,N_4144);
and U4246 (N_4246,N_4167,N_4147);
xnor U4247 (N_4247,N_4142,N_4160);
nor U4248 (N_4248,N_4113,N_4143);
and U4249 (N_4249,N_4136,N_4166);
xor U4250 (N_4250,N_4132,N_4143);
and U4251 (N_4251,N_4135,N_4149);
xnor U4252 (N_4252,N_4146,N_4142);
and U4253 (N_4253,N_4166,N_4167);
nand U4254 (N_4254,N_4133,N_4176);
nor U4255 (N_4255,N_4198,N_4142);
or U4256 (N_4256,N_4109,N_4146);
nor U4257 (N_4257,N_4118,N_4109);
or U4258 (N_4258,N_4158,N_4190);
xor U4259 (N_4259,N_4162,N_4105);
nand U4260 (N_4260,N_4137,N_4194);
or U4261 (N_4261,N_4142,N_4158);
nor U4262 (N_4262,N_4179,N_4191);
nor U4263 (N_4263,N_4163,N_4122);
and U4264 (N_4264,N_4154,N_4177);
nand U4265 (N_4265,N_4110,N_4188);
and U4266 (N_4266,N_4198,N_4106);
or U4267 (N_4267,N_4109,N_4112);
xnor U4268 (N_4268,N_4197,N_4194);
nor U4269 (N_4269,N_4101,N_4134);
and U4270 (N_4270,N_4127,N_4176);
or U4271 (N_4271,N_4195,N_4141);
xnor U4272 (N_4272,N_4169,N_4173);
nand U4273 (N_4273,N_4194,N_4135);
or U4274 (N_4274,N_4186,N_4137);
and U4275 (N_4275,N_4195,N_4134);
or U4276 (N_4276,N_4126,N_4131);
or U4277 (N_4277,N_4115,N_4141);
and U4278 (N_4278,N_4182,N_4181);
xor U4279 (N_4279,N_4193,N_4152);
nand U4280 (N_4280,N_4168,N_4130);
or U4281 (N_4281,N_4137,N_4196);
nand U4282 (N_4282,N_4150,N_4136);
and U4283 (N_4283,N_4129,N_4195);
and U4284 (N_4284,N_4171,N_4121);
or U4285 (N_4285,N_4131,N_4182);
nor U4286 (N_4286,N_4103,N_4195);
nor U4287 (N_4287,N_4175,N_4115);
nand U4288 (N_4288,N_4164,N_4151);
and U4289 (N_4289,N_4153,N_4186);
and U4290 (N_4290,N_4161,N_4150);
and U4291 (N_4291,N_4198,N_4151);
nand U4292 (N_4292,N_4166,N_4152);
and U4293 (N_4293,N_4167,N_4199);
or U4294 (N_4294,N_4181,N_4163);
nor U4295 (N_4295,N_4127,N_4182);
or U4296 (N_4296,N_4142,N_4152);
xnor U4297 (N_4297,N_4160,N_4141);
or U4298 (N_4298,N_4197,N_4176);
xor U4299 (N_4299,N_4186,N_4125);
nand U4300 (N_4300,N_4242,N_4240);
xor U4301 (N_4301,N_4270,N_4215);
and U4302 (N_4302,N_4287,N_4296);
or U4303 (N_4303,N_4221,N_4241);
nand U4304 (N_4304,N_4204,N_4294);
nand U4305 (N_4305,N_4274,N_4214);
nor U4306 (N_4306,N_4254,N_4276);
nand U4307 (N_4307,N_4228,N_4299);
and U4308 (N_4308,N_4236,N_4277);
and U4309 (N_4309,N_4283,N_4208);
and U4310 (N_4310,N_4249,N_4206);
or U4311 (N_4311,N_4278,N_4268);
or U4312 (N_4312,N_4225,N_4293);
nor U4313 (N_4313,N_4253,N_4265);
xnor U4314 (N_4314,N_4269,N_4262);
and U4315 (N_4315,N_4224,N_4203);
nor U4316 (N_4316,N_4280,N_4210);
or U4317 (N_4317,N_4211,N_4251);
xor U4318 (N_4318,N_4267,N_4288);
and U4319 (N_4319,N_4229,N_4271);
or U4320 (N_4320,N_4233,N_4201);
nor U4321 (N_4321,N_4218,N_4220);
and U4322 (N_4322,N_4272,N_4266);
xor U4323 (N_4323,N_4295,N_4258);
nor U4324 (N_4324,N_4235,N_4226);
or U4325 (N_4325,N_4244,N_4264);
nor U4326 (N_4326,N_4222,N_4216);
or U4327 (N_4327,N_4246,N_4292);
nor U4328 (N_4328,N_4217,N_4291);
xnor U4329 (N_4329,N_4237,N_4261);
nand U4330 (N_4330,N_4243,N_4232);
and U4331 (N_4331,N_4248,N_4239);
nor U4332 (N_4332,N_4257,N_4207);
or U4333 (N_4333,N_4285,N_4290);
xnor U4334 (N_4334,N_4238,N_4223);
nand U4335 (N_4335,N_4205,N_4209);
nor U4336 (N_4336,N_4252,N_4213);
nand U4337 (N_4337,N_4212,N_4260);
nand U4338 (N_4338,N_4250,N_4230);
nand U4339 (N_4339,N_4202,N_4247);
or U4340 (N_4340,N_4275,N_4219);
or U4341 (N_4341,N_4282,N_4298);
nand U4342 (N_4342,N_4259,N_4227);
nor U4343 (N_4343,N_4256,N_4245);
and U4344 (N_4344,N_4286,N_4263);
or U4345 (N_4345,N_4200,N_4234);
xor U4346 (N_4346,N_4255,N_4297);
xnor U4347 (N_4347,N_4231,N_4273);
nand U4348 (N_4348,N_4284,N_4279);
and U4349 (N_4349,N_4281,N_4289);
and U4350 (N_4350,N_4297,N_4269);
nor U4351 (N_4351,N_4204,N_4291);
nand U4352 (N_4352,N_4232,N_4218);
xor U4353 (N_4353,N_4269,N_4245);
nand U4354 (N_4354,N_4201,N_4281);
nand U4355 (N_4355,N_4206,N_4286);
or U4356 (N_4356,N_4274,N_4239);
nand U4357 (N_4357,N_4240,N_4213);
and U4358 (N_4358,N_4245,N_4218);
and U4359 (N_4359,N_4288,N_4253);
xnor U4360 (N_4360,N_4212,N_4283);
nor U4361 (N_4361,N_4208,N_4267);
or U4362 (N_4362,N_4276,N_4252);
or U4363 (N_4363,N_4263,N_4250);
or U4364 (N_4364,N_4211,N_4281);
or U4365 (N_4365,N_4270,N_4236);
xnor U4366 (N_4366,N_4267,N_4210);
or U4367 (N_4367,N_4267,N_4253);
xnor U4368 (N_4368,N_4289,N_4207);
nand U4369 (N_4369,N_4267,N_4246);
nor U4370 (N_4370,N_4261,N_4221);
nor U4371 (N_4371,N_4230,N_4271);
or U4372 (N_4372,N_4216,N_4251);
and U4373 (N_4373,N_4208,N_4235);
nor U4374 (N_4374,N_4277,N_4262);
and U4375 (N_4375,N_4286,N_4282);
xor U4376 (N_4376,N_4218,N_4277);
nand U4377 (N_4377,N_4209,N_4283);
or U4378 (N_4378,N_4232,N_4284);
or U4379 (N_4379,N_4262,N_4234);
and U4380 (N_4380,N_4206,N_4207);
xnor U4381 (N_4381,N_4290,N_4225);
xor U4382 (N_4382,N_4294,N_4202);
and U4383 (N_4383,N_4254,N_4251);
nand U4384 (N_4384,N_4279,N_4239);
xor U4385 (N_4385,N_4212,N_4211);
nor U4386 (N_4386,N_4231,N_4268);
and U4387 (N_4387,N_4294,N_4285);
nor U4388 (N_4388,N_4287,N_4254);
nand U4389 (N_4389,N_4223,N_4276);
nand U4390 (N_4390,N_4201,N_4248);
or U4391 (N_4391,N_4227,N_4201);
or U4392 (N_4392,N_4206,N_4256);
nand U4393 (N_4393,N_4293,N_4268);
nand U4394 (N_4394,N_4295,N_4283);
or U4395 (N_4395,N_4287,N_4294);
nand U4396 (N_4396,N_4204,N_4251);
nor U4397 (N_4397,N_4229,N_4274);
or U4398 (N_4398,N_4276,N_4248);
and U4399 (N_4399,N_4237,N_4218);
nand U4400 (N_4400,N_4381,N_4356);
nor U4401 (N_4401,N_4303,N_4376);
nand U4402 (N_4402,N_4305,N_4331);
or U4403 (N_4403,N_4384,N_4363);
or U4404 (N_4404,N_4369,N_4340);
nand U4405 (N_4405,N_4396,N_4385);
nor U4406 (N_4406,N_4316,N_4313);
and U4407 (N_4407,N_4374,N_4332);
nand U4408 (N_4408,N_4368,N_4373);
or U4409 (N_4409,N_4353,N_4317);
nand U4410 (N_4410,N_4338,N_4329);
nand U4411 (N_4411,N_4318,N_4386);
xor U4412 (N_4412,N_4304,N_4383);
or U4413 (N_4413,N_4394,N_4351);
xnor U4414 (N_4414,N_4314,N_4310);
nand U4415 (N_4415,N_4342,N_4359);
xor U4416 (N_4416,N_4336,N_4311);
or U4417 (N_4417,N_4308,N_4354);
xnor U4418 (N_4418,N_4377,N_4387);
or U4419 (N_4419,N_4350,N_4378);
xnor U4420 (N_4420,N_4388,N_4301);
and U4421 (N_4421,N_4325,N_4371);
nand U4422 (N_4422,N_4333,N_4343);
xor U4423 (N_4423,N_4328,N_4339);
or U4424 (N_4424,N_4393,N_4346);
or U4425 (N_4425,N_4380,N_4307);
nor U4426 (N_4426,N_4365,N_4352);
nor U4427 (N_4427,N_4399,N_4321);
nor U4428 (N_4428,N_4366,N_4344);
nor U4429 (N_4429,N_4355,N_4361);
or U4430 (N_4430,N_4390,N_4389);
nand U4431 (N_4431,N_4364,N_4322);
and U4432 (N_4432,N_4392,N_4372);
xnor U4433 (N_4433,N_4347,N_4312);
or U4434 (N_4434,N_4315,N_4391);
xnor U4435 (N_4435,N_4323,N_4362);
nor U4436 (N_4436,N_4335,N_4379);
xnor U4437 (N_4437,N_4306,N_4324);
xor U4438 (N_4438,N_4334,N_4375);
nor U4439 (N_4439,N_4319,N_4345);
or U4440 (N_4440,N_4357,N_4367);
or U4441 (N_4441,N_4326,N_4341);
nand U4442 (N_4442,N_4330,N_4349);
xor U4443 (N_4443,N_4320,N_4382);
xnor U4444 (N_4444,N_4300,N_4397);
nor U4445 (N_4445,N_4337,N_4302);
or U4446 (N_4446,N_4348,N_4395);
nand U4447 (N_4447,N_4370,N_4360);
nand U4448 (N_4448,N_4398,N_4327);
or U4449 (N_4449,N_4309,N_4358);
or U4450 (N_4450,N_4321,N_4328);
nor U4451 (N_4451,N_4392,N_4349);
and U4452 (N_4452,N_4301,N_4377);
and U4453 (N_4453,N_4385,N_4393);
or U4454 (N_4454,N_4331,N_4378);
xnor U4455 (N_4455,N_4334,N_4360);
and U4456 (N_4456,N_4398,N_4356);
xnor U4457 (N_4457,N_4388,N_4328);
or U4458 (N_4458,N_4368,N_4398);
xnor U4459 (N_4459,N_4362,N_4326);
and U4460 (N_4460,N_4350,N_4377);
and U4461 (N_4461,N_4381,N_4340);
nor U4462 (N_4462,N_4323,N_4393);
xnor U4463 (N_4463,N_4386,N_4341);
and U4464 (N_4464,N_4307,N_4363);
nor U4465 (N_4465,N_4349,N_4379);
xor U4466 (N_4466,N_4306,N_4335);
and U4467 (N_4467,N_4300,N_4395);
or U4468 (N_4468,N_4398,N_4314);
and U4469 (N_4469,N_4303,N_4391);
nand U4470 (N_4470,N_4396,N_4359);
nor U4471 (N_4471,N_4378,N_4307);
nor U4472 (N_4472,N_4333,N_4380);
or U4473 (N_4473,N_4354,N_4376);
nand U4474 (N_4474,N_4314,N_4386);
nand U4475 (N_4475,N_4357,N_4315);
nor U4476 (N_4476,N_4323,N_4353);
nor U4477 (N_4477,N_4382,N_4367);
nand U4478 (N_4478,N_4305,N_4378);
and U4479 (N_4479,N_4399,N_4322);
xnor U4480 (N_4480,N_4363,N_4364);
or U4481 (N_4481,N_4306,N_4353);
nand U4482 (N_4482,N_4338,N_4337);
xnor U4483 (N_4483,N_4370,N_4374);
and U4484 (N_4484,N_4396,N_4301);
xor U4485 (N_4485,N_4345,N_4368);
and U4486 (N_4486,N_4347,N_4356);
nor U4487 (N_4487,N_4348,N_4341);
nor U4488 (N_4488,N_4302,N_4335);
and U4489 (N_4489,N_4365,N_4392);
and U4490 (N_4490,N_4393,N_4301);
or U4491 (N_4491,N_4313,N_4356);
and U4492 (N_4492,N_4355,N_4362);
nand U4493 (N_4493,N_4334,N_4356);
nand U4494 (N_4494,N_4367,N_4340);
or U4495 (N_4495,N_4305,N_4388);
or U4496 (N_4496,N_4336,N_4393);
and U4497 (N_4497,N_4308,N_4345);
and U4498 (N_4498,N_4357,N_4394);
or U4499 (N_4499,N_4341,N_4303);
xor U4500 (N_4500,N_4406,N_4489);
or U4501 (N_4501,N_4484,N_4494);
or U4502 (N_4502,N_4416,N_4434);
and U4503 (N_4503,N_4499,N_4462);
nor U4504 (N_4504,N_4471,N_4476);
nor U4505 (N_4505,N_4419,N_4411);
xnor U4506 (N_4506,N_4437,N_4480);
or U4507 (N_4507,N_4415,N_4467);
nand U4508 (N_4508,N_4474,N_4426);
nor U4509 (N_4509,N_4403,N_4496);
nand U4510 (N_4510,N_4483,N_4478);
nand U4511 (N_4511,N_4427,N_4400);
nor U4512 (N_4512,N_4409,N_4430);
nand U4513 (N_4513,N_4444,N_4488);
xor U4514 (N_4514,N_4468,N_4482);
or U4515 (N_4515,N_4459,N_4413);
nand U4516 (N_4516,N_4423,N_4442);
xnor U4517 (N_4517,N_4420,N_4418);
nor U4518 (N_4518,N_4448,N_4487);
and U4519 (N_4519,N_4402,N_4431);
and U4520 (N_4520,N_4449,N_4455);
nand U4521 (N_4521,N_4473,N_4470);
xor U4522 (N_4522,N_4405,N_4410);
or U4523 (N_4523,N_4491,N_4446);
xor U4524 (N_4524,N_4486,N_4485);
nand U4525 (N_4525,N_4408,N_4441);
nand U4526 (N_4526,N_4439,N_4479);
and U4527 (N_4527,N_4477,N_4433);
and U4528 (N_4528,N_4464,N_4452);
xnor U4529 (N_4529,N_4414,N_4425);
nand U4530 (N_4530,N_4401,N_4466);
and U4531 (N_4531,N_4461,N_4492);
nor U4532 (N_4532,N_4428,N_4497);
nor U4533 (N_4533,N_4465,N_4404);
and U4534 (N_4534,N_4443,N_4438);
and U4535 (N_4535,N_4429,N_4436);
or U4536 (N_4536,N_4490,N_4424);
or U4537 (N_4537,N_4454,N_4440);
or U4538 (N_4538,N_4475,N_4481);
nand U4539 (N_4539,N_4412,N_4456);
nand U4540 (N_4540,N_4417,N_4460);
xnor U4541 (N_4541,N_4458,N_4498);
xnor U4542 (N_4542,N_4453,N_4457);
and U4543 (N_4543,N_4451,N_4472);
and U4544 (N_4544,N_4469,N_4421);
nand U4545 (N_4545,N_4447,N_4407);
xor U4546 (N_4546,N_4495,N_4435);
xor U4547 (N_4547,N_4445,N_4422);
and U4548 (N_4548,N_4432,N_4450);
xor U4549 (N_4549,N_4493,N_4463);
nor U4550 (N_4550,N_4461,N_4421);
nor U4551 (N_4551,N_4450,N_4415);
or U4552 (N_4552,N_4468,N_4403);
and U4553 (N_4553,N_4494,N_4481);
or U4554 (N_4554,N_4459,N_4404);
nand U4555 (N_4555,N_4454,N_4494);
or U4556 (N_4556,N_4436,N_4491);
and U4557 (N_4557,N_4449,N_4439);
and U4558 (N_4558,N_4408,N_4475);
and U4559 (N_4559,N_4408,N_4437);
nor U4560 (N_4560,N_4461,N_4494);
xor U4561 (N_4561,N_4479,N_4460);
and U4562 (N_4562,N_4452,N_4422);
or U4563 (N_4563,N_4470,N_4490);
nor U4564 (N_4564,N_4496,N_4426);
nor U4565 (N_4565,N_4469,N_4496);
nor U4566 (N_4566,N_4459,N_4400);
nor U4567 (N_4567,N_4462,N_4442);
nor U4568 (N_4568,N_4407,N_4493);
or U4569 (N_4569,N_4427,N_4459);
nor U4570 (N_4570,N_4450,N_4491);
and U4571 (N_4571,N_4442,N_4477);
nor U4572 (N_4572,N_4401,N_4445);
nor U4573 (N_4573,N_4434,N_4438);
and U4574 (N_4574,N_4481,N_4448);
nor U4575 (N_4575,N_4449,N_4426);
or U4576 (N_4576,N_4431,N_4437);
nand U4577 (N_4577,N_4489,N_4402);
and U4578 (N_4578,N_4436,N_4467);
and U4579 (N_4579,N_4449,N_4496);
and U4580 (N_4580,N_4411,N_4468);
nand U4581 (N_4581,N_4421,N_4440);
or U4582 (N_4582,N_4485,N_4482);
xnor U4583 (N_4583,N_4433,N_4488);
xnor U4584 (N_4584,N_4419,N_4492);
nor U4585 (N_4585,N_4493,N_4462);
or U4586 (N_4586,N_4427,N_4454);
or U4587 (N_4587,N_4457,N_4452);
nor U4588 (N_4588,N_4429,N_4480);
and U4589 (N_4589,N_4406,N_4417);
or U4590 (N_4590,N_4413,N_4487);
nor U4591 (N_4591,N_4419,N_4427);
xor U4592 (N_4592,N_4414,N_4438);
and U4593 (N_4593,N_4419,N_4445);
xnor U4594 (N_4594,N_4491,N_4495);
nand U4595 (N_4595,N_4498,N_4445);
and U4596 (N_4596,N_4408,N_4442);
nand U4597 (N_4597,N_4488,N_4418);
nand U4598 (N_4598,N_4424,N_4400);
xnor U4599 (N_4599,N_4401,N_4485);
nor U4600 (N_4600,N_4581,N_4586);
nand U4601 (N_4601,N_4584,N_4582);
and U4602 (N_4602,N_4598,N_4564);
or U4603 (N_4603,N_4592,N_4530);
nand U4604 (N_4604,N_4557,N_4572);
and U4605 (N_4605,N_4569,N_4541);
nand U4606 (N_4606,N_4590,N_4507);
xor U4607 (N_4607,N_4567,N_4548);
or U4608 (N_4608,N_4501,N_4558);
xnor U4609 (N_4609,N_4596,N_4540);
and U4610 (N_4610,N_4543,N_4510);
and U4611 (N_4611,N_4579,N_4553);
nor U4612 (N_4612,N_4528,N_4517);
or U4613 (N_4613,N_4515,N_4594);
and U4614 (N_4614,N_4589,N_4538);
or U4615 (N_4615,N_4576,N_4570);
nand U4616 (N_4616,N_4580,N_4568);
xor U4617 (N_4617,N_4560,N_4516);
nand U4618 (N_4618,N_4574,N_4591);
or U4619 (N_4619,N_4518,N_4512);
nor U4620 (N_4620,N_4542,N_4559);
or U4621 (N_4621,N_4513,N_4545);
nand U4622 (N_4622,N_4531,N_4539);
nand U4623 (N_4623,N_4504,N_4593);
and U4624 (N_4624,N_4523,N_4566);
or U4625 (N_4625,N_4522,N_4521);
nor U4626 (N_4626,N_4561,N_4527);
nor U4627 (N_4627,N_4571,N_4503);
nor U4628 (N_4628,N_4555,N_4599);
or U4629 (N_4629,N_4597,N_4502);
xor U4630 (N_4630,N_4583,N_4500);
and U4631 (N_4631,N_4595,N_4549);
or U4632 (N_4632,N_4573,N_4550);
and U4633 (N_4633,N_4575,N_4533);
nand U4634 (N_4634,N_4556,N_4544);
or U4635 (N_4635,N_4534,N_4519);
xor U4636 (N_4636,N_4511,N_4562);
and U4637 (N_4637,N_4546,N_4578);
nand U4638 (N_4638,N_4588,N_4514);
nor U4639 (N_4639,N_4535,N_4506);
nand U4640 (N_4640,N_4532,N_4509);
nand U4641 (N_4641,N_4508,N_4520);
nor U4642 (N_4642,N_4536,N_4537);
xnor U4643 (N_4643,N_4505,N_4585);
xnor U4644 (N_4644,N_4525,N_4526);
or U4645 (N_4645,N_4551,N_4565);
xnor U4646 (N_4646,N_4529,N_4587);
and U4647 (N_4647,N_4563,N_4552);
nor U4648 (N_4648,N_4524,N_4577);
nand U4649 (N_4649,N_4554,N_4547);
xor U4650 (N_4650,N_4582,N_4528);
and U4651 (N_4651,N_4500,N_4577);
nor U4652 (N_4652,N_4530,N_4540);
nand U4653 (N_4653,N_4521,N_4571);
nand U4654 (N_4654,N_4510,N_4554);
and U4655 (N_4655,N_4535,N_4564);
and U4656 (N_4656,N_4593,N_4563);
nand U4657 (N_4657,N_4557,N_4517);
xnor U4658 (N_4658,N_4512,N_4555);
or U4659 (N_4659,N_4580,N_4556);
xor U4660 (N_4660,N_4560,N_4542);
and U4661 (N_4661,N_4520,N_4559);
xnor U4662 (N_4662,N_4533,N_4512);
nand U4663 (N_4663,N_4565,N_4579);
xnor U4664 (N_4664,N_4570,N_4537);
or U4665 (N_4665,N_4554,N_4539);
or U4666 (N_4666,N_4511,N_4590);
xnor U4667 (N_4667,N_4522,N_4513);
or U4668 (N_4668,N_4589,N_4568);
nor U4669 (N_4669,N_4506,N_4505);
xnor U4670 (N_4670,N_4508,N_4512);
and U4671 (N_4671,N_4520,N_4541);
nor U4672 (N_4672,N_4574,N_4534);
nor U4673 (N_4673,N_4525,N_4574);
xor U4674 (N_4674,N_4504,N_4518);
and U4675 (N_4675,N_4575,N_4591);
and U4676 (N_4676,N_4540,N_4585);
xnor U4677 (N_4677,N_4556,N_4520);
or U4678 (N_4678,N_4525,N_4556);
nor U4679 (N_4679,N_4504,N_4557);
or U4680 (N_4680,N_4562,N_4528);
or U4681 (N_4681,N_4513,N_4502);
xnor U4682 (N_4682,N_4540,N_4570);
xnor U4683 (N_4683,N_4597,N_4581);
xor U4684 (N_4684,N_4565,N_4506);
xor U4685 (N_4685,N_4503,N_4567);
nor U4686 (N_4686,N_4574,N_4528);
and U4687 (N_4687,N_4543,N_4592);
xor U4688 (N_4688,N_4548,N_4539);
and U4689 (N_4689,N_4510,N_4548);
nand U4690 (N_4690,N_4507,N_4597);
xnor U4691 (N_4691,N_4594,N_4578);
nor U4692 (N_4692,N_4541,N_4585);
nor U4693 (N_4693,N_4596,N_4579);
nor U4694 (N_4694,N_4574,N_4539);
nor U4695 (N_4695,N_4544,N_4557);
nand U4696 (N_4696,N_4558,N_4550);
nand U4697 (N_4697,N_4562,N_4559);
or U4698 (N_4698,N_4523,N_4506);
or U4699 (N_4699,N_4527,N_4591);
and U4700 (N_4700,N_4646,N_4620);
nand U4701 (N_4701,N_4666,N_4695);
xor U4702 (N_4702,N_4625,N_4655);
or U4703 (N_4703,N_4665,N_4652);
nand U4704 (N_4704,N_4696,N_4673);
nand U4705 (N_4705,N_4692,N_4686);
xor U4706 (N_4706,N_4670,N_4662);
xor U4707 (N_4707,N_4647,N_4632);
xor U4708 (N_4708,N_4649,N_4667);
and U4709 (N_4709,N_4609,N_4699);
nand U4710 (N_4710,N_4641,N_4683);
nand U4711 (N_4711,N_4657,N_4614);
and U4712 (N_4712,N_4691,N_4656);
nand U4713 (N_4713,N_4644,N_4677);
xnor U4714 (N_4714,N_4602,N_4610);
nand U4715 (N_4715,N_4659,N_4611);
nand U4716 (N_4716,N_4690,N_4629);
nand U4717 (N_4717,N_4613,N_4674);
xnor U4718 (N_4718,N_4622,N_4619);
nor U4719 (N_4719,N_4668,N_4605);
xnor U4720 (N_4720,N_4661,N_4616);
xor U4721 (N_4721,N_4628,N_4624);
nor U4722 (N_4722,N_4643,N_4697);
xnor U4723 (N_4723,N_4604,N_4664);
and U4724 (N_4724,N_4617,N_4679);
or U4725 (N_4725,N_4689,N_4698);
and U4726 (N_4726,N_4653,N_4603);
or U4727 (N_4727,N_4678,N_4694);
and U4728 (N_4728,N_4636,N_4658);
and U4729 (N_4729,N_4654,N_4672);
xor U4730 (N_4730,N_4601,N_4627);
or U4731 (N_4731,N_4680,N_4612);
or U4732 (N_4732,N_4650,N_4693);
nand U4733 (N_4733,N_4633,N_4634);
nor U4734 (N_4734,N_4621,N_4631);
and U4735 (N_4735,N_4635,N_4642);
nand U4736 (N_4736,N_4600,N_4687);
nor U4737 (N_4737,N_4618,N_4630);
or U4738 (N_4738,N_4645,N_4663);
or U4739 (N_4739,N_4623,N_4637);
or U4740 (N_4740,N_4626,N_4638);
nand U4741 (N_4741,N_4688,N_4640);
or U4742 (N_4742,N_4639,N_4660);
xor U4743 (N_4743,N_4606,N_4648);
xnor U4744 (N_4744,N_4682,N_4676);
nor U4745 (N_4745,N_4671,N_4608);
nor U4746 (N_4746,N_4684,N_4607);
and U4747 (N_4747,N_4651,N_4681);
nand U4748 (N_4748,N_4675,N_4615);
nor U4749 (N_4749,N_4685,N_4669);
nand U4750 (N_4750,N_4615,N_4686);
nand U4751 (N_4751,N_4603,N_4612);
nand U4752 (N_4752,N_4609,N_4664);
xnor U4753 (N_4753,N_4605,N_4613);
and U4754 (N_4754,N_4647,N_4650);
nand U4755 (N_4755,N_4643,N_4665);
nand U4756 (N_4756,N_4698,N_4688);
or U4757 (N_4757,N_4611,N_4667);
nor U4758 (N_4758,N_4623,N_4604);
xor U4759 (N_4759,N_4606,N_4650);
and U4760 (N_4760,N_4608,N_4690);
and U4761 (N_4761,N_4688,N_4658);
or U4762 (N_4762,N_4669,N_4651);
nor U4763 (N_4763,N_4651,N_4629);
xor U4764 (N_4764,N_4603,N_4622);
xnor U4765 (N_4765,N_4674,N_4685);
xnor U4766 (N_4766,N_4695,N_4687);
and U4767 (N_4767,N_4604,N_4684);
or U4768 (N_4768,N_4673,N_4620);
or U4769 (N_4769,N_4625,N_4614);
nand U4770 (N_4770,N_4623,N_4656);
nor U4771 (N_4771,N_4699,N_4601);
or U4772 (N_4772,N_4685,N_4651);
or U4773 (N_4773,N_4665,N_4623);
or U4774 (N_4774,N_4614,N_4676);
nor U4775 (N_4775,N_4693,N_4647);
xor U4776 (N_4776,N_4614,N_4689);
or U4777 (N_4777,N_4608,N_4625);
nor U4778 (N_4778,N_4686,N_4654);
nor U4779 (N_4779,N_4662,N_4629);
nand U4780 (N_4780,N_4608,N_4691);
or U4781 (N_4781,N_4635,N_4669);
or U4782 (N_4782,N_4642,N_4634);
nor U4783 (N_4783,N_4621,N_4617);
and U4784 (N_4784,N_4625,N_4681);
xor U4785 (N_4785,N_4601,N_4671);
or U4786 (N_4786,N_4687,N_4668);
nand U4787 (N_4787,N_4664,N_4622);
nand U4788 (N_4788,N_4650,N_4646);
nand U4789 (N_4789,N_4644,N_4681);
and U4790 (N_4790,N_4640,N_4699);
and U4791 (N_4791,N_4684,N_4694);
or U4792 (N_4792,N_4632,N_4626);
xnor U4793 (N_4793,N_4607,N_4651);
xor U4794 (N_4794,N_4686,N_4641);
xor U4795 (N_4795,N_4649,N_4619);
nand U4796 (N_4796,N_4606,N_4605);
nor U4797 (N_4797,N_4643,N_4623);
nor U4798 (N_4798,N_4629,N_4633);
nor U4799 (N_4799,N_4631,N_4609);
nand U4800 (N_4800,N_4776,N_4763);
and U4801 (N_4801,N_4795,N_4762);
nand U4802 (N_4802,N_4787,N_4773);
and U4803 (N_4803,N_4724,N_4738);
or U4804 (N_4804,N_4735,N_4718);
nand U4805 (N_4805,N_4717,N_4708);
and U4806 (N_4806,N_4769,N_4722);
nor U4807 (N_4807,N_4714,N_4719);
nand U4808 (N_4808,N_4755,N_4706);
xnor U4809 (N_4809,N_4732,N_4752);
or U4810 (N_4810,N_4729,N_4782);
nor U4811 (N_4811,N_4705,N_4734);
xnor U4812 (N_4812,N_4702,N_4785);
nand U4813 (N_4813,N_4778,N_4771);
xnor U4814 (N_4814,N_4737,N_4703);
or U4815 (N_4815,N_4767,N_4748);
or U4816 (N_4816,N_4749,N_4726);
xor U4817 (N_4817,N_4790,N_4794);
xnor U4818 (N_4818,N_4730,N_4704);
or U4819 (N_4819,N_4774,N_4789);
nor U4820 (N_4820,N_4770,N_4709);
and U4821 (N_4821,N_4742,N_4798);
or U4822 (N_4822,N_4700,N_4751);
xnor U4823 (N_4823,N_4759,N_4747);
nand U4824 (N_4824,N_4739,N_4736);
nor U4825 (N_4825,N_4710,N_4757);
or U4826 (N_4826,N_4741,N_4746);
nor U4827 (N_4827,N_4723,N_4733);
and U4828 (N_4828,N_4791,N_4701);
xor U4829 (N_4829,N_4780,N_4799);
xor U4830 (N_4830,N_4797,N_4766);
xor U4831 (N_4831,N_4753,N_4792);
nor U4832 (N_4832,N_4775,N_4758);
nor U4833 (N_4833,N_4764,N_4750);
or U4834 (N_4834,N_4743,N_4772);
and U4835 (N_4835,N_4712,N_4779);
xor U4836 (N_4836,N_4728,N_4756);
or U4837 (N_4837,N_4796,N_4754);
and U4838 (N_4838,N_4784,N_4727);
nor U4839 (N_4839,N_4715,N_4786);
nor U4840 (N_4840,N_4777,N_4711);
xnor U4841 (N_4841,N_4793,N_4761);
nand U4842 (N_4842,N_4765,N_4707);
and U4843 (N_4843,N_4783,N_4721);
nand U4844 (N_4844,N_4788,N_4781);
nor U4845 (N_4845,N_4745,N_4725);
and U4846 (N_4846,N_4744,N_4768);
or U4847 (N_4847,N_4713,N_4716);
or U4848 (N_4848,N_4760,N_4731);
or U4849 (N_4849,N_4740,N_4720);
nand U4850 (N_4850,N_4701,N_4751);
xnor U4851 (N_4851,N_4722,N_4707);
xor U4852 (N_4852,N_4784,N_4711);
nor U4853 (N_4853,N_4775,N_4703);
xor U4854 (N_4854,N_4784,N_4796);
or U4855 (N_4855,N_4769,N_4785);
xnor U4856 (N_4856,N_4727,N_4717);
nor U4857 (N_4857,N_4772,N_4735);
nor U4858 (N_4858,N_4762,N_4769);
or U4859 (N_4859,N_4793,N_4715);
nor U4860 (N_4860,N_4761,N_4792);
nor U4861 (N_4861,N_4786,N_4783);
nor U4862 (N_4862,N_4712,N_4781);
nor U4863 (N_4863,N_4709,N_4728);
xnor U4864 (N_4864,N_4787,N_4742);
nand U4865 (N_4865,N_4756,N_4772);
nand U4866 (N_4866,N_4712,N_4730);
and U4867 (N_4867,N_4759,N_4703);
nor U4868 (N_4868,N_4714,N_4727);
nor U4869 (N_4869,N_4787,N_4729);
nand U4870 (N_4870,N_4701,N_4797);
xnor U4871 (N_4871,N_4701,N_4798);
or U4872 (N_4872,N_4733,N_4762);
nor U4873 (N_4873,N_4745,N_4751);
nand U4874 (N_4874,N_4736,N_4771);
or U4875 (N_4875,N_4723,N_4707);
xnor U4876 (N_4876,N_4746,N_4712);
or U4877 (N_4877,N_4784,N_4708);
and U4878 (N_4878,N_4722,N_4799);
or U4879 (N_4879,N_4798,N_4739);
and U4880 (N_4880,N_4790,N_4735);
and U4881 (N_4881,N_4796,N_4733);
or U4882 (N_4882,N_4735,N_4788);
xor U4883 (N_4883,N_4763,N_4730);
nor U4884 (N_4884,N_4787,N_4765);
xnor U4885 (N_4885,N_4706,N_4773);
xnor U4886 (N_4886,N_4787,N_4751);
and U4887 (N_4887,N_4763,N_4705);
nor U4888 (N_4888,N_4731,N_4785);
nor U4889 (N_4889,N_4764,N_4732);
or U4890 (N_4890,N_4707,N_4755);
nand U4891 (N_4891,N_4720,N_4705);
xnor U4892 (N_4892,N_4765,N_4788);
nor U4893 (N_4893,N_4754,N_4741);
nand U4894 (N_4894,N_4733,N_4716);
nand U4895 (N_4895,N_4749,N_4776);
xor U4896 (N_4896,N_4786,N_4769);
and U4897 (N_4897,N_4765,N_4726);
nor U4898 (N_4898,N_4748,N_4711);
nor U4899 (N_4899,N_4772,N_4713);
and U4900 (N_4900,N_4818,N_4831);
nand U4901 (N_4901,N_4853,N_4866);
xnor U4902 (N_4902,N_4800,N_4841);
nor U4903 (N_4903,N_4809,N_4858);
nor U4904 (N_4904,N_4806,N_4870);
nand U4905 (N_4905,N_4843,N_4896);
and U4906 (N_4906,N_4852,N_4857);
nand U4907 (N_4907,N_4836,N_4885);
nor U4908 (N_4908,N_4849,N_4862);
nand U4909 (N_4909,N_4838,N_4807);
xor U4910 (N_4910,N_4863,N_4815);
and U4911 (N_4911,N_4868,N_4899);
and U4912 (N_4912,N_4802,N_4822);
xor U4913 (N_4913,N_4842,N_4840);
nand U4914 (N_4914,N_4829,N_4875);
nand U4915 (N_4915,N_4869,N_4883);
or U4916 (N_4916,N_4887,N_4828);
nand U4917 (N_4917,N_4861,N_4879);
and U4918 (N_4918,N_4882,N_4808);
and U4919 (N_4919,N_4894,N_4845);
and U4920 (N_4920,N_4873,N_4837);
or U4921 (N_4921,N_4881,N_4892);
nor U4922 (N_4922,N_4859,N_4893);
nor U4923 (N_4923,N_4889,N_4803);
and U4924 (N_4924,N_4827,N_4805);
xnor U4925 (N_4925,N_4874,N_4884);
nand U4926 (N_4926,N_4891,N_4865);
and U4927 (N_4927,N_4816,N_4804);
nand U4928 (N_4928,N_4830,N_4819);
and U4929 (N_4929,N_4851,N_4832);
xor U4930 (N_4930,N_4820,N_4878);
and U4931 (N_4931,N_4847,N_4897);
and U4932 (N_4932,N_4864,N_4880);
xor U4933 (N_4933,N_4821,N_4826);
or U4934 (N_4934,N_4890,N_4833);
or U4935 (N_4935,N_4898,N_4813);
nand U4936 (N_4936,N_4854,N_4834);
xor U4937 (N_4937,N_4824,N_4846);
xnor U4938 (N_4938,N_4855,N_4812);
nand U4939 (N_4939,N_4817,N_4850);
nand U4940 (N_4940,N_4876,N_4801);
nor U4941 (N_4941,N_4860,N_4895);
or U4942 (N_4942,N_4871,N_4877);
and U4943 (N_4943,N_4844,N_4867);
xnor U4944 (N_4944,N_4839,N_4848);
xnor U4945 (N_4945,N_4888,N_4825);
xnor U4946 (N_4946,N_4886,N_4835);
xnor U4947 (N_4947,N_4872,N_4823);
nor U4948 (N_4948,N_4810,N_4814);
nor U4949 (N_4949,N_4811,N_4856);
and U4950 (N_4950,N_4894,N_4832);
nand U4951 (N_4951,N_4862,N_4853);
and U4952 (N_4952,N_4849,N_4851);
nor U4953 (N_4953,N_4836,N_4859);
or U4954 (N_4954,N_4811,N_4807);
nor U4955 (N_4955,N_4873,N_4890);
xnor U4956 (N_4956,N_4881,N_4813);
nand U4957 (N_4957,N_4811,N_4828);
xor U4958 (N_4958,N_4885,N_4841);
and U4959 (N_4959,N_4846,N_4814);
nor U4960 (N_4960,N_4838,N_4850);
and U4961 (N_4961,N_4853,N_4898);
nand U4962 (N_4962,N_4896,N_4829);
nor U4963 (N_4963,N_4855,N_4886);
xnor U4964 (N_4964,N_4823,N_4835);
nor U4965 (N_4965,N_4888,N_4805);
or U4966 (N_4966,N_4805,N_4842);
nand U4967 (N_4967,N_4866,N_4832);
nor U4968 (N_4968,N_4836,N_4889);
nor U4969 (N_4969,N_4818,N_4883);
xor U4970 (N_4970,N_4835,N_4859);
xor U4971 (N_4971,N_4806,N_4818);
or U4972 (N_4972,N_4856,N_4880);
nor U4973 (N_4973,N_4837,N_4808);
or U4974 (N_4974,N_4888,N_4868);
xnor U4975 (N_4975,N_4869,N_4855);
and U4976 (N_4976,N_4827,N_4866);
nand U4977 (N_4977,N_4852,N_4886);
nor U4978 (N_4978,N_4809,N_4825);
or U4979 (N_4979,N_4849,N_4829);
xor U4980 (N_4980,N_4850,N_4824);
and U4981 (N_4981,N_4845,N_4885);
and U4982 (N_4982,N_4861,N_4899);
xnor U4983 (N_4983,N_4865,N_4889);
nand U4984 (N_4984,N_4846,N_4875);
and U4985 (N_4985,N_4828,N_4872);
nand U4986 (N_4986,N_4898,N_4891);
nor U4987 (N_4987,N_4827,N_4842);
nor U4988 (N_4988,N_4886,N_4859);
nor U4989 (N_4989,N_4888,N_4897);
or U4990 (N_4990,N_4840,N_4848);
nor U4991 (N_4991,N_4879,N_4871);
nor U4992 (N_4992,N_4836,N_4814);
nand U4993 (N_4993,N_4887,N_4863);
nand U4994 (N_4994,N_4816,N_4878);
or U4995 (N_4995,N_4857,N_4873);
nand U4996 (N_4996,N_4858,N_4815);
xnor U4997 (N_4997,N_4883,N_4820);
xor U4998 (N_4998,N_4880,N_4884);
xor U4999 (N_4999,N_4815,N_4896);
or UO_0 (O_0,N_4982,N_4986);
nor UO_1 (O_1,N_4959,N_4938);
nand UO_2 (O_2,N_4958,N_4978);
xor UO_3 (O_3,N_4931,N_4924);
nand UO_4 (O_4,N_4972,N_4969);
nor UO_5 (O_5,N_4943,N_4964);
nor UO_6 (O_6,N_4976,N_4920);
nor UO_7 (O_7,N_4928,N_4904);
nor UO_8 (O_8,N_4905,N_4935);
xor UO_9 (O_9,N_4990,N_4911);
nand UO_10 (O_10,N_4917,N_4902);
nor UO_11 (O_11,N_4901,N_4979);
or UO_12 (O_12,N_4965,N_4949);
xor UO_13 (O_13,N_4908,N_4974);
nor UO_14 (O_14,N_4910,N_4980);
or UO_15 (O_15,N_4988,N_4983);
or UO_16 (O_16,N_4925,N_4952);
nor UO_17 (O_17,N_4916,N_4984);
and UO_18 (O_18,N_4957,N_4973);
xor UO_19 (O_19,N_4921,N_4947);
nand UO_20 (O_20,N_4971,N_4926);
nand UO_21 (O_21,N_4975,N_4927);
xor UO_22 (O_22,N_4946,N_4906);
nor UO_23 (O_23,N_4989,N_4951);
nand UO_24 (O_24,N_4950,N_4941);
nand UO_25 (O_25,N_4963,N_4914);
nand UO_26 (O_26,N_4934,N_4942);
xor UO_27 (O_27,N_4987,N_4915);
nand UO_28 (O_28,N_4944,N_4977);
and UO_29 (O_29,N_4903,N_4907);
nand UO_30 (O_30,N_4936,N_4918);
and UO_31 (O_31,N_4998,N_4997);
and UO_32 (O_32,N_4996,N_4991);
or UO_33 (O_33,N_4961,N_4930);
xor UO_34 (O_34,N_4970,N_4900);
xnor UO_35 (O_35,N_4999,N_4919);
xor UO_36 (O_36,N_4985,N_4995);
nand UO_37 (O_37,N_4966,N_4933);
nor UO_38 (O_38,N_4994,N_4981);
nand UO_39 (O_39,N_4960,N_4953);
and UO_40 (O_40,N_4948,N_4923);
nor UO_41 (O_41,N_4939,N_4962);
nor UO_42 (O_42,N_4932,N_4945);
or UO_43 (O_43,N_4967,N_4929);
or UO_44 (O_44,N_4912,N_4940);
or UO_45 (O_45,N_4968,N_4909);
and UO_46 (O_46,N_4955,N_4992);
or UO_47 (O_47,N_4937,N_4922);
nor UO_48 (O_48,N_4956,N_4993);
xnor UO_49 (O_49,N_4913,N_4954);
and UO_50 (O_50,N_4933,N_4946);
and UO_51 (O_51,N_4900,N_4993);
or UO_52 (O_52,N_4940,N_4928);
nand UO_53 (O_53,N_4924,N_4959);
nor UO_54 (O_54,N_4917,N_4922);
or UO_55 (O_55,N_4916,N_4955);
nand UO_56 (O_56,N_4994,N_4997);
nor UO_57 (O_57,N_4939,N_4938);
or UO_58 (O_58,N_4938,N_4954);
nand UO_59 (O_59,N_4921,N_4992);
and UO_60 (O_60,N_4908,N_4976);
and UO_61 (O_61,N_4987,N_4964);
xnor UO_62 (O_62,N_4950,N_4946);
and UO_63 (O_63,N_4919,N_4960);
or UO_64 (O_64,N_4945,N_4969);
or UO_65 (O_65,N_4916,N_4921);
nand UO_66 (O_66,N_4942,N_4981);
nand UO_67 (O_67,N_4966,N_4943);
xnor UO_68 (O_68,N_4947,N_4974);
or UO_69 (O_69,N_4922,N_4984);
nor UO_70 (O_70,N_4971,N_4900);
xor UO_71 (O_71,N_4966,N_4999);
xnor UO_72 (O_72,N_4956,N_4978);
nand UO_73 (O_73,N_4910,N_4940);
xnor UO_74 (O_74,N_4941,N_4943);
and UO_75 (O_75,N_4972,N_4927);
or UO_76 (O_76,N_4997,N_4966);
nand UO_77 (O_77,N_4949,N_4902);
nand UO_78 (O_78,N_4956,N_4974);
xnor UO_79 (O_79,N_4993,N_4951);
or UO_80 (O_80,N_4969,N_4988);
nor UO_81 (O_81,N_4908,N_4903);
and UO_82 (O_82,N_4923,N_4907);
nor UO_83 (O_83,N_4904,N_4906);
and UO_84 (O_84,N_4937,N_4917);
xnor UO_85 (O_85,N_4950,N_4940);
xor UO_86 (O_86,N_4944,N_4914);
or UO_87 (O_87,N_4988,N_4929);
nor UO_88 (O_88,N_4982,N_4910);
nor UO_89 (O_89,N_4959,N_4905);
nor UO_90 (O_90,N_4948,N_4918);
and UO_91 (O_91,N_4904,N_4939);
or UO_92 (O_92,N_4923,N_4911);
and UO_93 (O_93,N_4979,N_4954);
or UO_94 (O_94,N_4945,N_4952);
nand UO_95 (O_95,N_4971,N_4984);
xor UO_96 (O_96,N_4964,N_4975);
and UO_97 (O_97,N_4967,N_4931);
and UO_98 (O_98,N_4995,N_4951);
nand UO_99 (O_99,N_4975,N_4953);
xnor UO_100 (O_100,N_4932,N_4938);
and UO_101 (O_101,N_4937,N_4900);
and UO_102 (O_102,N_4905,N_4963);
or UO_103 (O_103,N_4926,N_4912);
and UO_104 (O_104,N_4907,N_4912);
xnor UO_105 (O_105,N_4957,N_4962);
xnor UO_106 (O_106,N_4957,N_4907);
or UO_107 (O_107,N_4931,N_4905);
xor UO_108 (O_108,N_4956,N_4905);
nand UO_109 (O_109,N_4946,N_4928);
nor UO_110 (O_110,N_4905,N_4934);
nand UO_111 (O_111,N_4914,N_4945);
nor UO_112 (O_112,N_4981,N_4965);
xor UO_113 (O_113,N_4921,N_4983);
or UO_114 (O_114,N_4911,N_4940);
xor UO_115 (O_115,N_4992,N_4904);
nand UO_116 (O_116,N_4904,N_4977);
and UO_117 (O_117,N_4985,N_4934);
nor UO_118 (O_118,N_4987,N_4918);
nor UO_119 (O_119,N_4980,N_4979);
or UO_120 (O_120,N_4980,N_4904);
or UO_121 (O_121,N_4937,N_4988);
xor UO_122 (O_122,N_4909,N_4932);
or UO_123 (O_123,N_4961,N_4926);
nor UO_124 (O_124,N_4920,N_4903);
or UO_125 (O_125,N_4944,N_4940);
nor UO_126 (O_126,N_4992,N_4906);
nand UO_127 (O_127,N_4960,N_4984);
xnor UO_128 (O_128,N_4945,N_4954);
or UO_129 (O_129,N_4970,N_4957);
and UO_130 (O_130,N_4935,N_4924);
nor UO_131 (O_131,N_4994,N_4968);
and UO_132 (O_132,N_4992,N_4928);
xnor UO_133 (O_133,N_4997,N_4951);
and UO_134 (O_134,N_4973,N_4996);
nor UO_135 (O_135,N_4963,N_4933);
xnor UO_136 (O_136,N_4926,N_4957);
nand UO_137 (O_137,N_4982,N_4919);
nand UO_138 (O_138,N_4977,N_4946);
nor UO_139 (O_139,N_4935,N_4915);
or UO_140 (O_140,N_4933,N_4919);
or UO_141 (O_141,N_4998,N_4936);
nor UO_142 (O_142,N_4950,N_4969);
xor UO_143 (O_143,N_4922,N_4934);
or UO_144 (O_144,N_4922,N_4956);
nor UO_145 (O_145,N_4982,N_4901);
and UO_146 (O_146,N_4939,N_4965);
xnor UO_147 (O_147,N_4911,N_4944);
nand UO_148 (O_148,N_4967,N_4973);
xnor UO_149 (O_149,N_4991,N_4937);
nor UO_150 (O_150,N_4991,N_4903);
xnor UO_151 (O_151,N_4970,N_4916);
or UO_152 (O_152,N_4972,N_4989);
or UO_153 (O_153,N_4930,N_4932);
and UO_154 (O_154,N_4931,N_4936);
or UO_155 (O_155,N_4949,N_4995);
nor UO_156 (O_156,N_4999,N_4906);
or UO_157 (O_157,N_4960,N_4935);
nand UO_158 (O_158,N_4968,N_4950);
xnor UO_159 (O_159,N_4961,N_4998);
or UO_160 (O_160,N_4948,N_4977);
nand UO_161 (O_161,N_4926,N_4915);
nor UO_162 (O_162,N_4928,N_4903);
nor UO_163 (O_163,N_4921,N_4953);
and UO_164 (O_164,N_4968,N_4978);
or UO_165 (O_165,N_4926,N_4976);
and UO_166 (O_166,N_4991,N_4905);
xor UO_167 (O_167,N_4990,N_4956);
nor UO_168 (O_168,N_4969,N_4983);
nand UO_169 (O_169,N_4903,N_4995);
nand UO_170 (O_170,N_4934,N_4926);
and UO_171 (O_171,N_4992,N_4967);
nand UO_172 (O_172,N_4957,N_4909);
nand UO_173 (O_173,N_4939,N_4934);
nor UO_174 (O_174,N_4913,N_4996);
or UO_175 (O_175,N_4995,N_4988);
xnor UO_176 (O_176,N_4987,N_4997);
and UO_177 (O_177,N_4977,N_4921);
xnor UO_178 (O_178,N_4991,N_4941);
or UO_179 (O_179,N_4949,N_4952);
xnor UO_180 (O_180,N_4906,N_4976);
nor UO_181 (O_181,N_4924,N_4933);
xnor UO_182 (O_182,N_4926,N_4972);
and UO_183 (O_183,N_4978,N_4910);
xor UO_184 (O_184,N_4958,N_4913);
nand UO_185 (O_185,N_4978,N_4988);
xnor UO_186 (O_186,N_4945,N_4917);
nor UO_187 (O_187,N_4946,N_4966);
nor UO_188 (O_188,N_4971,N_4979);
nor UO_189 (O_189,N_4911,N_4946);
and UO_190 (O_190,N_4951,N_4980);
nand UO_191 (O_191,N_4947,N_4946);
or UO_192 (O_192,N_4928,N_4966);
nand UO_193 (O_193,N_4960,N_4921);
xnor UO_194 (O_194,N_4958,N_4919);
and UO_195 (O_195,N_4928,N_4997);
and UO_196 (O_196,N_4918,N_4940);
xor UO_197 (O_197,N_4937,N_4956);
xnor UO_198 (O_198,N_4973,N_4932);
nand UO_199 (O_199,N_4973,N_4940);
and UO_200 (O_200,N_4949,N_4940);
and UO_201 (O_201,N_4949,N_4937);
or UO_202 (O_202,N_4994,N_4962);
or UO_203 (O_203,N_4989,N_4925);
nand UO_204 (O_204,N_4979,N_4976);
or UO_205 (O_205,N_4926,N_4997);
nand UO_206 (O_206,N_4985,N_4958);
xor UO_207 (O_207,N_4953,N_4998);
nor UO_208 (O_208,N_4923,N_4941);
and UO_209 (O_209,N_4976,N_4916);
xor UO_210 (O_210,N_4931,N_4950);
xor UO_211 (O_211,N_4932,N_4982);
nor UO_212 (O_212,N_4972,N_4965);
xor UO_213 (O_213,N_4960,N_4979);
or UO_214 (O_214,N_4983,N_4992);
xnor UO_215 (O_215,N_4953,N_4969);
xor UO_216 (O_216,N_4935,N_4929);
nor UO_217 (O_217,N_4952,N_4921);
or UO_218 (O_218,N_4990,N_4997);
and UO_219 (O_219,N_4933,N_4938);
nand UO_220 (O_220,N_4995,N_4996);
or UO_221 (O_221,N_4918,N_4950);
or UO_222 (O_222,N_4997,N_4947);
nor UO_223 (O_223,N_4958,N_4982);
and UO_224 (O_224,N_4979,N_4992);
or UO_225 (O_225,N_4971,N_4976);
and UO_226 (O_226,N_4941,N_4933);
or UO_227 (O_227,N_4975,N_4935);
nand UO_228 (O_228,N_4907,N_4979);
nand UO_229 (O_229,N_4905,N_4971);
nand UO_230 (O_230,N_4966,N_4907);
or UO_231 (O_231,N_4956,N_4945);
or UO_232 (O_232,N_4919,N_4942);
xnor UO_233 (O_233,N_4961,N_4907);
or UO_234 (O_234,N_4900,N_4948);
nand UO_235 (O_235,N_4994,N_4973);
or UO_236 (O_236,N_4913,N_4940);
xor UO_237 (O_237,N_4982,N_4917);
nand UO_238 (O_238,N_4925,N_4931);
xor UO_239 (O_239,N_4915,N_4914);
xor UO_240 (O_240,N_4929,N_4970);
and UO_241 (O_241,N_4915,N_4974);
and UO_242 (O_242,N_4964,N_4950);
and UO_243 (O_243,N_4915,N_4977);
and UO_244 (O_244,N_4930,N_4966);
xnor UO_245 (O_245,N_4902,N_4972);
and UO_246 (O_246,N_4997,N_4989);
nand UO_247 (O_247,N_4932,N_4924);
and UO_248 (O_248,N_4995,N_4994);
and UO_249 (O_249,N_4995,N_4939);
or UO_250 (O_250,N_4990,N_4945);
xor UO_251 (O_251,N_4931,N_4992);
and UO_252 (O_252,N_4964,N_4973);
and UO_253 (O_253,N_4987,N_4961);
and UO_254 (O_254,N_4934,N_4962);
nand UO_255 (O_255,N_4995,N_4947);
or UO_256 (O_256,N_4919,N_4996);
or UO_257 (O_257,N_4926,N_4918);
xnor UO_258 (O_258,N_4933,N_4983);
and UO_259 (O_259,N_4934,N_4965);
and UO_260 (O_260,N_4970,N_4953);
or UO_261 (O_261,N_4919,N_4988);
nor UO_262 (O_262,N_4912,N_4991);
xnor UO_263 (O_263,N_4960,N_4934);
nand UO_264 (O_264,N_4921,N_4924);
or UO_265 (O_265,N_4969,N_4986);
or UO_266 (O_266,N_4960,N_4988);
nand UO_267 (O_267,N_4927,N_4924);
nor UO_268 (O_268,N_4900,N_4962);
xor UO_269 (O_269,N_4957,N_4940);
or UO_270 (O_270,N_4998,N_4938);
nand UO_271 (O_271,N_4968,N_4951);
nand UO_272 (O_272,N_4909,N_4921);
nand UO_273 (O_273,N_4967,N_4982);
or UO_274 (O_274,N_4991,N_4904);
nor UO_275 (O_275,N_4999,N_4984);
xor UO_276 (O_276,N_4926,N_4927);
or UO_277 (O_277,N_4980,N_4989);
nor UO_278 (O_278,N_4945,N_4999);
nor UO_279 (O_279,N_4980,N_4948);
xor UO_280 (O_280,N_4900,N_4973);
or UO_281 (O_281,N_4909,N_4920);
and UO_282 (O_282,N_4970,N_4974);
and UO_283 (O_283,N_4933,N_4943);
or UO_284 (O_284,N_4938,N_4912);
xor UO_285 (O_285,N_4901,N_4927);
or UO_286 (O_286,N_4919,N_4925);
nand UO_287 (O_287,N_4986,N_4925);
nor UO_288 (O_288,N_4970,N_4996);
xor UO_289 (O_289,N_4984,N_4924);
nor UO_290 (O_290,N_4991,N_4949);
nor UO_291 (O_291,N_4935,N_4936);
nor UO_292 (O_292,N_4921,N_4942);
or UO_293 (O_293,N_4931,N_4984);
nor UO_294 (O_294,N_4994,N_4939);
xor UO_295 (O_295,N_4943,N_4945);
xnor UO_296 (O_296,N_4925,N_4901);
and UO_297 (O_297,N_4950,N_4938);
or UO_298 (O_298,N_4949,N_4903);
xnor UO_299 (O_299,N_4946,N_4959);
nand UO_300 (O_300,N_4977,N_4947);
nand UO_301 (O_301,N_4956,N_4985);
nand UO_302 (O_302,N_4946,N_4914);
or UO_303 (O_303,N_4943,N_4965);
nand UO_304 (O_304,N_4950,N_4943);
or UO_305 (O_305,N_4902,N_4960);
and UO_306 (O_306,N_4991,N_4957);
and UO_307 (O_307,N_4905,N_4909);
xnor UO_308 (O_308,N_4961,N_4984);
nand UO_309 (O_309,N_4944,N_4950);
xnor UO_310 (O_310,N_4913,N_4915);
xor UO_311 (O_311,N_4978,N_4902);
nand UO_312 (O_312,N_4990,N_4920);
nor UO_313 (O_313,N_4959,N_4902);
nor UO_314 (O_314,N_4940,N_4948);
nor UO_315 (O_315,N_4928,N_4988);
or UO_316 (O_316,N_4961,N_4995);
nand UO_317 (O_317,N_4959,N_4954);
nand UO_318 (O_318,N_4947,N_4954);
nand UO_319 (O_319,N_4931,N_4954);
xor UO_320 (O_320,N_4965,N_4994);
nand UO_321 (O_321,N_4976,N_4917);
xnor UO_322 (O_322,N_4921,N_4978);
or UO_323 (O_323,N_4980,N_4970);
nor UO_324 (O_324,N_4955,N_4960);
and UO_325 (O_325,N_4964,N_4977);
xor UO_326 (O_326,N_4963,N_4917);
nand UO_327 (O_327,N_4925,N_4963);
nor UO_328 (O_328,N_4993,N_4990);
xnor UO_329 (O_329,N_4915,N_4958);
or UO_330 (O_330,N_4938,N_4997);
and UO_331 (O_331,N_4900,N_4953);
and UO_332 (O_332,N_4998,N_4930);
nand UO_333 (O_333,N_4954,N_4928);
nor UO_334 (O_334,N_4929,N_4985);
nor UO_335 (O_335,N_4946,N_4903);
xor UO_336 (O_336,N_4969,N_4940);
xnor UO_337 (O_337,N_4926,N_4980);
nand UO_338 (O_338,N_4948,N_4905);
and UO_339 (O_339,N_4962,N_4963);
nand UO_340 (O_340,N_4918,N_4977);
nor UO_341 (O_341,N_4918,N_4941);
nand UO_342 (O_342,N_4908,N_4951);
or UO_343 (O_343,N_4940,N_4934);
and UO_344 (O_344,N_4937,N_4942);
or UO_345 (O_345,N_4909,N_4987);
xnor UO_346 (O_346,N_4975,N_4976);
xor UO_347 (O_347,N_4943,N_4984);
and UO_348 (O_348,N_4949,N_4918);
xor UO_349 (O_349,N_4901,N_4967);
nand UO_350 (O_350,N_4978,N_4949);
and UO_351 (O_351,N_4962,N_4983);
and UO_352 (O_352,N_4951,N_4913);
or UO_353 (O_353,N_4996,N_4961);
or UO_354 (O_354,N_4918,N_4956);
nor UO_355 (O_355,N_4991,N_4952);
nand UO_356 (O_356,N_4911,N_4915);
and UO_357 (O_357,N_4940,N_4970);
nand UO_358 (O_358,N_4974,N_4919);
nand UO_359 (O_359,N_4974,N_4948);
and UO_360 (O_360,N_4942,N_4954);
or UO_361 (O_361,N_4914,N_4982);
nor UO_362 (O_362,N_4922,N_4977);
nor UO_363 (O_363,N_4945,N_4931);
nor UO_364 (O_364,N_4998,N_4939);
or UO_365 (O_365,N_4955,N_4994);
nand UO_366 (O_366,N_4908,N_4940);
xor UO_367 (O_367,N_4916,N_4979);
nand UO_368 (O_368,N_4942,N_4932);
nor UO_369 (O_369,N_4962,N_4975);
or UO_370 (O_370,N_4905,N_4947);
or UO_371 (O_371,N_4968,N_4941);
or UO_372 (O_372,N_4997,N_4996);
and UO_373 (O_373,N_4989,N_4943);
and UO_374 (O_374,N_4975,N_4998);
nand UO_375 (O_375,N_4904,N_4998);
and UO_376 (O_376,N_4984,N_4981);
nand UO_377 (O_377,N_4907,N_4978);
nor UO_378 (O_378,N_4939,N_4996);
nand UO_379 (O_379,N_4953,N_4974);
or UO_380 (O_380,N_4939,N_4912);
or UO_381 (O_381,N_4973,N_4917);
nor UO_382 (O_382,N_4974,N_4927);
nor UO_383 (O_383,N_4900,N_4940);
nor UO_384 (O_384,N_4995,N_4942);
nand UO_385 (O_385,N_4929,N_4977);
nor UO_386 (O_386,N_4985,N_4967);
and UO_387 (O_387,N_4959,N_4989);
nand UO_388 (O_388,N_4914,N_4902);
and UO_389 (O_389,N_4909,N_4989);
or UO_390 (O_390,N_4908,N_4929);
nand UO_391 (O_391,N_4904,N_4935);
and UO_392 (O_392,N_4971,N_4903);
or UO_393 (O_393,N_4928,N_4980);
xor UO_394 (O_394,N_4986,N_4941);
and UO_395 (O_395,N_4915,N_4973);
nor UO_396 (O_396,N_4964,N_4904);
nand UO_397 (O_397,N_4980,N_4988);
nand UO_398 (O_398,N_4962,N_4973);
nand UO_399 (O_399,N_4993,N_4927);
nor UO_400 (O_400,N_4941,N_4936);
and UO_401 (O_401,N_4918,N_4931);
and UO_402 (O_402,N_4917,N_4997);
and UO_403 (O_403,N_4945,N_4979);
nor UO_404 (O_404,N_4987,N_4982);
xor UO_405 (O_405,N_4990,N_4972);
xor UO_406 (O_406,N_4906,N_4927);
nor UO_407 (O_407,N_4916,N_4988);
and UO_408 (O_408,N_4963,N_4980);
nand UO_409 (O_409,N_4909,N_4967);
nor UO_410 (O_410,N_4982,N_4943);
or UO_411 (O_411,N_4931,N_4923);
and UO_412 (O_412,N_4978,N_4901);
nand UO_413 (O_413,N_4971,N_4930);
and UO_414 (O_414,N_4957,N_4922);
nand UO_415 (O_415,N_4909,N_4961);
or UO_416 (O_416,N_4970,N_4914);
xnor UO_417 (O_417,N_4996,N_4977);
xnor UO_418 (O_418,N_4969,N_4967);
nor UO_419 (O_419,N_4977,N_4998);
or UO_420 (O_420,N_4918,N_4933);
xnor UO_421 (O_421,N_4925,N_4993);
nand UO_422 (O_422,N_4966,N_4922);
xnor UO_423 (O_423,N_4906,N_4901);
and UO_424 (O_424,N_4905,N_4961);
xnor UO_425 (O_425,N_4933,N_4972);
or UO_426 (O_426,N_4973,N_4931);
nor UO_427 (O_427,N_4904,N_4927);
or UO_428 (O_428,N_4919,N_4948);
or UO_429 (O_429,N_4953,N_4950);
or UO_430 (O_430,N_4965,N_4992);
or UO_431 (O_431,N_4932,N_4996);
nor UO_432 (O_432,N_4925,N_4910);
xor UO_433 (O_433,N_4900,N_4987);
nand UO_434 (O_434,N_4999,N_4996);
and UO_435 (O_435,N_4957,N_4910);
nand UO_436 (O_436,N_4948,N_4960);
nor UO_437 (O_437,N_4965,N_4962);
or UO_438 (O_438,N_4911,N_4945);
or UO_439 (O_439,N_4906,N_4979);
and UO_440 (O_440,N_4941,N_4914);
or UO_441 (O_441,N_4926,N_4942);
and UO_442 (O_442,N_4993,N_4952);
and UO_443 (O_443,N_4994,N_4910);
or UO_444 (O_444,N_4950,N_4955);
and UO_445 (O_445,N_4906,N_4905);
and UO_446 (O_446,N_4986,N_4970);
nand UO_447 (O_447,N_4981,N_4932);
and UO_448 (O_448,N_4937,N_4952);
nor UO_449 (O_449,N_4961,N_4973);
and UO_450 (O_450,N_4994,N_4946);
or UO_451 (O_451,N_4973,N_4924);
and UO_452 (O_452,N_4934,N_4959);
xor UO_453 (O_453,N_4974,N_4935);
xor UO_454 (O_454,N_4938,N_4957);
xor UO_455 (O_455,N_4938,N_4926);
xnor UO_456 (O_456,N_4922,N_4981);
nand UO_457 (O_457,N_4911,N_4901);
nor UO_458 (O_458,N_4916,N_4941);
xnor UO_459 (O_459,N_4949,N_4910);
or UO_460 (O_460,N_4951,N_4966);
nor UO_461 (O_461,N_4997,N_4953);
nand UO_462 (O_462,N_4908,N_4969);
xnor UO_463 (O_463,N_4938,N_4961);
nor UO_464 (O_464,N_4962,N_4958);
nor UO_465 (O_465,N_4968,N_4903);
nand UO_466 (O_466,N_4937,N_4947);
xor UO_467 (O_467,N_4920,N_4963);
or UO_468 (O_468,N_4917,N_4920);
nand UO_469 (O_469,N_4929,N_4922);
nor UO_470 (O_470,N_4908,N_4924);
xnor UO_471 (O_471,N_4970,N_4903);
or UO_472 (O_472,N_4970,N_4948);
xor UO_473 (O_473,N_4929,N_4971);
nor UO_474 (O_474,N_4923,N_4963);
and UO_475 (O_475,N_4939,N_4935);
nor UO_476 (O_476,N_4977,N_4979);
and UO_477 (O_477,N_4944,N_4959);
nor UO_478 (O_478,N_4902,N_4927);
xor UO_479 (O_479,N_4967,N_4927);
xnor UO_480 (O_480,N_4964,N_4981);
nand UO_481 (O_481,N_4986,N_4922);
xor UO_482 (O_482,N_4975,N_4908);
or UO_483 (O_483,N_4987,N_4983);
nor UO_484 (O_484,N_4948,N_4952);
xnor UO_485 (O_485,N_4951,N_4900);
xor UO_486 (O_486,N_4926,N_4959);
xor UO_487 (O_487,N_4965,N_4951);
and UO_488 (O_488,N_4906,N_4912);
nand UO_489 (O_489,N_4945,N_4975);
and UO_490 (O_490,N_4945,N_4991);
nand UO_491 (O_491,N_4958,N_4960);
nand UO_492 (O_492,N_4917,N_4946);
nor UO_493 (O_493,N_4985,N_4989);
nand UO_494 (O_494,N_4946,N_4916);
and UO_495 (O_495,N_4936,N_4902);
or UO_496 (O_496,N_4910,N_4941);
or UO_497 (O_497,N_4981,N_4901);
xor UO_498 (O_498,N_4972,N_4940);
or UO_499 (O_499,N_4990,N_4917);
nand UO_500 (O_500,N_4987,N_4941);
nor UO_501 (O_501,N_4980,N_4915);
or UO_502 (O_502,N_4983,N_4970);
xnor UO_503 (O_503,N_4945,N_4960);
xor UO_504 (O_504,N_4907,N_4902);
and UO_505 (O_505,N_4996,N_4979);
or UO_506 (O_506,N_4992,N_4943);
or UO_507 (O_507,N_4900,N_4939);
and UO_508 (O_508,N_4986,N_4990);
xor UO_509 (O_509,N_4921,N_4966);
and UO_510 (O_510,N_4920,N_4997);
or UO_511 (O_511,N_4946,N_4973);
and UO_512 (O_512,N_4963,N_4977);
and UO_513 (O_513,N_4906,N_4953);
and UO_514 (O_514,N_4948,N_4929);
xor UO_515 (O_515,N_4969,N_4901);
nand UO_516 (O_516,N_4971,N_4912);
and UO_517 (O_517,N_4926,N_4958);
xor UO_518 (O_518,N_4908,N_4916);
xnor UO_519 (O_519,N_4972,N_4915);
xor UO_520 (O_520,N_4929,N_4914);
xnor UO_521 (O_521,N_4933,N_4950);
or UO_522 (O_522,N_4938,N_4931);
xnor UO_523 (O_523,N_4974,N_4946);
nand UO_524 (O_524,N_4991,N_4976);
nand UO_525 (O_525,N_4935,N_4940);
xor UO_526 (O_526,N_4903,N_4972);
nor UO_527 (O_527,N_4971,N_4923);
xnor UO_528 (O_528,N_4988,N_4963);
and UO_529 (O_529,N_4962,N_4921);
or UO_530 (O_530,N_4910,N_4943);
nand UO_531 (O_531,N_4973,N_4921);
nand UO_532 (O_532,N_4954,N_4901);
nand UO_533 (O_533,N_4910,N_4971);
or UO_534 (O_534,N_4973,N_4941);
xnor UO_535 (O_535,N_4963,N_4939);
or UO_536 (O_536,N_4908,N_4971);
nand UO_537 (O_537,N_4966,N_4959);
xnor UO_538 (O_538,N_4971,N_4941);
nor UO_539 (O_539,N_4930,N_4913);
nor UO_540 (O_540,N_4989,N_4913);
nand UO_541 (O_541,N_4994,N_4925);
and UO_542 (O_542,N_4930,N_4994);
xor UO_543 (O_543,N_4941,N_4924);
nor UO_544 (O_544,N_4967,N_4906);
and UO_545 (O_545,N_4990,N_4955);
and UO_546 (O_546,N_4997,N_4980);
nor UO_547 (O_547,N_4907,N_4960);
and UO_548 (O_548,N_4952,N_4917);
or UO_549 (O_549,N_4999,N_4907);
nand UO_550 (O_550,N_4915,N_4962);
and UO_551 (O_551,N_4964,N_4930);
xnor UO_552 (O_552,N_4971,N_4928);
nand UO_553 (O_553,N_4973,N_4947);
and UO_554 (O_554,N_4942,N_4952);
nor UO_555 (O_555,N_4909,N_4943);
xnor UO_556 (O_556,N_4940,N_4983);
nand UO_557 (O_557,N_4944,N_4986);
xnor UO_558 (O_558,N_4947,N_4922);
nand UO_559 (O_559,N_4956,N_4910);
nor UO_560 (O_560,N_4900,N_4991);
xnor UO_561 (O_561,N_4939,N_4975);
xnor UO_562 (O_562,N_4905,N_4936);
and UO_563 (O_563,N_4962,N_4904);
nand UO_564 (O_564,N_4949,N_4938);
and UO_565 (O_565,N_4930,N_4939);
xnor UO_566 (O_566,N_4984,N_4966);
and UO_567 (O_567,N_4972,N_4952);
nand UO_568 (O_568,N_4925,N_4996);
nand UO_569 (O_569,N_4945,N_4986);
nand UO_570 (O_570,N_4977,N_4909);
nor UO_571 (O_571,N_4904,N_4945);
and UO_572 (O_572,N_4916,N_4997);
or UO_573 (O_573,N_4980,N_4914);
nand UO_574 (O_574,N_4982,N_4931);
and UO_575 (O_575,N_4961,N_4914);
nand UO_576 (O_576,N_4947,N_4906);
xor UO_577 (O_577,N_4968,N_4986);
nor UO_578 (O_578,N_4901,N_4918);
xor UO_579 (O_579,N_4973,N_4922);
nand UO_580 (O_580,N_4925,N_4941);
and UO_581 (O_581,N_4994,N_4938);
xor UO_582 (O_582,N_4970,N_4973);
nor UO_583 (O_583,N_4932,N_4931);
nand UO_584 (O_584,N_4966,N_4977);
xnor UO_585 (O_585,N_4988,N_4902);
and UO_586 (O_586,N_4987,N_4974);
nand UO_587 (O_587,N_4960,N_4983);
or UO_588 (O_588,N_4998,N_4973);
nand UO_589 (O_589,N_4918,N_4994);
nand UO_590 (O_590,N_4936,N_4952);
and UO_591 (O_591,N_4933,N_4911);
nand UO_592 (O_592,N_4949,N_4928);
nor UO_593 (O_593,N_4977,N_4940);
or UO_594 (O_594,N_4985,N_4960);
xor UO_595 (O_595,N_4945,N_4934);
nand UO_596 (O_596,N_4988,N_4925);
or UO_597 (O_597,N_4991,N_4953);
nand UO_598 (O_598,N_4907,N_4975);
xor UO_599 (O_599,N_4937,N_4932);
xnor UO_600 (O_600,N_4987,N_4908);
xor UO_601 (O_601,N_4984,N_4968);
or UO_602 (O_602,N_4994,N_4970);
nand UO_603 (O_603,N_4957,N_4955);
nor UO_604 (O_604,N_4931,N_4920);
nand UO_605 (O_605,N_4941,N_4932);
nor UO_606 (O_606,N_4973,N_4968);
xor UO_607 (O_607,N_4913,N_4957);
xnor UO_608 (O_608,N_4946,N_4910);
nand UO_609 (O_609,N_4998,N_4944);
and UO_610 (O_610,N_4912,N_4958);
and UO_611 (O_611,N_4982,N_4909);
and UO_612 (O_612,N_4930,N_4963);
nor UO_613 (O_613,N_4910,N_4926);
or UO_614 (O_614,N_4998,N_4943);
xnor UO_615 (O_615,N_4960,N_4939);
and UO_616 (O_616,N_4925,N_4908);
xnor UO_617 (O_617,N_4929,N_4951);
xnor UO_618 (O_618,N_4936,N_4948);
nand UO_619 (O_619,N_4902,N_4948);
or UO_620 (O_620,N_4909,N_4911);
or UO_621 (O_621,N_4993,N_4959);
and UO_622 (O_622,N_4969,N_4971);
nor UO_623 (O_623,N_4968,N_4913);
and UO_624 (O_624,N_4963,N_4989);
xnor UO_625 (O_625,N_4991,N_4974);
and UO_626 (O_626,N_4958,N_4933);
xnor UO_627 (O_627,N_4947,N_4941);
or UO_628 (O_628,N_4931,N_4922);
xor UO_629 (O_629,N_4927,N_4951);
and UO_630 (O_630,N_4906,N_4998);
and UO_631 (O_631,N_4955,N_4956);
nand UO_632 (O_632,N_4931,N_4937);
nand UO_633 (O_633,N_4979,N_4925);
or UO_634 (O_634,N_4941,N_4915);
nor UO_635 (O_635,N_4932,N_4965);
xnor UO_636 (O_636,N_4921,N_4945);
nor UO_637 (O_637,N_4903,N_4957);
or UO_638 (O_638,N_4906,N_4932);
or UO_639 (O_639,N_4961,N_4985);
and UO_640 (O_640,N_4997,N_4942);
or UO_641 (O_641,N_4990,N_4981);
or UO_642 (O_642,N_4983,N_4953);
nor UO_643 (O_643,N_4982,N_4993);
nor UO_644 (O_644,N_4907,N_4993);
xor UO_645 (O_645,N_4984,N_4911);
or UO_646 (O_646,N_4966,N_4910);
xnor UO_647 (O_647,N_4906,N_4980);
nor UO_648 (O_648,N_4937,N_4957);
xor UO_649 (O_649,N_4980,N_4964);
nor UO_650 (O_650,N_4920,N_4916);
or UO_651 (O_651,N_4901,N_4961);
or UO_652 (O_652,N_4914,N_4906);
xor UO_653 (O_653,N_4921,N_4987);
or UO_654 (O_654,N_4910,N_4979);
nor UO_655 (O_655,N_4937,N_4905);
or UO_656 (O_656,N_4999,N_4982);
and UO_657 (O_657,N_4901,N_4929);
nor UO_658 (O_658,N_4974,N_4992);
xnor UO_659 (O_659,N_4919,N_4946);
nor UO_660 (O_660,N_4948,N_4913);
nor UO_661 (O_661,N_4983,N_4997);
and UO_662 (O_662,N_4946,N_4982);
nand UO_663 (O_663,N_4965,N_4923);
or UO_664 (O_664,N_4912,N_4966);
nor UO_665 (O_665,N_4904,N_4985);
or UO_666 (O_666,N_4912,N_4936);
or UO_667 (O_667,N_4928,N_4956);
or UO_668 (O_668,N_4922,N_4959);
or UO_669 (O_669,N_4998,N_4959);
or UO_670 (O_670,N_4950,N_4922);
and UO_671 (O_671,N_4923,N_4973);
or UO_672 (O_672,N_4900,N_4905);
nor UO_673 (O_673,N_4913,N_4999);
nor UO_674 (O_674,N_4911,N_4967);
or UO_675 (O_675,N_4933,N_4995);
nor UO_676 (O_676,N_4956,N_4976);
nand UO_677 (O_677,N_4943,N_4937);
or UO_678 (O_678,N_4956,N_4900);
or UO_679 (O_679,N_4912,N_4948);
and UO_680 (O_680,N_4983,N_4900);
nand UO_681 (O_681,N_4943,N_4952);
nand UO_682 (O_682,N_4942,N_4936);
nor UO_683 (O_683,N_4956,N_4968);
or UO_684 (O_684,N_4944,N_4941);
nor UO_685 (O_685,N_4983,N_4955);
nor UO_686 (O_686,N_4927,N_4986);
or UO_687 (O_687,N_4990,N_4969);
xnor UO_688 (O_688,N_4914,N_4950);
nor UO_689 (O_689,N_4916,N_4927);
nor UO_690 (O_690,N_4934,N_4938);
or UO_691 (O_691,N_4952,N_4928);
and UO_692 (O_692,N_4987,N_4954);
nand UO_693 (O_693,N_4941,N_4970);
and UO_694 (O_694,N_4967,N_4910);
xnor UO_695 (O_695,N_4981,N_4993);
and UO_696 (O_696,N_4979,N_4923);
xor UO_697 (O_697,N_4988,N_4936);
or UO_698 (O_698,N_4932,N_4913);
nand UO_699 (O_699,N_4938,N_4963);
xor UO_700 (O_700,N_4910,N_4928);
and UO_701 (O_701,N_4974,N_4981);
or UO_702 (O_702,N_4999,N_4998);
or UO_703 (O_703,N_4937,N_4910);
nand UO_704 (O_704,N_4919,N_4927);
nor UO_705 (O_705,N_4919,N_4944);
and UO_706 (O_706,N_4931,N_4935);
xnor UO_707 (O_707,N_4996,N_4968);
nand UO_708 (O_708,N_4960,N_4916);
nand UO_709 (O_709,N_4957,N_4998);
and UO_710 (O_710,N_4926,N_4932);
nand UO_711 (O_711,N_4960,N_4905);
or UO_712 (O_712,N_4948,N_4931);
xor UO_713 (O_713,N_4938,N_4979);
and UO_714 (O_714,N_4923,N_4901);
xnor UO_715 (O_715,N_4901,N_4965);
xnor UO_716 (O_716,N_4938,N_4917);
and UO_717 (O_717,N_4948,N_4971);
or UO_718 (O_718,N_4968,N_4958);
nand UO_719 (O_719,N_4979,N_4970);
or UO_720 (O_720,N_4981,N_4958);
nand UO_721 (O_721,N_4988,N_4967);
xnor UO_722 (O_722,N_4983,N_4999);
and UO_723 (O_723,N_4916,N_4934);
or UO_724 (O_724,N_4999,N_4997);
xor UO_725 (O_725,N_4900,N_4938);
xnor UO_726 (O_726,N_4913,N_4974);
xnor UO_727 (O_727,N_4941,N_4907);
xor UO_728 (O_728,N_4936,N_4913);
xnor UO_729 (O_729,N_4943,N_4931);
nand UO_730 (O_730,N_4986,N_4964);
nor UO_731 (O_731,N_4999,N_4921);
nand UO_732 (O_732,N_4964,N_4903);
nand UO_733 (O_733,N_4957,N_4999);
xor UO_734 (O_734,N_4956,N_4999);
or UO_735 (O_735,N_4999,N_4953);
xor UO_736 (O_736,N_4975,N_4952);
and UO_737 (O_737,N_4951,N_4932);
nand UO_738 (O_738,N_4998,N_4948);
or UO_739 (O_739,N_4987,N_4969);
and UO_740 (O_740,N_4952,N_4964);
nor UO_741 (O_741,N_4993,N_4931);
xor UO_742 (O_742,N_4909,N_4906);
nor UO_743 (O_743,N_4940,N_4996);
or UO_744 (O_744,N_4952,N_4971);
nand UO_745 (O_745,N_4901,N_4916);
or UO_746 (O_746,N_4909,N_4916);
and UO_747 (O_747,N_4998,N_4984);
xnor UO_748 (O_748,N_4971,N_4959);
nand UO_749 (O_749,N_4922,N_4972);
xor UO_750 (O_750,N_4902,N_4921);
xor UO_751 (O_751,N_4913,N_4900);
and UO_752 (O_752,N_4973,N_4914);
nand UO_753 (O_753,N_4921,N_4969);
nand UO_754 (O_754,N_4941,N_4906);
and UO_755 (O_755,N_4926,N_4987);
and UO_756 (O_756,N_4912,N_4922);
nand UO_757 (O_757,N_4943,N_4927);
xnor UO_758 (O_758,N_4962,N_4987);
and UO_759 (O_759,N_4994,N_4941);
nor UO_760 (O_760,N_4909,N_4969);
nand UO_761 (O_761,N_4943,N_4916);
or UO_762 (O_762,N_4974,N_4901);
xor UO_763 (O_763,N_4926,N_4930);
nand UO_764 (O_764,N_4964,N_4970);
xnor UO_765 (O_765,N_4903,N_4936);
or UO_766 (O_766,N_4923,N_4900);
xnor UO_767 (O_767,N_4916,N_4968);
xnor UO_768 (O_768,N_4989,N_4903);
or UO_769 (O_769,N_4969,N_4934);
and UO_770 (O_770,N_4983,N_4944);
xor UO_771 (O_771,N_4953,N_4912);
nand UO_772 (O_772,N_4997,N_4967);
xor UO_773 (O_773,N_4970,N_4913);
nor UO_774 (O_774,N_4901,N_4932);
nor UO_775 (O_775,N_4916,N_4936);
and UO_776 (O_776,N_4972,N_4923);
and UO_777 (O_777,N_4989,N_4969);
xor UO_778 (O_778,N_4959,N_4927);
or UO_779 (O_779,N_4988,N_4981);
xnor UO_780 (O_780,N_4989,N_4953);
or UO_781 (O_781,N_4980,N_4955);
xor UO_782 (O_782,N_4967,N_4925);
nor UO_783 (O_783,N_4908,N_4910);
nand UO_784 (O_784,N_4911,N_4966);
and UO_785 (O_785,N_4932,N_4993);
or UO_786 (O_786,N_4940,N_4946);
nand UO_787 (O_787,N_4967,N_4948);
xnor UO_788 (O_788,N_4965,N_4914);
nor UO_789 (O_789,N_4908,N_4962);
or UO_790 (O_790,N_4921,N_4922);
or UO_791 (O_791,N_4922,N_4989);
nor UO_792 (O_792,N_4915,N_4946);
nand UO_793 (O_793,N_4964,N_4969);
and UO_794 (O_794,N_4984,N_4942);
and UO_795 (O_795,N_4977,N_4937);
nor UO_796 (O_796,N_4992,N_4941);
xor UO_797 (O_797,N_4985,N_4988);
xor UO_798 (O_798,N_4905,N_4986);
nand UO_799 (O_799,N_4903,N_4961);
and UO_800 (O_800,N_4982,N_4981);
nand UO_801 (O_801,N_4905,N_4992);
or UO_802 (O_802,N_4928,N_4925);
or UO_803 (O_803,N_4911,N_4937);
nor UO_804 (O_804,N_4997,N_4986);
and UO_805 (O_805,N_4918,N_4924);
xnor UO_806 (O_806,N_4957,N_4945);
or UO_807 (O_807,N_4973,N_4955);
nand UO_808 (O_808,N_4917,N_4972);
xor UO_809 (O_809,N_4915,N_4917);
nor UO_810 (O_810,N_4904,N_4942);
or UO_811 (O_811,N_4991,N_4909);
nand UO_812 (O_812,N_4953,N_4915);
nand UO_813 (O_813,N_4932,N_4991);
or UO_814 (O_814,N_4966,N_4989);
nand UO_815 (O_815,N_4939,N_4999);
nor UO_816 (O_816,N_4929,N_4911);
or UO_817 (O_817,N_4946,N_4907);
and UO_818 (O_818,N_4972,N_4959);
and UO_819 (O_819,N_4920,N_4955);
xor UO_820 (O_820,N_4920,N_4982);
xnor UO_821 (O_821,N_4969,N_4981);
nand UO_822 (O_822,N_4929,N_4954);
and UO_823 (O_823,N_4992,N_4910);
nor UO_824 (O_824,N_4948,N_4906);
nand UO_825 (O_825,N_4917,N_4904);
nor UO_826 (O_826,N_4939,N_4923);
xnor UO_827 (O_827,N_4933,N_4973);
and UO_828 (O_828,N_4914,N_4936);
or UO_829 (O_829,N_4973,N_4938);
or UO_830 (O_830,N_4931,N_4944);
or UO_831 (O_831,N_4987,N_4960);
nor UO_832 (O_832,N_4938,N_4968);
nand UO_833 (O_833,N_4919,N_4987);
xnor UO_834 (O_834,N_4939,N_4913);
and UO_835 (O_835,N_4908,N_4979);
xnor UO_836 (O_836,N_4949,N_4982);
and UO_837 (O_837,N_4957,N_4935);
nor UO_838 (O_838,N_4970,N_4937);
nand UO_839 (O_839,N_4900,N_4915);
nor UO_840 (O_840,N_4933,N_4979);
xnor UO_841 (O_841,N_4964,N_4927);
or UO_842 (O_842,N_4984,N_4962);
nor UO_843 (O_843,N_4925,N_4940);
nor UO_844 (O_844,N_4977,N_4989);
or UO_845 (O_845,N_4943,N_4971);
or UO_846 (O_846,N_4984,N_4996);
or UO_847 (O_847,N_4981,N_4972);
xor UO_848 (O_848,N_4961,N_4954);
nand UO_849 (O_849,N_4906,N_4918);
xnor UO_850 (O_850,N_4924,N_4977);
and UO_851 (O_851,N_4935,N_4925);
and UO_852 (O_852,N_4909,N_4958);
xor UO_853 (O_853,N_4912,N_4997);
and UO_854 (O_854,N_4947,N_4958);
and UO_855 (O_855,N_4931,N_4949);
or UO_856 (O_856,N_4926,N_4902);
and UO_857 (O_857,N_4965,N_4950);
or UO_858 (O_858,N_4926,N_4913);
nor UO_859 (O_859,N_4967,N_4951);
xor UO_860 (O_860,N_4915,N_4976);
nand UO_861 (O_861,N_4954,N_4955);
nand UO_862 (O_862,N_4918,N_4985);
or UO_863 (O_863,N_4946,N_4953);
nand UO_864 (O_864,N_4934,N_4987);
xor UO_865 (O_865,N_4994,N_4999);
and UO_866 (O_866,N_4907,N_4938);
or UO_867 (O_867,N_4990,N_4921);
or UO_868 (O_868,N_4914,N_4940);
nor UO_869 (O_869,N_4923,N_4983);
nor UO_870 (O_870,N_4991,N_4948);
nor UO_871 (O_871,N_4940,N_4956);
xor UO_872 (O_872,N_4935,N_4953);
or UO_873 (O_873,N_4919,N_4923);
nand UO_874 (O_874,N_4925,N_4944);
or UO_875 (O_875,N_4954,N_4903);
or UO_876 (O_876,N_4914,N_4968);
or UO_877 (O_877,N_4955,N_4914);
nand UO_878 (O_878,N_4935,N_4909);
nand UO_879 (O_879,N_4911,N_4994);
nand UO_880 (O_880,N_4947,N_4993);
xor UO_881 (O_881,N_4922,N_4930);
nand UO_882 (O_882,N_4951,N_4955);
nor UO_883 (O_883,N_4953,N_4977);
nor UO_884 (O_884,N_4960,N_4998);
xor UO_885 (O_885,N_4952,N_4976);
and UO_886 (O_886,N_4926,N_4973);
or UO_887 (O_887,N_4970,N_4936);
nor UO_888 (O_888,N_4904,N_4933);
nand UO_889 (O_889,N_4950,N_4984);
or UO_890 (O_890,N_4985,N_4923);
xor UO_891 (O_891,N_4991,N_4950);
or UO_892 (O_892,N_4991,N_4990);
xnor UO_893 (O_893,N_4989,N_4932);
or UO_894 (O_894,N_4940,N_4961);
or UO_895 (O_895,N_4948,N_4903);
nand UO_896 (O_896,N_4963,N_4936);
and UO_897 (O_897,N_4948,N_4921);
nor UO_898 (O_898,N_4986,N_4992);
xor UO_899 (O_899,N_4945,N_4902);
xnor UO_900 (O_900,N_4951,N_4901);
or UO_901 (O_901,N_4907,N_4919);
or UO_902 (O_902,N_4950,N_4936);
nor UO_903 (O_903,N_4936,N_4926);
and UO_904 (O_904,N_4960,N_4917);
nand UO_905 (O_905,N_4952,N_4906);
or UO_906 (O_906,N_4937,N_4913);
nand UO_907 (O_907,N_4906,N_4931);
or UO_908 (O_908,N_4915,N_4928);
and UO_909 (O_909,N_4908,N_4943);
nor UO_910 (O_910,N_4995,N_4910);
nand UO_911 (O_911,N_4908,N_4947);
or UO_912 (O_912,N_4940,N_4943);
and UO_913 (O_913,N_4923,N_4981);
or UO_914 (O_914,N_4916,N_4962);
xnor UO_915 (O_915,N_4938,N_4972);
and UO_916 (O_916,N_4906,N_4997);
and UO_917 (O_917,N_4912,N_4973);
nand UO_918 (O_918,N_4973,N_4975);
nand UO_919 (O_919,N_4945,N_4910);
xnor UO_920 (O_920,N_4902,N_4947);
and UO_921 (O_921,N_4999,N_4949);
nor UO_922 (O_922,N_4959,N_4931);
and UO_923 (O_923,N_4954,N_4965);
xnor UO_924 (O_924,N_4968,N_4940);
nor UO_925 (O_925,N_4971,N_4936);
nor UO_926 (O_926,N_4981,N_4936);
or UO_927 (O_927,N_4916,N_4951);
and UO_928 (O_928,N_4979,N_4918);
and UO_929 (O_929,N_4937,N_4990);
or UO_930 (O_930,N_4910,N_4944);
nor UO_931 (O_931,N_4929,N_4973);
nand UO_932 (O_932,N_4975,N_4933);
nand UO_933 (O_933,N_4915,N_4945);
or UO_934 (O_934,N_4922,N_4900);
nor UO_935 (O_935,N_4994,N_4991);
and UO_936 (O_936,N_4998,N_4947);
xnor UO_937 (O_937,N_4950,N_4927);
and UO_938 (O_938,N_4953,N_4981);
or UO_939 (O_939,N_4969,N_4956);
xnor UO_940 (O_940,N_4992,N_4948);
xnor UO_941 (O_941,N_4907,N_4947);
or UO_942 (O_942,N_4940,N_4945);
nand UO_943 (O_943,N_4985,N_4983);
or UO_944 (O_944,N_4935,N_4999);
and UO_945 (O_945,N_4924,N_4979);
nand UO_946 (O_946,N_4917,N_4967);
or UO_947 (O_947,N_4904,N_4937);
nand UO_948 (O_948,N_4949,N_4934);
xor UO_949 (O_949,N_4979,N_4926);
nor UO_950 (O_950,N_4946,N_4995);
or UO_951 (O_951,N_4951,N_4902);
xnor UO_952 (O_952,N_4955,N_4947);
nand UO_953 (O_953,N_4994,N_4924);
and UO_954 (O_954,N_4903,N_4994);
nand UO_955 (O_955,N_4902,N_4952);
or UO_956 (O_956,N_4989,N_4967);
xnor UO_957 (O_957,N_4947,N_4996);
xnor UO_958 (O_958,N_4908,N_4922);
or UO_959 (O_959,N_4986,N_4971);
xor UO_960 (O_960,N_4908,N_4957);
nand UO_961 (O_961,N_4998,N_4952);
nand UO_962 (O_962,N_4948,N_4950);
nor UO_963 (O_963,N_4956,N_4906);
nor UO_964 (O_964,N_4966,N_4975);
and UO_965 (O_965,N_4945,N_4923);
nand UO_966 (O_966,N_4980,N_4990);
nand UO_967 (O_967,N_4959,N_4932);
nor UO_968 (O_968,N_4937,N_4978);
xnor UO_969 (O_969,N_4916,N_4942);
xor UO_970 (O_970,N_4991,N_4982);
and UO_971 (O_971,N_4983,N_4924);
and UO_972 (O_972,N_4975,N_4925);
nor UO_973 (O_973,N_4933,N_4955);
nand UO_974 (O_974,N_4960,N_4954);
or UO_975 (O_975,N_4970,N_4971);
or UO_976 (O_976,N_4974,N_4988);
or UO_977 (O_977,N_4998,N_4924);
nand UO_978 (O_978,N_4957,N_4987);
nand UO_979 (O_979,N_4947,N_4917);
xnor UO_980 (O_980,N_4919,N_4918);
nand UO_981 (O_981,N_4905,N_4984);
nand UO_982 (O_982,N_4944,N_4901);
nor UO_983 (O_983,N_4956,N_4923);
nor UO_984 (O_984,N_4923,N_4966);
nand UO_985 (O_985,N_4925,N_4936);
nand UO_986 (O_986,N_4961,N_4999);
nor UO_987 (O_987,N_4965,N_4971);
nor UO_988 (O_988,N_4981,N_4931);
nand UO_989 (O_989,N_4932,N_4963);
or UO_990 (O_990,N_4978,N_4954);
xor UO_991 (O_991,N_4934,N_4935);
or UO_992 (O_992,N_4984,N_4933);
and UO_993 (O_993,N_4976,N_4996);
or UO_994 (O_994,N_4953,N_4934);
and UO_995 (O_995,N_4912,N_4999);
nor UO_996 (O_996,N_4968,N_4980);
and UO_997 (O_997,N_4915,N_4918);
xor UO_998 (O_998,N_4914,N_4959);
xor UO_999 (O_999,N_4966,N_4952);
endmodule