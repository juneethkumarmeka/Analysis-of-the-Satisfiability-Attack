module basic_2500_25000_3000_10_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_1392,In_1338);
or U1 (N_1,In_750,In_1051);
or U2 (N_2,In_2021,In_2282);
xnor U3 (N_3,In_1684,In_935);
xnor U4 (N_4,In_709,In_627);
nor U5 (N_5,In_1048,In_2475);
nor U6 (N_6,In_1029,In_190);
xnor U7 (N_7,In_2054,In_224);
and U8 (N_8,In_2161,In_1756);
nor U9 (N_9,In_2123,In_426);
nand U10 (N_10,In_1495,In_468);
xnor U11 (N_11,In_1373,In_2395);
xnor U12 (N_12,In_1843,In_1409);
nor U13 (N_13,In_759,In_1537);
xnor U14 (N_14,In_1199,In_1266);
or U15 (N_15,In_570,In_204);
xor U16 (N_16,In_409,In_1907);
nand U17 (N_17,In_1844,In_332);
nand U18 (N_18,In_1948,In_1660);
or U19 (N_19,In_1476,In_1092);
nand U20 (N_20,In_1846,In_425);
nand U21 (N_21,In_1312,In_2292);
nor U22 (N_22,In_2426,In_303);
and U23 (N_23,In_92,In_1551);
xor U24 (N_24,In_1608,In_1977);
nor U25 (N_25,In_1404,In_690);
xnor U26 (N_26,In_670,In_1172);
nand U27 (N_27,In_1541,In_1545);
or U28 (N_28,In_135,In_2470);
or U29 (N_29,In_677,In_209);
xnor U30 (N_30,In_1261,In_2219);
nor U31 (N_31,In_835,In_316);
or U32 (N_32,In_581,In_1938);
nor U33 (N_33,In_1847,In_1664);
and U34 (N_34,In_1787,In_1091);
nand U35 (N_35,In_557,In_1748);
xnor U36 (N_36,In_624,In_1354);
xor U37 (N_37,In_2402,In_2250);
and U38 (N_38,In_885,In_233);
and U39 (N_39,In_648,In_1694);
and U40 (N_40,In_2447,In_519);
and U41 (N_41,In_685,In_622);
nand U42 (N_42,In_1336,In_1220);
and U43 (N_43,In_857,In_75);
and U44 (N_44,In_2370,In_1350);
or U45 (N_45,In_1211,In_762);
nand U46 (N_46,In_27,In_1362);
xnor U47 (N_47,In_503,In_2129);
nand U48 (N_48,In_516,In_285);
nand U49 (N_49,In_1127,In_949);
nand U50 (N_50,In_1877,In_587);
nor U51 (N_51,In_873,In_609);
xor U52 (N_52,In_1702,In_1695);
and U53 (N_53,In_108,In_1281);
xnor U54 (N_54,In_2163,In_239);
nor U55 (N_55,In_1866,In_1654);
and U56 (N_56,In_1621,In_811);
nor U57 (N_57,In_459,In_1529);
or U58 (N_58,In_1449,In_321);
nand U59 (N_59,In_2483,In_1469);
xnor U60 (N_60,In_371,In_905);
xor U61 (N_61,In_1945,In_1254);
xor U62 (N_62,In_572,In_260);
xnor U63 (N_63,In_283,In_1921);
xor U64 (N_64,In_1982,In_132);
nand U65 (N_65,In_346,In_1600);
nor U66 (N_66,In_124,In_952);
and U67 (N_67,In_1275,In_252);
or U68 (N_68,In_1596,In_2325);
and U69 (N_69,In_131,In_1980);
xnor U70 (N_70,In_2328,In_819);
nor U71 (N_71,In_1810,In_289);
or U72 (N_72,In_152,In_76);
and U73 (N_73,In_480,In_118);
nand U74 (N_74,In_445,In_1284);
and U75 (N_75,In_1902,In_2059);
nor U76 (N_76,In_592,In_2258);
nor U77 (N_77,In_880,In_1652);
nand U78 (N_78,In_848,In_2376);
nor U79 (N_79,In_80,In_126);
or U80 (N_80,In_2225,In_481);
xnor U81 (N_81,In_2154,In_1082);
or U82 (N_82,In_1322,In_632);
xor U83 (N_83,In_254,In_1221);
or U84 (N_84,In_416,In_1166);
nor U85 (N_85,In_38,In_1549);
or U86 (N_86,In_1042,In_333);
nor U87 (N_87,In_1317,In_921);
or U88 (N_88,In_993,In_395);
or U89 (N_89,In_1944,In_2084);
and U90 (N_90,In_20,In_2201);
or U91 (N_91,In_653,In_1258);
or U92 (N_92,In_1732,In_2087);
and U93 (N_93,In_1739,In_2198);
or U94 (N_94,In_298,In_317);
nand U95 (N_95,In_1868,In_2007);
xor U96 (N_96,In_793,In_2037);
nand U97 (N_97,In_598,In_628);
nand U98 (N_98,In_1288,In_79);
or U99 (N_99,In_2236,In_1471);
and U100 (N_100,In_53,In_422);
nand U101 (N_101,In_1738,In_744);
or U102 (N_102,In_2126,In_944);
nand U103 (N_103,In_1767,In_2091);
nand U104 (N_104,In_1401,In_1713);
or U105 (N_105,In_697,In_1458);
xor U106 (N_106,In_1862,In_1396);
nor U107 (N_107,In_1052,In_218);
nand U108 (N_108,In_1524,In_774);
xnor U109 (N_109,In_2348,In_389);
nand U110 (N_110,In_57,In_573);
xor U111 (N_111,In_2436,In_1544);
nand U112 (N_112,In_403,In_2003);
and U113 (N_113,In_1780,In_585);
nor U114 (N_114,In_2389,In_658);
and U115 (N_115,In_896,In_121);
and U116 (N_116,In_443,In_2260);
or U117 (N_117,In_2031,In_286);
or U118 (N_118,In_216,In_2090);
and U119 (N_119,In_1849,In_1936);
nor U120 (N_120,In_339,In_2377);
and U121 (N_121,In_117,In_1501);
nor U122 (N_122,In_1192,In_326);
nor U123 (N_123,In_498,In_542);
nand U124 (N_124,In_24,In_2298);
nor U125 (N_125,In_1807,In_1771);
or U126 (N_126,In_977,In_1917);
or U127 (N_127,In_1260,In_2423);
and U128 (N_128,In_1132,In_1962);
nor U129 (N_129,In_2439,In_1644);
and U130 (N_130,In_1975,In_97);
xnor U131 (N_131,In_1487,In_1090);
and U132 (N_132,In_1467,In_193);
nor U133 (N_133,In_1834,In_1589);
xnor U134 (N_134,In_2013,In_1062);
nor U135 (N_135,In_248,In_1889);
xor U136 (N_136,In_353,In_1910);
and U137 (N_137,In_976,In_1958);
or U138 (N_138,In_1263,In_2092);
nor U139 (N_139,In_297,In_827);
and U140 (N_140,In_219,In_1900);
or U141 (N_141,In_1747,In_1295);
xnor U142 (N_142,In_1235,In_1195);
nor U143 (N_143,In_114,In_164);
nand U144 (N_144,In_143,In_915);
or U145 (N_145,In_2148,In_349);
nand U146 (N_146,In_1395,In_1525);
and U147 (N_147,In_579,In_2272);
nor U148 (N_148,In_494,In_2323);
xnor U149 (N_149,In_2467,In_510);
xnor U150 (N_150,In_2456,In_243);
or U151 (N_151,In_381,In_2243);
nor U152 (N_152,In_1286,In_236);
nand U153 (N_153,In_2297,In_1460);
nor U154 (N_154,In_1277,In_2138);
nor U155 (N_155,In_2019,In_633);
nor U156 (N_156,In_2246,In_476);
nand U157 (N_157,In_967,In_1138);
or U158 (N_158,In_895,In_1432);
nand U159 (N_159,In_1233,In_681);
nor U160 (N_160,In_734,In_1297);
or U161 (N_161,In_1207,In_464);
xor U162 (N_162,In_1,In_1247);
nand U163 (N_163,In_360,In_675);
nor U164 (N_164,In_50,In_2188);
nand U165 (N_165,In_382,In_1113);
xnor U166 (N_166,In_1878,In_1858);
nand U167 (N_167,In_2190,In_642);
nor U168 (N_168,In_2215,In_110);
nand U169 (N_169,In_52,In_2155);
or U170 (N_170,In_1802,In_1499);
and U171 (N_171,In_305,In_1214);
and U172 (N_172,In_467,In_1431);
and U173 (N_173,In_953,In_2081);
nand U174 (N_174,In_1223,In_733);
and U175 (N_175,In_2030,In_119);
nand U176 (N_176,In_745,In_1405);
xor U177 (N_177,In_1011,In_1349);
nor U178 (N_178,In_407,In_2079);
and U179 (N_179,In_1470,In_2070);
nand U180 (N_180,In_417,In_45);
and U181 (N_181,In_2329,In_2118);
xnor U182 (N_182,In_1358,In_525);
xor U183 (N_183,In_974,In_723);
or U184 (N_184,In_1319,In_1800);
nor U185 (N_185,In_414,In_350);
xor U186 (N_186,In_1604,In_2127);
and U187 (N_187,In_12,In_483);
and U188 (N_188,In_1988,In_2335);
xor U189 (N_189,In_1427,In_1264);
and U190 (N_190,In_1055,In_870);
nand U191 (N_191,In_761,In_829);
nor U192 (N_192,In_4,In_1402);
nor U193 (N_193,In_1150,In_2180);
and U194 (N_194,In_172,In_253);
and U195 (N_195,In_1506,In_641);
and U196 (N_196,In_1558,In_964);
xnor U197 (N_197,In_899,In_1759);
nor U198 (N_198,In_2427,In_44);
xnor U199 (N_199,In_2101,In_777);
and U200 (N_200,In_357,In_694);
nor U201 (N_201,In_461,In_918);
xnor U202 (N_202,In_597,In_1566);
or U203 (N_203,In_2100,In_1947);
and U204 (N_204,In_10,In_1946);
or U205 (N_205,In_2487,In_2386);
xor U206 (N_206,In_984,In_732);
nand U207 (N_207,In_826,In_13);
nand U208 (N_208,In_1490,In_2134);
nand U209 (N_209,In_1851,In_1163);
xor U210 (N_210,In_1033,In_262);
or U211 (N_211,In_191,In_1512);
or U212 (N_212,In_250,In_1368);
nor U213 (N_213,In_1193,In_2493);
nand U214 (N_214,In_563,In_2274);
nand U215 (N_215,In_85,In_1594);
and U216 (N_216,In_1996,In_2152);
nand U217 (N_217,In_308,In_2097);
or U218 (N_218,In_1316,In_2305);
and U219 (N_219,In_1581,In_238);
or U220 (N_220,In_1956,In_612);
xnor U221 (N_221,In_1611,In_2312);
and U222 (N_222,In_1578,In_2361);
and U223 (N_223,In_2318,In_63);
nor U224 (N_224,In_217,In_1197);
or U225 (N_225,In_813,In_1813);
nand U226 (N_226,In_824,In_725);
nor U227 (N_227,In_67,In_499);
nor U228 (N_228,In_1561,In_1175);
xnor U229 (N_229,In_1842,In_2414);
or U230 (N_230,In_1991,In_1840);
xor U231 (N_231,In_719,In_2355);
nor U232 (N_232,In_1606,In_1072);
nand U233 (N_233,In_1085,In_2041);
or U234 (N_234,In_1229,In_1880);
and U235 (N_235,In_814,In_374);
nand U236 (N_236,In_1194,In_2045);
nor U237 (N_237,In_2429,In_712);
nor U238 (N_238,In_1942,In_1287);
nand U239 (N_239,In_784,In_2227);
and U240 (N_240,In_916,In_2232);
or U241 (N_241,In_501,In_1446);
nor U242 (N_242,In_344,In_182);
or U243 (N_243,In_1179,In_771);
and U244 (N_244,In_828,In_2194);
or U245 (N_245,In_1721,In_306);
nor U246 (N_246,In_2327,In_2096);
xor U247 (N_247,In_1743,In_99);
xnor U248 (N_248,In_2284,In_2075);
or U249 (N_249,In_742,In_1355);
or U250 (N_250,In_1930,In_1273);
or U251 (N_251,In_738,In_1546);
nand U252 (N_252,In_1750,In_1775);
nand U253 (N_253,In_724,In_577);
nand U254 (N_254,In_1965,In_1334);
nand U255 (N_255,In_767,In_2463);
or U256 (N_256,In_1474,In_2162);
or U257 (N_257,In_2481,In_1839);
nand U258 (N_258,In_477,In_87);
nor U259 (N_259,In_715,In_865);
nand U260 (N_260,In_2207,In_2345);
xor U261 (N_261,In_1050,In_1579);
nor U262 (N_262,In_795,In_1379);
and U263 (N_263,In_1887,In_1200);
nor U264 (N_264,In_2202,In_1265);
nor U265 (N_265,In_769,In_199);
and U266 (N_266,In_1299,In_590);
xor U267 (N_267,In_1879,In_1827);
xnor U268 (N_268,In_1829,In_9);
nor U269 (N_269,In_89,In_688);
nor U270 (N_270,In_882,In_300);
or U271 (N_271,In_1937,In_2492);
nor U272 (N_272,In_1803,In_336);
xnor U273 (N_273,In_2050,In_1278);
xor U274 (N_274,In_1315,In_1259);
nand U275 (N_275,In_554,In_939);
xor U276 (N_276,In_1661,In_235);
nand U277 (N_277,In_809,In_1693);
and U278 (N_278,In_2094,In_1078);
or U279 (N_279,In_454,In_1502);
and U280 (N_280,In_904,In_1662);
nand U281 (N_281,In_208,In_1539);
and U282 (N_282,In_2151,In_666);
nand U283 (N_283,In_1765,In_2491);
nor U284 (N_284,In_1369,In_834);
or U285 (N_285,In_1382,In_1423);
and U286 (N_286,In_799,In_386);
or U287 (N_287,In_230,In_1871);
xor U288 (N_288,In_2185,In_1370);
or U289 (N_289,In_1522,In_1613);
xor U290 (N_290,In_1145,In_906);
or U291 (N_291,In_2358,In_1773);
or U292 (N_292,In_983,In_926);
nand U293 (N_293,In_740,In_2399);
and U294 (N_294,In_2497,In_574);
and U295 (N_295,In_620,In_676);
xor U296 (N_296,In_1384,In_1054);
nand U297 (N_297,In_2294,In_1215);
or U298 (N_298,In_2257,In_1933);
and U299 (N_299,In_1105,In_1129);
xor U300 (N_300,In_2109,In_1568);
xor U301 (N_301,In_1485,In_207);
or U302 (N_302,In_765,In_1450);
xor U303 (N_303,In_2472,In_1912);
xor U304 (N_304,In_1659,In_1651);
nor U305 (N_305,In_189,In_802);
xor U306 (N_306,In_49,In_457);
nand U307 (N_307,In_2145,In_1791);
and U308 (N_308,In_1285,In_307);
nor U309 (N_309,In_1068,In_2012);
or U310 (N_310,In_35,In_660);
nand U311 (N_311,In_1407,In_792);
nand U312 (N_312,In_534,In_874);
xor U313 (N_313,In_1711,In_1832);
nand U314 (N_314,In_643,In_328);
and U315 (N_315,In_469,In_269);
and U316 (N_316,In_631,In_1511);
nand U317 (N_317,In_441,In_16);
nand U318 (N_318,In_1023,In_1619);
xnor U319 (N_319,In_575,In_361);
xnor U320 (N_320,In_1083,In_1734);
or U321 (N_321,In_324,In_113);
nor U322 (N_322,In_1073,In_1292);
nand U323 (N_323,In_1805,In_26);
and U324 (N_324,In_736,In_615);
xor U325 (N_325,In_1974,In_1208);
nand U326 (N_326,In_2025,In_1952);
nor U327 (N_327,In_710,In_225);
and U328 (N_328,In_2052,In_2286);
nor U329 (N_329,In_900,In_28);
xnor U330 (N_330,In_807,In_544);
nand U331 (N_331,In_2000,In_1308);
or U332 (N_332,In_2344,In_1904);
xor U333 (N_333,In_2093,In_2428);
nand U334 (N_334,In_739,In_428);
or U335 (N_335,In_1815,In_2166);
nand U336 (N_336,In_334,In_1935);
or U337 (N_337,In_1624,In_2060);
and U338 (N_338,In_1157,In_936);
and U339 (N_339,In_2381,In_198);
xnor U340 (N_340,In_2105,In_523);
and U341 (N_341,In_1509,In_1184);
and U342 (N_342,In_2222,In_442);
nor U343 (N_343,In_1714,In_1557);
nor U344 (N_344,In_315,In_84);
or U345 (N_345,In_755,In_621);
nor U346 (N_346,In_86,In_2254);
nor U347 (N_347,In_2380,In_2224);
and U348 (N_348,In_1038,In_2432);
nor U349 (N_349,In_1472,In_1420);
nand U350 (N_350,In_2178,In_583);
xnor U351 (N_351,In_2149,In_1478);
or U352 (N_352,In_163,In_1547);
nor U353 (N_353,In_1473,In_2208);
nor U354 (N_354,In_475,In_39);
nand U355 (N_355,In_2339,In_1622);
nor U356 (N_356,In_279,In_1607);
xor U357 (N_357,In_810,In_1015);
nand U358 (N_358,In_1508,In_2150);
nand U359 (N_359,In_661,In_613);
xnor U360 (N_360,In_2285,In_1393);
nand U361 (N_361,In_120,In_1462);
xor U362 (N_362,In_1436,In_355);
nand U363 (N_363,In_1928,In_384);
xor U364 (N_364,In_1057,In_1479);
xnor U365 (N_365,In_825,In_111);
and U366 (N_366,In_1770,In_1171);
and U367 (N_367,In_251,In_2276);
xor U368 (N_368,In_1676,In_90);
and U369 (N_369,In_1484,In_18);
nor U370 (N_370,In_276,In_2437);
xor U371 (N_371,In_166,In_1893);
nand U372 (N_372,In_1990,In_1680);
nand U373 (N_373,In_1480,In_1481);
nand U374 (N_374,In_956,In_2357);
and U375 (N_375,In_971,In_2157);
and U376 (N_376,In_656,In_786);
and U377 (N_377,In_401,In_1272);
and U378 (N_378,In_611,In_484);
and U379 (N_379,In_1914,In_1642);
or U380 (N_380,In_907,In_2401);
xnor U381 (N_381,In_1086,In_1383);
and U382 (N_382,In_1210,In_460);
xor U383 (N_383,In_908,In_2369);
nand U384 (N_384,In_541,In_452);
nor U385 (N_385,In_2113,In_128);
xor U386 (N_386,In_955,In_1516);
or U387 (N_387,In_1030,In_5);
nor U388 (N_388,In_1656,In_379);
nand U389 (N_389,In_2065,In_1003);
or U390 (N_390,In_1911,In_2156);
and U391 (N_391,In_1181,In_1726);
and U392 (N_392,In_1328,In_133);
or U393 (N_393,In_803,In_1044);
xnor U394 (N_394,In_134,In_986);
nor U395 (N_395,In_854,In_1205);
or U396 (N_396,In_1874,In_1823);
and U397 (N_397,In_2363,In_748);
and U398 (N_398,In_782,In_539);
xnor U399 (N_399,In_1768,In_515);
nor U400 (N_400,In_497,In_954);
or U401 (N_401,In_638,In_2262);
nand U402 (N_402,In_1359,In_1709);
xor U403 (N_403,In_2032,In_2375);
nor U404 (N_404,In_2042,In_797);
xnor U405 (N_405,In_46,In_1919);
nand U406 (N_406,In_940,In_2210);
xnor U407 (N_407,In_1897,In_1735);
nor U408 (N_408,In_1682,In_402);
xnor U409 (N_409,In_1201,In_8);
nor U410 (N_410,In_1576,In_1898);
nor U411 (N_411,In_1754,In_1616);
nor U412 (N_412,In_836,In_2213);
nor U413 (N_413,In_830,In_1951);
xnor U414 (N_414,In_453,In_1097);
or U415 (N_415,In_1673,In_2387);
xor U416 (N_416,In_157,In_1999);
and U417 (N_417,In_2024,In_2314);
or U418 (N_418,In_2076,In_342);
xnor U419 (N_419,In_527,In_1239);
nand U420 (N_420,In_812,In_1095);
xor U421 (N_421,In_1523,In_2132);
nor U422 (N_422,In_2283,In_2119);
xor U423 (N_423,In_1888,In_1209);
nor U424 (N_424,In_2307,In_589);
nor U425 (N_425,In_2471,In_1027);
xor U426 (N_426,In_514,In_1135);
xnor U427 (N_427,In_1556,In_2136);
xnor U428 (N_428,In_1553,In_1961);
nand U429 (N_429,In_1045,In_48);
and U430 (N_430,In_1836,In_549);
nor U431 (N_431,In_352,In_268);
and U432 (N_432,In_1894,In_427);
or U433 (N_433,In_2016,In_1189);
nand U434 (N_434,In_168,In_1535);
and U435 (N_435,In_200,In_909);
xnor U436 (N_436,In_1416,In_385);
and U437 (N_437,In_702,In_1032);
nand U438 (N_438,In_214,In_2137);
or U439 (N_439,In_140,In_2383);
and U440 (N_440,In_816,In_2416);
nor U441 (N_441,In_1825,In_1587);
nor U442 (N_442,In_1468,In_1043);
or U443 (N_443,In_1675,In_1004);
nand U444 (N_444,In_107,In_2171);
and U445 (N_445,In_787,In_535);
nand U446 (N_446,In_2303,In_623);
nand U447 (N_447,In_1752,In_2261);
or U448 (N_448,In_1024,In_1067);
nor U449 (N_449,In_2400,In_569);
or U450 (N_450,In_1153,In_778);
nand U451 (N_451,In_1703,In_1635);
nand U452 (N_452,In_1463,In_862);
xnor U453 (N_453,In_2488,In_282);
xor U454 (N_454,In_337,In_910);
nand U455 (N_455,In_822,In_720);
or U456 (N_456,In_245,In_1447);
or U457 (N_457,In_1216,In_327);
nor U458 (N_458,In_1809,In_437);
xor U459 (N_459,In_1683,In_1941);
xnor U460 (N_460,In_844,In_1835);
nand U461 (N_461,In_1424,In_1021);
nor U462 (N_462,In_637,In_843);
and U463 (N_463,In_1385,In_1131);
xor U464 (N_464,In_1257,In_1300);
and U465 (N_465,In_2214,In_683);
and U466 (N_466,In_249,In_2068);
nor U467 (N_467,In_640,In_2099);
xnor U468 (N_468,In_506,In_1453);
nor U469 (N_469,In_1433,In_727);
and U470 (N_470,In_2264,In_897);
nand U471 (N_471,In_1001,In_1360);
nor U472 (N_472,In_1093,In_749);
xor U473 (N_473,In_2004,In_2067);
nor U474 (N_474,In_1830,In_2451);
xor U475 (N_475,In_2242,In_1357);
xnor U476 (N_476,In_2212,In_789);
and U477 (N_477,In_1390,In_1364);
nor U478 (N_478,In_619,In_2122);
or U479 (N_479,In_794,In_1203);
xor U480 (N_480,In_1301,In_1270);
and U481 (N_481,In_1710,In_1310);
nand U482 (N_482,In_275,In_1663);
nand U483 (N_483,In_1758,In_2495);
nand U484 (N_484,In_1324,In_891);
or U485 (N_485,In_1649,In_1995);
or U486 (N_486,In_2332,In_455);
and U487 (N_487,In_2352,In_398);
xor U488 (N_488,In_1326,In_1147);
xnor U489 (N_489,In_1012,In_2071);
nand U490 (N_490,In_487,In_1230);
xor U491 (N_491,In_1451,In_1018);
and U492 (N_492,In_991,In_2462);
nor U493 (N_493,In_2130,In_2479);
xnor U494 (N_494,In_1908,In_1824);
nand U495 (N_495,In_1969,In_1669);
nand U496 (N_496,In_1950,In_2182);
nor U497 (N_497,In_772,In_730);
and U498 (N_498,In_1442,In_482);
and U499 (N_499,In_318,In_1009);
or U500 (N_500,In_183,In_731);
nand U501 (N_501,In_1114,In_173);
or U502 (N_502,In_410,In_538);
nand U503 (N_503,In_2,In_2365);
nor U504 (N_504,In_992,In_2115);
nor U505 (N_505,In_1188,In_2478);
and U506 (N_506,In_212,In_171);
xor U507 (N_507,In_465,In_1586);
nor U508 (N_508,In_1108,In_71);
xnor U509 (N_509,In_540,In_66);
xor U510 (N_510,In_617,In_345);
and U511 (N_511,In_711,In_1896);
and U512 (N_512,In_942,In_432);
nor U513 (N_513,In_1954,In_1906);
or U514 (N_514,In_2005,In_1130);
nand U515 (N_515,In_729,In_1010);
and U516 (N_516,In_73,In_2058);
and U517 (N_517,In_528,In_576);
and U518 (N_518,In_911,In_2023);
xor U519 (N_519,In_1356,In_821);
and U520 (N_520,In_1049,In_2398);
or U521 (N_521,In_37,In_1020);
and U522 (N_522,In_1121,In_1926);
and U523 (N_523,In_1833,In_2160);
or U524 (N_524,In_41,In_1218);
and U525 (N_525,In_30,In_1144);
or U526 (N_526,In_1069,In_1744);
nor U527 (N_527,In_378,In_923);
or U528 (N_528,In_1242,In_1872);
nor U529 (N_529,In_489,In_451);
xor U530 (N_530,In_1388,In_1025);
nand U531 (N_531,In_1439,In_2098);
xnor U532 (N_532,In_2393,In_1425);
nor U533 (N_533,In_278,In_2438);
and U534 (N_534,In_931,In_2191);
nand U535 (N_535,In_40,In_33);
and U536 (N_536,In_682,In_1972);
nor U537 (N_537,In_2112,In_1267);
nand U538 (N_538,In_958,In_1161);
nand U539 (N_539,In_3,In_330);
xor U540 (N_540,In_875,In_14);
xor U541 (N_541,In_2281,In_994);
or U542 (N_542,In_917,In_1855);
or U543 (N_543,In_2265,In_878);
nand U544 (N_544,In_1741,In_625);
xor U545 (N_545,In_59,In_933);
xnor U546 (N_546,In_1968,In_2351);
and U547 (N_547,In_2244,In_1776);
or U548 (N_548,In_1294,In_743);
xnor U549 (N_549,In_1323,In_1548);
nand U550 (N_550,In_860,In_1614);
nor U551 (N_551,In_989,In_2234);
nor U552 (N_552,In_429,In_165);
or U553 (N_553,In_864,In_1477);
xor U554 (N_554,In_2397,In_1859);
and U555 (N_555,In_1101,In_969);
and U556 (N_556,In_1232,In_1040);
nor U557 (N_557,In_1348,In_51);
xnor U558 (N_558,In_2186,In_508);
or U559 (N_559,In_2267,In_922);
nand U560 (N_560,In_1876,In_1440);
nor U561 (N_561,In_1592,In_560);
xor U562 (N_562,In_366,In_2165);
and U563 (N_563,In_2110,In_1380);
nor U564 (N_564,In_657,In_2230);
nand U565 (N_565,In_602,In_495);
or U566 (N_566,In_752,In_421);
xor U567 (N_567,In_1913,In_561);
nor U568 (N_568,In_2026,In_1112);
or U569 (N_569,In_1647,In_1643);
and U570 (N_570,In_56,In_96);
or U571 (N_571,In_1099,In_1367);
or U572 (N_572,In_903,In_1140);
nand U573 (N_573,In_446,In_1096);
or U574 (N_574,In_2382,In_479);
xor U575 (N_575,In_438,In_237);
nor U576 (N_576,In_500,In_2141);
and U577 (N_577,In_1005,In_1376);
nand U578 (N_578,In_999,In_125);
nor U579 (N_579,In_1707,In_2310);
nor U580 (N_580,In_1857,In_1638);
and U581 (N_581,In_2342,In_684);
and U582 (N_582,In_1279,In_188);
or U583 (N_583,In_277,In_1155);
xor U584 (N_584,In_1372,In_737);
nor U585 (N_585,In_698,In_1677);
or U586 (N_586,In_2330,In_1971);
nand U587 (N_587,In_1252,In_1895);
nor U588 (N_588,In_1870,In_1339);
xor U589 (N_589,In_639,In_2174);
and U590 (N_590,In_1918,In_1891);
nor U591 (N_591,In_202,In_2346);
nor U592 (N_592,In_91,In_1753);
nand U593 (N_593,In_1627,In_302);
or U594 (N_594,In_473,In_707);
nand U595 (N_595,In_1430,In_879);
xor U596 (N_596,In_1881,In_1305);
or U597 (N_597,In_2268,In_58);
nor U598 (N_598,In_1814,In_1489);
nand U599 (N_599,In_1191,In_6);
nor U600 (N_600,In_1690,In_1959);
nor U601 (N_601,In_1136,In_2144);
and U602 (N_602,In_2120,In_1497);
nor U603 (N_603,In_380,In_1142);
nand U604 (N_604,In_2302,In_1346);
nand U605 (N_605,In_1250,In_2403);
nor U606 (N_606,In_507,In_902);
or U607 (N_607,In_2378,In_841);
or U608 (N_608,In_2295,In_678);
or U609 (N_609,In_881,In_383);
nand U610 (N_610,In_2354,In_1213);
or U611 (N_611,In_849,In_2116);
or U612 (N_612,In_1786,In_2425);
or U613 (N_613,In_2204,In_883);
nand U614 (N_614,In_1925,In_1408);
xor U615 (N_615,In_2206,In_2433);
and U616 (N_616,In_1345,In_272);
xnor U617 (N_617,In_1665,In_373);
and U618 (N_618,In_1679,In_2489);
and U619 (N_619,In_818,In_1796);
nor U620 (N_620,In_591,In_1778);
xnor U621 (N_621,In_2367,In_1014);
or U622 (N_622,In_1645,In_1426);
nor U623 (N_623,In_1922,In_2419);
and U624 (N_624,In_1289,In_444);
nand U625 (N_625,In_2104,In_287);
xor U626 (N_626,In_2418,In_2080);
xnor U627 (N_627,In_1955,In_1366);
nand U628 (N_628,In_559,In_392);
xnor U629 (N_629,In_1283,In_1059);
or U630 (N_630,In_932,In_1779);
and U631 (N_631,In_431,In_756);
xor U632 (N_632,In_1492,In_1046);
or U633 (N_633,In_901,In_449);
or U634 (N_634,In_1429,In_323);
nor U635 (N_635,In_2147,In_1903);
xor U636 (N_636,In_696,In_162);
xnor U637 (N_637,In_55,In_2290);
xor U638 (N_638,In_699,In_2229);
nor U639 (N_639,In_2324,In_1641);
and U640 (N_640,In_1251,In_1443);
nand U641 (N_641,In_914,In_2106);
and U642 (N_642,In_706,In_359);
xnor U643 (N_643,In_288,In_1573);
or U644 (N_644,In_726,In_1183);
and U645 (N_645,In_2288,In_673);
xor U646 (N_646,In_1811,In_753);
and U647 (N_647,In_1630,In_773);
nand U648 (N_648,In_466,In_257);
and U649 (N_649,In_1314,In_15);
and U650 (N_650,In_1792,In_1022);
and U651 (N_651,In_301,In_194);
or U652 (N_652,In_1901,In_1650);
and U653 (N_653,In_331,In_980);
and U654 (N_654,In_2033,In_735);
xnor U655 (N_655,In_979,In_687);
and U656 (N_656,In_545,In_2228);
nand U657 (N_657,In_1963,In_1798);
and U658 (N_658,In_713,In_1640);
xnor U659 (N_659,In_2072,In_70);
nor U660 (N_660,In_1386,In_309);
or U661 (N_661,In_871,In_1993);
nor U662 (N_662,In_404,In_1731);
or U663 (N_663,In_806,In_663);
nor U664 (N_664,In_192,In_798);
and U665 (N_665,In_390,In_610);
nor U666 (N_666,In_941,In_1164);
xor U667 (N_667,In_1111,In_2089);
xnor U668 (N_668,In_861,In_2280);
xnor U669 (N_669,In_169,In_1180);
nor U670 (N_670,In_2009,In_1330);
and U671 (N_671,In_470,In_2063);
xnor U672 (N_672,In_1056,In_2197);
nand U673 (N_673,In_2474,In_1219);
or U674 (N_674,In_1167,In_1417);
nand U675 (N_675,In_1625,In_2331);
xor U676 (N_676,In_505,In_2049);
xor U677 (N_677,In_88,In_1760);
xor U678 (N_678,In_1075,In_605);
or U679 (N_679,In_596,In_2069);
nor U680 (N_680,In_1822,In_1636);
nand U681 (N_681,In_158,In_858);
and U682 (N_682,In_680,In_161);
or U683 (N_683,In_531,In_2226);
or U684 (N_684,In_929,In_718);
nor U685 (N_685,In_1618,In_652);
or U686 (N_686,In_1533,In_1321);
nor U687 (N_687,In_270,In_1152);
xor U688 (N_688,In_512,In_820);
nor U689 (N_689,In_1720,In_292);
and U690 (N_690,In_1931,In_2095);
and U691 (N_691,In_716,In_1320);
nand U692 (N_692,In_1574,In_1146);
xnor U693 (N_693,In_1583,In_1733);
and U694 (N_694,In_1637,In_1063);
and U695 (N_695,In_588,In_2340);
or U696 (N_696,In_1986,In_1340);
nor U697 (N_697,In_1176,In_1884);
nand U698 (N_698,In_2457,In_1378);
and U699 (N_699,In_291,In_170);
and U700 (N_700,In_808,In_2017);
and U701 (N_701,In_2034,In_223);
xnor U702 (N_702,In_1565,In_293);
and U703 (N_703,In_550,In_100);
or U704 (N_704,In_1845,In_1841);
and U705 (N_705,In_1559,In_1742);
xor U706 (N_706,In_1343,In_195);
xor U707 (N_707,In_1749,In_1764);
nor U708 (N_708,In_1331,In_1528);
xor U709 (N_709,In_1118,In_2048);
or U710 (N_710,In_433,In_123);
or U711 (N_711,In_1875,In_1406);
nand U712 (N_712,In_1280,In_913);
nor U713 (N_713,In_1909,In_1860);
and U714 (N_714,In_2356,In_1500);
or U715 (N_715,In_116,In_630);
and U716 (N_716,In_1035,In_2394);
nand U717 (N_717,In_2164,In_367);
nor U718 (N_718,In_2193,In_833);
nor U719 (N_719,In_2300,In_2235);
or U720 (N_720,In_594,In_178);
xnor U721 (N_721,In_636,In_1667);
or U722 (N_722,In_68,In_536);
nor U723 (N_723,In_1282,In_400);
or U724 (N_724,In_78,In_448);
or U725 (N_725,In_1632,In_1751);
nand U726 (N_726,In_2349,In_2187);
and U727 (N_727,In_281,In_634);
xnor U728 (N_728,In_31,In_296);
xnor U729 (N_729,In_553,In_747);
xnor U730 (N_730,In_2249,In_187);
nand U731 (N_731,In_370,In_1507);
xnor U732 (N_732,In_148,In_1718);
xnor U733 (N_733,In_430,In_1577);
nor U734 (N_734,In_21,In_1400);
nor U735 (N_735,In_405,In_1957);
nor U736 (N_736,In_1098,In_1819);
xnor U737 (N_737,In_1784,In_1514);
xor U738 (N_738,In_1527,In_754);
xnor U739 (N_739,In_2482,In_267);
nand U740 (N_740,In_1949,In_1699);
or U741 (N_741,In_1785,In_1797);
nand U742 (N_742,In_1966,In_149);
or U743 (N_743,In_1352,In_1120);
and U744 (N_744,In_2111,In_496);
or U745 (N_745,In_271,In_1198);
and U746 (N_746,In_456,In_997);
xor U747 (N_747,In_36,In_205);
nand U748 (N_748,In_186,In_2053);
and U749 (N_749,In_1585,In_1353);
or U750 (N_750,In_1943,In_436);
and U751 (N_751,In_672,In_1498);
and U752 (N_752,In_693,In_2082);
or U753 (N_753,In_43,In_650);
nand U754 (N_754,In_144,In_1526);
nand U755 (N_755,In_1724,In_943);
and U756 (N_756,In_1795,In_2006);
or U757 (N_757,In_354,In_2279);
nor U758 (N_758,In_491,In_1728);
xor U759 (N_759,In_1705,In_185);
or U760 (N_760,In_1422,In_1240);
nand U761 (N_761,In_2074,In_1412);
or U762 (N_762,In_1570,In_2203);
xnor U763 (N_763,In_179,In_2269);
nor U764 (N_764,In_1542,In_1629);
nand U765 (N_765,In_1873,In_1591);
nand U766 (N_766,In_1882,In_1994);
nor U767 (N_767,In_1173,In_1757);
xnor U768 (N_768,In_2368,In_946);
or U769 (N_769,In_462,In_950);
xor U770 (N_770,In_1304,In_717);
and U771 (N_771,In_965,In_1543);
xnor U772 (N_772,In_669,In_1562);
nand U773 (N_773,In_2107,In_1555);
or U774 (N_774,In_1452,In_2189);
and U775 (N_775,In_1104,In_2044);
nand U776 (N_776,In_790,In_1041);
xor U777 (N_777,In_478,In_109);
nand U778 (N_778,In_1244,In_1831);
and U779 (N_779,In_2291,In_112);
nand U780 (N_780,In_651,In_406);
or U781 (N_781,In_2404,In_1671);
or U782 (N_782,In_1701,In_529);
xor U783 (N_783,In_518,In_17);
nand U784 (N_784,In_2396,In_788);
xor U785 (N_785,In_667,In_708);
nor U786 (N_786,In_2406,In_358);
and U787 (N_787,In_2392,In_1766);
and U788 (N_788,In_290,In_695);
xor U789 (N_789,In_1311,In_2360);
or U790 (N_790,In_1762,In_142);
xnor U791 (N_791,In_599,In_975);
nor U792 (N_792,In_2241,In_889);
nor U793 (N_793,In_227,In_937);
xor U794 (N_794,In_1139,In_1729);
nor U795 (N_795,In_2379,In_1806);
or U796 (N_796,In_1602,In_2454);
or U797 (N_797,In_396,In_1245);
xnor U798 (N_798,In_1290,In_2440);
nor U799 (N_799,In_146,In_504);
nand U800 (N_800,In_60,In_1413);
nor U801 (N_801,In_1291,In_852);
and U802 (N_802,In_804,In_1329);
nand U803 (N_803,In_2248,In_930);
and U804 (N_804,In_800,In_985);
nand U805 (N_805,In_102,In_115);
and U806 (N_806,In_2311,In_2442);
or U807 (N_807,In_266,In_766);
and U808 (N_808,In_471,In_2131);
nor U809 (N_809,In_783,In_665);
nor U810 (N_810,In_1979,In_2421);
or U811 (N_811,In_1620,In_1231);
nand U812 (N_812,In_2022,In_654);
nand U813 (N_813,In_1808,In_785);
and U814 (N_814,In_2499,In_945);
and U815 (N_815,In_1293,In_578);
xnor U816 (N_816,In_1826,In_1670);
or U817 (N_817,In_1115,In_1394);
and U818 (N_818,In_2011,In_2486);
and U819 (N_819,In_884,In_388);
or U820 (N_820,In_1371,In_2468);
and U821 (N_821,In_1598,In_509);
or U822 (N_822,In_423,In_2321);
or U823 (N_823,In_2240,In_184);
nor U824 (N_824,In_2496,In_393);
nand U825 (N_825,In_2480,In_1182);
nor U826 (N_826,In_662,In_957);
or U827 (N_827,In_580,In_760);
and U828 (N_828,In_548,In_197);
and U829 (N_829,In_530,In_1134);
and U830 (N_830,In_1170,In_1116);
nand U831 (N_831,In_1206,In_280);
and U832 (N_832,In_988,In_1374);
xnor U833 (N_833,In_1399,In_1486);
nor U834 (N_834,In_568,In_1517);
nand U835 (N_835,In_348,In_368);
nand U836 (N_836,In_990,In_616);
or U837 (N_837,In_95,In_1126);
nand U838 (N_838,In_832,In_127);
nand U839 (N_839,In_679,In_1212);
nor U840 (N_840,In_2108,In_1657);
nand U841 (N_841,In_1818,In_1123);
and U842 (N_842,In_701,In_2103);
nor U843 (N_843,In_556,In_961);
and U844 (N_844,In_1019,In_312);
nor U845 (N_845,In_919,In_1325);
or U846 (N_846,In_1639,In_1071);
nand U847 (N_847,In_1927,In_1580);
or U848 (N_848,In_412,In_555);
or U849 (N_849,In_2256,In_2014);
xnor U850 (N_850,In_1493,In_1569);
nand U851 (N_851,In_1998,In_1332);
and U852 (N_852,In_1079,In_2231);
xor U853 (N_853,In_1363,In_2293);
nor U854 (N_854,In_1309,In_1599);
or U855 (N_855,In_2062,In_64);
nand U856 (N_856,In_2114,In_1000);
or U857 (N_857,In_25,In_363);
nand U858 (N_858,In_2028,In_1706);
nor U859 (N_859,In_54,In_1939);
and U860 (N_860,In_1790,In_1494);
and U861 (N_861,In_1100,In_1668);
xnor U862 (N_862,In_1466,In_1435);
nand U863 (N_863,In_1154,In_1335);
nor U864 (N_864,In_105,In_831);
xnor U865 (N_865,In_492,In_129);
and U866 (N_866,In_147,In_770);
nor U867 (N_867,In_912,In_894);
and U868 (N_868,In_1838,In_1187);
xnor U869 (N_869,In_1674,In_2010);
or U870 (N_870,In_104,In_1588);
nor U871 (N_871,In_1448,In_1503);
nand U872 (N_872,In_2494,In_261);
and U873 (N_873,In_2047,In_1421);
xor U874 (N_874,In_1989,In_313);
xnor U875 (N_875,In_1603,In_2435);
xor U876 (N_876,In_1464,In_1740);
and U877 (N_877,In_1687,In_1564);
and U878 (N_878,In_1076,In_1865);
nand U879 (N_879,In_2177,In_365);
nand U880 (N_880,In_2056,In_2461);
nor U881 (N_881,In_2446,In_1454);
xor U882 (N_882,In_1563,In_1064);
nand U883 (N_883,In_2453,In_1722);
nor U884 (N_884,In_2449,In_2452);
xnor U885 (N_885,In_2015,In_2064);
nand U886 (N_886,In_600,In_2445);
xnor U887 (N_887,In_1536,In_2018);
xnor U888 (N_888,In_703,In_1821);
and U889 (N_889,In_2477,In_2443);
xor U890 (N_890,In_2422,In_851);
nand U891 (N_891,In_2088,In_341);
and U892 (N_892,In_751,In_2181);
nor U893 (N_893,In_22,In_1418);
or U894 (N_894,In_973,In_1236);
nor U895 (N_895,In_106,In_2200);
nand U896 (N_896,In_213,In_1337);
and U897 (N_897,In_325,In_1445);
and U898 (N_898,In_842,In_1031);
nand U899 (N_899,In_635,In_2469);
or U900 (N_900,In_274,In_888);
xnor U901 (N_901,In_256,In_2417);
nor U902 (N_902,In_1061,In_2371);
and U903 (N_903,In_1691,In_1915);
nand U904 (N_904,In_2159,In_2313);
and U905 (N_905,In_1028,In_817);
or U906 (N_906,In_1269,In_2450);
xnor U907 (N_907,In_145,In_1716);
xnor U908 (N_908,In_2167,In_1110);
xor U909 (N_909,In_1375,In_391);
and U910 (N_910,In_1804,In_618);
nor U911 (N_911,In_928,In_1848);
or U912 (N_912,In_2066,In_2085);
or U913 (N_913,In_1920,In_2253);
xnor U914 (N_914,In_2476,In_626);
nor U915 (N_915,In_565,In_866);
or U916 (N_916,In_1274,In_2390);
nand U917 (N_917,In_82,In_1697);
nor U918 (N_918,In_1534,In_566);
or U919 (N_919,In_1692,In_335);
xnor U920 (N_920,In_1008,In_1976);
xor U921 (N_921,In_122,In_299);
xnor U922 (N_922,In_966,In_859);
or U923 (N_923,In_938,In_1248);
xor U924 (N_924,In_1970,In_1016);
xor U925 (N_925,In_1725,In_319);
nand U926 (N_926,In_607,In_2046);
nor U927 (N_927,In_1595,In_397);
nand U928 (N_928,In_1717,In_2040);
or U929 (N_929,In_242,In_1863);
or U930 (N_930,In_920,In_1241);
and U931 (N_931,In_154,In_2195);
nand U932 (N_932,In_2223,In_2319);
xor U933 (N_933,In_2247,In_1307);
or U934 (N_934,In_2139,In_1678);
nor U935 (N_935,In_968,In_1916);
nand U936 (N_936,In_2385,In_2315);
and U937 (N_937,In_1973,In_1812);
and U938 (N_938,In_2384,In_674);
nor U939 (N_939,In_1246,In_1610);
xnor U940 (N_940,In_776,In_241);
or U941 (N_941,In_1037,In_2273);
xnor U942 (N_942,In_564,In_1053);
or U943 (N_943,In_2441,In_1793);
or U944 (N_944,In_1243,In_763);
and U945 (N_945,In_1411,In_1080);
nor U946 (N_946,In_1601,In_2142);
or U947 (N_947,In_791,In_898);
or U948 (N_948,In_2266,In_2278);
nor U949 (N_949,In_2405,In_2343);
and U950 (N_950,In_2408,In_1854);
nor U951 (N_951,In_2464,In_562);
nand U952 (N_952,In_1475,In_2407);
xnor U953 (N_953,In_340,In_1107);
or U954 (N_954,In_686,In_1255);
nor U955 (N_955,In_2043,In_1137);
xor U956 (N_956,In_659,In_2073);
and U957 (N_957,In_869,In_138);
or U958 (N_958,In_959,In_1852);
or U959 (N_959,In_1222,In_2336);
nand U960 (N_960,In_2036,In_2196);
xor U961 (N_961,In_1886,In_2170);
nor U962 (N_962,In_1781,In_1820);
xnor U963 (N_963,In_1799,In_603);
and U964 (N_964,In_419,In_1387);
xor U965 (N_965,In_606,In_714);
nor U966 (N_966,In_2301,In_2372);
and U967 (N_967,In_181,In_671);
and U968 (N_968,In_1065,In_1666);
nor U969 (N_969,In_764,In_61);
and U970 (N_970,In_2484,In_329);
xnor U971 (N_971,In_2263,In_2415);
xnor U972 (N_972,In_1217,In_1117);
xor U973 (N_973,In_604,In_987);
and U974 (N_974,In_1415,In_240);
and U975 (N_975,In_1983,In_1185);
nor U976 (N_976,In_850,In_1538);
xnor U977 (N_977,In_1612,In_1124);
nor U978 (N_978,In_2199,In_1002);
nor U979 (N_979,In_1929,In_310);
xor U980 (N_980,In_1837,In_1584);
xnor U981 (N_981,In_2077,In_311);
and U982 (N_982,In_2338,In_644);
nand U983 (N_983,In_246,In_1715);
and U984 (N_984,In_524,In_376);
or U985 (N_985,In_823,In_153);
nor U986 (N_986,In_258,In_2179);
or U987 (N_987,In_244,In_2259);
xnor U988 (N_988,In_1978,In_1892);
xnor U989 (N_989,In_963,In_215);
and U990 (N_990,In_1590,In_1626);
or U991 (N_991,In_1262,In_1794);
or U992 (N_992,In_0,In_136);
and U993 (N_993,In_1036,In_704);
nand U994 (N_994,In_1165,In_839);
and U995 (N_995,In_485,In_1159);
nand U996 (N_996,In_424,In_2366);
and U997 (N_997,In_1817,In_1026);
and U998 (N_998,In_1238,In_1597);
xnor U999 (N_999,In_1646,In_1923);
nor U1000 (N_1000,In_847,In_1997);
xor U1001 (N_1001,In_2209,In_180);
xor U1002 (N_1002,In_65,In_552);
xor U1003 (N_1003,In_815,In_1960);
xnor U1004 (N_1004,In_263,In_1341);
xor U1005 (N_1005,In_2458,In_1615);
and U1006 (N_1006,In_1782,In_1531);
nand U1007 (N_1007,In_1940,In_1438);
nor U1008 (N_1008,In_1389,In_2029);
nand U1009 (N_1009,In_1237,In_1457);
xor U1010 (N_1010,In_1225,In_2239);
nand U1011 (N_1011,In_265,In_757);
nor U1012 (N_1012,In_1459,In_2078);
nand U1013 (N_1013,In_537,In_322);
or U1014 (N_1014,In_486,In_1482);
nand U1015 (N_1015,In_855,In_2173);
nand U1016 (N_1016,In_1700,In_1017);
and U1017 (N_1017,In_1303,In_141);
and U1018 (N_1018,In_1039,In_629);
xor U1019 (N_1019,In_567,In_2473);
and U1020 (N_1020,In_1521,In_210);
or U1021 (N_1021,In_2359,In_1306);
or U1022 (N_1022,In_2374,In_746);
xnor U1023 (N_1023,In_758,In_375);
and U1024 (N_1024,In_174,In_2333);
or U1025 (N_1025,In_1510,In_1504);
and U1026 (N_1026,In_1333,In_1133);
nand U1027 (N_1027,In_394,In_2238);
and U1028 (N_1028,In_2362,In_845);
xor U1029 (N_1029,In_1532,In_2237);
xnor U1030 (N_1030,In_947,In_1391);
nand U1031 (N_1031,In_2326,In_2083);
or U1032 (N_1032,In_1774,In_1623);
nand U1033 (N_1033,In_877,In_62);
xnor U1034 (N_1034,In_511,In_356);
xor U1035 (N_1035,In_1730,In_925);
and U1036 (N_1036,In_779,In_47);
nand U1037 (N_1037,In_2169,In_226);
nand U1038 (N_1038,In_440,In_130);
nand U1039 (N_1039,In_1672,In_586);
or U1040 (N_1040,In_1365,In_1103);
nor U1041 (N_1041,In_1992,In_1128);
nor U1042 (N_1042,In_982,In_2255);
xor U1043 (N_1043,In_2061,In_2102);
nor U1044 (N_1044,In_705,In_1094);
xnor U1045 (N_1045,In_264,In_1361);
xor U1046 (N_1046,In_1605,In_1932);
xor U1047 (N_1047,In_2490,In_1719);
nand U1048 (N_1048,In_1727,In_255);
or U1049 (N_1049,In_1109,In_692);
nand U1050 (N_1050,In_2183,In_2289);
and U1051 (N_1051,In_372,In_351);
nor U1052 (N_1052,In_1351,In_837);
nor U1053 (N_1053,In_101,In_196);
nand U1054 (N_1054,In_94,In_582);
and U1055 (N_1055,In_11,In_1658);
and U1056 (N_1056,In_304,In_1685);
and U1057 (N_1057,In_1746,In_1772);
xnor U1058 (N_1058,In_1761,In_408);
nand U1059 (N_1059,In_608,In_1084);
nor U1060 (N_1060,In_320,In_1419);
nand U1061 (N_1061,In_1788,In_1967);
nand U1062 (N_1062,In_2498,In_2121);
and U1063 (N_1063,In_876,In_1634);
nor U1064 (N_1064,In_34,In_1783);
nand U1065 (N_1065,In_1655,In_1441);
nor U1066 (N_1066,In_543,In_2270);
or U1067 (N_1067,In_77,In_722);
or U1068 (N_1068,In_2035,In_1410);
nor U1069 (N_1069,In_176,In_1227);
and U1070 (N_1070,In_1987,In_655);
and U1071 (N_1071,In_1828,In_2002);
and U1072 (N_1072,In_1609,In_1867);
nand U1073 (N_1073,In_418,In_458);
xor U1074 (N_1074,In_649,In_1006);
xnor U1075 (N_1075,In_863,In_1196);
xor U1076 (N_1076,In_2287,In_1853);
and U1077 (N_1077,In_273,In_2306);
or U1078 (N_1078,In_1081,In_175);
nor U1079 (N_1079,In_1151,In_892);
xnor U1080 (N_1080,In_1461,In_934);
and U1081 (N_1081,In_415,In_1515);
nor U1082 (N_1082,In_1554,In_551);
xor U1083 (N_1083,In_1149,In_2039);
and U1084 (N_1084,In_2218,In_890);
nand U1085 (N_1085,In_1572,In_1850);
and U1086 (N_1086,In_1397,In_1186);
or U1087 (N_1087,In_893,In_1455);
xor U1088 (N_1088,In_2411,In_2460);
xnor U1089 (N_1089,In_2153,In_1190);
or U1090 (N_1090,In_1228,In_886);
nor U1091 (N_1091,In_951,In_231);
nor U1092 (N_1092,In_1177,In_137);
and U1093 (N_1093,In_768,In_2140);
nor U1094 (N_1094,In_1088,In_159);
nand U1095 (N_1095,In_490,In_1377);
nor U1096 (N_1096,In_1953,In_98);
xor U1097 (N_1097,In_411,In_2353);
nor U1098 (N_1098,In_156,In_1934);
xnor U1099 (N_1099,In_2388,In_2211);
xor U1100 (N_1100,In_532,In_1593);
xnor U1101 (N_1101,In_558,In_1582);
xnor U1102 (N_1102,In_1256,In_970);
nor U1103 (N_1103,In_2444,In_1414);
and U1104 (N_1104,In_228,In_522);
xor U1105 (N_1105,In_1034,In_1296);
or U1106 (N_1106,In_2412,In_1704);
or U1107 (N_1107,In_2001,In_201);
or U1108 (N_1108,In_995,In_347);
xnor U1109 (N_1109,In_1465,In_2217);
and U1110 (N_1110,In_1518,In_972);
and U1111 (N_1111,In_927,In_29);
nand U1112 (N_1112,In_1488,In_203);
or U1113 (N_1113,In_780,In_924);
nor U1114 (N_1114,In_2252,In_234);
and U1115 (N_1115,In_1736,In_846);
nor U1116 (N_1116,In_2420,In_1087);
and U1117 (N_1117,In_2055,In_1696);
and U1118 (N_1118,In_1964,In_295);
xor U1119 (N_1119,In_1342,In_1347);
and U1120 (N_1120,In_362,In_2008);
and U1121 (N_1121,In_520,In_1302);
xnor U1122 (N_1122,In_595,In_1869);
nor U1123 (N_1123,In_1763,In_103);
xnor U1124 (N_1124,In_2168,In_1143);
nand U1125 (N_1125,In_93,In_948);
and U1126 (N_1126,In_434,In_2410);
nor U1127 (N_1127,In_868,In_1883);
nor U1128 (N_1128,In_593,In_2430);
and U1129 (N_1129,In_7,In_2158);
and U1130 (N_1130,In_1890,In_2143);
nor U1131 (N_1131,In_2391,In_1403);
nand U1132 (N_1132,In_1520,In_1249);
xor U1133 (N_1133,In_2220,In_1160);
nand U1134 (N_1134,In_2135,In_1505);
xor U1135 (N_1135,In_338,In_867);
and U1136 (N_1136,In_1648,In_1571);
and U1137 (N_1137,In_646,In_1074);
nand U1138 (N_1138,In_83,In_1428);
xor U1139 (N_1139,In_571,In_2434);
or U1140 (N_1140,In_1712,In_488);
and U1141 (N_1141,In_1483,In_1125);
nand U1142 (N_1142,In_81,In_2216);
xnor U1143 (N_1143,In_463,In_221);
nor U1144 (N_1144,In_364,In_1899);
or U1145 (N_1145,In_1202,In_1755);
or U1146 (N_1146,In_741,In_728);
or U1147 (N_1147,In_1513,In_1801);
nor U1148 (N_1148,In_2184,In_206);
nand U1149 (N_1149,In_139,In_2431);
and U1150 (N_1150,In_1856,In_450);
or U1151 (N_1151,In_2172,In_447);
nand U1152 (N_1152,In_2455,In_547);
or U1153 (N_1153,In_2320,In_700);
xnor U1154 (N_1154,In_1816,In_1984);
nor U1155 (N_1155,In_1575,In_502);
nor U1156 (N_1156,In_2086,In_2347);
xor U1157 (N_1157,In_1007,In_2038);
and U1158 (N_1158,In_2322,In_1437);
nand U1159 (N_1159,In_2364,In_284);
xnor U1160 (N_1160,In_1633,In_1496);
and U1161 (N_1161,In_2128,In_2057);
xnor U1162 (N_1162,In_2125,In_1047);
nor U1163 (N_1163,In_19,In_840);
nand U1164 (N_1164,In_2192,In_2459);
or U1165 (N_1165,In_377,In_177);
and U1166 (N_1166,In_796,In_2117);
nor U1167 (N_1167,In_664,In_160);
or U1168 (N_1168,In_1148,In_601);
nand U1169 (N_1169,In_1985,In_998);
and U1170 (N_1170,In_584,In_1204);
nor U1171 (N_1171,In_689,In_155);
nand U1172 (N_1172,In_856,In_72);
nor U1173 (N_1173,In_420,In_1681);
or U1174 (N_1174,In_2413,In_1271);
xor U1175 (N_1175,In_2316,In_1276);
and U1176 (N_1176,In_222,In_1122);
nor U1177 (N_1177,In_1631,In_2299);
and U1178 (N_1178,In_781,In_1737);
xor U1179 (N_1179,In_1253,In_1106);
nand U1180 (N_1180,In_1234,In_1313);
and U1181 (N_1181,In_1861,In_1102);
and U1182 (N_1182,In_2350,In_1560);
or U1183 (N_1183,In_259,In_1905);
or U1184 (N_1184,In_1060,In_472);
and U1185 (N_1185,In_1158,In_2424);
nor U1186 (N_1186,In_691,In_838);
xor U1187 (N_1187,In_42,In_1885);
or U1188 (N_1188,In_294,In_2221);
and U1189 (N_1189,In_978,In_1617);
and U1190 (N_1190,In_2334,In_413);
nand U1191 (N_1191,In_1141,In_387);
nor U1192 (N_1192,In_32,In_721);
xnor U1193 (N_1193,In_211,In_2020);
or U1194 (N_1194,In_2271,In_1344);
and U1195 (N_1195,In_1174,In_1327);
nor U1196 (N_1196,In_2205,In_1769);
xor U1197 (N_1197,In_69,In_1540);
and U1198 (N_1198,In_1156,In_526);
nor U1199 (N_1199,In_1550,In_645);
and U1200 (N_1200,In_521,In_2466);
xor U1201 (N_1201,In_2296,In_2448);
xnor U1202 (N_1202,In_1708,In_1318);
xor U1203 (N_1203,In_1789,In_2304);
nor U1204 (N_1204,In_1169,In_2124);
xor U1205 (N_1205,In_1777,In_668);
xnor U1206 (N_1206,In_2051,In_2341);
nand U1207 (N_1207,In_805,In_1981);
nor U1208 (N_1208,In_1723,In_1070);
or U1209 (N_1209,In_314,In_1552);
nor U1210 (N_1210,In_2373,In_647);
or U1211 (N_1211,In_1119,In_343);
nor U1212 (N_1212,In_533,In_1567);
nand U1213 (N_1213,In_1444,In_1686);
nor U1214 (N_1214,In_1530,In_1168);
and U1215 (N_1215,In_2337,In_1298);
nor U1216 (N_1216,In_2233,In_1077);
xor U1217 (N_1217,In_1226,In_1519);
nand U1218 (N_1218,In_2485,In_2275);
nor U1219 (N_1219,In_2176,In_1491);
nand U1220 (N_1220,In_439,In_1058);
xor U1221 (N_1221,In_887,In_1698);
nor U1222 (N_1222,In_2465,In_150);
nand U1223 (N_1223,In_513,In_1689);
and U1224 (N_1224,In_1066,In_493);
nor U1225 (N_1225,In_435,In_872);
and U1226 (N_1226,In_614,In_2027);
and U1227 (N_1227,In_399,In_2409);
nor U1228 (N_1228,In_2175,In_1398);
nand U1229 (N_1229,In_220,In_996);
and U1230 (N_1230,In_2146,In_1178);
xnor U1231 (N_1231,In_2308,In_775);
xor U1232 (N_1232,In_801,In_1089);
or U1233 (N_1233,In_962,In_474);
xnor U1234 (N_1234,In_1268,In_2277);
and U1235 (N_1235,In_369,In_1224);
and U1236 (N_1236,In_853,In_2309);
or U1237 (N_1237,In_2317,In_247);
and U1238 (N_1238,In_167,In_23);
or U1239 (N_1239,In_1653,In_229);
nor U1240 (N_1240,In_1013,In_74);
xor U1241 (N_1241,In_546,In_2133);
or U1242 (N_1242,In_1864,In_1745);
xor U1243 (N_1243,In_1434,In_1162);
nor U1244 (N_1244,In_151,In_1628);
and U1245 (N_1245,In_1688,In_517);
nor U1246 (N_1246,In_2251,In_981);
nand U1247 (N_1247,In_960,In_1381);
xnor U1248 (N_1248,In_1924,In_2245);
nor U1249 (N_1249,In_1456,In_232);
or U1250 (N_1250,In_815,In_1946);
xnor U1251 (N_1251,In_942,In_224);
nand U1252 (N_1252,In_1417,In_18);
nand U1253 (N_1253,In_1240,In_176);
or U1254 (N_1254,In_1514,In_1061);
xor U1255 (N_1255,In_1768,In_2333);
and U1256 (N_1256,In_1726,In_1164);
nor U1257 (N_1257,In_282,In_2347);
xnor U1258 (N_1258,In_2449,In_1866);
or U1259 (N_1259,In_2317,In_336);
or U1260 (N_1260,In_1635,In_839);
xor U1261 (N_1261,In_1045,In_518);
and U1262 (N_1262,In_602,In_1050);
xnor U1263 (N_1263,In_250,In_1239);
and U1264 (N_1264,In_1180,In_215);
or U1265 (N_1265,In_305,In_1111);
or U1266 (N_1266,In_1393,In_261);
or U1267 (N_1267,In_525,In_945);
nand U1268 (N_1268,In_1692,In_7);
xnor U1269 (N_1269,In_206,In_641);
and U1270 (N_1270,In_1802,In_1761);
xor U1271 (N_1271,In_2474,In_988);
xor U1272 (N_1272,In_739,In_582);
and U1273 (N_1273,In_80,In_1816);
xor U1274 (N_1274,In_2426,In_2142);
or U1275 (N_1275,In_454,In_2433);
or U1276 (N_1276,In_2475,In_1524);
xor U1277 (N_1277,In_895,In_158);
nand U1278 (N_1278,In_568,In_646);
nand U1279 (N_1279,In_2282,In_2154);
xor U1280 (N_1280,In_2161,In_1751);
and U1281 (N_1281,In_1857,In_2116);
nor U1282 (N_1282,In_270,In_1110);
nor U1283 (N_1283,In_387,In_1382);
xor U1284 (N_1284,In_1089,In_91);
and U1285 (N_1285,In_1577,In_263);
nand U1286 (N_1286,In_2266,In_206);
xnor U1287 (N_1287,In_498,In_1137);
or U1288 (N_1288,In_1312,In_246);
or U1289 (N_1289,In_2479,In_392);
nand U1290 (N_1290,In_1429,In_1698);
xnor U1291 (N_1291,In_1170,In_505);
or U1292 (N_1292,In_752,In_216);
or U1293 (N_1293,In_848,In_1020);
nor U1294 (N_1294,In_2317,In_1294);
xor U1295 (N_1295,In_1183,In_1938);
and U1296 (N_1296,In_2292,In_2426);
or U1297 (N_1297,In_2386,In_2226);
and U1298 (N_1298,In_141,In_2254);
nand U1299 (N_1299,In_858,In_2093);
nand U1300 (N_1300,In_989,In_926);
nand U1301 (N_1301,In_2014,In_1455);
or U1302 (N_1302,In_1603,In_1446);
and U1303 (N_1303,In_1770,In_2179);
nor U1304 (N_1304,In_1704,In_514);
nor U1305 (N_1305,In_1312,In_1944);
nand U1306 (N_1306,In_1848,In_1208);
nor U1307 (N_1307,In_477,In_833);
xor U1308 (N_1308,In_2064,In_146);
and U1309 (N_1309,In_1979,In_349);
xor U1310 (N_1310,In_537,In_43);
xor U1311 (N_1311,In_1491,In_835);
xor U1312 (N_1312,In_641,In_1508);
or U1313 (N_1313,In_2463,In_583);
nand U1314 (N_1314,In_730,In_1080);
and U1315 (N_1315,In_1996,In_331);
nor U1316 (N_1316,In_1844,In_163);
and U1317 (N_1317,In_661,In_270);
or U1318 (N_1318,In_278,In_1628);
and U1319 (N_1319,In_1713,In_1679);
nor U1320 (N_1320,In_1441,In_1584);
xnor U1321 (N_1321,In_1199,In_63);
nor U1322 (N_1322,In_188,In_1747);
nor U1323 (N_1323,In_966,In_2257);
or U1324 (N_1324,In_292,In_2188);
nor U1325 (N_1325,In_915,In_302);
xnor U1326 (N_1326,In_1369,In_333);
xor U1327 (N_1327,In_2387,In_273);
nand U1328 (N_1328,In_457,In_1293);
and U1329 (N_1329,In_2340,In_1190);
nor U1330 (N_1330,In_2439,In_856);
xnor U1331 (N_1331,In_1271,In_2408);
and U1332 (N_1332,In_415,In_1047);
nor U1333 (N_1333,In_964,In_1662);
xnor U1334 (N_1334,In_2446,In_2438);
nor U1335 (N_1335,In_1424,In_1859);
xor U1336 (N_1336,In_2197,In_1757);
xnor U1337 (N_1337,In_396,In_200);
nor U1338 (N_1338,In_398,In_1037);
nand U1339 (N_1339,In_897,In_365);
nand U1340 (N_1340,In_1174,In_1598);
nand U1341 (N_1341,In_735,In_1895);
or U1342 (N_1342,In_1168,In_701);
xor U1343 (N_1343,In_2436,In_1155);
and U1344 (N_1344,In_1619,In_1312);
and U1345 (N_1345,In_925,In_54);
nor U1346 (N_1346,In_1040,In_524);
nor U1347 (N_1347,In_41,In_1541);
xnor U1348 (N_1348,In_1578,In_1280);
xor U1349 (N_1349,In_1932,In_1297);
nor U1350 (N_1350,In_2065,In_2280);
or U1351 (N_1351,In_1099,In_454);
or U1352 (N_1352,In_443,In_2118);
xnor U1353 (N_1353,In_1103,In_1973);
and U1354 (N_1354,In_1062,In_425);
nor U1355 (N_1355,In_244,In_680);
nor U1356 (N_1356,In_423,In_507);
nand U1357 (N_1357,In_487,In_2063);
nand U1358 (N_1358,In_92,In_1107);
and U1359 (N_1359,In_1570,In_2198);
nand U1360 (N_1360,In_559,In_703);
or U1361 (N_1361,In_480,In_725);
nor U1362 (N_1362,In_30,In_864);
xor U1363 (N_1363,In_1324,In_1628);
and U1364 (N_1364,In_1536,In_1841);
nor U1365 (N_1365,In_2055,In_2036);
nor U1366 (N_1366,In_479,In_1209);
xor U1367 (N_1367,In_366,In_1868);
or U1368 (N_1368,In_393,In_2400);
or U1369 (N_1369,In_761,In_462);
nand U1370 (N_1370,In_0,In_2207);
nor U1371 (N_1371,In_1330,In_2034);
and U1372 (N_1372,In_1096,In_1986);
nor U1373 (N_1373,In_2122,In_640);
xor U1374 (N_1374,In_836,In_251);
nand U1375 (N_1375,In_2293,In_2297);
nand U1376 (N_1376,In_316,In_1938);
nor U1377 (N_1377,In_184,In_2472);
nand U1378 (N_1378,In_2412,In_1749);
nor U1379 (N_1379,In_2236,In_1118);
and U1380 (N_1380,In_1473,In_2361);
or U1381 (N_1381,In_1344,In_432);
and U1382 (N_1382,In_1198,In_560);
xnor U1383 (N_1383,In_1652,In_1101);
nand U1384 (N_1384,In_486,In_92);
nand U1385 (N_1385,In_2311,In_103);
and U1386 (N_1386,In_1416,In_1588);
and U1387 (N_1387,In_1404,In_1317);
nand U1388 (N_1388,In_215,In_1927);
or U1389 (N_1389,In_1813,In_400);
nor U1390 (N_1390,In_249,In_1171);
nor U1391 (N_1391,In_515,In_2340);
or U1392 (N_1392,In_509,In_1472);
xnor U1393 (N_1393,In_2444,In_1469);
and U1394 (N_1394,In_204,In_2294);
nor U1395 (N_1395,In_1224,In_943);
nor U1396 (N_1396,In_2018,In_174);
and U1397 (N_1397,In_324,In_2152);
xor U1398 (N_1398,In_973,In_794);
xor U1399 (N_1399,In_1928,In_795);
and U1400 (N_1400,In_1679,In_1599);
nor U1401 (N_1401,In_1584,In_2394);
xnor U1402 (N_1402,In_252,In_1528);
or U1403 (N_1403,In_808,In_699);
nand U1404 (N_1404,In_2274,In_1503);
and U1405 (N_1405,In_271,In_2119);
nor U1406 (N_1406,In_933,In_2002);
nand U1407 (N_1407,In_1098,In_2369);
nand U1408 (N_1408,In_2210,In_583);
or U1409 (N_1409,In_1672,In_845);
nand U1410 (N_1410,In_522,In_1846);
nor U1411 (N_1411,In_1236,In_1830);
nor U1412 (N_1412,In_1355,In_872);
nand U1413 (N_1413,In_1858,In_1093);
and U1414 (N_1414,In_2343,In_1962);
nand U1415 (N_1415,In_681,In_1528);
xor U1416 (N_1416,In_1156,In_1284);
and U1417 (N_1417,In_1635,In_1083);
and U1418 (N_1418,In_1931,In_737);
nor U1419 (N_1419,In_1060,In_1953);
nor U1420 (N_1420,In_2356,In_1462);
and U1421 (N_1421,In_2304,In_613);
nand U1422 (N_1422,In_845,In_1666);
nand U1423 (N_1423,In_1928,In_1684);
or U1424 (N_1424,In_2125,In_558);
nand U1425 (N_1425,In_1517,In_62);
or U1426 (N_1426,In_1424,In_891);
and U1427 (N_1427,In_724,In_1775);
and U1428 (N_1428,In_1393,In_11);
and U1429 (N_1429,In_103,In_461);
and U1430 (N_1430,In_696,In_842);
nor U1431 (N_1431,In_2341,In_2271);
nor U1432 (N_1432,In_622,In_2332);
xor U1433 (N_1433,In_854,In_2266);
nor U1434 (N_1434,In_1000,In_2175);
nor U1435 (N_1435,In_1211,In_2477);
xor U1436 (N_1436,In_678,In_1372);
or U1437 (N_1437,In_2187,In_698);
nand U1438 (N_1438,In_282,In_630);
nand U1439 (N_1439,In_438,In_1437);
or U1440 (N_1440,In_2272,In_578);
nor U1441 (N_1441,In_698,In_1905);
nand U1442 (N_1442,In_1020,In_651);
nand U1443 (N_1443,In_722,In_447);
nor U1444 (N_1444,In_9,In_2355);
nand U1445 (N_1445,In_2471,In_262);
or U1446 (N_1446,In_1339,In_1633);
and U1447 (N_1447,In_2291,In_1921);
nor U1448 (N_1448,In_2259,In_1131);
and U1449 (N_1449,In_1136,In_946);
and U1450 (N_1450,In_866,In_1292);
nor U1451 (N_1451,In_383,In_301);
or U1452 (N_1452,In_583,In_1902);
and U1453 (N_1453,In_1188,In_1214);
and U1454 (N_1454,In_2176,In_1632);
nor U1455 (N_1455,In_471,In_980);
nor U1456 (N_1456,In_727,In_574);
and U1457 (N_1457,In_397,In_2184);
or U1458 (N_1458,In_1653,In_1140);
xor U1459 (N_1459,In_1844,In_692);
xnor U1460 (N_1460,In_1626,In_429);
nand U1461 (N_1461,In_658,In_723);
xor U1462 (N_1462,In_1792,In_2179);
nor U1463 (N_1463,In_512,In_816);
nor U1464 (N_1464,In_522,In_870);
xor U1465 (N_1465,In_2134,In_1322);
nand U1466 (N_1466,In_1135,In_1709);
xor U1467 (N_1467,In_1461,In_931);
nand U1468 (N_1468,In_2109,In_1262);
nand U1469 (N_1469,In_1375,In_995);
xnor U1470 (N_1470,In_714,In_1799);
nand U1471 (N_1471,In_410,In_1446);
or U1472 (N_1472,In_2284,In_1965);
xor U1473 (N_1473,In_1150,In_111);
nor U1474 (N_1474,In_931,In_1468);
nor U1475 (N_1475,In_440,In_1513);
nor U1476 (N_1476,In_2204,In_1171);
nand U1477 (N_1477,In_529,In_1953);
xor U1478 (N_1478,In_1963,In_1557);
or U1479 (N_1479,In_1157,In_2357);
and U1480 (N_1480,In_1441,In_1404);
and U1481 (N_1481,In_2002,In_1556);
nand U1482 (N_1482,In_738,In_1772);
nand U1483 (N_1483,In_1608,In_1590);
or U1484 (N_1484,In_60,In_190);
or U1485 (N_1485,In_577,In_1570);
and U1486 (N_1486,In_1430,In_845);
nor U1487 (N_1487,In_1042,In_2080);
nand U1488 (N_1488,In_696,In_628);
xnor U1489 (N_1489,In_2034,In_397);
nor U1490 (N_1490,In_1264,In_915);
nor U1491 (N_1491,In_1151,In_1307);
or U1492 (N_1492,In_1904,In_560);
or U1493 (N_1493,In_2486,In_434);
nand U1494 (N_1494,In_1806,In_2327);
xor U1495 (N_1495,In_2271,In_2024);
nor U1496 (N_1496,In_726,In_971);
xnor U1497 (N_1497,In_302,In_1694);
or U1498 (N_1498,In_1285,In_65);
or U1499 (N_1499,In_2255,In_712);
nand U1500 (N_1500,In_1906,In_47);
or U1501 (N_1501,In_1316,In_1766);
and U1502 (N_1502,In_2498,In_287);
or U1503 (N_1503,In_2118,In_1245);
nor U1504 (N_1504,In_569,In_1772);
nor U1505 (N_1505,In_1041,In_1860);
and U1506 (N_1506,In_334,In_1259);
or U1507 (N_1507,In_1814,In_1256);
xnor U1508 (N_1508,In_445,In_1934);
xnor U1509 (N_1509,In_1317,In_330);
nor U1510 (N_1510,In_979,In_517);
nand U1511 (N_1511,In_1713,In_2293);
or U1512 (N_1512,In_1641,In_1404);
nor U1513 (N_1513,In_2455,In_1091);
xor U1514 (N_1514,In_408,In_1658);
nand U1515 (N_1515,In_2109,In_2338);
and U1516 (N_1516,In_2440,In_1276);
nor U1517 (N_1517,In_1803,In_377);
and U1518 (N_1518,In_798,In_2414);
xor U1519 (N_1519,In_607,In_797);
or U1520 (N_1520,In_1002,In_1718);
or U1521 (N_1521,In_2278,In_2151);
nor U1522 (N_1522,In_1104,In_745);
and U1523 (N_1523,In_2002,In_1511);
and U1524 (N_1524,In_1744,In_1060);
nor U1525 (N_1525,In_538,In_1265);
or U1526 (N_1526,In_207,In_1307);
or U1527 (N_1527,In_1606,In_950);
nand U1528 (N_1528,In_169,In_2220);
nor U1529 (N_1529,In_281,In_295);
nor U1530 (N_1530,In_733,In_1545);
and U1531 (N_1531,In_967,In_340);
or U1532 (N_1532,In_2169,In_1817);
or U1533 (N_1533,In_246,In_1904);
xor U1534 (N_1534,In_1925,In_7);
nor U1535 (N_1535,In_791,In_1606);
nor U1536 (N_1536,In_1766,In_456);
nor U1537 (N_1537,In_2116,In_2145);
and U1538 (N_1538,In_2078,In_1360);
and U1539 (N_1539,In_1952,In_431);
and U1540 (N_1540,In_692,In_1789);
xnor U1541 (N_1541,In_30,In_821);
and U1542 (N_1542,In_744,In_1483);
xor U1543 (N_1543,In_199,In_1481);
nor U1544 (N_1544,In_1498,In_149);
nand U1545 (N_1545,In_822,In_2260);
nor U1546 (N_1546,In_1549,In_1211);
and U1547 (N_1547,In_394,In_877);
nor U1548 (N_1548,In_1288,In_554);
xnor U1549 (N_1549,In_2187,In_1331);
xnor U1550 (N_1550,In_779,In_883);
nor U1551 (N_1551,In_269,In_1265);
and U1552 (N_1552,In_797,In_2452);
nor U1553 (N_1553,In_795,In_617);
and U1554 (N_1554,In_2365,In_1500);
xor U1555 (N_1555,In_1535,In_902);
xnor U1556 (N_1556,In_2150,In_2053);
nor U1557 (N_1557,In_2335,In_683);
nor U1558 (N_1558,In_1620,In_187);
xnor U1559 (N_1559,In_765,In_2349);
nand U1560 (N_1560,In_558,In_1662);
nand U1561 (N_1561,In_2360,In_613);
nor U1562 (N_1562,In_339,In_873);
and U1563 (N_1563,In_527,In_2092);
nand U1564 (N_1564,In_2359,In_2393);
nand U1565 (N_1565,In_901,In_1516);
xor U1566 (N_1566,In_446,In_266);
or U1567 (N_1567,In_1584,In_2080);
nand U1568 (N_1568,In_2190,In_227);
xor U1569 (N_1569,In_1993,In_1706);
and U1570 (N_1570,In_163,In_1753);
or U1571 (N_1571,In_1810,In_1200);
or U1572 (N_1572,In_1751,In_862);
nor U1573 (N_1573,In_360,In_247);
and U1574 (N_1574,In_1045,In_1990);
xor U1575 (N_1575,In_1503,In_66);
or U1576 (N_1576,In_2365,In_575);
and U1577 (N_1577,In_34,In_240);
nand U1578 (N_1578,In_399,In_1135);
nand U1579 (N_1579,In_444,In_1564);
or U1580 (N_1580,In_1357,In_1666);
and U1581 (N_1581,In_1954,In_2218);
and U1582 (N_1582,In_907,In_2002);
and U1583 (N_1583,In_605,In_631);
nor U1584 (N_1584,In_2208,In_2472);
nand U1585 (N_1585,In_1929,In_1104);
nand U1586 (N_1586,In_719,In_277);
nor U1587 (N_1587,In_195,In_650);
nor U1588 (N_1588,In_1483,In_2498);
nand U1589 (N_1589,In_891,In_207);
nor U1590 (N_1590,In_700,In_1711);
or U1591 (N_1591,In_183,In_819);
xor U1592 (N_1592,In_2472,In_989);
and U1593 (N_1593,In_1620,In_941);
nor U1594 (N_1594,In_1840,In_36);
nor U1595 (N_1595,In_2072,In_2153);
nor U1596 (N_1596,In_1540,In_186);
nand U1597 (N_1597,In_91,In_1783);
nand U1598 (N_1598,In_171,In_1373);
xor U1599 (N_1599,In_521,In_848);
and U1600 (N_1600,In_1323,In_1411);
xor U1601 (N_1601,In_1757,In_2125);
and U1602 (N_1602,In_110,In_1421);
nor U1603 (N_1603,In_2237,In_1261);
nand U1604 (N_1604,In_2484,In_1014);
nand U1605 (N_1605,In_578,In_2156);
nor U1606 (N_1606,In_2345,In_834);
nand U1607 (N_1607,In_2441,In_1048);
xor U1608 (N_1608,In_1306,In_1672);
xnor U1609 (N_1609,In_1422,In_125);
and U1610 (N_1610,In_2103,In_1580);
nor U1611 (N_1611,In_899,In_1760);
nand U1612 (N_1612,In_169,In_2456);
and U1613 (N_1613,In_1129,In_1487);
nor U1614 (N_1614,In_1231,In_1713);
and U1615 (N_1615,In_1685,In_2045);
or U1616 (N_1616,In_1520,In_793);
and U1617 (N_1617,In_2474,In_2452);
and U1618 (N_1618,In_2198,In_549);
and U1619 (N_1619,In_764,In_1742);
and U1620 (N_1620,In_845,In_941);
nand U1621 (N_1621,In_1269,In_827);
nand U1622 (N_1622,In_2157,In_885);
and U1623 (N_1623,In_1597,In_15);
xor U1624 (N_1624,In_884,In_1079);
nand U1625 (N_1625,In_356,In_995);
or U1626 (N_1626,In_1608,In_2185);
nor U1627 (N_1627,In_832,In_2133);
and U1628 (N_1628,In_857,In_1296);
nor U1629 (N_1629,In_552,In_2211);
nor U1630 (N_1630,In_2297,In_2225);
and U1631 (N_1631,In_173,In_639);
or U1632 (N_1632,In_2354,In_1910);
nand U1633 (N_1633,In_2063,In_1465);
xnor U1634 (N_1634,In_423,In_2329);
and U1635 (N_1635,In_1062,In_175);
nand U1636 (N_1636,In_1751,In_1670);
xnor U1637 (N_1637,In_1370,In_374);
xnor U1638 (N_1638,In_2423,In_1651);
or U1639 (N_1639,In_2289,In_108);
xor U1640 (N_1640,In_1174,In_18);
or U1641 (N_1641,In_151,In_512);
nand U1642 (N_1642,In_1167,In_2318);
nand U1643 (N_1643,In_964,In_616);
xor U1644 (N_1644,In_855,In_1735);
or U1645 (N_1645,In_1155,In_991);
or U1646 (N_1646,In_2207,In_275);
or U1647 (N_1647,In_2273,In_1822);
nor U1648 (N_1648,In_482,In_894);
nand U1649 (N_1649,In_2162,In_30);
or U1650 (N_1650,In_950,In_2004);
nor U1651 (N_1651,In_218,In_342);
or U1652 (N_1652,In_470,In_447);
nand U1653 (N_1653,In_810,In_1531);
nand U1654 (N_1654,In_2359,In_2376);
nand U1655 (N_1655,In_1855,In_1442);
xor U1656 (N_1656,In_2051,In_2468);
or U1657 (N_1657,In_208,In_1265);
nand U1658 (N_1658,In_956,In_1516);
nand U1659 (N_1659,In_2128,In_1286);
nand U1660 (N_1660,In_1944,In_580);
nand U1661 (N_1661,In_1618,In_932);
or U1662 (N_1662,In_638,In_128);
and U1663 (N_1663,In_2150,In_531);
nand U1664 (N_1664,In_1016,In_1018);
and U1665 (N_1665,In_523,In_1026);
and U1666 (N_1666,In_1056,In_910);
nor U1667 (N_1667,In_2297,In_25);
nand U1668 (N_1668,In_1107,In_1466);
nor U1669 (N_1669,In_355,In_1733);
xor U1670 (N_1670,In_914,In_1195);
or U1671 (N_1671,In_270,In_790);
and U1672 (N_1672,In_1504,In_73);
nand U1673 (N_1673,In_2305,In_2047);
or U1674 (N_1674,In_2016,In_2450);
and U1675 (N_1675,In_1887,In_835);
or U1676 (N_1676,In_671,In_1489);
and U1677 (N_1677,In_1504,In_1654);
or U1678 (N_1678,In_526,In_2007);
nand U1679 (N_1679,In_1223,In_229);
xnor U1680 (N_1680,In_1323,In_904);
nor U1681 (N_1681,In_225,In_1166);
nand U1682 (N_1682,In_4,In_2102);
nand U1683 (N_1683,In_837,In_1622);
or U1684 (N_1684,In_422,In_1697);
nor U1685 (N_1685,In_2439,In_317);
nor U1686 (N_1686,In_9,In_939);
nand U1687 (N_1687,In_678,In_670);
nand U1688 (N_1688,In_678,In_1323);
and U1689 (N_1689,In_1585,In_1075);
or U1690 (N_1690,In_1552,In_2185);
nand U1691 (N_1691,In_1615,In_1461);
or U1692 (N_1692,In_13,In_269);
and U1693 (N_1693,In_861,In_1921);
or U1694 (N_1694,In_2198,In_630);
or U1695 (N_1695,In_278,In_723);
nand U1696 (N_1696,In_1596,In_180);
or U1697 (N_1697,In_1653,In_1743);
nand U1698 (N_1698,In_90,In_1388);
nor U1699 (N_1699,In_268,In_928);
nand U1700 (N_1700,In_2200,In_970);
nor U1701 (N_1701,In_703,In_90);
nor U1702 (N_1702,In_1028,In_765);
nand U1703 (N_1703,In_2250,In_1783);
nand U1704 (N_1704,In_1324,In_1141);
nor U1705 (N_1705,In_713,In_859);
and U1706 (N_1706,In_700,In_1257);
and U1707 (N_1707,In_1942,In_152);
or U1708 (N_1708,In_2096,In_2209);
and U1709 (N_1709,In_1059,In_27);
nand U1710 (N_1710,In_959,In_2147);
xor U1711 (N_1711,In_341,In_1336);
or U1712 (N_1712,In_2125,In_2449);
nand U1713 (N_1713,In_2289,In_608);
or U1714 (N_1714,In_1620,In_1158);
and U1715 (N_1715,In_1485,In_2426);
nor U1716 (N_1716,In_107,In_52);
xor U1717 (N_1717,In_2279,In_1086);
nand U1718 (N_1718,In_1297,In_1953);
or U1719 (N_1719,In_1650,In_498);
nand U1720 (N_1720,In_1974,In_1869);
or U1721 (N_1721,In_264,In_618);
nor U1722 (N_1722,In_1441,In_1145);
or U1723 (N_1723,In_1541,In_2075);
nand U1724 (N_1724,In_425,In_2231);
nand U1725 (N_1725,In_603,In_1530);
and U1726 (N_1726,In_1198,In_2228);
or U1727 (N_1727,In_1123,In_1399);
nand U1728 (N_1728,In_828,In_1845);
and U1729 (N_1729,In_1753,In_751);
nor U1730 (N_1730,In_2310,In_98);
and U1731 (N_1731,In_2053,In_2067);
nand U1732 (N_1732,In_1628,In_1644);
and U1733 (N_1733,In_2405,In_1742);
nor U1734 (N_1734,In_1032,In_459);
nand U1735 (N_1735,In_1763,In_907);
and U1736 (N_1736,In_1722,In_198);
xnor U1737 (N_1737,In_505,In_2381);
and U1738 (N_1738,In_368,In_1211);
and U1739 (N_1739,In_1573,In_352);
nor U1740 (N_1740,In_2317,In_1803);
nand U1741 (N_1741,In_593,In_1655);
and U1742 (N_1742,In_1818,In_1934);
xor U1743 (N_1743,In_1200,In_773);
xor U1744 (N_1744,In_2133,In_1528);
nand U1745 (N_1745,In_1324,In_744);
and U1746 (N_1746,In_1243,In_1903);
nand U1747 (N_1747,In_2196,In_1018);
or U1748 (N_1748,In_1735,In_1779);
nor U1749 (N_1749,In_679,In_269);
nor U1750 (N_1750,In_2125,In_707);
nor U1751 (N_1751,In_1085,In_2255);
or U1752 (N_1752,In_274,In_1384);
xor U1753 (N_1753,In_237,In_920);
xor U1754 (N_1754,In_2063,In_1332);
xnor U1755 (N_1755,In_574,In_1585);
nor U1756 (N_1756,In_549,In_1399);
and U1757 (N_1757,In_869,In_2248);
nand U1758 (N_1758,In_775,In_2244);
or U1759 (N_1759,In_1598,In_1513);
and U1760 (N_1760,In_2058,In_547);
nor U1761 (N_1761,In_1112,In_644);
and U1762 (N_1762,In_164,In_2465);
nand U1763 (N_1763,In_296,In_1802);
or U1764 (N_1764,In_2282,In_309);
nand U1765 (N_1765,In_809,In_1759);
or U1766 (N_1766,In_1220,In_1037);
nor U1767 (N_1767,In_367,In_1569);
xnor U1768 (N_1768,In_2430,In_1071);
xnor U1769 (N_1769,In_827,In_1743);
xnor U1770 (N_1770,In_670,In_2424);
nand U1771 (N_1771,In_1830,In_1661);
or U1772 (N_1772,In_2488,In_1459);
and U1773 (N_1773,In_1525,In_2179);
nor U1774 (N_1774,In_1865,In_1969);
nand U1775 (N_1775,In_2400,In_66);
or U1776 (N_1776,In_398,In_510);
nor U1777 (N_1777,In_926,In_226);
and U1778 (N_1778,In_795,In_1224);
xnor U1779 (N_1779,In_713,In_663);
or U1780 (N_1780,In_2201,In_204);
xnor U1781 (N_1781,In_669,In_2395);
nand U1782 (N_1782,In_2464,In_1505);
and U1783 (N_1783,In_2241,In_563);
xor U1784 (N_1784,In_1745,In_1749);
and U1785 (N_1785,In_1017,In_1834);
xor U1786 (N_1786,In_1026,In_1200);
and U1787 (N_1787,In_1915,In_1530);
xor U1788 (N_1788,In_1073,In_544);
and U1789 (N_1789,In_1792,In_377);
and U1790 (N_1790,In_87,In_1265);
nor U1791 (N_1791,In_736,In_747);
nor U1792 (N_1792,In_1497,In_565);
or U1793 (N_1793,In_1816,In_1339);
nor U1794 (N_1794,In_1014,In_2084);
xor U1795 (N_1795,In_1014,In_187);
and U1796 (N_1796,In_1573,In_1053);
and U1797 (N_1797,In_1515,In_2000);
and U1798 (N_1798,In_2371,In_2318);
or U1799 (N_1799,In_2337,In_329);
or U1800 (N_1800,In_143,In_2194);
xnor U1801 (N_1801,In_2425,In_552);
nand U1802 (N_1802,In_1227,In_610);
and U1803 (N_1803,In_845,In_1328);
nand U1804 (N_1804,In_380,In_2174);
or U1805 (N_1805,In_2196,In_1475);
nand U1806 (N_1806,In_890,In_90);
xor U1807 (N_1807,In_619,In_2191);
xor U1808 (N_1808,In_1372,In_1035);
or U1809 (N_1809,In_1379,In_1332);
and U1810 (N_1810,In_860,In_2335);
or U1811 (N_1811,In_1793,In_2213);
and U1812 (N_1812,In_2340,In_1);
nor U1813 (N_1813,In_2083,In_1135);
nor U1814 (N_1814,In_2421,In_2150);
and U1815 (N_1815,In_1429,In_490);
and U1816 (N_1816,In_1799,In_1955);
nor U1817 (N_1817,In_1254,In_151);
and U1818 (N_1818,In_1233,In_347);
xor U1819 (N_1819,In_435,In_777);
or U1820 (N_1820,In_922,In_323);
nor U1821 (N_1821,In_964,In_995);
or U1822 (N_1822,In_118,In_1561);
and U1823 (N_1823,In_804,In_497);
nand U1824 (N_1824,In_1187,In_1908);
or U1825 (N_1825,In_1994,In_1729);
or U1826 (N_1826,In_1008,In_1770);
or U1827 (N_1827,In_1626,In_1065);
nor U1828 (N_1828,In_1688,In_173);
and U1829 (N_1829,In_1061,In_1473);
nand U1830 (N_1830,In_1300,In_124);
and U1831 (N_1831,In_150,In_1575);
or U1832 (N_1832,In_2384,In_30);
nand U1833 (N_1833,In_1495,In_1030);
and U1834 (N_1834,In_146,In_1223);
or U1835 (N_1835,In_802,In_616);
or U1836 (N_1836,In_493,In_475);
xor U1837 (N_1837,In_2499,In_777);
and U1838 (N_1838,In_2389,In_1714);
nor U1839 (N_1839,In_1709,In_1790);
nand U1840 (N_1840,In_599,In_1695);
nor U1841 (N_1841,In_795,In_1974);
or U1842 (N_1842,In_2086,In_2247);
nor U1843 (N_1843,In_1336,In_1534);
xnor U1844 (N_1844,In_895,In_275);
nand U1845 (N_1845,In_219,In_2346);
nor U1846 (N_1846,In_188,In_1985);
nor U1847 (N_1847,In_624,In_273);
nand U1848 (N_1848,In_1512,In_2463);
or U1849 (N_1849,In_1077,In_1044);
or U1850 (N_1850,In_1789,In_2370);
xnor U1851 (N_1851,In_721,In_1533);
or U1852 (N_1852,In_593,In_1220);
and U1853 (N_1853,In_1175,In_2352);
xor U1854 (N_1854,In_1367,In_2468);
nand U1855 (N_1855,In_2369,In_507);
or U1856 (N_1856,In_2113,In_1516);
and U1857 (N_1857,In_2457,In_1674);
or U1858 (N_1858,In_1476,In_1266);
and U1859 (N_1859,In_794,In_1808);
or U1860 (N_1860,In_563,In_1677);
or U1861 (N_1861,In_61,In_1544);
nand U1862 (N_1862,In_944,In_1577);
nand U1863 (N_1863,In_2334,In_1583);
and U1864 (N_1864,In_1082,In_976);
or U1865 (N_1865,In_1595,In_1133);
nor U1866 (N_1866,In_1036,In_2392);
or U1867 (N_1867,In_547,In_115);
or U1868 (N_1868,In_1873,In_709);
and U1869 (N_1869,In_1858,In_643);
and U1870 (N_1870,In_1564,In_1563);
xor U1871 (N_1871,In_1505,In_1913);
and U1872 (N_1872,In_2031,In_1587);
xnor U1873 (N_1873,In_1838,In_618);
and U1874 (N_1874,In_2159,In_2356);
nand U1875 (N_1875,In_561,In_214);
and U1876 (N_1876,In_1753,In_264);
nand U1877 (N_1877,In_109,In_769);
nand U1878 (N_1878,In_639,In_1105);
xnor U1879 (N_1879,In_1003,In_1508);
xor U1880 (N_1880,In_1225,In_452);
xnor U1881 (N_1881,In_1042,In_2095);
and U1882 (N_1882,In_4,In_515);
xnor U1883 (N_1883,In_786,In_546);
or U1884 (N_1884,In_160,In_83);
and U1885 (N_1885,In_2463,In_2303);
xor U1886 (N_1886,In_1370,In_1264);
and U1887 (N_1887,In_820,In_818);
xor U1888 (N_1888,In_2380,In_1480);
and U1889 (N_1889,In_2018,In_507);
or U1890 (N_1890,In_884,In_2335);
xor U1891 (N_1891,In_454,In_632);
or U1892 (N_1892,In_229,In_89);
and U1893 (N_1893,In_1162,In_753);
and U1894 (N_1894,In_754,In_600);
nand U1895 (N_1895,In_1960,In_497);
or U1896 (N_1896,In_925,In_2223);
nor U1897 (N_1897,In_2065,In_2012);
nor U1898 (N_1898,In_85,In_1597);
nor U1899 (N_1899,In_769,In_1457);
nor U1900 (N_1900,In_2119,In_556);
nand U1901 (N_1901,In_119,In_1075);
or U1902 (N_1902,In_759,In_2239);
or U1903 (N_1903,In_1246,In_1496);
xor U1904 (N_1904,In_726,In_678);
nor U1905 (N_1905,In_1880,In_2021);
nand U1906 (N_1906,In_664,In_585);
nand U1907 (N_1907,In_1888,In_2219);
and U1908 (N_1908,In_1444,In_985);
nand U1909 (N_1909,In_1209,In_738);
or U1910 (N_1910,In_1278,In_2151);
or U1911 (N_1911,In_871,In_1174);
xor U1912 (N_1912,In_1349,In_2313);
and U1913 (N_1913,In_1867,In_1939);
xor U1914 (N_1914,In_2079,In_2413);
xnor U1915 (N_1915,In_539,In_2004);
nor U1916 (N_1916,In_2439,In_2135);
nand U1917 (N_1917,In_1158,In_1994);
xor U1918 (N_1918,In_2093,In_1504);
or U1919 (N_1919,In_1,In_1978);
and U1920 (N_1920,In_110,In_2469);
nor U1921 (N_1921,In_2114,In_2029);
nand U1922 (N_1922,In_1522,In_987);
nand U1923 (N_1923,In_44,In_981);
nand U1924 (N_1924,In_200,In_1274);
nand U1925 (N_1925,In_460,In_1988);
xor U1926 (N_1926,In_1400,In_2024);
and U1927 (N_1927,In_1010,In_1541);
or U1928 (N_1928,In_2409,In_190);
nand U1929 (N_1929,In_1559,In_1041);
nor U1930 (N_1930,In_2388,In_668);
and U1931 (N_1931,In_269,In_1253);
or U1932 (N_1932,In_33,In_674);
xor U1933 (N_1933,In_1245,In_2234);
and U1934 (N_1934,In_2394,In_2335);
or U1935 (N_1935,In_2102,In_1325);
nor U1936 (N_1936,In_1423,In_1829);
xor U1937 (N_1937,In_2359,In_1080);
and U1938 (N_1938,In_793,In_1137);
and U1939 (N_1939,In_2456,In_723);
xnor U1940 (N_1940,In_1274,In_964);
xor U1941 (N_1941,In_1032,In_2200);
xnor U1942 (N_1942,In_1572,In_486);
xor U1943 (N_1943,In_900,In_877);
xnor U1944 (N_1944,In_1658,In_2319);
nor U1945 (N_1945,In_2461,In_1682);
xnor U1946 (N_1946,In_466,In_164);
and U1947 (N_1947,In_909,In_1968);
and U1948 (N_1948,In_458,In_477);
nor U1949 (N_1949,In_1262,In_143);
and U1950 (N_1950,In_441,In_2167);
or U1951 (N_1951,In_888,In_404);
nor U1952 (N_1952,In_2068,In_1975);
xnor U1953 (N_1953,In_1884,In_1089);
and U1954 (N_1954,In_0,In_1245);
xor U1955 (N_1955,In_1149,In_1577);
nand U1956 (N_1956,In_708,In_1469);
and U1957 (N_1957,In_1281,In_1771);
nand U1958 (N_1958,In_276,In_154);
or U1959 (N_1959,In_1693,In_1966);
nor U1960 (N_1960,In_22,In_1922);
nor U1961 (N_1961,In_184,In_1683);
and U1962 (N_1962,In_1624,In_1218);
and U1963 (N_1963,In_643,In_1074);
xor U1964 (N_1964,In_2393,In_468);
nand U1965 (N_1965,In_472,In_1094);
xor U1966 (N_1966,In_1345,In_301);
and U1967 (N_1967,In_1129,In_153);
nand U1968 (N_1968,In_1772,In_1238);
or U1969 (N_1969,In_2038,In_445);
or U1970 (N_1970,In_2311,In_213);
and U1971 (N_1971,In_50,In_2335);
and U1972 (N_1972,In_2175,In_399);
and U1973 (N_1973,In_912,In_1948);
nor U1974 (N_1974,In_475,In_1618);
or U1975 (N_1975,In_1219,In_2039);
nor U1976 (N_1976,In_1886,In_757);
or U1977 (N_1977,In_1946,In_1264);
xnor U1978 (N_1978,In_1815,In_99);
and U1979 (N_1979,In_1966,In_2444);
xnor U1980 (N_1980,In_2030,In_2217);
and U1981 (N_1981,In_506,In_599);
or U1982 (N_1982,In_476,In_1175);
nor U1983 (N_1983,In_1479,In_1454);
nand U1984 (N_1984,In_2318,In_1824);
xor U1985 (N_1985,In_1391,In_836);
xnor U1986 (N_1986,In_1144,In_769);
nor U1987 (N_1987,In_2363,In_1295);
or U1988 (N_1988,In_169,In_191);
or U1989 (N_1989,In_126,In_1237);
xor U1990 (N_1990,In_467,In_1302);
or U1991 (N_1991,In_375,In_1391);
or U1992 (N_1992,In_691,In_678);
nand U1993 (N_1993,In_1090,In_1095);
nor U1994 (N_1994,In_1735,In_2262);
nor U1995 (N_1995,In_1236,In_55);
xor U1996 (N_1996,In_599,In_609);
nand U1997 (N_1997,In_805,In_54);
and U1998 (N_1998,In_588,In_2019);
xnor U1999 (N_1999,In_114,In_873);
xnor U2000 (N_2000,In_1865,In_721);
nor U2001 (N_2001,In_1040,In_2030);
or U2002 (N_2002,In_1392,In_800);
or U2003 (N_2003,In_1444,In_2054);
xnor U2004 (N_2004,In_1506,In_1591);
nand U2005 (N_2005,In_2191,In_22);
and U2006 (N_2006,In_2301,In_1528);
or U2007 (N_2007,In_1832,In_43);
and U2008 (N_2008,In_1217,In_1046);
xor U2009 (N_2009,In_1020,In_1120);
xnor U2010 (N_2010,In_384,In_2034);
nor U2011 (N_2011,In_1517,In_1013);
and U2012 (N_2012,In_156,In_2357);
nand U2013 (N_2013,In_1631,In_1766);
nor U2014 (N_2014,In_135,In_547);
or U2015 (N_2015,In_2049,In_528);
nor U2016 (N_2016,In_579,In_2491);
or U2017 (N_2017,In_401,In_969);
xnor U2018 (N_2018,In_2083,In_1951);
xor U2019 (N_2019,In_606,In_69);
or U2020 (N_2020,In_2374,In_794);
or U2021 (N_2021,In_2386,In_25);
nor U2022 (N_2022,In_1539,In_2331);
xor U2023 (N_2023,In_2411,In_605);
xnor U2024 (N_2024,In_1929,In_2154);
and U2025 (N_2025,In_333,In_1321);
xor U2026 (N_2026,In_158,In_1041);
nand U2027 (N_2027,In_689,In_1144);
nand U2028 (N_2028,In_1621,In_797);
and U2029 (N_2029,In_1506,In_919);
nor U2030 (N_2030,In_294,In_1137);
and U2031 (N_2031,In_2135,In_2290);
nand U2032 (N_2032,In_1741,In_334);
nand U2033 (N_2033,In_2349,In_1638);
or U2034 (N_2034,In_1833,In_1240);
nor U2035 (N_2035,In_690,In_289);
nor U2036 (N_2036,In_911,In_2128);
xnor U2037 (N_2037,In_1741,In_2459);
or U2038 (N_2038,In_971,In_1106);
nor U2039 (N_2039,In_1402,In_1558);
xor U2040 (N_2040,In_40,In_346);
and U2041 (N_2041,In_1031,In_2028);
xor U2042 (N_2042,In_1959,In_430);
or U2043 (N_2043,In_2034,In_2142);
nand U2044 (N_2044,In_871,In_2109);
xnor U2045 (N_2045,In_2313,In_1424);
nand U2046 (N_2046,In_901,In_1306);
xnor U2047 (N_2047,In_1497,In_1355);
nor U2048 (N_2048,In_1724,In_1850);
xor U2049 (N_2049,In_727,In_1677);
nor U2050 (N_2050,In_1542,In_1057);
xnor U2051 (N_2051,In_1983,In_1839);
nor U2052 (N_2052,In_878,In_1835);
nor U2053 (N_2053,In_1614,In_116);
and U2054 (N_2054,In_2458,In_2291);
nor U2055 (N_2055,In_1427,In_384);
nor U2056 (N_2056,In_1433,In_1613);
xor U2057 (N_2057,In_1884,In_948);
or U2058 (N_2058,In_563,In_2006);
nor U2059 (N_2059,In_2122,In_441);
and U2060 (N_2060,In_1000,In_1204);
and U2061 (N_2061,In_82,In_571);
and U2062 (N_2062,In_1688,In_508);
xnor U2063 (N_2063,In_1629,In_1194);
nand U2064 (N_2064,In_2450,In_1669);
nor U2065 (N_2065,In_862,In_1216);
nor U2066 (N_2066,In_1713,In_668);
nand U2067 (N_2067,In_2283,In_1846);
nor U2068 (N_2068,In_284,In_2402);
and U2069 (N_2069,In_2112,In_473);
and U2070 (N_2070,In_1226,In_161);
or U2071 (N_2071,In_1861,In_2142);
nor U2072 (N_2072,In_1047,In_1615);
nand U2073 (N_2073,In_2110,In_2425);
xor U2074 (N_2074,In_501,In_914);
xor U2075 (N_2075,In_2344,In_615);
xnor U2076 (N_2076,In_1421,In_2496);
nor U2077 (N_2077,In_1146,In_2374);
and U2078 (N_2078,In_1864,In_2023);
nor U2079 (N_2079,In_1912,In_839);
xor U2080 (N_2080,In_1706,In_552);
and U2081 (N_2081,In_1126,In_1339);
xnor U2082 (N_2082,In_730,In_766);
and U2083 (N_2083,In_622,In_2333);
nand U2084 (N_2084,In_784,In_2351);
and U2085 (N_2085,In_1686,In_1008);
nand U2086 (N_2086,In_1527,In_1529);
nor U2087 (N_2087,In_1433,In_1693);
or U2088 (N_2088,In_2161,In_2370);
nand U2089 (N_2089,In_249,In_1565);
nor U2090 (N_2090,In_769,In_2134);
and U2091 (N_2091,In_115,In_573);
xor U2092 (N_2092,In_856,In_2419);
and U2093 (N_2093,In_1114,In_2423);
nor U2094 (N_2094,In_1254,In_512);
nor U2095 (N_2095,In_1952,In_177);
or U2096 (N_2096,In_758,In_506);
xor U2097 (N_2097,In_12,In_1254);
and U2098 (N_2098,In_762,In_968);
and U2099 (N_2099,In_2084,In_31);
nand U2100 (N_2100,In_1856,In_755);
nor U2101 (N_2101,In_669,In_2226);
or U2102 (N_2102,In_1218,In_950);
nand U2103 (N_2103,In_853,In_1866);
xnor U2104 (N_2104,In_1836,In_49);
nor U2105 (N_2105,In_2230,In_1623);
and U2106 (N_2106,In_2021,In_1014);
nor U2107 (N_2107,In_620,In_2452);
xor U2108 (N_2108,In_2084,In_1252);
xor U2109 (N_2109,In_1892,In_2347);
and U2110 (N_2110,In_1293,In_1930);
nor U2111 (N_2111,In_1100,In_1149);
nand U2112 (N_2112,In_455,In_2011);
xnor U2113 (N_2113,In_401,In_41);
or U2114 (N_2114,In_1740,In_784);
and U2115 (N_2115,In_2008,In_1621);
nor U2116 (N_2116,In_2157,In_615);
xor U2117 (N_2117,In_688,In_1607);
nor U2118 (N_2118,In_2411,In_2295);
xor U2119 (N_2119,In_1191,In_1719);
xnor U2120 (N_2120,In_1609,In_2351);
and U2121 (N_2121,In_2200,In_685);
xor U2122 (N_2122,In_316,In_2365);
and U2123 (N_2123,In_2283,In_1147);
nand U2124 (N_2124,In_2421,In_1287);
and U2125 (N_2125,In_921,In_1777);
and U2126 (N_2126,In_820,In_903);
and U2127 (N_2127,In_302,In_2477);
xnor U2128 (N_2128,In_2215,In_1398);
or U2129 (N_2129,In_1020,In_230);
nand U2130 (N_2130,In_1239,In_2469);
nand U2131 (N_2131,In_1864,In_2371);
nor U2132 (N_2132,In_2172,In_523);
nand U2133 (N_2133,In_642,In_1675);
nor U2134 (N_2134,In_881,In_49);
or U2135 (N_2135,In_138,In_1041);
xor U2136 (N_2136,In_456,In_1324);
or U2137 (N_2137,In_502,In_451);
or U2138 (N_2138,In_139,In_1496);
xnor U2139 (N_2139,In_438,In_348);
or U2140 (N_2140,In_1890,In_2421);
and U2141 (N_2141,In_1552,In_1932);
nor U2142 (N_2142,In_69,In_543);
or U2143 (N_2143,In_1967,In_2323);
nor U2144 (N_2144,In_2278,In_1606);
nor U2145 (N_2145,In_2132,In_294);
nor U2146 (N_2146,In_1966,In_209);
xor U2147 (N_2147,In_2199,In_225);
nor U2148 (N_2148,In_71,In_2397);
xor U2149 (N_2149,In_902,In_1466);
xor U2150 (N_2150,In_1649,In_493);
nand U2151 (N_2151,In_1434,In_279);
nand U2152 (N_2152,In_1480,In_1158);
or U2153 (N_2153,In_1887,In_1286);
nor U2154 (N_2154,In_959,In_810);
nand U2155 (N_2155,In_1550,In_1067);
nor U2156 (N_2156,In_371,In_1897);
nor U2157 (N_2157,In_1623,In_922);
nand U2158 (N_2158,In_2479,In_2119);
xnor U2159 (N_2159,In_1887,In_1199);
or U2160 (N_2160,In_1938,In_1846);
and U2161 (N_2161,In_1748,In_1200);
and U2162 (N_2162,In_2403,In_113);
or U2163 (N_2163,In_2278,In_1291);
and U2164 (N_2164,In_1139,In_649);
nor U2165 (N_2165,In_390,In_1809);
xor U2166 (N_2166,In_1243,In_1440);
xor U2167 (N_2167,In_263,In_1486);
nand U2168 (N_2168,In_1780,In_2265);
nor U2169 (N_2169,In_1304,In_246);
xnor U2170 (N_2170,In_2155,In_1564);
or U2171 (N_2171,In_1703,In_1363);
and U2172 (N_2172,In_1162,In_1031);
xor U2173 (N_2173,In_894,In_1783);
xor U2174 (N_2174,In_1500,In_1874);
nand U2175 (N_2175,In_1664,In_1154);
xor U2176 (N_2176,In_339,In_2392);
nor U2177 (N_2177,In_250,In_2114);
or U2178 (N_2178,In_2295,In_531);
nor U2179 (N_2179,In_2131,In_1858);
xor U2180 (N_2180,In_2281,In_381);
nand U2181 (N_2181,In_469,In_401);
and U2182 (N_2182,In_1261,In_726);
nor U2183 (N_2183,In_693,In_1932);
nor U2184 (N_2184,In_886,In_541);
or U2185 (N_2185,In_1970,In_1793);
nor U2186 (N_2186,In_2325,In_1908);
nand U2187 (N_2187,In_832,In_2206);
and U2188 (N_2188,In_1776,In_1272);
xnor U2189 (N_2189,In_854,In_619);
and U2190 (N_2190,In_490,In_749);
nor U2191 (N_2191,In_1155,In_24);
nor U2192 (N_2192,In_1840,In_2223);
xor U2193 (N_2193,In_1673,In_1853);
and U2194 (N_2194,In_1644,In_242);
or U2195 (N_2195,In_1052,In_1207);
xnor U2196 (N_2196,In_2273,In_1031);
and U2197 (N_2197,In_2312,In_760);
nor U2198 (N_2198,In_177,In_1449);
and U2199 (N_2199,In_1474,In_1596);
xor U2200 (N_2200,In_118,In_1125);
or U2201 (N_2201,In_307,In_717);
nand U2202 (N_2202,In_758,In_1055);
nor U2203 (N_2203,In_2214,In_754);
or U2204 (N_2204,In_1542,In_240);
nor U2205 (N_2205,In_2174,In_432);
nand U2206 (N_2206,In_1282,In_512);
and U2207 (N_2207,In_1854,In_1893);
nor U2208 (N_2208,In_806,In_1902);
nor U2209 (N_2209,In_1624,In_865);
nand U2210 (N_2210,In_2398,In_1832);
xnor U2211 (N_2211,In_1503,In_2188);
or U2212 (N_2212,In_386,In_2337);
and U2213 (N_2213,In_45,In_702);
and U2214 (N_2214,In_650,In_228);
or U2215 (N_2215,In_1754,In_411);
xnor U2216 (N_2216,In_2181,In_818);
nand U2217 (N_2217,In_2306,In_2232);
xor U2218 (N_2218,In_2103,In_1710);
nand U2219 (N_2219,In_1216,In_1008);
nand U2220 (N_2220,In_2239,In_487);
nor U2221 (N_2221,In_1758,In_1523);
nor U2222 (N_2222,In_901,In_1983);
and U2223 (N_2223,In_1665,In_1802);
or U2224 (N_2224,In_959,In_2145);
nor U2225 (N_2225,In_2145,In_1566);
and U2226 (N_2226,In_1864,In_2418);
and U2227 (N_2227,In_141,In_380);
nand U2228 (N_2228,In_564,In_886);
or U2229 (N_2229,In_1474,In_1762);
or U2230 (N_2230,In_587,In_1815);
or U2231 (N_2231,In_600,In_429);
nand U2232 (N_2232,In_749,In_2355);
nand U2233 (N_2233,In_998,In_1053);
nand U2234 (N_2234,In_2172,In_2262);
nand U2235 (N_2235,In_2102,In_2384);
nor U2236 (N_2236,In_1038,In_2163);
nor U2237 (N_2237,In_1844,In_2295);
or U2238 (N_2238,In_438,In_919);
and U2239 (N_2239,In_1614,In_809);
nand U2240 (N_2240,In_2183,In_2324);
nor U2241 (N_2241,In_1921,In_210);
nand U2242 (N_2242,In_620,In_2457);
nand U2243 (N_2243,In_1334,In_1270);
xor U2244 (N_2244,In_2307,In_2297);
nor U2245 (N_2245,In_860,In_687);
and U2246 (N_2246,In_1138,In_152);
xor U2247 (N_2247,In_2037,In_1111);
xnor U2248 (N_2248,In_287,In_2106);
and U2249 (N_2249,In_1204,In_600);
nand U2250 (N_2250,In_96,In_2401);
xnor U2251 (N_2251,In_1433,In_23);
xnor U2252 (N_2252,In_2049,In_117);
xor U2253 (N_2253,In_1941,In_553);
nand U2254 (N_2254,In_1634,In_3);
nand U2255 (N_2255,In_210,In_363);
nor U2256 (N_2256,In_768,In_962);
nand U2257 (N_2257,In_1920,In_2275);
and U2258 (N_2258,In_2122,In_1825);
and U2259 (N_2259,In_2283,In_2459);
xnor U2260 (N_2260,In_1998,In_1944);
and U2261 (N_2261,In_2391,In_1003);
or U2262 (N_2262,In_2144,In_963);
or U2263 (N_2263,In_1688,In_2450);
xor U2264 (N_2264,In_1247,In_1514);
and U2265 (N_2265,In_1183,In_1292);
xor U2266 (N_2266,In_1841,In_336);
nor U2267 (N_2267,In_1843,In_1486);
xor U2268 (N_2268,In_128,In_2496);
nor U2269 (N_2269,In_33,In_908);
or U2270 (N_2270,In_1604,In_2370);
nor U2271 (N_2271,In_2159,In_956);
nor U2272 (N_2272,In_637,In_756);
and U2273 (N_2273,In_1796,In_1967);
and U2274 (N_2274,In_1348,In_1482);
and U2275 (N_2275,In_402,In_1106);
nor U2276 (N_2276,In_2331,In_1920);
nand U2277 (N_2277,In_2408,In_611);
nand U2278 (N_2278,In_417,In_1970);
xnor U2279 (N_2279,In_1889,In_2011);
nor U2280 (N_2280,In_885,In_2431);
xor U2281 (N_2281,In_1374,In_2048);
or U2282 (N_2282,In_1055,In_1812);
or U2283 (N_2283,In_2044,In_930);
nor U2284 (N_2284,In_2092,In_89);
nand U2285 (N_2285,In_361,In_205);
nor U2286 (N_2286,In_35,In_895);
xnor U2287 (N_2287,In_1849,In_2056);
nor U2288 (N_2288,In_2174,In_283);
xnor U2289 (N_2289,In_2174,In_1157);
nand U2290 (N_2290,In_234,In_854);
nand U2291 (N_2291,In_1748,In_1939);
and U2292 (N_2292,In_1547,In_1688);
or U2293 (N_2293,In_1612,In_1412);
nor U2294 (N_2294,In_496,In_1144);
and U2295 (N_2295,In_777,In_717);
or U2296 (N_2296,In_1731,In_134);
nor U2297 (N_2297,In_1077,In_819);
xor U2298 (N_2298,In_2388,In_2356);
nand U2299 (N_2299,In_1533,In_1823);
nand U2300 (N_2300,In_292,In_2169);
and U2301 (N_2301,In_1320,In_420);
nor U2302 (N_2302,In_1331,In_1890);
nand U2303 (N_2303,In_1165,In_1338);
nor U2304 (N_2304,In_1612,In_1475);
or U2305 (N_2305,In_210,In_402);
and U2306 (N_2306,In_996,In_1803);
nor U2307 (N_2307,In_706,In_246);
or U2308 (N_2308,In_52,In_2288);
nor U2309 (N_2309,In_1580,In_831);
or U2310 (N_2310,In_198,In_1000);
nand U2311 (N_2311,In_2193,In_1344);
nor U2312 (N_2312,In_681,In_1945);
xor U2313 (N_2313,In_765,In_1314);
nand U2314 (N_2314,In_253,In_1080);
or U2315 (N_2315,In_2385,In_1850);
nand U2316 (N_2316,In_1014,In_1634);
or U2317 (N_2317,In_2084,In_452);
or U2318 (N_2318,In_530,In_2008);
or U2319 (N_2319,In_1813,In_955);
xor U2320 (N_2320,In_2424,In_726);
xnor U2321 (N_2321,In_2232,In_2092);
and U2322 (N_2322,In_448,In_1794);
or U2323 (N_2323,In_627,In_243);
and U2324 (N_2324,In_821,In_1409);
xor U2325 (N_2325,In_1238,In_701);
and U2326 (N_2326,In_1391,In_2158);
xnor U2327 (N_2327,In_2185,In_2495);
xor U2328 (N_2328,In_1838,In_2012);
nor U2329 (N_2329,In_1496,In_657);
nand U2330 (N_2330,In_514,In_2226);
and U2331 (N_2331,In_1169,In_673);
and U2332 (N_2332,In_2208,In_789);
and U2333 (N_2333,In_435,In_32);
xor U2334 (N_2334,In_2235,In_1318);
nor U2335 (N_2335,In_193,In_1682);
or U2336 (N_2336,In_1308,In_342);
nor U2337 (N_2337,In_2090,In_535);
and U2338 (N_2338,In_798,In_2162);
nor U2339 (N_2339,In_1440,In_1912);
xor U2340 (N_2340,In_1941,In_1036);
or U2341 (N_2341,In_2165,In_532);
or U2342 (N_2342,In_2066,In_1863);
nand U2343 (N_2343,In_785,In_2039);
or U2344 (N_2344,In_1144,In_1890);
nor U2345 (N_2345,In_2449,In_561);
xor U2346 (N_2346,In_726,In_929);
and U2347 (N_2347,In_787,In_624);
nand U2348 (N_2348,In_500,In_1319);
or U2349 (N_2349,In_309,In_2042);
or U2350 (N_2350,In_1296,In_1166);
nand U2351 (N_2351,In_668,In_2360);
or U2352 (N_2352,In_1821,In_1048);
nor U2353 (N_2353,In_2074,In_820);
or U2354 (N_2354,In_618,In_734);
nand U2355 (N_2355,In_181,In_764);
xnor U2356 (N_2356,In_2463,In_807);
nand U2357 (N_2357,In_1653,In_1712);
and U2358 (N_2358,In_539,In_1060);
nand U2359 (N_2359,In_1860,In_1465);
or U2360 (N_2360,In_1393,In_2136);
nor U2361 (N_2361,In_1943,In_1744);
nor U2362 (N_2362,In_880,In_632);
or U2363 (N_2363,In_1188,In_2226);
nor U2364 (N_2364,In_982,In_2439);
nand U2365 (N_2365,In_1016,In_1267);
and U2366 (N_2366,In_1611,In_1123);
or U2367 (N_2367,In_1953,In_1913);
or U2368 (N_2368,In_274,In_1163);
nor U2369 (N_2369,In_1348,In_1333);
nor U2370 (N_2370,In_642,In_570);
or U2371 (N_2371,In_1012,In_2003);
nand U2372 (N_2372,In_1777,In_1662);
nand U2373 (N_2373,In_941,In_2107);
nor U2374 (N_2374,In_1499,In_1329);
or U2375 (N_2375,In_1017,In_79);
xnor U2376 (N_2376,In_1542,In_910);
nand U2377 (N_2377,In_646,In_1010);
and U2378 (N_2378,In_90,In_1398);
nand U2379 (N_2379,In_1192,In_2038);
xnor U2380 (N_2380,In_678,In_1009);
nand U2381 (N_2381,In_1015,In_133);
nor U2382 (N_2382,In_1140,In_2287);
nand U2383 (N_2383,In_86,In_656);
nor U2384 (N_2384,In_2448,In_1660);
nand U2385 (N_2385,In_2275,In_104);
or U2386 (N_2386,In_1593,In_2008);
or U2387 (N_2387,In_1488,In_30);
and U2388 (N_2388,In_2341,In_1875);
nor U2389 (N_2389,In_833,In_2353);
nor U2390 (N_2390,In_954,In_1736);
nor U2391 (N_2391,In_1489,In_1305);
nand U2392 (N_2392,In_217,In_93);
nor U2393 (N_2393,In_295,In_537);
or U2394 (N_2394,In_2162,In_2392);
nor U2395 (N_2395,In_567,In_538);
and U2396 (N_2396,In_581,In_511);
xor U2397 (N_2397,In_282,In_1610);
nor U2398 (N_2398,In_1987,In_1300);
and U2399 (N_2399,In_1297,In_639);
or U2400 (N_2400,In_67,In_2199);
or U2401 (N_2401,In_1749,In_1378);
nor U2402 (N_2402,In_482,In_1562);
and U2403 (N_2403,In_1706,In_748);
nand U2404 (N_2404,In_461,In_253);
nand U2405 (N_2405,In_149,In_1407);
nor U2406 (N_2406,In_819,In_1310);
xor U2407 (N_2407,In_2375,In_584);
nor U2408 (N_2408,In_2451,In_1856);
xor U2409 (N_2409,In_2171,In_41);
xnor U2410 (N_2410,In_1174,In_171);
or U2411 (N_2411,In_1650,In_679);
nand U2412 (N_2412,In_120,In_1497);
and U2413 (N_2413,In_77,In_238);
xor U2414 (N_2414,In_1170,In_2369);
xor U2415 (N_2415,In_131,In_137);
xor U2416 (N_2416,In_990,In_341);
nand U2417 (N_2417,In_554,In_526);
xnor U2418 (N_2418,In_71,In_29);
nand U2419 (N_2419,In_390,In_1115);
xnor U2420 (N_2420,In_1942,In_489);
nand U2421 (N_2421,In_70,In_1626);
or U2422 (N_2422,In_1994,In_1193);
xor U2423 (N_2423,In_1353,In_1603);
or U2424 (N_2424,In_980,In_1468);
and U2425 (N_2425,In_1503,In_483);
and U2426 (N_2426,In_2295,In_1381);
xor U2427 (N_2427,In_576,In_951);
and U2428 (N_2428,In_1101,In_630);
xnor U2429 (N_2429,In_1290,In_885);
or U2430 (N_2430,In_362,In_1380);
and U2431 (N_2431,In_844,In_813);
or U2432 (N_2432,In_525,In_2471);
xnor U2433 (N_2433,In_1174,In_491);
and U2434 (N_2434,In_1259,In_977);
nand U2435 (N_2435,In_1269,In_524);
nand U2436 (N_2436,In_2483,In_350);
or U2437 (N_2437,In_256,In_2076);
and U2438 (N_2438,In_685,In_718);
xor U2439 (N_2439,In_2072,In_2204);
nand U2440 (N_2440,In_1663,In_2429);
xor U2441 (N_2441,In_1532,In_1392);
or U2442 (N_2442,In_423,In_2173);
nor U2443 (N_2443,In_2439,In_680);
and U2444 (N_2444,In_863,In_2035);
and U2445 (N_2445,In_1313,In_1220);
and U2446 (N_2446,In_2304,In_686);
or U2447 (N_2447,In_161,In_1531);
nor U2448 (N_2448,In_1764,In_518);
nor U2449 (N_2449,In_697,In_2235);
or U2450 (N_2450,In_1722,In_867);
or U2451 (N_2451,In_1979,In_316);
nor U2452 (N_2452,In_511,In_933);
xor U2453 (N_2453,In_39,In_308);
nor U2454 (N_2454,In_487,In_1527);
nor U2455 (N_2455,In_671,In_773);
and U2456 (N_2456,In_1555,In_691);
nor U2457 (N_2457,In_2345,In_887);
xnor U2458 (N_2458,In_2281,In_1812);
xnor U2459 (N_2459,In_2416,In_1423);
nor U2460 (N_2460,In_2016,In_1865);
nand U2461 (N_2461,In_81,In_1480);
nand U2462 (N_2462,In_276,In_1089);
nor U2463 (N_2463,In_2207,In_799);
and U2464 (N_2464,In_991,In_1256);
or U2465 (N_2465,In_824,In_979);
or U2466 (N_2466,In_2497,In_1287);
xnor U2467 (N_2467,In_2164,In_1464);
or U2468 (N_2468,In_1089,In_1316);
or U2469 (N_2469,In_881,In_185);
nand U2470 (N_2470,In_280,In_2396);
and U2471 (N_2471,In_761,In_343);
nand U2472 (N_2472,In_2356,In_290);
xor U2473 (N_2473,In_1814,In_634);
and U2474 (N_2474,In_82,In_2350);
nor U2475 (N_2475,In_2104,In_865);
xor U2476 (N_2476,In_2471,In_543);
nand U2477 (N_2477,In_1186,In_1740);
nor U2478 (N_2478,In_252,In_458);
and U2479 (N_2479,In_596,In_281);
nand U2480 (N_2480,In_1796,In_1496);
nand U2481 (N_2481,In_26,In_2120);
nor U2482 (N_2482,In_70,In_722);
and U2483 (N_2483,In_728,In_1166);
and U2484 (N_2484,In_1958,In_592);
or U2485 (N_2485,In_19,In_2360);
nor U2486 (N_2486,In_88,In_80);
nand U2487 (N_2487,In_709,In_1944);
or U2488 (N_2488,In_1190,In_2488);
nor U2489 (N_2489,In_40,In_1469);
nor U2490 (N_2490,In_426,In_1191);
and U2491 (N_2491,In_565,In_94);
xnor U2492 (N_2492,In_195,In_173);
xnor U2493 (N_2493,In_1280,In_1899);
and U2494 (N_2494,In_2316,In_2260);
or U2495 (N_2495,In_1869,In_1819);
and U2496 (N_2496,In_86,In_2343);
and U2497 (N_2497,In_959,In_1863);
xnor U2498 (N_2498,In_1315,In_1667);
and U2499 (N_2499,In_58,In_1152);
nand U2500 (N_2500,N_1152,N_643);
xnor U2501 (N_2501,N_557,N_943);
xor U2502 (N_2502,N_1901,N_2426);
or U2503 (N_2503,N_444,N_1523);
and U2504 (N_2504,N_1237,N_145);
xor U2505 (N_2505,N_1082,N_604);
or U2506 (N_2506,N_2470,N_1483);
or U2507 (N_2507,N_1013,N_302);
and U2508 (N_2508,N_2499,N_914);
and U2509 (N_2509,N_2276,N_285);
nor U2510 (N_2510,N_1987,N_365);
nand U2511 (N_2511,N_1073,N_1413);
nor U2512 (N_2512,N_1709,N_2031);
xnor U2513 (N_2513,N_1321,N_63);
and U2514 (N_2514,N_693,N_793);
nand U2515 (N_2515,N_1398,N_1912);
nand U2516 (N_2516,N_927,N_2270);
or U2517 (N_2517,N_2479,N_1031);
xnor U2518 (N_2518,N_1316,N_1384);
xor U2519 (N_2519,N_695,N_610);
and U2520 (N_2520,N_1388,N_300);
and U2521 (N_2521,N_1324,N_1971);
and U2522 (N_2522,N_458,N_235);
and U2523 (N_2523,N_1042,N_2446);
xor U2524 (N_2524,N_192,N_470);
and U2525 (N_2525,N_1501,N_1207);
or U2526 (N_2526,N_1184,N_280);
xor U2527 (N_2527,N_2045,N_709);
and U2528 (N_2528,N_1105,N_1012);
nand U2529 (N_2529,N_577,N_369);
nand U2530 (N_2530,N_2219,N_1559);
and U2531 (N_2531,N_407,N_2221);
or U2532 (N_2532,N_1880,N_772);
xor U2533 (N_2533,N_1286,N_176);
xor U2534 (N_2534,N_1740,N_2016);
nor U2535 (N_2535,N_1532,N_892);
xor U2536 (N_2536,N_1599,N_1077);
or U2537 (N_2537,N_1728,N_1203);
xnor U2538 (N_2538,N_2356,N_1010);
or U2539 (N_2539,N_651,N_1179);
xor U2540 (N_2540,N_2493,N_583);
or U2541 (N_2541,N_483,N_74);
nor U2542 (N_2542,N_1186,N_1940);
nand U2543 (N_2543,N_1490,N_1036);
xnor U2544 (N_2544,N_1339,N_1638);
xnor U2545 (N_2545,N_1691,N_479);
nor U2546 (N_2546,N_716,N_159);
xnor U2547 (N_2547,N_1109,N_212);
nand U2548 (N_2548,N_1270,N_449);
nor U2549 (N_2549,N_489,N_231);
nand U2550 (N_2550,N_2013,N_2110);
nor U2551 (N_2551,N_826,N_1580);
or U2552 (N_2552,N_1498,N_1762);
and U2553 (N_2553,N_2268,N_2393);
or U2554 (N_2554,N_298,N_805);
xor U2555 (N_2555,N_1431,N_1208);
and U2556 (N_2556,N_1141,N_2108);
nor U2557 (N_2557,N_572,N_1120);
nand U2558 (N_2558,N_2142,N_971);
nand U2559 (N_2559,N_1056,N_388);
nand U2560 (N_2560,N_509,N_1524);
nor U2561 (N_2561,N_527,N_1887);
nand U2562 (N_2562,N_59,N_1255);
and U2563 (N_2563,N_893,N_2107);
nand U2564 (N_2564,N_1342,N_201);
and U2565 (N_2565,N_1725,N_2069);
and U2566 (N_2566,N_1656,N_1061);
nor U2567 (N_2567,N_1153,N_99);
and U2568 (N_2568,N_871,N_2321);
and U2569 (N_2569,N_579,N_901);
nand U2570 (N_2570,N_129,N_2434);
xor U2571 (N_2571,N_1845,N_800);
and U2572 (N_2572,N_206,N_1275);
nand U2573 (N_2573,N_1832,N_1333);
xor U2574 (N_2574,N_658,N_4);
xnor U2575 (N_2575,N_202,N_1983);
or U2576 (N_2576,N_416,N_2329);
or U2577 (N_2577,N_1145,N_1889);
nand U2578 (N_2578,N_561,N_1586);
nor U2579 (N_2579,N_267,N_2036);
and U2580 (N_2580,N_511,N_1747);
xnor U2581 (N_2581,N_1755,N_1235);
or U2582 (N_2582,N_1942,N_714);
and U2583 (N_2583,N_1347,N_382);
or U2584 (N_2584,N_2012,N_398);
and U2585 (N_2585,N_44,N_1516);
and U2586 (N_2586,N_2291,N_406);
xnor U2587 (N_2587,N_1076,N_2309);
and U2588 (N_2588,N_1817,N_379);
xnor U2589 (N_2589,N_1276,N_2299);
nor U2590 (N_2590,N_1200,N_2156);
nand U2591 (N_2591,N_466,N_1063);
and U2592 (N_2592,N_1415,N_214);
nor U2593 (N_2593,N_763,N_1598);
xor U2594 (N_2594,N_1915,N_908);
nand U2595 (N_2595,N_1329,N_1807);
nor U2596 (N_2596,N_316,N_440);
nand U2597 (N_2597,N_1773,N_834);
xnor U2598 (N_2598,N_543,N_1188);
nor U2599 (N_2599,N_784,N_592);
nand U2600 (N_2600,N_143,N_215);
nor U2601 (N_2601,N_1542,N_2055);
xnor U2602 (N_2602,N_838,N_1245);
nor U2603 (N_2603,N_2189,N_2227);
and U2604 (N_2604,N_2430,N_1039);
and U2605 (N_2605,N_749,N_701);
and U2606 (N_2606,N_1164,N_183);
or U2607 (N_2607,N_1630,N_498);
or U2608 (N_2608,N_1812,N_865);
nand U2609 (N_2609,N_1615,N_736);
and U2610 (N_2610,N_1739,N_1119);
nor U2611 (N_2611,N_802,N_1970);
xor U2612 (N_2612,N_1367,N_2303);
or U2613 (N_2613,N_545,N_127);
xnor U2614 (N_2614,N_1225,N_2275);
xnor U2615 (N_2615,N_2497,N_80);
or U2616 (N_2616,N_153,N_955);
or U2617 (N_2617,N_353,N_912);
and U2618 (N_2618,N_2226,N_2178);
or U2619 (N_2619,N_1953,N_2200);
or U2620 (N_2620,N_1272,N_1440);
nand U2621 (N_2621,N_2491,N_1204);
xnor U2622 (N_2622,N_1634,N_1167);
and U2623 (N_2623,N_1209,N_2067);
and U2624 (N_2624,N_1143,N_173);
nor U2625 (N_2625,N_1512,N_376);
and U2626 (N_2626,N_1287,N_1304);
nor U2627 (N_2627,N_1657,N_2486);
nor U2628 (N_2628,N_372,N_1219);
xor U2629 (N_2629,N_1420,N_491);
nor U2630 (N_2630,N_890,N_524);
and U2631 (N_2631,N_616,N_2205);
nand U2632 (N_2632,N_1863,N_1642);
nor U2633 (N_2633,N_593,N_1414);
and U2634 (N_2634,N_197,N_2377);
and U2635 (N_2635,N_712,N_20);
and U2636 (N_2636,N_619,N_2338);
nor U2637 (N_2637,N_1531,N_245);
xnor U2638 (N_2638,N_1262,N_875);
or U2639 (N_2639,N_1961,N_98);
xnor U2640 (N_2640,N_84,N_144);
or U2641 (N_2641,N_1266,N_375);
nand U2642 (N_2642,N_69,N_1635);
nor U2643 (N_2643,N_645,N_1867);
xnor U2644 (N_2644,N_2024,N_2111);
or U2645 (N_2645,N_623,N_2139);
or U2646 (N_2646,N_1273,N_1350);
nand U2647 (N_2647,N_1995,N_2168);
nor U2648 (N_2648,N_420,N_1711);
xor U2649 (N_2649,N_433,N_1375);
or U2650 (N_2650,N_1001,N_526);
xor U2651 (N_2651,N_1791,N_2021);
nor U2652 (N_2652,N_226,N_66);
xnor U2653 (N_2653,N_964,N_2266);
nand U2654 (N_2654,N_1162,N_669);
xnor U2655 (N_2655,N_175,N_1707);
nand U2656 (N_2656,N_2467,N_442);
or U2657 (N_2657,N_1803,N_568);
or U2658 (N_2658,N_881,N_2346);
xor U2659 (N_2659,N_2458,N_502);
or U2660 (N_2660,N_752,N_1299);
xor U2661 (N_2661,N_1944,N_2402);
nand U2662 (N_2662,N_2089,N_2084);
xor U2663 (N_2663,N_1301,N_1972);
and U2664 (N_2664,N_2176,N_1538);
xnor U2665 (N_2665,N_1232,N_2043);
xor U2666 (N_2666,N_1969,N_2245);
or U2667 (N_2667,N_1328,N_1144);
or U2668 (N_2668,N_1959,N_1752);
nor U2669 (N_2669,N_724,N_625);
nor U2670 (N_2670,N_1006,N_29);
or U2671 (N_2671,N_295,N_1268);
or U2672 (N_2672,N_163,N_778);
nand U2673 (N_2673,N_2201,N_90);
nor U2674 (N_2674,N_1871,N_1462);
xnor U2675 (N_2675,N_270,N_564);
or U2676 (N_2676,N_1651,N_2415);
and U2677 (N_2677,N_1704,N_965);
nor U2678 (N_2678,N_149,N_2392);
nor U2679 (N_2679,N_2004,N_166);
xnor U2680 (N_2680,N_473,N_942);
or U2681 (N_2681,N_1756,N_2416);
and U2682 (N_2682,N_2397,N_2048);
xor U2683 (N_2683,N_1341,N_620);
xor U2684 (N_2684,N_2241,N_138);
nor U2685 (N_2685,N_1916,N_797);
or U2686 (N_2686,N_2026,N_2459);
nor U2687 (N_2687,N_1500,N_726);
or U2688 (N_2688,N_1424,N_1850);
xor U2689 (N_2689,N_182,N_1543);
nor U2690 (N_2690,N_1362,N_899);
or U2691 (N_2691,N_707,N_1908);
or U2692 (N_2692,N_2421,N_1662);
nor U2693 (N_2693,N_142,N_2059);
nor U2694 (N_2694,N_409,N_1734);
nor U2695 (N_2695,N_1379,N_1406);
or U2696 (N_2696,N_451,N_56);
xnor U2697 (N_2697,N_2032,N_886);
or U2698 (N_2698,N_1477,N_827);
and U2699 (N_2699,N_294,N_1693);
and U2700 (N_2700,N_1975,N_1596);
nand U2701 (N_2701,N_6,N_1508);
and U2702 (N_2702,N_1359,N_1592);
xor U2703 (N_2703,N_638,N_1802);
and U2704 (N_2704,N_363,N_1996);
xnor U2705 (N_2705,N_244,N_2382);
nand U2706 (N_2706,N_552,N_600);
nand U2707 (N_2707,N_1781,N_2222);
or U2708 (N_2708,N_2097,N_759);
or U2709 (N_2709,N_576,N_2487);
xnor U2710 (N_2710,N_1800,N_1148);
xnor U2711 (N_2711,N_1027,N_1553);
and U2712 (N_2712,N_612,N_1757);
xnor U2713 (N_2713,N_405,N_1421);
and U2714 (N_2714,N_2071,N_782);
nand U2715 (N_2715,N_377,N_1400);
and U2716 (N_2716,N_342,N_373);
xor U2717 (N_2717,N_246,N_515);
nand U2718 (N_2718,N_1327,N_1569);
and U2719 (N_2719,N_229,N_428);
nand U2720 (N_2720,N_2234,N_1236);
nand U2721 (N_2721,N_1552,N_2453);
nor U2722 (N_2722,N_1821,N_1385);
or U2723 (N_2723,N_1718,N_2160);
nand U2724 (N_2724,N_2370,N_949);
or U2725 (N_2725,N_1899,N_1730);
nor U2726 (N_2726,N_2436,N_476);
nor U2727 (N_2727,N_824,N_789);
nor U2728 (N_2728,N_1218,N_1713);
nor U2729 (N_2729,N_856,N_1924);
xor U2730 (N_2730,N_977,N_49);
or U2731 (N_2731,N_2450,N_866);
xnor U2732 (N_2732,N_1973,N_1425);
nor U2733 (N_2733,N_550,N_2283);
and U2734 (N_2734,N_1074,N_1550);
nand U2735 (N_2735,N_715,N_191);
nor U2736 (N_2736,N_1790,N_2420);
nand U2737 (N_2737,N_554,N_2064);
or U2738 (N_2738,N_837,N_457);
or U2739 (N_2739,N_1891,N_396);
nand U2740 (N_2740,N_1558,N_1842);
xnor U2741 (N_2741,N_1976,N_1412);
nor U2742 (N_2742,N_321,N_2288);
xor U2743 (N_2743,N_1044,N_2088);
or U2744 (N_2744,N_1234,N_412);
xnor U2745 (N_2745,N_351,N_1585);
or U2746 (N_2746,N_2468,N_1607);
and U2747 (N_2747,N_492,N_1066);
and U2748 (N_2748,N_340,N_1652);
or U2749 (N_2749,N_1374,N_931);
nor U2750 (N_2750,N_1295,N_2293);
and U2751 (N_2751,N_2239,N_87);
nand U2752 (N_2752,N_1606,N_2195);
nand U2753 (N_2753,N_381,N_2127);
xor U2754 (N_2754,N_1214,N_0);
nand U2755 (N_2755,N_953,N_1720);
nor U2756 (N_2756,N_522,N_2376);
or U2757 (N_2757,N_1934,N_1526);
nor U2758 (N_2758,N_2040,N_2058);
xnor U2759 (N_2759,N_888,N_265);
xnor U2760 (N_2760,N_1841,N_2247);
nor U2761 (N_2761,N_2118,N_1834);
nor U2762 (N_2762,N_77,N_534);
nand U2763 (N_2763,N_767,N_934);
nand U2764 (N_2764,N_2286,N_336);
nand U2765 (N_2765,N_1833,N_1838);
or U2766 (N_2766,N_1396,N_1920);
or U2767 (N_2767,N_1496,N_1018);
or U2768 (N_2768,N_739,N_504);
nand U2769 (N_2769,N_989,N_779);
nor U2770 (N_2770,N_217,N_464);
or U2771 (N_2771,N_380,N_1170);
nor U2772 (N_2772,N_2072,N_1175);
nor U2773 (N_2773,N_1460,N_1765);
and U2774 (N_2774,N_1069,N_1622);
and U2775 (N_2775,N_2070,N_401);
and U2776 (N_2776,N_627,N_1556);
and U2777 (N_2777,N_11,N_1226);
xor U2778 (N_2778,N_2049,N_291);
or U2779 (N_2779,N_1741,N_1933);
nand U2780 (N_2780,N_1659,N_1360);
and U2781 (N_2781,N_1482,N_536);
and U2782 (N_2782,N_975,N_2061);
nor U2783 (N_2783,N_279,N_1767);
nand U2784 (N_2784,N_776,N_94);
xnor U2785 (N_2785,N_1977,N_1932);
or U2786 (N_2786,N_939,N_952);
xor U2787 (N_2787,N_2271,N_454);
nand U2788 (N_2788,N_417,N_1719);
xor U2789 (N_2789,N_1768,N_874);
nand U2790 (N_2790,N_1928,N_1795);
and U2791 (N_2791,N_1305,N_1563);
and U2792 (N_2792,N_25,N_1411);
or U2793 (N_2793,N_2334,N_1437);
or U2794 (N_2794,N_105,N_835);
and U2795 (N_2795,N_165,N_1665);
xnor U2796 (N_2796,N_879,N_944);
nor U2797 (N_2797,N_2335,N_1052);
nor U2798 (N_2798,N_867,N_791);
or U2799 (N_2799,N_2137,N_1468);
or U2800 (N_2800,N_1690,N_303);
or U2801 (N_2801,N_747,N_366);
or U2802 (N_2802,N_637,N_281);
nor U2803 (N_2803,N_1610,N_653);
and U2804 (N_2804,N_521,N_1947);
xnor U2805 (N_2805,N_113,N_589);
xnor U2806 (N_2806,N_1211,N_1518);
or U2807 (N_2807,N_1670,N_51);
xnor U2808 (N_2808,N_1878,N_474);
or U2809 (N_2809,N_1830,N_690);
nor U2810 (N_2810,N_859,N_773);
xnor U2811 (N_2811,N_1094,N_1522);
and U2812 (N_2812,N_2123,N_1548);
nand U2813 (N_2813,N_1993,N_553);
nor U2814 (N_2814,N_8,N_1794);
and U2815 (N_2815,N_755,N_555);
nor U2816 (N_2816,N_43,N_1216);
or U2817 (N_2817,N_574,N_1856);
and U2818 (N_2818,N_2203,N_2355);
and U2819 (N_2819,N_2010,N_1163);
xnor U2820 (N_2820,N_2431,N_787);
nor U2821 (N_2821,N_2481,N_825);
xnor U2822 (N_2822,N_50,N_2399);
nand U2823 (N_2823,N_146,N_426);
or U2824 (N_2824,N_2180,N_2437);
nor U2825 (N_2825,N_1603,N_1687);
nor U2826 (N_2826,N_1250,N_210);
and U2827 (N_2827,N_1637,N_851);
nor U2828 (N_2828,N_21,N_1363);
xor U2829 (N_2829,N_1435,N_1353);
xnor U2830 (N_2830,N_2462,N_180);
and U2831 (N_2831,N_887,N_904);
nor U2832 (N_2832,N_410,N_558);
xnor U2833 (N_2833,N_2375,N_82);
nand U2834 (N_2834,N_2051,N_1849);
or U2835 (N_2835,N_1815,N_199);
nand U2836 (N_2836,N_1241,N_1729);
or U2837 (N_2837,N_1102,N_394);
nand U2838 (N_2838,N_1862,N_41);
nor U2839 (N_2839,N_1682,N_1963);
and U2840 (N_2840,N_1988,N_560);
nand U2841 (N_2841,N_2102,N_2406);
and U2842 (N_2842,N_1159,N_1269);
and U2843 (N_2843,N_2361,N_2225);
nand U2844 (N_2844,N_2007,N_2378);
nor U2845 (N_2845,N_2100,N_1540);
nand U2846 (N_2846,N_648,N_367);
or U2847 (N_2847,N_775,N_1007);
and U2848 (N_2848,N_1660,N_1681);
nand U2849 (N_2849,N_1195,N_1311);
or U2850 (N_2850,N_869,N_967);
and U2851 (N_2851,N_1716,N_1138);
xnor U2852 (N_2852,N_313,N_1857);
nor U2853 (N_2853,N_537,N_882);
xnor U2854 (N_2854,N_950,N_806);
or U2855 (N_2855,N_1161,N_2207);
nor U2856 (N_2856,N_518,N_1140);
and U2857 (N_2857,N_501,N_2383);
xnor U2858 (N_2858,N_453,N_2065);
xor U2859 (N_2859,N_2220,N_626);
or U2860 (N_2860,N_757,N_885);
nand U2861 (N_2861,N_894,N_2365);
or U2862 (N_2862,N_441,N_1894);
nor U2863 (N_2863,N_2318,N_2196);
xor U2864 (N_2864,N_1189,N_1294);
nand U2865 (N_2865,N_1537,N_2223);
or U2866 (N_2866,N_131,N_1277);
nand U2867 (N_2867,N_1777,N_208);
and U2868 (N_2868,N_2216,N_2279);
nor U2869 (N_2869,N_1893,N_1723);
or U2870 (N_2870,N_1905,N_2344);
and U2871 (N_2871,N_2407,N_2348);
or U2872 (N_2872,N_1191,N_30);
nor U2873 (N_2873,N_1703,N_1187);
or U2874 (N_2874,N_1217,N_982);
or U2875 (N_2875,N_1626,N_275);
nand U2876 (N_2876,N_2232,N_902);
or U2877 (N_2877,N_355,N_39);
nand U2878 (N_2878,N_3,N_706);
xor U2879 (N_2879,N_1283,N_1583);
and U2880 (N_2880,N_2103,N_1562);
xor U2881 (N_2881,N_1067,N_532);
and U2882 (N_2882,N_897,N_1405);
or U2883 (N_2883,N_1647,N_76);
or U2884 (N_2884,N_2091,N_1366);
nor U2885 (N_2885,N_2155,N_988);
nand U2886 (N_2886,N_929,N_384);
nor U2887 (N_2887,N_1493,N_970);
nor U2888 (N_2888,N_2498,N_1679);
or U2889 (N_2889,N_718,N_644);
nand U2890 (N_2890,N_186,N_1065);
and U2891 (N_2891,N_843,N_346);
nand U2892 (N_2892,N_2454,N_530);
nand U2893 (N_2893,N_1124,N_469);
xor U2894 (N_2894,N_811,N_1779);
or U2895 (N_2895,N_2244,N_1594);
or U2896 (N_2896,N_1183,N_661);
or U2897 (N_2897,N_1697,N_959);
nand U2898 (N_2898,N_2256,N_263);
xnor U2899 (N_2899,N_1605,N_597);
xnor U2900 (N_2900,N_1395,N_218);
nor U2901 (N_2901,N_672,N_1265);
and U2902 (N_2902,N_2248,N_660);
nor U2903 (N_2903,N_109,N_1865);
or U2904 (N_2904,N_110,N_986);
nand U2905 (N_2905,N_1037,N_1688);
nor U2906 (N_2906,N_287,N_247);
nor U2907 (N_2907,N_2238,N_195);
nand U2908 (N_2908,N_2255,N_1858);
and U2909 (N_2909,N_1248,N_692);
nand U2910 (N_2910,N_753,N_134);
or U2911 (N_2911,N_1097,N_2442);
xor U2912 (N_2912,N_679,N_1735);
nor U2913 (N_2913,N_1019,N_60);
nand U2914 (N_2914,N_1151,N_92);
and U2915 (N_2915,N_1520,N_2077);
xnor U2916 (N_2916,N_2443,N_1368);
xor U2917 (N_2917,N_1877,N_503);
nand U2918 (N_2918,N_1576,N_531);
xor U2919 (N_2919,N_2099,N_663);
nand U2920 (N_2920,N_960,N_352);
nand U2921 (N_2921,N_1409,N_758);
nor U2922 (N_2922,N_1989,N_1882);
and U2923 (N_2923,N_1616,N_1567);
nor U2924 (N_2924,N_68,N_1201);
or U2925 (N_2925,N_1632,N_562);
xor U2926 (N_2926,N_1123,N_203);
or U2927 (N_2927,N_1478,N_228);
xnor U2928 (N_2928,N_1701,N_1261);
nand U2929 (N_2929,N_849,N_1966);
xor U2930 (N_2930,N_2068,N_1048);
or U2931 (N_2931,N_650,N_1499);
nor U2932 (N_2932,N_1075,N_1957);
nor U2933 (N_2933,N_2472,N_1999);
nand U2934 (N_2934,N_1212,N_2224);
nand U2935 (N_2935,N_288,N_1369);
nand U2936 (N_2936,N_386,N_1106);
xnor U2937 (N_2937,N_499,N_1149);
nor U2938 (N_2938,N_1199,N_383);
or U2939 (N_2939,N_614,N_546);
xnor U2940 (N_2940,N_2433,N_1320);
and U2941 (N_2941,N_617,N_2164);
nor U2942 (N_2942,N_820,N_2152);
nor U2943 (N_2943,N_1020,N_222);
xor U2944 (N_2944,N_12,N_2085);
nor U2945 (N_2945,N_488,N_538);
nor U2946 (N_2946,N_204,N_387);
nand U2947 (N_2947,N_1564,N_936);
nor U2948 (N_2948,N_2186,N_1177);
or U2949 (N_2949,N_1215,N_1264);
or U2950 (N_2950,N_602,N_2320);
nor U2951 (N_2951,N_116,N_1387);
nand U2952 (N_2952,N_1323,N_1060);
xor U2953 (N_2953,N_2237,N_320);
nand U2954 (N_2954,N_721,N_731);
nand U2955 (N_2955,N_2405,N_2157);
and U2956 (N_2956,N_1093,N_547);
and U2957 (N_2957,N_2466,N_1588);
nor U2958 (N_2958,N_2285,N_2367);
xnor U2959 (N_2959,N_1608,N_1474);
and U2960 (N_2960,N_72,N_2120);
nand U2961 (N_2961,N_659,N_2126);
xnor U2962 (N_2962,N_400,N_2418);
nor U2963 (N_2963,N_1011,N_1238);
xor U2964 (N_2964,N_1917,N_1091);
nand U2965 (N_2965,N_2253,N_86);
nor U2966 (N_2966,N_1130,N_24);
or U2967 (N_2967,N_722,N_1443);
nor U2968 (N_2968,N_1668,N_705);
xnor U2969 (N_2969,N_850,N_1813);
nor U2970 (N_2970,N_1355,N_1612);
nand U2971 (N_2971,N_896,N_1965);
nor U2972 (N_2972,N_2265,N_1487);
and U2973 (N_2973,N_2212,N_1103);
xnor U2974 (N_2974,N_1945,N_284);
or U2975 (N_2975,N_1373,N_2423);
or U2976 (N_2976,N_1246,N_1620);
or U2977 (N_2977,N_1939,N_1686);
nand U2978 (N_2978,N_831,N_680);
or U2979 (N_2979,N_1986,N_1736);
nand U2980 (N_2980,N_1278,N_31);
nor U2981 (N_2981,N_64,N_2166);
xor U2982 (N_2982,N_1879,N_2116);
xor U2983 (N_2983,N_937,N_306);
nor U2984 (N_2984,N_2341,N_1213);
or U2985 (N_2985,N_1633,N_2083);
xnor U2986 (N_2986,N_704,N_467);
and U2987 (N_2987,N_2428,N_973);
or U2988 (N_2988,N_2047,N_2485);
xnor U2989 (N_2989,N_1169,N_2363);
or U2990 (N_2990,N_1913,N_1764);
and U2991 (N_2991,N_487,N_326);
and U2992 (N_2992,N_2122,N_2417);
or U2993 (N_2993,N_1371,N_1297);
and U2994 (N_2994,N_2243,N_2389);
nand U2995 (N_2995,N_2448,N_2027);
nor U2996 (N_2996,N_1104,N_1337);
and U2997 (N_2997,N_2175,N_2394);
xnor U2998 (N_2998,N_533,N_1445);
xor U2999 (N_2999,N_2317,N_359);
or U3000 (N_3000,N_2327,N_2337);
xor U3001 (N_3001,N_697,N_1875);
xor U3002 (N_3002,N_1835,N_675);
xnor U3003 (N_3003,N_1244,N_1551);
nor U3004 (N_3004,N_1423,N_2259);
xnor U3005 (N_3005,N_2184,N_1991);
nand U3006 (N_3006,N_1904,N_1290);
xnor U3007 (N_3007,N_1197,N_780);
nor U3008 (N_3008,N_630,N_2194);
xor U3009 (N_3009,N_994,N_1621);
or U3010 (N_3010,N_2198,N_666);
nor U3011 (N_3011,N_271,N_932);
xnor U3012 (N_3012,N_2336,N_297);
nand U3013 (N_3013,N_2304,N_2432);
nand U3014 (N_3014,N_1705,N_1582);
nand U3015 (N_3015,N_1092,N_877);
nand U3016 (N_3016,N_19,N_729);
and U3017 (N_3017,N_1041,N_2213);
or U3018 (N_3018,N_423,N_1450);
xor U3019 (N_3019,N_980,N_2424);
or U3020 (N_3020,N_2105,N_1165);
xor U3021 (N_3021,N_1125,N_1925);
and U3022 (N_3022,N_817,N_350);
nand U3023 (N_3023,N_331,N_282);
or U3024 (N_3024,N_829,N_1291);
xnor U3025 (N_3025,N_588,N_974);
or U3026 (N_3026,N_1121,N_870);
xor U3027 (N_3027,N_1157,N_155);
or U3028 (N_3028,N_1534,N_1536);
nor U3029 (N_3029,N_1726,N_1658);
xnor U3030 (N_3030,N_2172,N_1113);
xnor U3031 (N_3031,N_801,N_1009);
nand U3032 (N_3032,N_1738,N_1386);
nor U3033 (N_3033,N_1410,N_2360);
xor U3034 (N_3034,N_946,N_765);
nand U3035 (N_3035,N_1804,N_2046);
and U3036 (N_3036,N_777,N_1611);
nor U3037 (N_3037,N_55,N_1579);
xnor U3038 (N_3038,N_2395,N_1661);
nand U3039 (N_3039,N_1628,N_239);
xnor U3040 (N_3040,N_1786,N_324);
xnor U3041 (N_3041,N_374,N_2119);
xor U3042 (N_3042,N_2075,N_430);
nor U3043 (N_3043,N_1340,N_2052);
nor U3044 (N_3044,N_1602,N_1968);
nand U3045 (N_3045,N_862,N_2000);
nor U3046 (N_3046,N_7,N_1809);
nand U3047 (N_3047,N_1310,N_2115);
and U3048 (N_3048,N_413,N_1528);
and U3049 (N_3049,N_719,N_238);
nand U3050 (N_3050,N_1014,N_830);
or U3051 (N_3051,N_1717,N_189);
nor U3052 (N_3052,N_513,N_566);
xor U3053 (N_3053,N_1086,N_478);
and U3054 (N_3054,N_951,N_1958);
nand U3055 (N_3055,N_1466,N_304);
and U3056 (N_3056,N_2006,N_456);
nand U3057 (N_3057,N_1846,N_1702);
nand U3058 (N_3058,N_1950,N_1038);
xor U3059 (N_3059,N_1308,N_1561);
and U3060 (N_3060,N_1792,N_2372);
xnor U3061 (N_3061,N_921,N_2235);
nand U3062 (N_3062,N_1072,N_961);
xnor U3063 (N_3063,N_2273,N_819);
xnor U3064 (N_3064,N_1743,N_1771);
or U3065 (N_3065,N_608,N_1003);
xor U3066 (N_3066,N_1122,N_1452);
nor U3067 (N_3067,N_259,N_2060);
or U3068 (N_3068,N_2173,N_1869);
or U3069 (N_3069,N_1114,N_1806);
and U3070 (N_3070,N_1180,N_140);
xor U3071 (N_3071,N_1128,N_2456);
and U3072 (N_3072,N_744,N_508);
and U3073 (N_3073,N_906,N_1541);
and U3074 (N_3074,N_1503,N_193);
nor U3075 (N_3075,N_286,N_236);
and U3076 (N_3076,N_1302,N_2440);
or U3077 (N_3077,N_65,N_1769);
and U3078 (N_3078,N_1910,N_992);
nor U3079 (N_3079,N_328,N_2483);
and U3080 (N_3080,N_575,N_237);
xnor U3081 (N_3081,N_2215,N_2187);
nor U3082 (N_3082,N_1100,N_22);
or U3083 (N_3083,N_1172,N_764);
and U3084 (N_3084,N_1874,N_633);
and U3085 (N_3085,N_1903,N_1332);
nand U3086 (N_3086,N_1814,N_861);
and U3087 (N_3087,N_256,N_2307);
or U3088 (N_3088,N_293,N_2345);
or U3089 (N_3089,N_1252,N_1573);
xnor U3090 (N_3090,N_1227,N_462);
nand U3091 (N_3091,N_673,N_1298);
nand U3092 (N_3092,N_120,N_1344);
nor U3093 (N_3093,N_1312,N_1046);
xnor U3094 (N_3094,N_2358,N_1058);
or U3095 (N_3095,N_1441,N_46);
and U3096 (N_3096,N_2351,N_1253);
or U3097 (N_3097,N_48,N_1673);
nor U3098 (N_3098,N_2204,N_305);
or U3099 (N_3099,N_839,N_924);
and U3100 (N_3100,N_2177,N_1021);
nor U3101 (N_3101,N_622,N_945);
and U3102 (N_3102,N_1967,N_1853);
or U3103 (N_3103,N_1233,N_2141);
nand U3104 (N_3104,N_853,N_807);
nor U3105 (N_3105,N_1285,N_925);
or U3106 (N_3106,N_1352,N_2310);
xor U3107 (N_3107,N_1818,N_685);
or U3108 (N_3108,N_2257,N_2278);
and U3109 (N_3109,N_1372,N_2267);
or U3110 (N_3110,N_1851,N_1282);
xor U3111 (N_3111,N_615,N_1313);
nand U3112 (N_3112,N_1597,N_1354);
nor U3113 (N_3113,N_118,N_985);
nor U3114 (N_3114,N_551,N_710);
or U3115 (N_3115,N_1111,N_1389);
nor U3116 (N_3116,N_356,N_1254);
nand U3117 (N_3117,N_2350,N_2410);
xnor U3118 (N_3118,N_70,N_649);
nand U3119 (N_3119,N_2014,N_1419);
and U3120 (N_3120,N_358,N_187);
nand U3121 (N_3121,N_1451,N_419);
xnor U3122 (N_3122,N_1979,N_813);
nand U3123 (N_3123,N_269,N_762);
nand U3124 (N_3124,N_1890,N_786);
xnor U3125 (N_3125,N_635,N_1584);
nor U3126 (N_3126,N_1418,N_2117);
or U3127 (N_3127,N_1787,N_1962);
or U3128 (N_3128,N_1870,N_913);
nor U3129 (N_3129,N_2182,N_2388);
or U3130 (N_3130,N_1085,N_681);
nor U3131 (N_3131,N_329,N_112);
nor U3132 (N_3132,N_520,N_1852);
nand U3133 (N_3133,N_1545,N_900);
or U3134 (N_3134,N_2413,N_408);
and U3135 (N_3135,N_580,N_100);
or U3136 (N_3136,N_683,N_1619);
or U3137 (N_3137,N_2368,N_917);
nand U3138 (N_3138,N_594,N_71);
or U3139 (N_3139,N_2435,N_242);
or U3140 (N_3140,N_1568,N_1514);
or U3141 (N_3141,N_1491,N_1724);
or U3142 (N_3142,N_2400,N_477);
and U3143 (N_3143,N_357,N_1810);
nand U3144 (N_3144,N_1326,N_563);
nor U3145 (N_3145,N_2231,N_1055);
nor U3146 (N_3146,N_266,N_923);
nor U3147 (N_3147,N_1049,N_1330);
or U3148 (N_3148,N_976,N_1098);
xnor U3149 (N_3149,N_2277,N_338);
nor U3150 (N_3150,N_1855,N_2332);
or U3151 (N_3151,N_947,N_1376);
nand U3152 (N_3152,N_262,N_345);
xor U3153 (N_3153,N_1549,N_2330);
xnor U3154 (N_3154,N_1645,N_840);
nand U3155 (N_3155,N_1456,N_2480);
or U3156 (N_3156,N_1289,N_1577);
nand U3157 (N_3157,N_1527,N_1392);
nor U3158 (N_3158,N_1416,N_940);
xnor U3159 (N_3159,N_2246,N_1954);
nor U3160 (N_3160,N_347,N_257);
nand U3161 (N_3161,N_1182,N_1799);
and U3162 (N_3162,N_1919,N_2030);
xnor U3163 (N_3163,N_111,N_1495);
nand U3164 (N_3164,N_2087,N_2092);
and U3165 (N_3165,N_1335,N_1883);
or U3166 (N_3166,N_2153,N_224);
or U3167 (N_3167,N_584,N_95);
or U3168 (N_3168,N_2101,N_1943);
nand U3169 (N_3169,N_1417,N_1343);
and U3170 (N_3170,N_1745,N_2066);
nor U3171 (N_3171,N_993,N_2419);
xor U3172 (N_3172,N_268,N_2038);
or U3173 (N_3173,N_1775,N_1178);
or U3174 (N_3174,N_1677,N_114);
or U3175 (N_3175,N_2008,N_1578);
xnor U3176 (N_3176,N_139,N_2076);
nand U3177 (N_3177,N_1751,N_828);
or U3178 (N_3178,N_1271,N_2146);
or U3179 (N_3179,N_2333,N_2094);
and U3180 (N_3180,N_1990,N_1763);
or U3181 (N_3181,N_2425,N_221);
nand U3182 (N_3182,N_2347,N_743);
nand U3183 (N_3183,N_1900,N_162);
or U3184 (N_3184,N_471,N_700);
or U3185 (N_3185,N_2414,N_2492);
and U3186 (N_3186,N_1955,N_1843);
xnor U3187 (N_3187,N_1080,N_2217);
nand U3188 (N_3188,N_548,N_2449);
nand U3189 (N_3189,N_641,N_2297);
nand U3190 (N_3190,N_655,N_1998);
nor U3191 (N_3191,N_948,N_1064);
nand U3192 (N_3192,N_1951,N_205);
nand U3193 (N_3193,N_1035,N_1222);
or U3194 (N_3194,N_1949,N_1488);
or U3195 (N_3195,N_1492,N_264);
nand U3196 (N_3196,N_686,N_200);
nor U3197 (N_3197,N_101,N_905);
nand U3198 (N_3198,N_1228,N_1486);
nor U3199 (N_3199,N_1546,N_103);
xnor U3200 (N_3200,N_1479,N_2322);
or U3201 (N_3201,N_2260,N_40);
nand U3202 (N_3202,N_301,N_1481);
and U3203 (N_3203,N_2474,N_2009);
nand U3204 (N_3204,N_855,N_337);
and U3205 (N_3205,N_1365,N_1439);
or U3206 (N_3206,N_1083,N_1808);
or U3207 (N_3207,N_385,N_1560);
nor U3208 (N_3208,N_915,N_1150);
and U3209 (N_3209,N_1455,N_2130);
nor U3210 (N_3210,N_1547,N_2121);
or U3211 (N_3211,N_2140,N_1744);
and U3212 (N_3212,N_437,N_997);
nand U3213 (N_3213,N_507,N_452);
and U3214 (N_3214,N_1793,N_211);
xor U3215 (N_3215,N_540,N_1507);
and U3216 (N_3216,N_1139,N_1257);
nand U3217 (N_3217,N_2019,N_586);
or U3218 (N_3218,N_174,N_1047);
nand U3219 (N_3219,N_1936,N_621);
and U3220 (N_3220,N_85,N_1627);
and U3221 (N_3221,N_1731,N_1453);
nand U3222 (N_3222,N_2003,N_96);
or U3223 (N_3223,N_147,N_343);
nand U3224 (N_3224,N_1087,N_2106);
or U3225 (N_3225,N_2455,N_1675);
xor U3226 (N_3226,N_1780,N_930);
xor U3227 (N_3227,N_1154,N_1727);
nor U3228 (N_3228,N_2090,N_984);
nor U3229 (N_3229,N_609,N_2022);
xnor U3230 (N_3230,N_968,N_309);
nor U3231 (N_3231,N_2352,N_770);
nor U3232 (N_3232,N_768,N_1158);
nand U3233 (N_3233,N_10,N_1117);
nor U3234 (N_3234,N_2294,N_1749);
or U3235 (N_3235,N_14,N_1938);
xor U3236 (N_3236,N_1378,N_1571);
nand U3237 (N_3237,N_1022,N_1695);
nor U3238 (N_3238,N_2369,N_2132);
nand U3239 (N_3239,N_783,N_2230);
and U3240 (N_3240,N_2353,N_570);
and U3241 (N_3241,N_170,N_429);
nand U3242 (N_3242,N_1930,N_2001);
nor U3243 (N_3243,N_1708,N_5);
nor U3244 (N_3244,N_2319,N_821);
or U3245 (N_3245,N_334,N_126);
and U3246 (N_3246,N_1517,N_2109);
nand U3247 (N_3247,N_1306,N_1000);
xor U3248 (N_3248,N_1732,N_814);
and U3249 (N_3249,N_2469,N_1084);
nand U3250 (N_3250,N_1485,N_196);
or U3251 (N_3251,N_991,N_2305);
or U3252 (N_3252,N_425,N_1404);
or U3253 (N_3253,N_1300,N_1683);
nor U3254 (N_3254,N_2281,N_788);
nor U3255 (N_3255,N_1314,N_2113);
nand U3256 (N_3256,N_678,N_1666);
nor U3257 (N_3257,N_123,N_422);
xnor U3258 (N_3258,N_2465,N_2039);
xnor U3259 (N_3259,N_1062,N_124);
or U3260 (N_3260,N_2484,N_711);
nor U3261 (N_3261,N_276,N_1267);
or U3262 (N_3262,N_581,N_809);
xnor U3263 (N_3263,N_1346,N_395);
nor U3264 (N_3264,N_1742,N_2098);
and U3265 (N_3265,N_1430,N_1315);
or U3266 (N_3266,N_591,N_1896);
or U3267 (N_3267,N_254,N_1349);
and U3268 (N_3268,N_995,N_1589);
nor U3269 (N_3269,N_1274,N_1442);
xor U3270 (N_3270,N_1676,N_393);
or U3271 (N_3271,N_1750,N_1772);
nand U3272 (N_3272,N_1922,N_1334);
nor U3273 (N_3273,N_1811,N_2249);
xnor U3274 (N_3274,N_158,N_694);
nand U3275 (N_3275,N_1079,N_2062);
nand U3276 (N_3276,N_1131,N_1357);
or U3277 (N_3277,N_89,N_402);
xor U3278 (N_3278,N_1040,N_823);
nor U3279 (N_3279,N_1694,N_1797);
nor U3280 (N_3280,N_1296,N_1698);
xnor U3281 (N_3281,N_2438,N_399);
and U3282 (N_3282,N_468,N_958);
xnor U3283 (N_3283,N_1733,N_794);
xnor U3284 (N_3284,N_1024,N_463);
nand U3285 (N_3285,N_2290,N_1692);
xor U3286 (N_3286,N_1618,N_455);
xnor U3287 (N_3287,N_260,N_790);
nand U3288 (N_3288,N_605,N_1317);
nor U3289 (N_3289,N_919,N_847);
and U3290 (N_3290,N_1715,N_1181);
or U3291 (N_3291,N_1088,N_42);
and U3292 (N_3292,N_482,N_1461);
nand U3293 (N_3293,N_1888,N_607);
nand U3294 (N_3294,N_1399,N_133);
or U3295 (N_3295,N_1515,N_1502);
and U3296 (N_3296,N_2020,N_181);
or U3297 (N_3297,N_2170,N_26);
xnor U3298 (N_3298,N_2029,N_327);
nand U3299 (N_3299,N_987,N_962);
or U3300 (N_3300,N_1721,N_1043);
xnor U3301 (N_3301,N_318,N_278);
xor U3302 (N_3302,N_2096,N_2340);
and U3303 (N_3303,N_361,N_220);
nand U3304 (N_3304,N_446,N_647);
or U3305 (N_3305,N_1489,N_2135);
or U3306 (N_3306,N_798,N_397);
nand U3307 (N_3307,N_415,N_569);
or U3308 (N_3308,N_2463,N_277);
and U3309 (N_3309,N_1230,N_1646);
xor U3310 (N_3310,N_1394,N_194);
and U3311 (N_3311,N_480,N_1674);
nand U3312 (N_3312,N_1240,N_325);
xor U3313 (N_3313,N_45,N_148);
nand U3314 (N_3314,N_1509,N_249);
nor U3315 (N_3315,N_2313,N_1118);
xor U3316 (N_3316,N_815,N_2403);
and U3317 (N_3317,N_2165,N_2229);
xnor U3318 (N_3318,N_447,N_1465);
nand U3319 (N_3319,N_1648,N_702);
and U3320 (N_3320,N_601,N_1631);
nand U3321 (N_3321,N_2411,N_1614);
nand U3322 (N_3322,N_2464,N_863);
and U3323 (N_3323,N_1383,N_1050);
and U3324 (N_3324,N_2017,N_1623);
or U3325 (N_3325,N_876,N_371);
nor U3326 (N_3326,N_852,N_541);
nor U3327 (N_3327,N_1859,N_514);
or U3328 (N_3328,N_639,N_1557);
xnor U3329 (N_3329,N_848,N_2387);
nor U3330 (N_3330,N_93,N_1525);
nand U3331 (N_3331,N_1408,N_634);
and U3332 (N_3332,N_1081,N_1005);
or U3333 (N_3333,N_438,N_2171);
nor U3334 (N_3334,N_2074,N_972);
xnor U3335 (N_3335,N_2079,N_115);
and U3336 (N_3336,N_1090,N_230);
xor U3337 (N_3337,N_13,N_2136);
nor U3338 (N_3338,N_1023,N_1663);
nor U3339 (N_3339,N_1820,N_1566);
nand U3340 (N_3340,N_2343,N_1263);
nand U3341 (N_3341,N_2181,N_519);
or U3342 (N_3342,N_2296,N_1754);
xor U3343 (N_3343,N_674,N_1223);
or U3344 (N_3344,N_667,N_1982);
nor U3345 (N_3345,N_935,N_2011);
nor U3346 (N_3346,N_1788,N_354);
xor U3347 (N_3347,N_32,N_251);
and U3348 (N_3348,N_1844,N_1643);
or U3349 (N_3349,N_969,N_1338);
nor U3350 (N_3350,N_1476,N_500);
and U3351 (N_3351,N_730,N_754);
or U3352 (N_3352,N_1873,N_2287);
xor U3353 (N_3353,N_1370,N_2452);
or U3354 (N_3354,N_571,N_227);
nand U3355 (N_3355,N_723,N_1828);
or U3356 (N_3356,N_1382,N_2295);
or U3357 (N_3357,N_662,N_1504);
xor U3358 (N_3358,N_559,N_857);
nand U3359 (N_3359,N_990,N_978);
or U3360 (N_3360,N_389,N_1448);
or U3361 (N_3361,N_1403,N_999);
nor U3362 (N_3362,N_822,N_1);
or U3363 (N_3363,N_1402,N_2095);
nand U3364 (N_3364,N_549,N_1664);
or U3365 (N_3365,N_1401,N_1776);
nor U3366 (N_3366,N_528,N_1581);
nor U3367 (N_3367,N_232,N_258);
nand U3368 (N_3368,N_2439,N_587);
xor U3369 (N_3369,N_535,N_2114);
xnor U3370 (N_3370,N_2134,N_2412);
nor U3371 (N_3371,N_1710,N_624);
nand U3372 (N_3372,N_78,N_1202);
xnor U3373 (N_3373,N_1176,N_154);
nor U3374 (N_3374,N_878,N_391);
xor U3375 (N_3375,N_1572,N_889);
nand U3376 (N_3376,N_274,N_2209);
xnor U3377 (N_3377,N_2289,N_1819);
nor U3378 (N_3378,N_252,N_1345);
nand U3379 (N_3379,N_708,N_1801);
xor U3380 (N_3380,N_198,N_2401);
nand U3381 (N_3381,N_73,N_785);
and U3382 (N_3382,N_104,N_1529);
nand U3383 (N_3383,N_585,N_864);
and U3384 (N_3384,N_1544,N_567);
nand U3385 (N_3385,N_2080,N_1876);
or U3386 (N_3386,N_404,N_1609);
nand U3387 (N_3387,N_1171,N_414);
nor U3388 (N_3388,N_2023,N_1281);
nor U3389 (N_3389,N_1591,N_2314);
nor U3390 (N_3390,N_2150,N_1847);
nand U3391 (N_3391,N_219,N_872);
and U3392 (N_3392,N_748,N_2477);
xnor U3393 (N_3393,N_1984,N_846);
xor U3394 (N_3394,N_1918,N_2385);
xor U3395 (N_3395,N_737,N_1892);
or U3396 (N_3396,N_1604,N_1436);
xnor U3397 (N_3397,N_1303,N_2489);
nor U3398 (N_3398,N_47,N_665);
and U3399 (N_3399,N_2041,N_1422);
and U3400 (N_3400,N_1758,N_2236);
and U3401 (N_3401,N_1135,N_1654);
xnor U3402 (N_3402,N_688,N_727);
nand U3403 (N_3403,N_954,N_1446);
nand U3404 (N_3404,N_1881,N_424);
or U3405 (N_3405,N_756,N_1669);
or U3406 (N_3406,N_1519,N_1307);
nor U3407 (N_3407,N_1737,N_1595);
or U3408 (N_3408,N_796,N_676);
xor U3409 (N_3409,N_1348,N_1016);
and U3410 (N_3410,N_738,N_734);
nand U3411 (N_3411,N_733,N_1826);
xor U3412 (N_3412,N_1351,N_370);
nor U3413 (N_3413,N_2325,N_2396);
nor U3414 (N_3414,N_640,N_1364);
xnor U3415 (N_3415,N_606,N_2323);
xnor U3416 (N_3416,N_2250,N_130);
or U3417 (N_3417,N_1239,N_2211);
nor U3418 (N_3418,N_2311,N_1484);
nor U3419 (N_3419,N_1356,N_792);
nor U3420 (N_3420,N_629,N_898);
and U3421 (N_3421,N_2471,N_717);
nor U3422 (N_3422,N_2359,N_1997);
nor U3423 (N_3423,N_496,N_79);
and U3424 (N_3424,N_2240,N_1377);
nor U3425 (N_3425,N_603,N_2292);
nor U3426 (N_3426,N_582,N_2282);
nor U3427 (N_3427,N_332,N_36);
nor U3428 (N_3428,N_1173,N_2357);
or U3429 (N_3429,N_2374,N_895);
nand U3430 (N_3430,N_1473,N_167);
nand U3431 (N_3431,N_233,N_1426);
and U3432 (N_3432,N_2381,N_2057);
nand U3433 (N_3433,N_1914,N_510);
and U3434 (N_3434,N_684,N_810);
xor U3435 (N_3435,N_1107,N_2188);
nand U3436 (N_3436,N_1680,N_1051);
nor U3437 (N_3437,N_2445,N_335);
or U3438 (N_3438,N_1133,N_216);
nand U3439 (N_3439,N_497,N_1361);
nand U3440 (N_3440,N_1671,N_289);
nor U3441 (N_3441,N_225,N_255);
nand U3442 (N_3442,N_2183,N_390);
xnor U3443 (N_3443,N_1259,N_1407);
and U3444 (N_3444,N_1288,N_137);
nand U3445 (N_3445,N_2163,N_2159);
nand U3446 (N_3446,N_1147,N_461);
or U3447 (N_3447,N_2478,N_296);
or U3448 (N_3448,N_241,N_836);
nand U3449 (N_3449,N_1570,N_1472);
or U3450 (N_3450,N_618,N_1782);
or U3451 (N_3451,N_539,N_1974);
or U3452 (N_3452,N_1895,N_1906);
nand U3453 (N_3453,N_1816,N_2082);
and U3454 (N_3454,N_689,N_54);
or U3455 (N_3455,N_1672,N_1206);
xor U3456 (N_3456,N_121,N_1057);
xor U3457 (N_3457,N_432,N_745);
nor U3458 (N_3458,N_884,N_1992);
nand U3459 (N_3459,N_1318,N_1590);
xnor U3460 (N_3460,N_135,N_348);
nor U3461 (N_3461,N_2490,N_907);
nor U3462 (N_3462,N_2133,N_322);
or U3463 (N_3463,N_2362,N_2429);
nand U3464 (N_3464,N_1837,N_1649);
or U3465 (N_3465,N_1868,N_2302);
nand U3466 (N_3466,N_315,N_2284);
xor U3467 (N_3467,N_1653,N_460);
nor U3468 (N_3468,N_1054,N_963);
or U3469 (N_3469,N_169,N_1132);
nand U3470 (N_3470,N_1429,N_2138);
nor U3471 (N_3471,N_611,N_1229);
nand U3472 (N_3472,N_2228,N_1438);
xor U3473 (N_3473,N_2005,N_436);
and U3474 (N_3474,N_188,N_2331);
xor U3475 (N_3475,N_37,N_2202);
xor U3476 (N_3476,N_933,N_490);
nor U3477 (N_3477,N_2308,N_1624);
xnor U3478 (N_3478,N_1956,N_1155);
and U3479 (N_3479,N_1381,N_646);
nand U3480 (N_3480,N_803,N_2124);
nor U3481 (N_3481,N_732,N_2391);
or U3482 (N_3482,N_1449,N_17);
nand U3483 (N_3483,N_1126,N_209);
or U3484 (N_3484,N_818,N_1070);
nor U3485 (N_3485,N_1640,N_494);
nor U3486 (N_3486,N_1937,N_1028);
and U3487 (N_3487,N_761,N_250);
nand U3488 (N_3488,N_2349,N_33);
and U3489 (N_3489,N_141,N_1714);
or U3490 (N_3490,N_1336,N_161);
nand U3491 (N_3491,N_2408,N_1644);
xor U3492 (N_3492,N_1108,N_746);
and U3493 (N_3493,N_2272,N_1101);
and U3494 (N_3494,N_107,N_1247);
or U3495 (N_3495,N_1839,N_1761);
or U3496 (N_3496,N_1463,N_108);
or U3497 (N_3497,N_956,N_698);
nor U3498 (N_3498,N_578,N_1174);
nand U3499 (N_3499,N_2054,N_922);
nand U3500 (N_3500,N_2104,N_842);
or U3501 (N_3501,N_2034,N_1078);
and U3502 (N_3502,N_1284,N_495);
or U3503 (N_3503,N_1480,N_2473);
and U3504 (N_3504,N_769,N_1196);
nand U3505 (N_3505,N_506,N_1127);
nand U3506 (N_3506,N_2404,N_1722);
nand U3507 (N_3507,N_1457,N_833);
or U3508 (N_3508,N_1641,N_27);
nor U3509 (N_3509,N_57,N_1866);
nor U3510 (N_3510,N_1475,N_2028);
xnor U3511 (N_3511,N_1243,N_1823);
nor U3512 (N_3512,N_760,N_529);
nor U3513 (N_3513,N_668,N_1136);
nor U3514 (N_3514,N_1510,N_2002);
nand U3515 (N_3515,N_243,N_1521);
xor U3516 (N_3516,N_2364,N_505);
nand U3517 (N_3517,N_1459,N_966);
nand U3518 (N_3518,N_2251,N_435);
nor U3519 (N_3519,N_595,N_1280);
nand U3520 (N_3520,N_1746,N_845);
or U3521 (N_3521,N_362,N_742);
xnor U3522 (N_3522,N_119,N_2191);
nor U3523 (N_3523,N_61,N_1980);
nor U3524 (N_3524,N_1554,N_1096);
xor U3525 (N_3525,N_2315,N_1696);
and U3526 (N_3526,N_1824,N_1712);
or U3527 (N_3527,N_1926,N_450);
or U3528 (N_3528,N_9,N_1864);
nand U3529 (N_3529,N_1242,N_2145);
nor U3530 (N_3530,N_699,N_207);
or U3531 (N_3531,N_481,N_687);
nor U3532 (N_3532,N_728,N_1778);
nand U3533 (N_3533,N_799,N_2301);
and U3534 (N_3534,N_18,N_2125);
xor U3535 (N_3535,N_1059,N_1593);
or U3536 (N_3536,N_1427,N_2326);
xor U3537 (N_3537,N_2316,N_916);
and U3538 (N_3538,N_1655,N_808);
and U3539 (N_3539,N_2,N_523);
xor U3540 (N_3540,N_1089,N_1909);
nor U3541 (N_3541,N_128,N_1840);
and U3542 (N_3542,N_2274,N_1256);
nand U3543 (N_3543,N_938,N_918);
nor U3544 (N_3544,N_125,N_1985);
nand U3545 (N_3545,N_1861,N_1471);
and U3546 (N_3546,N_1390,N_1454);
and U3547 (N_3547,N_1325,N_1497);
or U3548 (N_3548,N_75,N_1116);
or U3549 (N_3549,N_439,N_1045);
xnor U3550 (N_3550,N_2242,N_240);
nor U3551 (N_3551,N_2373,N_771);
nor U3552 (N_3552,N_150,N_160);
or U3553 (N_3553,N_411,N_2143);
nand U3554 (N_3554,N_725,N_1539);
xor U3555 (N_3555,N_1952,N_234);
or U3556 (N_3556,N_766,N_983);
nand U3557 (N_3557,N_431,N_1166);
and U3558 (N_3558,N_330,N_190);
nor U3559 (N_3559,N_136,N_418);
or U3560 (N_3560,N_2148,N_590);
nor U3561 (N_3561,N_542,N_2206);
nor U3562 (N_3562,N_2161,N_1805);
nor U3563 (N_3563,N_2447,N_2044);
xnor U3564 (N_3564,N_2018,N_2073);
and U3565 (N_3565,N_475,N_1785);
nor U3566 (N_3566,N_2258,N_1190);
or U3567 (N_3567,N_1533,N_1115);
and U3568 (N_3568,N_1494,N_2482);
or U3569 (N_3569,N_860,N_2174);
nand U3570 (N_3570,N_378,N_2269);
and U3571 (N_3571,N_1322,N_996);
nor U3572 (N_3572,N_1829,N_213);
nand U3573 (N_3573,N_599,N_2384);
or U3574 (N_3574,N_1002,N_1836);
or U3575 (N_3575,N_310,N_1293);
nor U3576 (N_3576,N_781,N_319);
xnor U3577 (N_3577,N_392,N_816);
and U3578 (N_3578,N_544,N_1774);
and U3579 (N_3579,N_841,N_854);
nor U3580 (N_3580,N_2154,N_485);
or U3581 (N_3581,N_2042,N_360);
or U3582 (N_3582,N_1796,N_2342);
nand U3583 (N_3583,N_903,N_1112);
xnor U3584 (N_3584,N_565,N_642);
or U3585 (N_3585,N_1260,N_1667);
xnor U3586 (N_3586,N_652,N_151);
and U3587 (N_3587,N_1393,N_1946);
or U3588 (N_3588,N_1160,N_323);
xor U3589 (N_3589,N_290,N_156);
xor U3590 (N_3590,N_750,N_459);
and U3591 (N_3591,N_184,N_333);
and U3592 (N_3592,N_2476,N_2193);
nor U3593 (N_3593,N_35,N_1231);
xnor U3594 (N_3594,N_891,N_1898);
and U3595 (N_3595,N_1331,N_465);
and U3596 (N_3596,N_177,N_1689);
or U3597 (N_3597,N_880,N_1513);
nand U3598 (N_3598,N_52,N_1684);
or U3599 (N_3599,N_1458,N_1617);
and U3600 (N_3600,N_1053,N_2210);
or U3601 (N_3601,N_2162,N_1251);
nor U3602 (N_3602,N_1129,N_1380);
or U3603 (N_3603,N_2261,N_1506);
xnor U3604 (N_3604,N_1029,N_339);
xor U3605 (N_3605,N_1146,N_613);
nor U3606 (N_3606,N_664,N_632);
and U3607 (N_3607,N_223,N_795);
nor U3608 (N_3608,N_307,N_873);
nand U3609 (N_3609,N_311,N_2300);
nor U3610 (N_3610,N_1210,N_448);
nor U3611 (N_3611,N_1574,N_832);
and U3612 (N_3612,N_2158,N_2093);
and U3613 (N_3613,N_272,N_67);
nor U3614 (N_3614,N_2147,N_1902);
nand U3615 (N_3615,N_2086,N_1142);
nand U3616 (N_3616,N_2233,N_1071);
and U3617 (N_3617,N_2306,N_1309);
and U3618 (N_3618,N_1025,N_2015);
nand U3619 (N_3619,N_1789,N_691);
and U3620 (N_3620,N_1827,N_883);
and U3621 (N_3621,N_1469,N_2179);
nand U3622 (N_3622,N_1220,N_2037);
nand U3623 (N_3623,N_2339,N_957);
or U3624 (N_3624,N_88,N_1613);
nor U3625 (N_3625,N_2264,N_164);
and U3626 (N_3626,N_1185,N_2422);
or U3627 (N_3627,N_740,N_1884);
and U3628 (N_3628,N_1699,N_1447);
or U3629 (N_3629,N_1759,N_1848);
or U3630 (N_3630,N_631,N_1636);
nand U3631 (N_3631,N_53,N_774);
xnor U3632 (N_3632,N_2379,N_1391);
nor U3633 (N_3633,N_2324,N_804);
or U3634 (N_3634,N_1921,N_1935);
and U3635 (N_3635,N_2199,N_172);
nor U3636 (N_3636,N_1639,N_1205);
xnor U3637 (N_3637,N_1748,N_2444);
or U3638 (N_3638,N_2214,N_812);
or U3639 (N_3639,N_1923,N_1555);
xor U3640 (N_3640,N_2252,N_696);
or U3641 (N_3641,N_1467,N_1030);
nor U3642 (N_3642,N_1587,N_910);
xor U3643 (N_3643,N_981,N_2033);
or U3644 (N_3644,N_2081,N_926);
and U3645 (N_3645,N_751,N_97);
nor U3646 (N_3646,N_1464,N_2328);
xor U3647 (N_3647,N_434,N_1198);
and U3648 (N_3648,N_1319,N_998);
and U3649 (N_3649,N_314,N_248);
nor U3650 (N_3650,N_1444,N_1964);
and U3651 (N_3651,N_1706,N_2254);
nor U3652 (N_3652,N_312,N_261);
nand U3653 (N_3653,N_2366,N_2218);
nor U3654 (N_3654,N_1897,N_349);
and U3655 (N_3655,N_2380,N_1831);
nor U3656 (N_3656,N_2063,N_2131);
or U3657 (N_3657,N_1575,N_2451);
or U3658 (N_3658,N_928,N_2078);
nand U3659 (N_3659,N_1432,N_1784);
nand U3660 (N_3660,N_81,N_1224);
and U3661 (N_3661,N_1279,N_670);
or U3662 (N_3662,N_341,N_1292);
or U3663 (N_3663,N_1960,N_1783);
and U3664 (N_3664,N_703,N_403);
xor U3665 (N_3665,N_525,N_2298);
nand U3666 (N_3666,N_2129,N_1193);
and U3667 (N_3667,N_486,N_941);
nand U3668 (N_3668,N_1565,N_62);
nand U3669 (N_3669,N_1929,N_1535);
or U3670 (N_3670,N_152,N_1192);
or U3671 (N_3671,N_2151,N_657);
nand U3672 (N_3672,N_443,N_628);
or U3673 (N_3673,N_1134,N_2185);
or U3674 (N_3674,N_23,N_1008);
and U3675 (N_3675,N_2460,N_2149);
nand U3676 (N_3676,N_1004,N_484);
nand U3677 (N_3677,N_1258,N_1033);
nor U3678 (N_3678,N_868,N_2050);
nor U3679 (N_3679,N_299,N_1034);
nor U3680 (N_3680,N_2441,N_2427);
xnor U3681 (N_3681,N_1249,N_2457);
nor U3682 (N_3682,N_1095,N_1927);
or U3683 (N_3683,N_2035,N_106);
nor U3684 (N_3684,N_445,N_253);
or U3685 (N_3685,N_2190,N_132);
nand U3686 (N_3686,N_920,N_493);
nand U3687 (N_3687,N_741,N_58);
nor U3688 (N_3688,N_2262,N_2112);
nand U3689 (N_3689,N_1931,N_1911);
nor U3690 (N_3690,N_517,N_171);
xnor U3691 (N_3691,N_1685,N_1885);
nand U3692 (N_3692,N_979,N_1428);
nand U3693 (N_3693,N_292,N_2398);
and U3694 (N_3694,N_91,N_1907);
and U3695 (N_3695,N_1530,N_1511);
and U3696 (N_3696,N_1860,N_2280);
and U3697 (N_3697,N_1221,N_1470);
xnor U3698 (N_3698,N_654,N_368);
or U3699 (N_3699,N_178,N_1650);
and U3700 (N_3700,N_273,N_2208);
or U3701 (N_3701,N_15,N_596);
nor U3702 (N_3702,N_102,N_1168);
xnor U3703 (N_3703,N_720,N_2488);
and U3704 (N_3704,N_636,N_1629);
nand U3705 (N_3705,N_2053,N_364);
xnor U3706 (N_3706,N_38,N_28);
nand U3707 (N_3707,N_2386,N_157);
nor U3708 (N_3708,N_1766,N_1798);
or U3709 (N_3709,N_2056,N_16);
or U3710 (N_3710,N_2495,N_1397);
or U3711 (N_3711,N_185,N_1601);
nand U3712 (N_3712,N_1015,N_1600);
and U3713 (N_3713,N_1770,N_713);
nand U3714 (N_3714,N_1872,N_122);
or U3715 (N_3715,N_858,N_1625);
nor U3716 (N_3716,N_1854,N_735);
nor U3717 (N_3717,N_1505,N_2409);
and U3718 (N_3718,N_512,N_682);
or U3719 (N_3719,N_179,N_2312);
nor U3720 (N_3720,N_1032,N_1194);
or U3721 (N_3721,N_1700,N_317);
nand U3722 (N_3722,N_1358,N_1156);
and U3723 (N_3723,N_1099,N_1434);
or U3724 (N_3724,N_427,N_1825);
and U3725 (N_3725,N_1433,N_573);
and U3726 (N_3726,N_1822,N_117);
nor U3727 (N_3727,N_909,N_844);
nand U3728 (N_3728,N_1026,N_1886);
nor U3729 (N_3729,N_421,N_283);
and U3730 (N_3730,N_344,N_1017);
nand U3731 (N_3731,N_2169,N_2128);
xor U3732 (N_3732,N_2025,N_556);
xnor U3733 (N_3733,N_34,N_1948);
xor U3734 (N_3734,N_2197,N_2461);
nor U3735 (N_3735,N_1678,N_2494);
nand U3736 (N_3736,N_1981,N_1753);
xor U3737 (N_3737,N_1978,N_2192);
nand U3738 (N_3738,N_83,N_598);
and U3739 (N_3739,N_168,N_2263);
nor U3740 (N_3740,N_1760,N_472);
xor U3741 (N_3741,N_677,N_1110);
nand U3742 (N_3742,N_1137,N_516);
nor U3743 (N_3743,N_2144,N_671);
xnor U3744 (N_3744,N_2390,N_1941);
nand U3745 (N_3745,N_656,N_911);
xor U3746 (N_3746,N_2371,N_1994);
and U3747 (N_3747,N_2496,N_308);
nand U3748 (N_3748,N_1068,N_2167);
nor U3749 (N_3749,N_2354,N_2475);
nor U3750 (N_3750,N_2089,N_107);
nor U3751 (N_3751,N_1024,N_1782);
xor U3752 (N_3752,N_988,N_1878);
xnor U3753 (N_3753,N_2315,N_1005);
and U3754 (N_3754,N_1655,N_928);
nor U3755 (N_3755,N_379,N_2355);
nand U3756 (N_3756,N_1533,N_729);
or U3757 (N_3757,N_867,N_828);
and U3758 (N_3758,N_927,N_2254);
nand U3759 (N_3759,N_274,N_749);
nor U3760 (N_3760,N_2448,N_424);
xor U3761 (N_3761,N_1466,N_1327);
and U3762 (N_3762,N_2348,N_286);
and U3763 (N_3763,N_2074,N_1092);
and U3764 (N_3764,N_675,N_848);
and U3765 (N_3765,N_1811,N_31);
or U3766 (N_3766,N_776,N_2069);
or U3767 (N_3767,N_181,N_1469);
or U3768 (N_3768,N_1824,N_1352);
nor U3769 (N_3769,N_71,N_2021);
and U3770 (N_3770,N_1137,N_823);
nor U3771 (N_3771,N_2194,N_615);
nor U3772 (N_3772,N_2234,N_1970);
nor U3773 (N_3773,N_648,N_23);
xnor U3774 (N_3774,N_1818,N_784);
or U3775 (N_3775,N_2382,N_2226);
and U3776 (N_3776,N_910,N_683);
and U3777 (N_3777,N_1419,N_1484);
nand U3778 (N_3778,N_1948,N_1823);
nor U3779 (N_3779,N_1670,N_1327);
nor U3780 (N_3780,N_119,N_116);
nor U3781 (N_3781,N_2434,N_1716);
and U3782 (N_3782,N_47,N_54);
nor U3783 (N_3783,N_951,N_1248);
nor U3784 (N_3784,N_166,N_2054);
and U3785 (N_3785,N_1844,N_1);
nor U3786 (N_3786,N_1881,N_1837);
nor U3787 (N_3787,N_2332,N_481);
and U3788 (N_3788,N_818,N_41);
nor U3789 (N_3789,N_379,N_1443);
xor U3790 (N_3790,N_1014,N_32);
nand U3791 (N_3791,N_907,N_5);
and U3792 (N_3792,N_1820,N_2145);
nor U3793 (N_3793,N_1198,N_515);
nand U3794 (N_3794,N_1888,N_1375);
or U3795 (N_3795,N_578,N_1168);
or U3796 (N_3796,N_2249,N_717);
nor U3797 (N_3797,N_1071,N_1643);
xnor U3798 (N_3798,N_1509,N_1159);
xor U3799 (N_3799,N_28,N_2468);
or U3800 (N_3800,N_1890,N_809);
and U3801 (N_3801,N_1514,N_514);
or U3802 (N_3802,N_2243,N_2202);
or U3803 (N_3803,N_2246,N_2277);
nor U3804 (N_3804,N_994,N_2090);
xnor U3805 (N_3805,N_900,N_941);
nor U3806 (N_3806,N_966,N_335);
and U3807 (N_3807,N_1236,N_447);
nand U3808 (N_3808,N_1473,N_1286);
nand U3809 (N_3809,N_768,N_424);
nor U3810 (N_3810,N_1812,N_2125);
nand U3811 (N_3811,N_2297,N_2199);
nand U3812 (N_3812,N_955,N_813);
or U3813 (N_3813,N_1531,N_738);
and U3814 (N_3814,N_158,N_744);
xnor U3815 (N_3815,N_1397,N_1193);
or U3816 (N_3816,N_691,N_2327);
or U3817 (N_3817,N_1754,N_476);
and U3818 (N_3818,N_1411,N_1292);
or U3819 (N_3819,N_1107,N_1877);
and U3820 (N_3820,N_34,N_628);
and U3821 (N_3821,N_868,N_2191);
nand U3822 (N_3822,N_1514,N_1028);
nor U3823 (N_3823,N_929,N_1425);
xor U3824 (N_3824,N_1086,N_2368);
xnor U3825 (N_3825,N_1593,N_1020);
and U3826 (N_3826,N_1253,N_1531);
xor U3827 (N_3827,N_1032,N_2217);
nand U3828 (N_3828,N_1154,N_548);
and U3829 (N_3829,N_1550,N_62);
and U3830 (N_3830,N_1170,N_1801);
xor U3831 (N_3831,N_233,N_1836);
nor U3832 (N_3832,N_511,N_2222);
and U3833 (N_3833,N_1188,N_1400);
nand U3834 (N_3834,N_1760,N_92);
or U3835 (N_3835,N_2456,N_906);
or U3836 (N_3836,N_1887,N_1378);
xnor U3837 (N_3837,N_510,N_2368);
xor U3838 (N_3838,N_2324,N_1752);
nor U3839 (N_3839,N_2409,N_2219);
nor U3840 (N_3840,N_10,N_709);
nor U3841 (N_3841,N_1103,N_2241);
nor U3842 (N_3842,N_1703,N_531);
or U3843 (N_3843,N_1847,N_2489);
nor U3844 (N_3844,N_89,N_859);
nor U3845 (N_3845,N_1153,N_2375);
and U3846 (N_3846,N_2405,N_355);
or U3847 (N_3847,N_2371,N_764);
and U3848 (N_3848,N_1035,N_1335);
nor U3849 (N_3849,N_1481,N_220);
xor U3850 (N_3850,N_243,N_244);
nand U3851 (N_3851,N_1227,N_2496);
nand U3852 (N_3852,N_751,N_257);
and U3853 (N_3853,N_2361,N_965);
xnor U3854 (N_3854,N_1335,N_1364);
xnor U3855 (N_3855,N_1413,N_1088);
nor U3856 (N_3856,N_911,N_1390);
nor U3857 (N_3857,N_987,N_1599);
nor U3858 (N_3858,N_2440,N_510);
xnor U3859 (N_3859,N_74,N_416);
xor U3860 (N_3860,N_761,N_1369);
xnor U3861 (N_3861,N_648,N_2037);
and U3862 (N_3862,N_32,N_1757);
nor U3863 (N_3863,N_1602,N_1420);
and U3864 (N_3864,N_1205,N_1896);
or U3865 (N_3865,N_774,N_1346);
and U3866 (N_3866,N_485,N_1193);
or U3867 (N_3867,N_367,N_1889);
xnor U3868 (N_3868,N_1701,N_2327);
and U3869 (N_3869,N_1229,N_1172);
or U3870 (N_3870,N_533,N_867);
and U3871 (N_3871,N_1027,N_339);
or U3872 (N_3872,N_1893,N_668);
xnor U3873 (N_3873,N_1762,N_1058);
xnor U3874 (N_3874,N_1743,N_396);
nand U3875 (N_3875,N_1470,N_955);
nand U3876 (N_3876,N_875,N_467);
xor U3877 (N_3877,N_328,N_1171);
and U3878 (N_3878,N_2378,N_421);
and U3879 (N_3879,N_577,N_1351);
nor U3880 (N_3880,N_284,N_2463);
or U3881 (N_3881,N_54,N_1862);
nand U3882 (N_3882,N_1552,N_1250);
xnor U3883 (N_3883,N_2473,N_1570);
and U3884 (N_3884,N_742,N_235);
and U3885 (N_3885,N_1913,N_138);
nand U3886 (N_3886,N_218,N_1821);
xor U3887 (N_3887,N_964,N_1036);
or U3888 (N_3888,N_885,N_1329);
xor U3889 (N_3889,N_1286,N_395);
and U3890 (N_3890,N_1431,N_476);
and U3891 (N_3891,N_421,N_639);
nand U3892 (N_3892,N_1672,N_887);
xor U3893 (N_3893,N_276,N_563);
or U3894 (N_3894,N_602,N_918);
or U3895 (N_3895,N_1309,N_1729);
and U3896 (N_3896,N_2445,N_183);
and U3897 (N_3897,N_2127,N_2496);
nand U3898 (N_3898,N_1923,N_2275);
and U3899 (N_3899,N_771,N_873);
nor U3900 (N_3900,N_1790,N_453);
nor U3901 (N_3901,N_2138,N_1249);
and U3902 (N_3902,N_1087,N_2420);
or U3903 (N_3903,N_193,N_1470);
nand U3904 (N_3904,N_1689,N_1369);
xor U3905 (N_3905,N_1291,N_1822);
nor U3906 (N_3906,N_1196,N_378);
or U3907 (N_3907,N_1473,N_1711);
nand U3908 (N_3908,N_749,N_454);
nor U3909 (N_3909,N_98,N_319);
or U3910 (N_3910,N_1751,N_2453);
or U3911 (N_3911,N_1145,N_1970);
nor U3912 (N_3912,N_2491,N_2066);
and U3913 (N_3913,N_553,N_2025);
nor U3914 (N_3914,N_1703,N_1328);
and U3915 (N_3915,N_1527,N_368);
or U3916 (N_3916,N_551,N_632);
nor U3917 (N_3917,N_495,N_987);
nand U3918 (N_3918,N_702,N_1039);
nor U3919 (N_3919,N_2272,N_611);
or U3920 (N_3920,N_1452,N_903);
and U3921 (N_3921,N_946,N_93);
or U3922 (N_3922,N_1595,N_22);
and U3923 (N_3923,N_2334,N_621);
or U3924 (N_3924,N_459,N_1202);
or U3925 (N_3925,N_485,N_1597);
or U3926 (N_3926,N_161,N_552);
xnor U3927 (N_3927,N_586,N_841);
and U3928 (N_3928,N_2332,N_525);
nor U3929 (N_3929,N_1010,N_2216);
or U3930 (N_3930,N_1006,N_1401);
nand U3931 (N_3931,N_398,N_497);
nor U3932 (N_3932,N_436,N_697);
xnor U3933 (N_3933,N_547,N_2008);
nand U3934 (N_3934,N_203,N_1530);
or U3935 (N_3935,N_1018,N_2159);
nor U3936 (N_3936,N_520,N_1462);
xnor U3937 (N_3937,N_572,N_1935);
nand U3938 (N_3938,N_754,N_1215);
or U3939 (N_3939,N_1892,N_1299);
and U3940 (N_3940,N_1345,N_8);
or U3941 (N_3941,N_1119,N_1868);
or U3942 (N_3942,N_1297,N_2361);
nor U3943 (N_3943,N_2433,N_1825);
nand U3944 (N_3944,N_1075,N_1707);
xor U3945 (N_3945,N_1321,N_1947);
nand U3946 (N_3946,N_1927,N_2340);
nor U3947 (N_3947,N_276,N_2205);
and U3948 (N_3948,N_185,N_616);
or U3949 (N_3949,N_2268,N_1709);
xor U3950 (N_3950,N_1996,N_1623);
nor U3951 (N_3951,N_1753,N_449);
and U3952 (N_3952,N_10,N_1707);
xnor U3953 (N_3953,N_2172,N_2143);
nor U3954 (N_3954,N_210,N_1924);
nor U3955 (N_3955,N_1778,N_2120);
nand U3956 (N_3956,N_6,N_10);
nor U3957 (N_3957,N_218,N_1902);
xnor U3958 (N_3958,N_398,N_423);
nand U3959 (N_3959,N_1001,N_2297);
xor U3960 (N_3960,N_558,N_548);
nand U3961 (N_3961,N_2114,N_1033);
nor U3962 (N_3962,N_1830,N_1263);
nand U3963 (N_3963,N_134,N_708);
nor U3964 (N_3964,N_103,N_2113);
and U3965 (N_3965,N_1263,N_898);
or U3966 (N_3966,N_1681,N_44);
or U3967 (N_3967,N_1299,N_125);
or U3968 (N_3968,N_1736,N_1679);
nor U3969 (N_3969,N_2125,N_572);
nor U3970 (N_3970,N_292,N_1808);
nor U3971 (N_3971,N_2130,N_1476);
or U3972 (N_3972,N_1762,N_2306);
nand U3973 (N_3973,N_1235,N_1177);
xnor U3974 (N_3974,N_1753,N_1792);
or U3975 (N_3975,N_856,N_915);
and U3976 (N_3976,N_1303,N_1805);
or U3977 (N_3977,N_1742,N_2466);
xnor U3978 (N_3978,N_1242,N_2255);
nor U3979 (N_3979,N_2397,N_2476);
and U3980 (N_3980,N_2377,N_2101);
and U3981 (N_3981,N_1323,N_1653);
xnor U3982 (N_3982,N_830,N_851);
nor U3983 (N_3983,N_623,N_177);
nand U3984 (N_3984,N_1779,N_188);
or U3985 (N_3985,N_1003,N_24);
nand U3986 (N_3986,N_2414,N_1434);
xor U3987 (N_3987,N_2459,N_2219);
or U3988 (N_3988,N_844,N_728);
or U3989 (N_3989,N_449,N_1953);
or U3990 (N_3990,N_1206,N_2165);
or U3991 (N_3991,N_2447,N_76);
and U3992 (N_3992,N_428,N_262);
xnor U3993 (N_3993,N_645,N_2451);
nor U3994 (N_3994,N_1256,N_1581);
xor U3995 (N_3995,N_398,N_312);
nand U3996 (N_3996,N_269,N_1095);
nand U3997 (N_3997,N_2491,N_2168);
nand U3998 (N_3998,N_445,N_950);
or U3999 (N_3999,N_1178,N_2070);
or U4000 (N_4000,N_2434,N_2398);
xnor U4001 (N_4001,N_1473,N_144);
and U4002 (N_4002,N_907,N_1441);
nor U4003 (N_4003,N_1360,N_561);
nand U4004 (N_4004,N_189,N_173);
or U4005 (N_4005,N_2294,N_1524);
and U4006 (N_4006,N_2001,N_1671);
nor U4007 (N_4007,N_534,N_2008);
nor U4008 (N_4008,N_1330,N_1522);
xor U4009 (N_4009,N_1587,N_1443);
or U4010 (N_4010,N_366,N_1574);
xor U4011 (N_4011,N_976,N_40);
and U4012 (N_4012,N_2139,N_1429);
nand U4013 (N_4013,N_1810,N_2410);
and U4014 (N_4014,N_2423,N_10);
xor U4015 (N_4015,N_618,N_1121);
or U4016 (N_4016,N_616,N_1042);
nand U4017 (N_4017,N_1310,N_1647);
or U4018 (N_4018,N_27,N_2158);
nand U4019 (N_4019,N_354,N_884);
nor U4020 (N_4020,N_1851,N_2145);
and U4021 (N_4021,N_1304,N_1954);
xor U4022 (N_4022,N_205,N_735);
xor U4023 (N_4023,N_491,N_2176);
or U4024 (N_4024,N_993,N_1883);
xnor U4025 (N_4025,N_281,N_1948);
nor U4026 (N_4026,N_2398,N_795);
xor U4027 (N_4027,N_2473,N_1318);
and U4028 (N_4028,N_1040,N_1761);
and U4029 (N_4029,N_2288,N_1368);
or U4030 (N_4030,N_2475,N_596);
nand U4031 (N_4031,N_396,N_1597);
and U4032 (N_4032,N_1724,N_2177);
or U4033 (N_4033,N_1449,N_1645);
xnor U4034 (N_4034,N_1788,N_2356);
or U4035 (N_4035,N_1523,N_1210);
and U4036 (N_4036,N_311,N_92);
nor U4037 (N_4037,N_855,N_223);
nand U4038 (N_4038,N_82,N_1773);
or U4039 (N_4039,N_1461,N_1615);
xnor U4040 (N_4040,N_1629,N_284);
xor U4041 (N_4041,N_2283,N_1311);
and U4042 (N_4042,N_286,N_2222);
xor U4043 (N_4043,N_2153,N_1589);
nor U4044 (N_4044,N_1681,N_295);
nor U4045 (N_4045,N_1105,N_795);
or U4046 (N_4046,N_1992,N_264);
xnor U4047 (N_4047,N_315,N_1929);
nand U4048 (N_4048,N_2347,N_766);
and U4049 (N_4049,N_691,N_630);
nand U4050 (N_4050,N_2028,N_1518);
and U4051 (N_4051,N_1373,N_853);
nand U4052 (N_4052,N_753,N_2127);
xnor U4053 (N_4053,N_1789,N_1825);
or U4054 (N_4054,N_157,N_926);
nor U4055 (N_4055,N_407,N_1581);
nand U4056 (N_4056,N_1268,N_1776);
or U4057 (N_4057,N_1656,N_478);
or U4058 (N_4058,N_393,N_1374);
and U4059 (N_4059,N_2222,N_2099);
or U4060 (N_4060,N_779,N_1775);
and U4061 (N_4061,N_2248,N_813);
and U4062 (N_4062,N_2078,N_1198);
and U4063 (N_4063,N_1309,N_1419);
or U4064 (N_4064,N_855,N_229);
nor U4065 (N_4065,N_1721,N_818);
nor U4066 (N_4066,N_2429,N_331);
nand U4067 (N_4067,N_1448,N_2210);
nor U4068 (N_4068,N_492,N_1039);
or U4069 (N_4069,N_2282,N_2188);
xnor U4070 (N_4070,N_2094,N_2349);
and U4071 (N_4071,N_2477,N_2156);
or U4072 (N_4072,N_1798,N_2204);
or U4073 (N_4073,N_1918,N_2395);
xnor U4074 (N_4074,N_556,N_2413);
and U4075 (N_4075,N_1852,N_2028);
nor U4076 (N_4076,N_358,N_1206);
or U4077 (N_4077,N_2214,N_1069);
xnor U4078 (N_4078,N_1608,N_2217);
and U4079 (N_4079,N_1040,N_2215);
or U4080 (N_4080,N_1585,N_1987);
nand U4081 (N_4081,N_1844,N_999);
or U4082 (N_4082,N_974,N_1593);
nand U4083 (N_4083,N_2150,N_1413);
nand U4084 (N_4084,N_1765,N_279);
xnor U4085 (N_4085,N_1508,N_1268);
nor U4086 (N_4086,N_1542,N_2253);
or U4087 (N_4087,N_1091,N_761);
and U4088 (N_4088,N_1792,N_2473);
or U4089 (N_4089,N_2422,N_34);
or U4090 (N_4090,N_2018,N_1325);
and U4091 (N_4091,N_1067,N_1253);
xnor U4092 (N_4092,N_910,N_666);
and U4093 (N_4093,N_2039,N_2420);
xor U4094 (N_4094,N_1081,N_607);
or U4095 (N_4095,N_2185,N_579);
or U4096 (N_4096,N_2183,N_2358);
nand U4097 (N_4097,N_2010,N_2091);
nor U4098 (N_4098,N_2458,N_85);
xnor U4099 (N_4099,N_304,N_1419);
or U4100 (N_4100,N_2243,N_89);
nor U4101 (N_4101,N_243,N_1451);
xnor U4102 (N_4102,N_1972,N_114);
or U4103 (N_4103,N_1103,N_766);
xnor U4104 (N_4104,N_76,N_1343);
nand U4105 (N_4105,N_1640,N_2038);
nor U4106 (N_4106,N_1844,N_1608);
nor U4107 (N_4107,N_59,N_734);
nor U4108 (N_4108,N_982,N_1449);
and U4109 (N_4109,N_1270,N_1242);
nor U4110 (N_4110,N_649,N_1222);
and U4111 (N_4111,N_2461,N_488);
nor U4112 (N_4112,N_1595,N_2348);
nand U4113 (N_4113,N_783,N_965);
xnor U4114 (N_4114,N_1244,N_396);
and U4115 (N_4115,N_562,N_788);
nor U4116 (N_4116,N_551,N_2254);
and U4117 (N_4117,N_1244,N_356);
or U4118 (N_4118,N_2475,N_1726);
nor U4119 (N_4119,N_1355,N_2396);
and U4120 (N_4120,N_102,N_646);
nand U4121 (N_4121,N_1852,N_88);
xnor U4122 (N_4122,N_2311,N_2267);
nor U4123 (N_4123,N_2420,N_2153);
xnor U4124 (N_4124,N_922,N_1524);
and U4125 (N_4125,N_1902,N_2441);
or U4126 (N_4126,N_135,N_1858);
nor U4127 (N_4127,N_2276,N_800);
xnor U4128 (N_4128,N_213,N_385);
or U4129 (N_4129,N_1282,N_663);
or U4130 (N_4130,N_1479,N_1296);
nand U4131 (N_4131,N_1667,N_1806);
nor U4132 (N_4132,N_847,N_2248);
or U4133 (N_4133,N_570,N_2399);
xnor U4134 (N_4134,N_1701,N_1832);
or U4135 (N_4135,N_854,N_1737);
xnor U4136 (N_4136,N_2136,N_2199);
or U4137 (N_4137,N_903,N_442);
xor U4138 (N_4138,N_1898,N_1292);
nand U4139 (N_4139,N_1073,N_1002);
and U4140 (N_4140,N_967,N_1316);
xor U4141 (N_4141,N_732,N_1762);
and U4142 (N_4142,N_1248,N_1985);
xnor U4143 (N_4143,N_1951,N_2316);
nor U4144 (N_4144,N_2332,N_1466);
and U4145 (N_4145,N_1910,N_1515);
or U4146 (N_4146,N_1743,N_1630);
and U4147 (N_4147,N_171,N_1944);
and U4148 (N_4148,N_2237,N_725);
nor U4149 (N_4149,N_1743,N_1265);
nand U4150 (N_4150,N_1480,N_1848);
and U4151 (N_4151,N_1578,N_799);
and U4152 (N_4152,N_1958,N_1638);
or U4153 (N_4153,N_965,N_297);
and U4154 (N_4154,N_1317,N_1176);
xor U4155 (N_4155,N_1823,N_241);
nor U4156 (N_4156,N_1330,N_2231);
xor U4157 (N_4157,N_688,N_1568);
nand U4158 (N_4158,N_1771,N_733);
or U4159 (N_4159,N_928,N_1423);
nand U4160 (N_4160,N_2409,N_2241);
xnor U4161 (N_4161,N_914,N_769);
and U4162 (N_4162,N_2044,N_2210);
or U4163 (N_4163,N_181,N_1650);
nor U4164 (N_4164,N_2365,N_1620);
or U4165 (N_4165,N_2491,N_312);
nor U4166 (N_4166,N_1101,N_1585);
nor U4167 (N_4167,N_1528,N_1901);
and U4168 (N_4168,N_1986,N_131);
and U4169 (N_4169,N_1366,N_1721);
and U4170 (N_4170,N_485,N_1092);
xor U4171 (N_4171,N_2094,N_697);
xnor U4172 (N_4172,N_1394,N_2366);
nand U4173 (N_4173,N_1709,N_2146);
and U4174 (N_4174,N_281,N_2144);
nand U4175 (N_4175,N_1648,N_626);
and U4176 (N_4176,N_1887,N_77);
nor U4177 (N_4177,N_1910,N_1407);
or U4178 (N_4178,N_719,N_92);
xor U4179 (N_4179,N_1364,N_183);
nand U4180 (N_4180,N_2494,N_527);
and U4181 (N_4181,N_2131,N_0);
nand U4182 (N_4182,N_1006,N_366);
or U4183 (N_4183,N_1601,N_1210);
nand U4184 (N_4184,N_994,N_2146);
and U4185 (N_4185,N_1030,N_1998);
nand U4186 (N_4186,N_1407,N_329);
and U4187 (N_4187,N_676,N_1908);
xor U4188 (N_4188,N_2499,N_1359);
and U4189 (N_4189,N_596,N_570);
and U4190 (N_4190,N_2146,N_1303);
and U4191 (N_4191,N_2395,N_793);
nor U4192 (N_4192,N_657,N_1419);
nor U4193 (N_4193,N_2173,N_1939);
nand U4194 (N_4194,N_2356,N_2015);
nand U4195 (N_4195,N_1412,N_1831);
nor U4196 (N_4196,N_1613,N_228);
and U4197 (N_4197,N_2066,N_2291);
nand U4198 (N_4198,N_2117,N_2158);
and U4199 (N_4199,N_2421,N_1921);
xor U4200 (N_4200,N_1522,N_195);
or U4201 (N_4201,N_638,N_2427);
or U4202 (N_4202,N_895,N_1190);
nor U4203 (N_4203,N_988,N_1407);
nor U4204 (N_4204,N_2443,N_989);
nor U4205 (N_4205,N_462,N_522);
nand U4206 (N_4206,N_494,N_2125);
nor U4207 (N_4207,N_2212,N_1859);
and U4208 (N_4208,N_560,N_2095);
or U4209 (N_4209,N_1814,N_109);
nor U4210 (N_4210,N_790,N_1652);
or U4211 (N_4211,N_1244,N_55);
or U4212 (N_4212,N_2034,N_1111);
or U4213 (N_4213,N_2004,N_313);
nand U4214 (N_4214,N_834,N_1941);
nor U4215 (N_4215,N_1920,N_980);
nand U4216 (N_4216,N_47,N_2159);
xnor U4217 (N_4217,N_778,N_898);
nor U4218 (N_4218,N_2078,N_649);
or U4219 (N_4219,N_1995,N_750);
xor U4220 (N_4220,N_74,N_987);
and U4221 (N_4221,N_836,N_706);
or U4222 (N_4222,N_111,N_178);
xor U4223 (N_4223,N_604,N_2155);
nand U4224 (N_4224,N_449,N_376);
nor U4225 (N_4225,N_2443,N_166);
or U4226 (N_4226,N_62,N_113);
xnor U4227 (N_4227,N_611,N_75);
or U4228 (N_4228,N_605,N_1211);
nor U4229 (N_4229,N_2124,N_617);
xor U4230 (N_4230,N_2431,N_128);
and U4231 (N_4231,N_507,N_377);
or U4232 (N_4232,N_701,N_232);
or U4233 (N_4233,N_698,N_1903);
or U4234 (N_4234,N_2094,N_2186);
and U4235 (N_4235,N_2473,N_54);
and U4236 (N_4236,N_1834,N_2410);
xor U4237 (N_4237,N_560,N_241);
or U4238 (N_4238,N_276,N_1222);
xor U4239 (N_4239,N_289,N_2391);
nand U4240 (N_4240,N_1221,N_768);
nor U4241 (N_4241,N_412,N_1072);
and U4242 (N_4242,N_278,N_1222);
and U4243 (N_4243,N_1823,N_263);
nor U4244 (N_4244,N_1831,N_1509);
nor U4245 (N_4245,N_872,N_984);
or U4246 (N_4246,N_22,N_2021);
xnor U4247 (N_4247,N_1028,N_2443);
nor U4248 (N_4248,N_559,N_198);
xor U4249 (N_4249,N_2292,N_2465);
nor U4250 (N_4250,N_311,N_148);
or U4251 (N_4251,N_2243,N_1392);
or U4252 (N_4252,N_2049,N_1618);
xor U4253 (N_4253,N_1237,N_652);
and U4254 (N_4254,N_265,N_1654);
xor U4255 (N_4255,N_1047,N_1139);
nor U4256 (N_4256,N_1760,N_1093);
and U4257 (N_4257,N_2444,N_1411);
and U4258 (N_4258,N_267,N_1315);
and U4259 (N_4259,N_2290,N_551);
nor U4260 (N_4260,N_2097,N_2015);
nand U4261 (N_4261,N_1045,N_2386);
and U4262 (N_4262,N_2467,N_2446);
xor U4263 (N_4263,N_1369,N_2283);
and U4264 (N_4264,N_131,N_1970);
nor U4265 (N_4265,N_2342,N_807);
or U4266 (N_4266,N_382,N_1061);
xnor U4267 (N_4267,N_339,N_1803);
nand U4268 (N_4268,N_315,N_932);
and U4269 (N_4269,N_190,N_456);
nand U4270 (N_4270,N_1702,N_132);
and U4271 (N_4271,N_2193,N_1386);
or U4272 (N_4272,N_824,N_1207);
and U4273 (N_4273,N_733,N_322);
nor U4274 (N_4274,N_1526,N_2148);
and U4275 (N_4275,N_903,N_2000);
or U4276 (N_4276,N_420,N_740);
and U4277 (N_4277,N_105,N_1278);
nand U4278 (N_4278,N_2238,N_2072);
and U4279 (N_4279,N_580,N_1089);
nor U4280 (N_4280,N_583,N_423);
nor U4281 (N_4281,N_2101,N_1104);
and U4282 (N_4282,N_1645,N_1881);
or U4283 (N_4283,N_1263,N_106);
xor U4284 (N_4284,N_2263,N_669);
nor U4285 (N_4285,N_2211,N_855);
nor U4286 (N_4286,N_1305,N_1127);
nor U4287 (N_4287,N_2208,N_1111);
nor U4288 (N_4288,N_1274,N_856);
or U4289 (N_4289,N_823,N_1161);
and U4290 (N_4290,N_952,N_488);
nand U4291 (N_4291,N_2301,N_1416);
and U4292 (N_4292,N_160,N_1524);
nand U4293 (N_4293,N_1702,N_378);
nand U4294 (N_4294,N_2055,N_1186);
and U4295 (N_4295,N_1787,N_2103);
or U4296 (N_4296,N_1717,N_583);
nor U4297 (N_4297,N_1705,N_277);
or U4298 (N_4298,N_798,N_1919);
nand U4299 (N_4299,N_554,N_917);
and U4300 (N_4300,N_1795,N_820);
and U4301 (N_4301,N_564,N_1454);
xor U4302 (N_4302,N_1273,N_1899);
and U4303 (N_4303,N_730,N_1302);
nor U4304 (N_4304,N_934,N_1616);
nand U4305 (N_4305,N_1702,N_1853);
nand U4306 (N_4306,N_1877,N_767);
xor U4307 (N_4307,N_1639,N_705);
nor U4308 (N_4308,N_486,N_1515);
xor U4309 (N_4309,N_138,N_995);
nor U4310 (N_4310,N_2166,N_2369);
nand U4311 (N_4311,N_1059,N_2422);
and U4312 (N_4312,N_2033,N_1337);
or U4313 (N_4313,N_764,N_1439);
nand U4314 (N_4314,N_831,N_51);
xnor U4315 (N_4315,N_1979,N_2242);
nand U4316 (N_4316,N_2006,N_24);
and U4317 (N_4317,N_1509,N_2330);
nor U4318 (N_4318,N_1837,N_1766);
and U4319 (N_4319,N_879,N_1008);
xnor U4320 (N_4320,N_1396,N_2425);
nor U4321 (N_4321,N_1230,N_2456);
or U4322 (N_4322,N_851,N_77);
nand U4323 (N_4323,N_2440,N_2343);
xor U4324 (N_4324,N_2463,N_1797);
xnor U4325 (N_4325,N_152,N_2464);
or U4326 (N_4326,N_291,N_1558);
nand U4327 (N_4327,N_1961,N_111);
and U4328 (N_4328,N_1060,N_1728);
or U4329 (N_4329,N_1671,N_1065);
nand U4330 (N_4330,N_1018,N_1142);
nor U4331 (N_4331,N_1992,N_1220);
xor U4332 (N_4332,N_2048,N_740);
nor U4333 (N_4333,N_1718,N_2055);
nand U4334 (N_4334,N_1752,N_2070);
nor U4335 (N_4335,N_2460,N_1291);
or U4336 (N_4336,N_2399,N_632);
xnor U4337 (N_4337,N_1703,N_346);
or U4338 (N_4338,N_221,N_300);
nand U4339 (N_4339,N_235,N_26);
nor U4340 (N_4340,N_1399,N_910);
nand U4341 (N_4341,N_2374,N_964);
and U4342 (N_4342,N_1519,N_2126);
nand U4343 (N_4343,N_441,N_489);
or U4344 (N_4344,N_1404,N_1389);
and U4345 (N_4345,N_365,N_2073);
or U4346 (N_4346,N_1192,N_1555);
or U4347 (N_4347,N_448,N_1999);
nand U4348 (N_4348,N_581,N_453);
or U4349 (N_4349,N_1543,N_312);
and U4350 (N_4350,N_2060,N_2145);
or U4351 (N_4351,N_1947,N_349);
nand U4352 (N_4352,N_1349,N_9);
and U4353 (N_4353,N_2223,N_1817);
nor U4354 (N_4354,N_2383,N_24);
nand U4355 (N_4355,N_1062,N_45);
or U4356 (N_4356,N_1635,N_2011);
nor U4357 (N_4357,N_1270,N_2094);
xnor U4358 (N_4358,N_2002,N_1218);
nor U4359 (N_4359,N_1796,N_2164);
nand U4360 (N_4360,N_118,N_554);
nand U4361 (N_4361,N_2238,N_1500);
and U4362 (N_4362,N_1144,N_93);
and U4363 (N_4363,N_146,N_81);
nand U4364 (N_4364,N_569,N_281);
or U4365 (N_4365,N_203,N_1452);
or U4366 (N_4366,N_2443,N_729);
and U4367 (N_4367,N_2047,N_262);
xnor U4368 (N_4368,N_1406,N_117);
or U4369 (N_4369,N_1240,N_893);
nor U4370 (N_4370,N_893,N_2237);
or U4371 (N_4371,N_309,N_1825);
nand U4372 (N_4372,N_1612,N_1738);
nand U4373 (N_4373,N_1375,N_882);
nor U4374 (N_4374,N_900,N_1729);
nor U4375 (N_4375,N_58,N_521);
and U4376 (N_4376,N_2248,N_1147);
nand U4377 (N_4377,N_766,N_1856);
or U4378 (N_4378,N_1194,N_1804);
or U4379 (N_4379,N_2179,N_148);
or U4380 (N_4380,N_1698,N_2480);
nor U4381 (N_4381,N_1022,N_1696);
nand U4382 (N_4382,N_291,N_418);
nand U4383 (N_4383,N_1696,N_2017);
nor U4384 (N_4384,N_661,N_1719);
and U4385 (N_4385,N_1133,N_1326);
and U4386 (N_4386,N_2218,N_1346);
and U4387 (N_4387,N_2290,N_839);
or U4388 (N_4388,N_2274,N_1294);
nand U4389 (N_4389,N_1607,N_2390);
and U4390 (N_4390,N_693,N_880);
nand U4391 (N_4391,N_1556,N_1635);
nand U4392 (N_4392,N_1196,N_438);
nand U4393 (N_4393,N_529,N_434);
nor U4394 (N_4394,N_842,N_905);
nor U4395 (N_4395,N_724,N_1893);
and U4396 (N_4396,N_276,N_624);
nand U4397 (N_4397,N_1026,N_1209);
nand U4398 (N_4398,N_2316,N_569);
nor U4399 (N_4399,N_54,N_2127);
or U4400 (N_4400,N_2275,N_1547);
or U4401 (N_4401,N_344,N_1353);
or U4402 (N_4402,N_399,N_528);
or U4403 (N_4403,N_462,N_1089);
xnor U4404 (N_4404,N_1009,N_1031);
or U4405 (N_4405,N_1766,N_1476);
nand U4406 (N_4406,N_1426,N_1058);
and U4407 (N_4407,N_2113,N_453);
nand U4408 (N_4408,N_406,N_545);
and U4409 (N_4409,N_1327,N_1276);
or U4410 (N_4410,N_1430,N_1062);
xnor U4411 (N_4411,N_1202,N_172);
or U4412 (N_4412,N_1036,N_1969);
or U4413 (N_4413,N_38,N_1200);
and U4414 (N_4414,N_251,N_1297);
or U4415 (N_4415,N_1612,N_489);
xnor U4416 (N_4416,N_1384,N_381);
nor U4417 (N_4417,N_2356,N_390);
or U4418 (N_4418,N_1653,N_950);
xor U4419 (N_4419,N_2153,N_1221);
and U4420 (N_4420,N_740,N_1234);
xor U4421 (N_4421,N_1653,N_1749);
nand U4422 (N_4422,N_1263,N_1443);
or U4423 (N_4423,N_1682,N_1047);
or U4424 (N_4424,N_386,N_1765);
or U4425 (N_4425,N_1138,N_1195);
nand U4426 (N_4426,N_752,N_2355);
nor U4427 (N_4427,N_669,N_1727);
xor U4428 (N_4428,N_978,N_173);
and U4429 (N_4429,N_860,N_997);
nor U4430 (N_4430,N_1756,N_2495);
and U4431 (N_4431,N_288,N_657);
nand U4432 (N_4432,N_23,N_292);
or U4433 (N_4433,N_505,N_783);
and U4434 (N_4434,N_978,N_234);
nor U4435 (N_4435,N_727,N_2262);
or U4436 (N_4436,N_278,N_2106);
xnor U4437 (N_4437,N_2431,N_885);
xor U4438 (N_4438,N_1524,N_957);
nand U4439 (N_4439,N_130,N_458);
xor U4440 (N_4440,N_2445,N_153);
or U4441 (N_4441,N_982,N_684);
nand U4442 (N_4442,N_1061,N_801);
xnor U4443 (N_4443,N_806,N_444);
or U4444 (N_4444,N_1599,N_1505);
xor U4445 (N_4445,N_1068,N_65);
and U4446 (N_4446,N_878,N_2139);
xnor U4447 (N_4447,N_834,N_1878);
nand U4448 (N_4448,N_332,N_1136);
xnor U4449 (N_4449,N_1017,N_2119);
xor U4450 (N_4450,N_57,N_862);
xor U4451 (N_4451,N_921,N_2366);
nand U4452 (N_4452,N_355,N_1953);
xor U4453 (N_4453,N_1202,N_1859);
and U4454 (N_4454,N_2348,N_1492);
or U4455 (N_4455,N_181,N_352);
nor U4456 (N_4456,N_765,N_254);
nand U4457 (N_4457,N_66,N_1583);
or U4458 (N_4458,N_1181,N_2000);
nor U4459 (N_4459,N_1634,N_73);
or U4460 (N_4460,N_1460,N_1961);
nor U4461 (N_4461,N_2334,N_520);
nor U4462 (N_4462,N_1186,N_2426);
xor U4463 (N_4463,N_173,N_454);
xnor U4464 (N_4464,N_289,N_2182);
or U4465 (N_4465,N_886,N_1789);
nand U4466 (N_4466,N_1987,N_2376);
nor U4467 (N_4467,N_2,N_2190);
nor U4468 (N_4468,N_1591,N_1040);
xor U4469 (N_4469,N_1371,N_1045);
and U4470 (N_4470,N_1650,N_796);
and U4471 (N_4471,N_841,N_2039);
or U4472 (N_4472,N_1727,N_889);
and U4473 (N_4473,N_1622,N_2102);
xnor U4474 (N_4474,N_102,N_373);
or U4475 (N_4475,N_569,N_1518);
xnor U4476 (N_4476,N_2218,N_1964);
xor U4477 (N_4477,N_1047,N_1650);
xnor U4478 (N_4478,N_336,N_2184);
nor U4479 (N_4479,N_294,N_339);
and U4480 (N_4480,N_1785,N_1466);
nor U4481 (N_4481,N_1172,N_97);
and U4482 (N_4482,N_2332,N_1804);
nand U4483 (N_4483,N_1984,N_901);
and U4484 (N_4484,N_1368,N_410);
or U4485 (N_4485,N_1396,N_1346);
nand U4486 (N_4486,N_269,N_671);
and U4487 (N_4487,N_936,N_1455);
nor U4488 (N_4488,N_541,N_1087);
and U4489 (N_4489,N_1987,N_450);
xor U4490 (N_4490,N_2181,N_2201);
and U4491 (N_4491,N_1803,N_1177);
or U4492 (N_4492,N_1438,N_1269);
and U4493 (N_4493,N_1790,N_1751);
xnor U4494 (N_4494,N_47,N_2409);
nand U4495 (N_4495,N_652,N_685);
nand U4496 (N_4496,N_1507,N_1141);
nor U4497 (N_4497,N_619,N_1621);
nor U4498 (N_4498,N_1257,N_2065);
nor U4499 (N_4499,N_2421,N_1354);
or U4500 (N_4500,N_1021,N_717);
and U4501 (N_4501,N_370,N_1802);
nor U4502 (N_4502,N_428,N_1024);
nand U4503 (N_4503,N_293,N_1768);
nand U4504 (N_4504,N_1418,N_2170);
and U4505 (N_4505,N_63,N_1839);
xnor U4506 (N_4506,N_711,N_1292);
nand U4507 (N_4507,N_146,N_1432);
nand U4508 (N_4508,N_551,N_2493);
nand U4509 (N_4509,N_2035,N_1529);
and U4510 (N_4510,N_896,N_2295);
and U4511 (N_4511,N_1785,N_935);
nand U4512 (N_4512,N_69,N_736);
nor U4513 (N_4513,N_1787,N_1748);
nor U4514 (N_4514,N_2203,N_2497);
xnor U4515 (N_4515,N_2329,N_499);
xor U4516 (N_4516,N_101,N_334);
xnor U4517 (N_4517,N_1934,N_61);
xor U4518 (N_4518,N_2440,N_61);
or U4519 (N_4519,N_1296,N_1555);
or U4520 (N_4520,N_2104,N_1278);
xnor U4521 (N_4521,N_1251,N_207);
or U4522 (N_4522,N_1731,N_2115);
and U4523 (N_4523,N_2196,N_433);
xnor U4524 (N_4524,N_1925,N_623);
xor U4525 (N_4525,N_1649,N_15);
nand U4526 (N_4526,N_283,N_1375);
nand U4527 (N_4527,N_798,N_1686);
or U4528 (N_4528,N_1144,N_1421);
and U4529 (N_4529,N_428,N_2406);
xnor U4530 (N_4530,N_1572,N_259);
or U4531 (N_4531,N_1223,N_2273);
or U4532 (N_4532,N_525,N_115);
nor U4533 (N_4533,N_1679,N_1708);
or U4534 (N_4534,N_257,N_921);
nand U4535 (N_4535,N_1021,N_1563);
and U4536 (N_4536,N_202,N_197);
nand U4537 (N_4537,N_877,N_1979);
nor U4538 (N_4538,N_1746,N_1810);
xor U4539 (N_4539,N_1907,N_1627);
or U4540 (N_4540,N_1336,N_940);
and U4541 (N_4541,N_1175,N_673);
xor U4542 (N_4542,N_819,N_1165);
and U4543 (N_4543,N_790,N_221);
nor U4544 (N_4544,N_145,N_1682);
xnor U4545 (N_4545,N_496,N_2105);
nand U4546 (N_4546,N_1960,N_371);
or U4547 (N_4547,N_1189,N_94);
and U4548 (N_4548,N_955,N_1727);
nor U4549 (N_4549,N_130,N_427);
nand U4550 (N_4550,N_2116,N_380);
nor U4551 (N_4551,N_392,N_1504);
nor U4552 (N_4552,N_2070,N_2041);
and U4553 (N_4553,N_1482,N_345);
and U4554 (N_4554,N_156,N_629);
and U4555 (N_4555,N_2024,N_1618);
or U4556 (N_4556,N_795,N_688);
nand U4557 (N_4557,N_2490,N_63);
xnor U4558 (N_4558,N_2133,N_199);
xor U4559 (N_4559,N_2182,N_1625);
nor U4560 (N_4560,N_668,N_2428);
nor U4561 (N_4561,N_675,N_1880);
nand U4562 (N_4562,N_314,N_1271);
or U4563 (N_4563,N_2035,N_1182);
and U4564 (N_4564,N_672,N_1356);
and U4565 (N_4565,N_932,N_1686);
xnor U4566 (N_4566,N_1900,N_115);
xor U4567 (N_4567,N_950,N_1369);
or U4568 (N_4568,N_2291,N_1870);
or U4569 (N_4569,N_400,N_2054);
xor U4570 (N_4570,N_2090,N_583);
or U4571 (N_4571,N_2232,N_1197);
nand U4572 (N_4572,N_31,N_992);
nor U4573 (N_4573,N_2309,N_953);
or U4574 (N_4574,N_325,N_1117);
nand U4575 (N_4575,N_2488,N_301);
or U4576 (N_4576,N_2366,N_940);
or U4577 (N_4577,N_1047,N_1469);
nor U4578 (N_4578,N_799,N_702);
or U4579 (N_4579,N_182,N_22);
and U4580 (N_4580,N_2279,N_262);
and U4581 (N_4581,N_1475,N_370);
nand U4582 (N_4582,N_353,N_2220);
or U4583 (N_4583,N_2446,N_947);
and U4584 (N_4584,N_1782,N_218);
nand U4585 (N_4585,N_2346,N_1482);
nor U4586 (N_4586,N_1597,N_9);
or U4587 (N_4587,N_1164,N_1274);
nand U4588 (N_4588,N_2430,N_257);
or U4589 (N_4589,N_2494,N_898);
xor U4590 (N_4590,N_904,N_1357);
and U4591 (N_4591,N_1179,N_2450);
and U4592 (N_4592,N_1896,N_2090);
xor U4593 (N_4593,N_1202,N_1482);
or U4594 (N_4594,N_267,N_776);
nand U4595 (N_4595,N_49,N_2451);
nand U4596 (N_4596,N_2165,N_1547);
xor U4597 (N_4597,N_641,N_692);
and U4598 (N_4598,N_2373,N_139);
and U4599 (N_4599,N_2328,N_2166);
nand U4600 (N_4600,N_1897,N_1121);
nand U4601 (N_4601,N_1487,N_1515);
xnor U4602 (N_4602,N_1913,N_1915);
or U4603 (N_4603,N_679,N_1172);
or U4604 (N_4604,N_1945,N_2041);
or U4605 (N_4605,N_1450,N_2444);
nor U4606 (N_4606,N_264,N_2235);
nor U4607 (N_4607,N_476,N_433);
nand U4608 (N_4608,N_2344,N_1425);
and U4609 (N_4609,N_997,N_2040);
nand U4610 (N_4610,N_1468,N_1130);
xnor U4611 (N_4611,N_697,N_1171);
nand U4612 (N_4612,N_1627,N_1403);
nand U4613 (N_4613,N_1105,N_819);
nor U4614 (N_4614,N_438,N_1580);
and U4615 (N_4615,N_444,N_1097);
nand U4616 (N_4616,N_1298,N_1744);
or U4617 (N_4617,N_2187,N_925);
nor U4618 (N_4618,N_233,N_1050);
and U4619 (N_4619,N_25,N_555);
nor U4620 (N_4620,N_984,N_862);
nor U4621 (N_4621,N_2223,N_1900);
nor U4622 (N_4622,N_2016,N_1781);
xnor U4623 (N_4623,N_1984,N_1465);
or U4624 (N_4624,N_1174,N_367);
xor U4625 (N_4625,N_1238,N_1094);
or U4626 (N_4626,N_1184,N_677);
nor U4627 (N_4627,N_1937,N_2260);
and U4628 (N_4628,N_1968,N_42);
and U4629 (N_4629,N_930,N_1454);
or U4630 (N_4630,N_509,N_985);
or U4631 (N_4631,N_1384,N_159);
or U4632 (N_4632,N_580,N_516);
nor U4633 (N_4633,N_1274,N_2286);
or U4634 (N_4634,N_1610,N_2209);
nor U4635 (N_4635,N_169,N_1696);
nor U4636 (N_4636,N_2081,N_1917);
nor U4637 (N_4637,N_867,N_2357);
xnor U4638 (N_4638,N_1313,N_323);
xor U4639 (N_4639,N_1886,N_2393);
nor U4640 (N_4640,N_540,N_525);
and U4641 (N_4641,N_90,N_1611);
nand U4642 (N_4642,N_2468,N_292);
nor U4643 (N_4643,N_251,N_888);
nor U4644 (N_4644,N_819,N_1869);
nand U4645 (N_4645,N_2084,N_522);
and U4646 (N_4646,N_2343,N_2388);
and U4647 (N_4647,N_1214,N_1519);
or U4648 (N_4648,N_438,N_1565);
xnor U4649 (N_4649,N_1668,N_497);
or U4650 (N_4650,N_1719,N_1118);
nand U4651 (N_4651,N_2455,N_1913);
nor U4652 (N_4652,N_1466,N_262);
and U4653 (N_4653,N_819,N_1856);
nor U4654 (N_4654,N_829,N_979);
nand U4655 (N_4655,N_472,N_1250);
or U4656 (N_4656,N_272,N_597);
or U4657 (N_4657,N_573,N_499);
xnor U4658 (N_4658,N_1681,N_844);
and U4659 (N_4659,N_2262,N_759);
and U4660 (N_4660,N_1337,N_925);
nor U4661 (N_4661,N_2273,N_7);
nor U4662 (N_4662,N_2393,N_1299);
nand U4663 (N_4663,N_2098,N_70);
and U4664 (N_4664,N_2256,N_2025);
or U4665 (N_4665,N_321,N_767);
xnor U4666 (N_4666,N_651,N_662);
nand U4667 (N_4667,N_2352,N_180);
nor U4668 (N_4668,N_832,N_1173);
and U4669 (N_4669,N_95,N_1314);
nor U4670 (N_4670,N_1174,N_1061);
nand U4671 (N_4671,N_184,N_1683);
and U4672 (N_4672,N_497,N_36);
nor U4673 (N_4673,N_2318,N_1084);
and U4674 (N_4674,N_1415,N_1754);
and U4675 (N_4675,N_2052,N_1783);
xor U4676 (N_4676,N_431,N_462);
xor U4677 (N_4677,N_1066,N_52);
nor U4678 (N_4678,N_145,N_1790);
xor U4679 (N_4679,N_198,N_194);
xor U4680 (N_4680,N_2253,N_2424);
nand U4681 (N_4681,N_608,N_21);
and U4682 (N_4682,N_799,N_4);
nand U4683 (N_4683,N_2340,N_1354);
nand U4684 (N_4684,N_1755,N_2096);
nand U4685 (N_4685,N_1400,N_316);
xor U4686 (N_4686,N_1851,N_442);
nand U4687 (N_4687,N_1886,N_2247);
or U4688 (N_4688,N_1404,N_2402);
xnor U4689 (N_4689,N_1074,N_45);
and U4690 (N_4690,N_2007,N_854);
nor U4691 (N_4691,N_1410,N_2064);
and U4692 (N_4692,N_709,N_924);
nor U4693 (N_4693,N_307,N_278);
or U4694 (N_4694,N_1400,N_1836);
nor U4695 (N_4695,N_1928,N_66);
nand U4696 (N_4696,N_1069,N_2009);
or U4697 (N_4697,N_375,N_1108);
and U4698 (N_4698,N_417,N_112);
nand U4699 (N_4699,N_2118,N_125);
and U4700 (N_4700,N_1733,N_2126);
nor U4701 (N_4701,N_1915,N_960);
or U4702 (N_4702,N_414,N_1827);
and U4703 (N_4703,N_2150,N_720);
or U4704 (N_4704,N_463,N_1912);
nor U4705 (N_4705,N_1019,N_2222);
nor U4706 (N_4706,N_696,N_743);
and U4707 (N_4707,N_1556,N_1562);
and U4708 (N_4708,N_1594,N_295);
and U4709 (N_4709,N_1609,N_405);
or U4710 (N_4710,N_305,N_1445);
and U4711 (N_4711,N_1599,N_2112);
xnor U4712 (N_4712,N_635,N_2476);
nand U4713 (N_4713,N_1348,N_543);
or U4714 (N_4714,N_2148,N_2404);
and U4715 (N_4715,N_1334,N_2495);
nand U4716 (N_4716,N_981,N_464);
nor U4717 (N_4717,N_2251,N_1101);
nor U4718 (N_4718,N_1314,N_623);
nand U4719 (N_4719,N_721,N_1637);
nor U4720 (N_4720,N_2278,N_2080);
nor U4721 (N_4721,N_1784,N_996);
xor U4722 (N_4722,N_2460,N_2399);
or U4723 (N_4723,N_885,N_2058);
or U4724 (N_4724,N_2425,N_2166);
and U4725 (N_4725,N_2052,N_897);
nor U4726 (N_4726,N_1948,N_877);
nor U4727 (N_4727,N_1623,N_2462);
nand U4728 (N_4728,N_1581,N_2294);
and U4729 (N_4729,N_1224,N_643);
xor U4730 (N_4730,N_2337,N_1647);
and U4731 (N_4731,N_1840,N_495);
or U4732 (N_4732,N_1613,N_1600);
or U4733 (N_4733,N_81,N_598);
or U4734 (N_4734,N_438,N_2326);
and U4735 (N_4735,N_1410,N_914);
or U4736 (N_4736,N_1118,N_734);
nand U4737 (N_4737,N_226,N_1309);
nor U4738 (N_4738,N_1896,N_1758);
xor U4739 (N_4739,N_1826,N_591);
or U4740 (N_4740,N_2481,N_918);
and U4741 (N_4741,N_1257,N_11);
and U4742 (N_4742,N_1641,N_892);
xnor U4743 (N_4743,N_148,N_2297);
nor U4744 (N_4744,N_2003,N_1534);
or U4745 (N_4745,N_668,N_614);
or U4746 (N_4746,N_1933,N_354);
xor U4747 (N_4747,N_291,N_1177);
nor U4748 (N_4748,N_9,N_581);
and U4749 (N_4749,N_1327,N_474);
and U4750 (N_4750,N_2334,N_1156);
and U4751 (N_4751,N_1103,N_228);
nor U4752 (N_4752,N_854,N_330);
and U4753 (N_4753,N_1132,N_534);
nand U4754 (N_4754,N_491,N_1776);
and U4755 (N_4755,N_2136,N_2162);
xnor U4756 (N_4756,N_339,N_2496);
xnor U4757 (N_4757,N_1615,N_245);
or U4758 (N_4758,N_1643,N_2301);
nor U4759 (N_4759,N_598,N_1397);
nand U4760 (N_4760,N_1241,N_2311);
or U4761 (N_4761,N_1899,N_685);
or U4762 (N_4762,N_1280,N_959);
nand U4763 (N_4763,N_679,N_1787);
nor U4764 (N_4764,N_32,N_2155);
nand U4765 (N_4765,N_895,N_2492);
and U4766 (N_4766,N_1253,N_2065);
nand U4767 (N_4767,N_2184,N_987);
nor U4768 (N_4768,N_2386,N_1428);
nor U4769 (N_4769,N_1206,N_1402);
xor U4770 (N_4770,N_667,N_1383);
nor U4771 (N_4771,N_1312,N_2317);
or U4772 (N_4772,N_271,N_1433);
xor U4773 (N_4773,N_1323,N_2426);
nor U4774 (N_4774,N_1878,N_797);
xor U4775 (N_4775,N_2303,N_691);
nor U4776 (N_4776,N_1341,N_2032);
nand U4777 (N_4777,N_943,N_1140);
or U4778 (N_4778,N_1260,N_817);
and U4779 (N_4779,N_1900,N_2100);
nor U4780 (N_4780,N_700,N_2162);
and U4781 (N_4781,N_581,N_1191);
or U4782 (N_4782,N_420,N_673);
nor U4783 (N_4783,N_94,N_465);
nand U4784 (N_4784,N_1607,N_1675);
and U4785 (N_4785,N_19,N_2028);
xnor U4786 (N_4786,N_777,N_1591);
nand U4787 (N_4787,N_2419,N_142);
xor U4788 (N_4788,N_1029,N_2091);
xnor U4789 (N_4789,N_2012,N_222);
xor U4790 (N_4790,N_1664,N_2307);
nor U4791 (N_4791,N_1157,N_398);
xor U4792 (N_4792,N_182,N_2021);
or U4793 (N_4793,N_1702,N_1767);
xor U4794 (N_4794,N_680,N_431);
xor U4795 (N_4795,N_1212,N_1843);
and U4796 (N_4796,N_1761,N_503);
or U4797 (N_4797,N_590,N_456);
nor U4798 (N_4798,N_1570,N_696);
xor U4799 (N_4799,N_2249,N_1600);
nand U4800 (N_4800,N_1757,N_497);
xnor U4801 (N_4801,N_47,N_1367);
xor U4802 (N_4802,N_2465,N_1975);
nor U4803 (N_4803,N_2487,N_2062);
and U4804 (N_4804,N_563,N_1642);
nand U4805 (N_4805,N_78,N_424);
and U4806 (N_4806,N_877,N_1635);
xnor U4807 (N_4807,N_663,N_186);
or U4808 (N_4808,N_1051,N_2391);
and U4809 (N_4809,N_2251,N_1202);
and U4810 (N_4810,N_1874,N_1061);
nand U4811 (N_4811,N_83,N_2315);
nand U4812 (N_4812,N_441,N_2199);
nand U4813 (N_4813,N_347,N_1483);
nor U4814 (N_4814,N_338,N_1845);
nor U4815 (N_4815,N_796,N_2112);
or U4816 (N_4816,N_1037,N_862);
nand U4817 (N_4817,N_353,N_1885);
or U4818 (N_4818,N_198,N_1078);
nor U4819 (N_4819,N_481,N_2095);
or U4820 (N_4820,N_1712,N_566);
nor U4821 (N_4821,N_9,N_108);
nor U4822 (N_4822,N_1812,N_2410);
nand U4823 (N_4823,N_2246,N_2019);
and U4824 (N_4824,N_207,N_2399);
or U4825 (N_4825,N_1494,N_2460);
xor U4826 (N_4826,N_9,N_2188);
and U4827 (N_4827,N_1950,N_1013);
nor U4828 (N_4828,N_1366,N_2093);
or U4829 (N_4829,N_2017,N_809);
or U4830 (N_4830,N_116,N_751);
nor U4831 (N_4831,N_90,N_2127);
nand U4832 (N_4832,N_1972,N_2133);
nand U4833 (N_4833,N_193,N_2028);
nand U4834 (N_4834,N_807,N_1602);
and U4835 (N_4835,N_2157,N_2440);
or U4836 (N_4836,N_384,N_410);
nor U4837 (N_4837,N_32,N_1632);
xnor U4838 (N_4838,N_2274,N_99);
nor U4839 (N_4839,N_56,N_1333);
and U4840 (N_4840,N_2083,N_479);
or U4841 (N_4841,N_2469,N_1527);
xnor U4842 (N_4842,N_2026,N_2257);
and U4843 (N_4843,N_245,N_21);
xor U4844 (N_4844,N_266,N_1634);
nand U4845 (N_4845,N_1114,N_1035);
or U4846 (N_4846,N_274,N_2094);
xnor U4847 (N_4847,N_238,N_293);
or U4848 (N_4848,N_957,N_2391);
and U4849 (N_4849,N_2274,N_373);
or U4850 (N_4850,N_1878,N_1121);
nor U4851 (N_4851,N_1502,N_427);
or U4852 (N_4852,N_1057,N_353);
nand U4853 (N_4853,N_398,N_1153);
and U4854 (N_4854,N_730,N_284);
or U4855 (N_4855,N_1652,N_1273);
or U4856 (N_4856,N_1054,N_1431);
or U4857 (N_4857,N_1132,N_960);
nor U4858 (N_4858,N_1780,N_463);
xnor U4859 (N_4859,N_2220,N_1120);
nand U4860 (N_4860,N_477,N_2203);
nand U4861 (N_4861,N_1038,N_1202);
and U4862 (N_4862,N_155,N_2173);
or U4863 (N_4863,N_676,N_1171);
or U4864 (N_4864,N_252,N_1181);
or U4865 (N_4865,N_313,N_1906);
or U4866 (N_4866,N_2093,N_2175);
xnor U4867 (N_4867,N_1279,N_1527);
xor U4868 (N_4868,N_1095,N_459);
or U4869 (N_4869,N_1347,N_854);
or U4870 (N_4870,N_92,N_600);
and U4871 (N_4871,N_206,N_1778);
and U4872 (N_4872,N_2131,N_113);
or U4873 (N_4873,N_2217,N_251);
xor U4874 (N_4874,N_172,N_1146);
nor U4875 (N_4875,N_1829,N_2147);
xnor U4876 (N_4876,N_1886,N_2382);
xnor U4877 (N_4877,N_2204,N_820);
or U4878 (N_4878,N_2336,N_250);
nor U4879 (N_4879,N_2145,N_920);
or U4880 (N_4880,N_2021,N_1034);
and U4881 (N_4881,N_413,N_569);
nand U4882 (N_4882,N_541,N_2421);
nand U4883 (N_4883,N_972,N_1153);
and U4884 (N_4884,N_1017,N_1023);
nand U4885 (N_4885,N_1898,N_8);
xnor U4886 (N_4886,N_1633,N_2432);
xor U4887 (N_4887,N_702,N_635);
nand U4888 (N_4888,N_2395,N_1280);
or U4889 (N_4889,N_1542,N_1521);
and U4890 (N_4890,N_2341,N_1569);
nor U4891 (N_4891,N_2066,N_781);
xor U4892 (N_4892,N_766,N_2272);
xnor U4893 (N_4893,N_860,N_2488);
nor U4894 (N_4894,N_832,N_1638);
xnor U4895 (N_4895,N_1054,N_1948);
nand U4896 (N_4896,N_1239,N_2103);
and U4897 (N_4897,N_357,N_2432);
and U4898 (N_4898,N_12,N_672);
xor U4899 (N_4899,N_364,N_1563);
xor U4900 (N_4900,N_1452,N_838);
nor U4901 (N_4901,N_2135,N_2108);
nor U4902 (N_4902,N_1949,N_1470);
nand U4903 (N_4903,N_619,N_1321);
nand U4904 (N_4904,N_1528,N_1383);
or U4905 (N_4905,N_661,N_1435);
or U4906 (N_4906,N_1442,N_342);
or U4907 (N_4907,N_644,N_1304);
nand U4908 (N_4908,N_1344,N_357);
xnor U4909 (N_4909,N_129,N_1574);
xnor U4910 (N_4910,N_1002,N_1161);
nand U4911 (N_4911,N_2426,N_1069);
nand U4912 (N_4912,N_1964,N_447);
xnor U4913 (N_4913,N_20,N_1801);
and U4914 (N_4914,N_538,N_2286);
xor U4915 (N_4915,N_1675,N_2358);
nor U4916 (N_4916,N_434,N_7);
nand U4917 (N_4917,N_249,N_1312);
and U4918 (N_4918,N_2325,N_539);
xnor U4919 (N_4919,N_1523,N_1023);
nand U4920 (N_4920,N_444,N_1333);
and U4921 (N_4921,N_596,N_2441);
and U4922 (N_4922,N_272,N_2260);
nor U4923 (N_4923,N_307,N_25);
and U4924 (N_4924,N_2248,N_393);
nand U4925 (N_4925,N_986,N_448);
xor U4926 (N_4926,N_1037,N_104);
xnor U4927 (N_4927,N_132,N_1634);
xor U4928 (N_4928,N_2192,N_1085);
nor U4929 (N_4929,N_1578,N_1418);
nand U4930 (N_4930,N_1619,N_2331);
nand U4931 (N_4931,N_1152,N_2020);
nor U4932 (N_4932,N_254,N_1844);
or U4933 (N_4933,N_1939,N_1423);
or U4934 (N_4934,N_1389,N_2361);
nand U4935 (N_4935,N_281,N_2006);
xnor U4936 (N_4936,N_1442,N_924);
and U4937 (N_4937,N_1163,N_1673);
and U4938 (N_4938,N_1735,N_1872);
nor U4939 (N_4939,N_544,N_518);
nor U4940 (N_4940,N_367,N_124);
and U4941 (N_4941,N_250,N_792);
or U4942 (N_4942,N_964,N_1383);
or U4943 (N_4943,N_786,N_1397);
nor U4944 (N_4944,N_70,N_1733);
nand U4945 (N_4945,N_1389,N_621);
nor U4946 (N_4946,N_1674,N_1681);
and U4947 (N_4947,N_2023,N_513);
nor U4948 (N_4948,N_337,N_905);
nand U4949 (N_4949,N_463,N_1141);
nor U4950 (N_4950,N_1403,N_330);
xor U4951 (N_4951,N_1093,N_1012);
and U4952 (N_4952,N_173,N_1996);
nor U4953 (N_4953,N_1180,N_1316);
xnor U4954 (N_4954,N_354,N_343);
nor U4955 (N_4955,N_1672,N_1708);
or U4956 (N_4956,N_546,N_960);
or U4957 (N_4957,N_1097,N_104);
or U4958 (N_4958,N_2088,N_1795);
nand U4959 (N_4959,N_2411,N_2331);
nand U4960 (N_4960,N_1539,N_2148);
and U4961 (N_4961,N_846,N_2203);
xnor U4962 (N_4962,N_329,N_1979);
and U4963 (N_4963,N_56,N_379);
nor U4964 (N_4964,N_1690,N_2440);
and U4965 (N_4965,N_216,N_2473);
nand U4966 (N_4966,N_695,N_2349);
or U4967 (N_4967,N_2481,N_407);
nand U4968 (N_4968,N_641,N_404);
or U4969 (N_4969,N_272,N_405);
xnor U4970 (N_4970,N_596,N_2285);
xor U4971 (N_4971,N_1974,N_852);
nor U4972 (N_4972,N_1048,N_423);
nor U4973 (N_4973,N_624,N_2269);
nand U4974 (N_4974,N_2488,N_737);
or U4975 (N_4975,N_2267,N_1788);
or U4976 (N_4976,N_725,N_1010);
nor U4977 (N_4977,N_961,N_1584);
xor U4978 (N_4978,N_721,N_829);
xor U4979 (N_4979,N_535,N_1428);
or U4980 (N_4980,N_1967,N_1684);
nor U4981 (N_4981,N_1580,N_2334);
and U4982 (N_4982,N_1463,N_612);
nand U4983 (N_4983,N_2253,N_2379);
or U4984 (N_4984,N_876,N_1021);
or U4985 (N_4985,N_682,N_1724);
xnor U4986 (N_4986,N_845,N_449);
nand U4987 (N_4987,N_884,N_1703);
and U4988 (N_4988,N_490,N_705);
nand U4989 (N_4989,N_395,N_2018);
nand U4990 (N_4990,N_2294,N_896);
and U4991 (N_4991,N_1399,N_1774);
nand U4992 (N_4992,N_638,N_128);
or U4993 (N_4993,N_1861,N_1924);
or U4994 (N_4994,N_1771,N_2145);
xnor U4995 (N_4995,N_2390,N_1654);
xor U4996 (N_4996,N_1462,N_2042);
nand U4997 (N_4997,N_2498,N_2227);
nor U4998 (N_4998,N_2263,N_2437);
or U4999 (N_4999,N_213,N_1600);
or U5000 (N_5000,N_4671,N_3938);
nor U5001 (N_5001,N_4179,N_3551);
and U5002 (N_5002,N_4077,N_3971);
and U5003 (N_5003,N_3552,N_3654);
and U5004 (N_5004,N_4468,N_4119);
nand U5005 (N_5005,N_4215,N_4349);
xor U5006 (N_5006,N_2999,N_3055);
and U5007 (N_5007,N_2655,N_3534);
nor U5008 (N_5008,N_2679,N_4780);
and U5009 (N_5009,N_4266,N_2928);
nand U5010 (N_5010,N_3924,N_2678);
nand U5011 (N_5011,N_3983,N_4348);
or U5012 (N_5012,N_3127,N_3724);
nor U5013 (N_5013,N_3350,N_4894);
and U5014 (N_5014,N_2686,N_3302);
nand U5015 (N_5015,N_4370,N_3521);
and U5016 (N_5016,N_2971,N_2908);
and U5017 (N_5017,N_4842,N_4421);
and U5018 (N_5018,N_4974,N_3524);
or U5019 (N_5019,N_4098,N_4422);
xor U5020 (N_5020,N_3992,N_2652);
and U5021 (N_5021,N_2550,N_4448);
nor U5022 (N_5022,N_3575,N_2761);
xor U5023 (N_5023,N_3297,N_3159);
xnor U5024 (N_5024,N_2977,N_4471);
nor U5025 (N_5025,N_4071,N_2855);
nor U5026 (N_5026,N_3199,N_4067);
or U5027 (N_5027,N_3123,N_4717);
nor U5028 (N_5028,N_4845,N_3639);
or U5029 (N_5029,N_2870,N_4714);
and U5030 (N_5030,N_4482,N_4764);
or U5031 (N_5031,N_4672,N_2903);
nand U5032 (N_5032,N_3970,N_4645);
or U5033 (N_5033,N_2738,N_2718);
or U5034 (N_5034,N_3816,N_4824);
and U5035 (N_5035,N_3641,N_2551);
nor U5036 (N_5036,N_2713,N_2683);
nand U5037 (N_5037,N_4698,N_4877);
and U5038 (N_5038,N_3894,N_4347);
nand U5039 (N_5039,N_2911,N_2882);
and U5040 (N_5040,N_2914,N_4641);
nor U5041 (N_5041,N_3996,N_3382);
or U5042 (N_5042,N_3266,N_4725);
or U5043 (N_5043,N_4913,N_3761);
and U5044 (N_5044,N_2974,N_4419);
xnor U5045 (N_5045,N_4802,N_4866);
xor U5046 (N_5046,N_4222,N_4752);
nand U5047 (N_5047,N_4689,N_4073);
xnor U5048 (N_5048,N_3206,N_4582);
xor U5049 (N_5049,N_3963,N_4490);
and U5050 (N_5050,N_3864,N_4408);
xor U5051 (N_5051,N_3481,N_3166);
or U5052 (N_5052,N_4008,N_3325);
and U5053 (N_5053,N_3445,N_3193);
xor U5054 (N_5054,N_4327,N_4898);
and U5055 (N_5055,N_4909,N_2622);
nor U5056 (N_5056,N_4839,N_2544);
nand U5057 (N_5057,N_2778,N_3932);
and U5058 (N_5058,N_4878,N_4001);
nor U5059 (N_5059,N_4973,N_4616);
nand U5060 (N_5060,N_3847,N_4190);
nor U5061 (N_5061,N_3071,N_2852);
or U5062 (N_5062,N_3453,N_4893);
or U5063 (N_5063,N_4628,N_4412);
or U5064 (N_5064,N_3516,N_4465);
nor U5065 (N_5065,N_3665,N_3929);
nor U5066 (N_5066,N_3042,N_2824);
nand U5067 (N_5067,N_4226,N_3743);
xnor U5068 (N_5068,N_3561,N_4522);
or U5069 (N_5069,N_4346,N_2577);
nor U5070 (N_5070,N_3897,N_4210);
and U5071 (N_5071,N_2917,N_3044);
nor U5072 (N_5072,N_4636,N_3340);
nor U5073 (N_5073,N_3269,N_3474);
or U5074 (N_5074,N_4384,N_3510);
xor U5075 (N_5075,N_3160,N_2641);
or U5076 (N_5076,N_4143,N_2990);
nand U5077 (N_5077,N_3492,N_4053);
and U5078 (N_5078,N_2647,N_4472);
xor U5079 (N_5079,N_4564,N_4508);
xnor U5080 (N_5080,N_3859,N_3263);
xor U5081 (N_5081,N_4286,N_3987);
and U5082 (N_5082,N_4665,N_3498);
and U5083 (N_5083,N_2827,N_2814);
nor U5084 (N_5084,N_4826,N_3262);
nor U5085 (N_5085,N_3241,N_3362);
or U5086 (N_5086,N_4278,N_2602);
nand U5087 (N_5087,N_4738,N_3046);
xnor U5088 (N_5088,N_2515,N_4682);
and U5089 (N_5089,N_2560,N_2630);
and U5090 (N_5090,N_3951,N_3935);
nor U5091 (N_5091,N_4528,N_4583);
or U5092 (N_5092,N_4830,N_4762);
nand U5093 (N_5093,N_3130,N_4763);
or U5094 (N_5094,N_4829,N_2751);
or U5095 (N_5095,N_3410,N_2811);
xnor U5096 (N_5096,N_2984,N_4542);
xor U5097 (N_5097,N_3997,N_3860);
nand U5098 (N_5098,N_3776,N_2846);
nor U5099 (N_5099,N_4673,N_4133);
and U5100 (N_5100,N_2813,N_2989);
xnor U5101 (N_5101,N_3694,N_3161);
nor U5102 (N_5102,N_3947,N_4706);
nor U5103 (N_5103,N_2708,N_2644);
xor U5104 (N_5104,N_3244,N_4275);
and U5105 (N_5105,N_3975,N_4051);
nor U5106 (N_5106,N_3030,N_3092);
nor U5107 (N_5107,N_3794,N_4825);
nand U5108 (N_5108,N_2609,N_2775);
nand U5109 (N_5109,N_3614,N_4467);
nor U5110 (N_5110,N_3178,N_4678);
nor U5111 (N_5111,N_4569,N_3733);
xnor U5112 (N_5112,N_4962,N_3381);
nor U5113 (N_5113,N_2754,N_3739);
nand U5114 (N_5114,N_2972,N_4655);
xnor U5115 (N_5115,N_4117,N_2621);
and U5116 (N_5116,N_4024,N_3687);
xor U5117 (N_5117,N_4799,N_4724);
nor U5118 (N_5118,N_3462,N_3829);
and U5119 (N_5119,N_3376,N_4161);
or U5120 (N_5120,N_3497,N_4021);
nor U5121 (N_5121,N_2753,N_4108);
xnor U5122 (N_5122,N_3818,N_2782);
or U5123 (N_5123,N_4201,N_3259);
and U5124 (N_5124,N_3905,N_3682);
nor U5125 (N_5125,N_4341,N_3307);
xnor U5126 (N_5126,N_2823,N_4708);
and U5127 (N_5127,N_3783,N_2514);
nor U5128 (N_5128,N_4933,N_3710);
nor U5129 (N_5129,N_2502,N_4459);
xor U5130 (N_5130,N_4722,N_2563);
or U5131 (N_5131,N_3502,N_2532);
xnor U5132 (N_5132,N_3260,N_3597);
nor U5133 (N_5133,N_4075,N_3045);
or U5134 (N_5134,N_3930,N_3334);
nor U5135 (N_5135,N_4262,N_4385);
nand U5136 (N_5136,N_2759,N_4103);
xnor U5137 (N_5137,N_3479,N_4506);
xor U5138 (N_5138,N_3770,N_4633);
nand U5139 (N_5139,N_3836,N_2840);
nand U5140 (N_5140,N_3383,N_4157);
or U5141 (N_5141,N_3642,N_3038);
or U5142 (N_5142,N_3448,N_4047);
xnor U5143 (N_5143,N_3495,N_4943);
and U5144 (N_5144,N_4081,N_3240);
nor U5145 (N_5145,N_4382,N_4978);
xor U5146 (N_5146,N_2832,N_4129);
nand U5147 (N_5147,N_4959,N_3143);
and U5148 (N_5148,N_3117,N_4018);
nand U5149 (N_5149,N_2777,N_3844);
and U5150 (N_5150,N_3728,N_4922);
and U5151 (N_5151,N_3039,N_2867);
and U5152 (N_5152,N_4595,N_4835);
and U5153 (N_5153,N_4777,N_3664);
xor U5154 (N_5154,N_4063,N_2534);
or U5155 (N_5155,N_3558,N_2715);
and U5156 (N_5156,N_3730,N_2547);
xor U5157 (N_5157,N_2921,N_2851);
xor U5158 (N_5158,N_4547,N_3564);
or U5159 (N_5159,N_4545,N_3407);
nand U5160 (N_5160,N_4934,N_3031);
or U5161 (N_5161,N_4365,N_2915);
nand U5162 (N_5162,N_3631,N_2739);
nor U5163 (N_5163,N_4086,N_3295);
or U5164 (N_5164,N_3406,N_4424);
xor U5165 (N_5165,N_3156,N_4167);
nand U5166 (N_5166,N_3218,N_3751);
nand U5167 (N_5167,N_3141,N_4277);
xor U5168 (N_5168,N_4991,N_2746);
xor U5169 (N_5169,N_4152,N_3572);
nor U5170 (N_5170,N_3686,N_3985);
nand U5171 (N_5171,N_3966,N_4876);
or U5172 (N_5172,N_4045,N_2604);
xor U5173 (N_5173,N_3484,N_3248);
and U5174 (N_5174,N_3135,N_3283);
xor U5175 (N_5175,N_4390,N_2830);
and U5176 (N_5176,N_4240,N_3726);
nor U5177 (N_5177,N_3979,N_3679);
and U5178 (N_5178,N_4709,N_3287);
or U5179 (N_5179,N_4526,N_3895);
xor U5180 (N_5180,N_3440,N_2537);
and U5181 (N_5181,N_4158,N_4435);
xnor U5182 (N_5182,N_3223,N_2626);
nor U5183 (N_5183,N_3347,N_3986);
xor U5184 (N_5184,N_2880,N_3934);
nor U5185 (N_5185,N_2815,N_3197);
nor U5186 (N_5186,N_4247,N_4366);
and U5187 (N_5187,N_3204,N_3111);
or U5188 (N_5188,N_3949,N_3870);
and U5189 (N_5189,N_4515,N_3662);
xor U5190 (N_5190,N_3667,N_2618);
nand U5191 (N_5191,N_4817,N_4410);
nand U5192 (N_5192,N_4165,N_3742);
xor U5193 (N_5193,N_3719,N_3183);
nand U5194 (N_5194,N_3936,N_4891);
and U5195 (N_5195,N_2520,N_4359);
xnor U5196 (N_5196,N_4666,N_4514);
nand U5197 (N_5197,N_2765,N_4213);
and U5198 (N_5198,N_2853,N_4242);
nand U5199 (N_5199,N_3465,N_3789);
and U5200 (N_5200,N_3621,N_3471);
or U5201 (N_5201,N_2740,N_3115);
and U5202 (N_5202,N_3539,N_3946);
or U5203 (N_5203,N_2669,N_4554);
nand U5204 (N_5204,N_4504,N_3529);
or U5205 (N_5205,N_2800,N_3467);
xnor U5206 (N_5206,N_3065,N_3624);
xor U5207 (N_5207,N_2504,N_3514);
or U5208 (N_5208,N_4439,N_4844);
or U5209 (N_5209,N_4355,N_4259);
nor U5210 (N_5210,N_3557,N_4010);
or U5211 (N_5211,N_4818,N_2579);
and U5212 (N_5212,N_3457,N_2877);
and U5213 (N_5213,N_3010,N_3923);
and U5214 (N_5214,N_4123,N_2654);
xor U5215 (N_5215,N_3250,N_3403);
and U5216 (N_5216,N_3139,N_2965);
nand U5217 (N_5217,N_3819,N_4224);
or U5218 (N_5218,N_2845,N_2897);
or U5219 (N_5219,N_3875,N_4172);
and U5220 (N_5220,N_4718,N_3268);
xor U5221 (N_5221,N_2817,N_2511);
or U5222 (N_5222,N_4897,N_4074);
nor U5223 (N_5223,N_3508,N_4606);
xnor U5224 (N_5224,N_2894,N_4142);
nor U5225 (N_5225,N_2764,N_3734);
nor U5226 (N_5226,N_3960,N_3443);
nand U5227 (N_5227,N_4649,N_3310);
xor U5228 (N_5228,N_4085,N_4772);
nor U5229 (N_5229,N_3242,N_4761);
or U5230 (N_5230,N_4062,N_4460);
nand U5231 (N_5231,N_4720,N_4100);
or U5232 (N_5232,N_4507,N_4579);
nand U5233 (N_5233,N_2844,N_2926);
nor U5234 (N_5234,N_4338,N_2970);
nand U5235 (N_5235,N_4039,N_3215);
xor U5236 (N_5236,N_4250,N_4106);
or U5237 (N_5237,N_2714,N_2909);
xnor U5238 (N_5238,N_3649,N_3792);
nor U5239 (N_5239,N_2549,N_3331);
xor U5240 (N_5240,N_4314,N_4336);
and U5241 (N_5241,N_3808,N_3332);
xnor U5242 (N_5242,N_4397,N_2501);
and U5243 (N_5243,N_2527,N_3814);
xor U5244 (N_5244,N_3736,N_3413);
and U5245 (N_5245,N_4193,N_4900);
nor U5246 (N_5246,N_2500,N_4216);
nor U5247 (N_5247,N_2969,N_4396);
nor U5248 (N_5248,N_3470,N_4011);
or U5249 (N_5249,N_4393,N_3893);
and U5250 (N_5250,N_4581,N_3834);
xnor U5251 (N_5251,N_4322,N_3221);
nand U5252 (N_5252,N_3790,N_4874);
nor U5253 (N_5253,N_2806,N_3757);
nand U5254 (N_5254,N_4319,N_4170);
or U5255 (N_5255,N_3314,N_3780);
or U5256 (N_5256,N_3764,N_4773);
or U5257 (N_5257,N_4065,N_2694);
xor U5258 (N_5258,N_3353,N_3607);
nor U5259 (N_5259,N_3021,N_3696);
nor U5260 (N_5260,N_2848,N_3933);
nand U5261 (N_5261,N_4070,N_4832);
xor U5262 (N_5262,N_3116,N_3638);
or U5263 (N_5263,N_2519,N_4475);
nand U5264 (N_5264,N_4050,N_3344);
nand U5265 (N_5265,N_2774,N_3646);
xor U5266 (N_5266,N_3758,N_3090);
nor U5267 (N_5267,N_3276,N_2783);
nand U5268 (N_5268,N_4776,N_3286);
nor U5269 (N_5269,N_4494,N_4759);
and U5270 (N_5270,N_4749,N_2750);
and U5271 (N_5271,N_4809,N_2810);
and U5272 (N_5272,N_4441,N_4036);
nand U5273 (N_5273,N_4668,N_3771);
nand U5274 (N_5274,N_3858,N_3831);
nand U5275 (N_5275,N_3252,N_3584);
nor U5276 (N_5276,N_3014,N_4623);
or U5277 (N_5277,N_3677,N_4187);
nand U5278 (N_5278,N_4169,N_3202);
nand U5279 (N_5279,N_3336,N_4942);
nor U5280 (N_5280,N_2963,N_3772);
nand U5281 (N_5281,N_4200,N_3527);
nor U5282 (N_5282,N_2996,N_4937);
xor U5283 (N_5283,N_2961,N_3873);
nand U5284 (N_5284,N_3404,N_3553);
nor U5285 (N_5285,N_2864,N_4034);
nor U5286 (N_5286,N_4091,N_3239);
and U5287 (N_5287,N_4303,N_2756);
and U5288 (N_5288,N_2930,N_4916);
xor U5289 (N_5289,N_3033,N_4171);
or U5290 (N_5290,N_4307,N_2820);
xor U5291 (N_5291,N_4518,N_4675);
nor U5292 (N_5292,N_3081,N_4821);
or U5293 (N_5293,N_3267,N_4713);
xnor U5294 (N_5294,N_3684,N_4395);
and U5295 (N_5295,N_3569,N_3568);
and U5296 (N_5296,N_2637,N_4093);
xnor U5297 (N_5297,N_3676,N_4992);
nor U5298 (N_5298,N_4434,N_3454);
xnor U5299 (N_5299,N_4095,N_2865);
nor U5300 (N_5300,N_4028,N_4363);
xor U5301 (N_5301,N_3522,N_2653);
nand U5302 (N_5302,N_4596,N_3586);
and U5303 (N_5303,N_4862,N_4638);
and U5304 (N_5304,N_2603,N_2842);
nand U5305 (N_5305,N_2868,N_2874);
and U5306 (N_5306,N_4220,N_2508);
and U5307 (N_5307,N_2606,N_3800);
and U5308 (N_5308,N_4492,N_3181);
nand U5309 (N_5309,N_4931,N_3591);
nor U5310 (N_5310,N_2925,N_4455);
and U5311 (N_5311,N_3530,N_3578);
xnor U5312 (N_5312,N_4651,N_2610);
and U5313 (N_5313,N_3673,N_4715);
nor U5314 (N_5314,N_2662,N_3709);
or U5315 (N_5315,N_2731,N_4911);
or U5316 (N_5316,N_4237,N_3812);
and U5317 (N_5317,N_2856,N_3309);
nor U5318 (N_5318,N_3965,N_3211);
xnor U5319 (N_5319,N_4430,N_3926);
xnor U5320 (N_5320,N_3412,N_2766);
nand U5321 (N_5321,N_4013,N_4228);
or U5322 (N_5322,N_4425,N_4159);
nand U5323 (N_5323,N_3000,N_4733);
nor U5324 (N_5324,N_3356,N_4400);
or U5325 (N_5325,N_2573,N_4107);
nand U5326 (N_5326,N_4532,N_3098);
nand U5327 (N_5327,N_4120,N_3617);
nor U5328 (N_5328,N_4640,N_2732);
xnor U5329 (N_5329,N_3388,N_3265);
or U5330 (N_5330,N_2985,N_3200);
or U5331 (N_5331,N_3653,N_4041);
and U5332 (N_5332,N_3571,N_4880);
nor U5333 (N_5333,N_4551,N_3366);
and U5334 (N_5334,N_4695,N_4189);
and U5335 (N_5335,N_4527,N_2676);
nand U5336 (N_5336,N_2734,N_3994);
nor U5337 (N_5337,N_2829,N_2681);
nor U5338 (N_5338,N_3918,N_3898);
nand U5339 (N_5339,N_4500,N_3121);
nor U5340 (N_5340,N_3999,N_4561);
nor U5341 (N_5341,N_3175,N_3149);
or U5342 (N_5342,N_4352,N_2617);
or U5343 (N_5343,N_4767,N_3627);
nor U5344 (N_5344,N_3881,N_3040);
and U5345 (N_5345,N_3243,N_4578);
nand U5346 (N_5346,N_3168,N_2854);
xor U5347 (N_5347,N_4339,N_4854);
and U5348 (N_5348,N_3026,N_3271);
xnor U5349 (N_5349,N_3424,N_3886);
nor U5350 (N_5350,N_2900,N_3230);
nand U5351 (N_5351,N_3773,N_2650);
nor U5352 (N_5352,N_4573,N_2831);
or U5353 (N_5353,N_3133,N_4163);
xnor U5354 (N_5354,N_3070,N_4949);
and U5355 (N_5355,N_2539,N_3393);
nand U5356 (N_5356,N_4615,N_3763);
xor U5357 (N_5357,N_3962,N_3798);
nand U5358 (N_5358,N_3174,N_4534);
or U5359 (N_5359,N_4519,N_2729);
nor U5360 (N_5360,N_4644,N_4234);
xor U5361 (N_5361,N_4334,N_4729);
nor U5362 (N_5362,N_4917,N_4361);
or U5363 (N_5363,N_3955,N_4588);
xor U5364 (N_5364,N_4146,N_4731);
nand U5365 (N_5365,N_3085,N_3803);
xnor U5366 (N_5366,N_3096,N_4840);
nor U5367 (N_5367,N_3351,N_3861);
or U5368 (N_5368,N_3172,N_4323);
xor U5369 (N_5369,N_4919,N_2956);
xnor U5370 (N_5370,N_4930,N_3632);
and U5371 (N_5371,N_3787,N_2932);
and U5372 (N_5372,N_3348,N_2656);
nor U5373 (N_5373,N_2742,N_3207);
and U5374 (N_5374,N_3043,N_2841);
xnor U5375 (N_5375,N_4403,N_2546);
nand U5376 (N_5376,N_3146,N_2808);
or U5377 (N_5377,N_3004,N_4076);
nand U5378 (N_5378,N_2727,N_3464);
or U5379 (N_5379,N_3235,N_4377);
nor U5380 (N_5380,N_4751,N_3488);
or U5381 (N_5381,N_4687,N_4971);
xnor U5382 (N_5382,N_2940,N_2803);
nor U5383 (N_5383,N_3746,N_4178);
nor U5384 (N_5384,N_3520,N_3176);
xnor U5385 (N_5385,N_3459,N_3852);
nand U5386 (N_5386,N_3827,N_3120);
xor U5387 (N_5387,N_4997,N_3279);
xnor U5388 (N_5388,N_3815,N_4203);
nor U5389 (N_5389,N_4865,N_2838);
xor U5390 (N_5390,N_3073,N_4639);
nand U5391 (N_5391,N_4122,N_3748);
and U5392 (N_5392,N_3328,N_2712);
or U5393 (N_5393,N_3018,N_3483);
nand U5394 (N_5394,N_3226,N_4806);
and U5395 (N_5395,N_2684,N_4868);
nor U5396 (N_5396,N_4479,N_2558);
nor U5397 (N_5397,N_2529,N_2860);
or U5398 (N_5398,N_3089,N_4654);
and U5399 (N_5399,N_3668,N_3846);
or U5400 (N_5400,N_3067,N_3112);
nand U5401 (N_5401,N_4061,N_2871);
nand U5402 (N_5402,N_3990,N_4032);
nand U5403 (N_5403,N_3107,N_4432);
nand U5404 (N_5404,N_2507,N_3035);
nor U5405 (N_5405,N_4022,N_3801);
and U5406 (N_5406,N_4501,N_3456);
nor U5407 (N_5407,N_4109,N_4691);
xnor U5408 (N_5408,N_3888,N_3194);
nor U5409 (N_5409,N_4092,N_4260);
or U5410 (N_5410,N_2625,N_4600);
and U5411 (N_5411,N_2862,N_4469);
xor U5412 (N_5412,N_3716,N_2667);
nor U5413 (N_5413,N_3854,N_3285);
nor U5414 (N_5414,N_4066,N_3830);
or U5415 (N_5415,N_3180,N_3084);
nor U5416 (N_5416,N_4052,N_3229);
and U5417 (N_5417,N_2705,N_4005);
or U5418 (N_5418,N_2665,N_3587);
xnor U5419 (N_5419,N_3173,N_4374);
xnor U5420 (N_5420,N_3610,N_2793);
or U5421 (N_5421,N_3187,N_3647);
nand U5422 (N_5422,N_3705,N_3455);
xnor U5423 (N_5423,N_3838,N_4498);
nor U5424 (N_5424,N_3486,N_4779);
nor U5425 (N_5425,N_4139,N_3750);
or U5426 (N_5426,N_4975,N_4181);
nor U5427 (N_5427,N_4711,N_2593);
nor U5428 (N_5428,N_4730,N_4483);
or U5429 (N_5429,N_2918,N_2680);
or U5430 (N_5430,N_4433,N_3738);
nor U5431 (N_5431,N_4755,N_3841);
and U5432 (N_5432,N_3273,N_3912);
and U5433 (N_5433,N_4788,N_4196);
xor U5434 (N_5434,N_2943,N_4279);
xor U5435 (N_5435,N_3950,N_4966);
xnor U5436 (N_5436,N_3540,N_2847);
and U5437 (N_5437,N_3320,N_3969);
xnor U5438 (N_5438,N_2920,N_4935);
nand U5439 (N_5439,N_2968,N_2649);
or U5440 (N_5440,N_4285,N_4114);
or U5441 (N_5441,N_4531,N_4183);
xnor U5442 (N_5442,N_3517,N_2540);
or U5443 (N_5443,N_4175,N_4619);
and U5444 (N_5444,N_3767,N_3024);
xnor U5445 (N_5445,N_4177,N_3601);
or U5446 (N_5446,N_3220,N_4552);
and U5447 (N_5447,N_3378,N_3012);
and U5448 (N_5448,N_4814,N_4924);
nand U5449 (N_5449,N_3482,N_3835);
nor U5450 (N_5450,N_3109,N_4128);
nand U5451 (N_5451,N_2993,N_3967);
nor U5452 (N_5452,N_3419,N_2752);
and U5453 (N_5453,N_3064,N_2976);
or U5454 (N_5454,N_4176,N_3784);
xnor U5455 (N_5455,N_4389,N_3057);
nor U5456 (N_5456,N_2671,N_2675);
xor U5457 (N_5457,N_4727,N_2640);
nor U5458 (N_5458,N_4321,N_2666);
and U5459 (N_5459,N_3909,N_3102);
nor U5460 (N_5460,N_3439,N_3397);
and U5461 (N_5461,N_3125,N_3721);
nand U5462 (N_5462,N_3543,N_4921);
xnor U5463 (N_5463,N_3634,N_3427);
nor U5464 (N_5464,N_4820,N_3217);
or U5465 (N_5465,N_3535,N_3349);
and U5466 (N_5466,N_4693,N_3670);
xor U5467 (N_5467,N_3164,N_2895);
nand U5468 (N_5468,N_4885,N_4446);
or U5469 (N_5469,N_4059,N_4778);
and U5470 (N_5470,N_3028,N_3681);
and U5471 (N_5471,N_2624,N_4020);
nand U5472 (N_5472,N_3525,N_4782);
nor U5473 (N_5473,N_2594,N_3755);
xor U5474 (N_5474,N_3203,N_3429);
xor U5475 (N_5475,N_3177,N_2589);
nand U5476 (N_5476,N_4127,N_4357);
and U5477 (N_5477,N_3872,N_3612);
nand U5478 (N_5478,N_2564,N_4317);
and U5479 (N_5479,N_3972,N_3329);
or U5480 (N_5480,N_4604,N_3536);
nand U5481 (N_5481,N_3671,N_4245);
xor U5482 (N_5482,N_2986,N_2693);
nand U5483 (N_5483,N_4512,N_2747);
and U5484 (N_5484,N_3956,N_4948);
xor U5485 (N_5485,N_3251,N_4529);
or U5486 (N_5486,N_3478,N_2706);
or U5487 (N_5487,N_3565,N_2720);
and U5488 (N_5488,N_4470,N_4340);
nand U5489 (N_5489,N_2931,N_3678);
xnor U5490 (N_5490,N_4701,N_4147);
xor U5491 (N_5491,N_3526,N_4669);
xor U5492 (N_5492,N_4822,N_4947);
nand U5493 (N_5493,N_4753,N_2799);
and U5494 (N_5494,N_3560,N_4792);
or U5495 (N_5495,N_2872,N_4986);
nand U5496 (N_5496,N_3450,N_4505);
nor U5497 (N_5497,N_3943,N_3228);
nand U5498 (N_5498,N_4575,N_3782);
and U5499 (N_5499,N_4783,N_4420);
nor U5500 (N_5500,N_3423,N_3840);
xor U5501 (N_5501,N_3785,N_3500);
nand U5502 (N_5502,N_4372,N_2634);
nor U5503 (N_5503,N_4741,N_3294);
and U5504 (N_5504,N_3910,N_4662);
and U5505 (N_5505,N_3321,N_4622);
nor U5506 (N_5506,N_4864,N_3629);
and U5507 (N_5507,N_4496,N_4392);
or U5508 (N_5508,N_3054,N_3915);
xnor U5509 (N_5509,N_2949,N_4710);
and U5510 (N_5510,N_3982,N_4153);
nor U5511 (N_5511,N_4236,N_4509);
xnor U5512 (N_5512,N_4756,N_4437);
nand U5513 (N_5513,N_3008,N_2839);
nand U5514 (N_5514,N_4684,N_4790);
or U5515 (N_5515,N_3145,N_3891);
and U5516 (N_5516,N_3184,N_3078);
nand U5517 (N_5517,N_3559,N_3280);
xor U5518 (N_5518,N_4069,N_3637);
or U5519 (N_5519,N_4476,N_3618);
nand U5520 (N_5520,N_2651,N_3887);
or U5521 (N_5521,N_3702,N_4110);
or U5522 (N_5522,N_3034,N_2924);
xnor U5523 (N_5523,N_4617,N_2888);
xnor U5524 (N_5524,N_4373,N_3741);
and U5525 (N_5525,N_4431,N_3952);
and U5526 (N_5526,N_2645,N_3606);
nor U5527 (N_5527,N_4436,N_2568);
xor U5528 (N_5528,N_2889,N_4386);
nand U5529 (N_5529,N_3623,N_2768);
or U5530 (N_5530,N_4810,N_3976);
or U5531 (N_5531,N_3515,N_2691);
nand U5532 (N_5532,N_3416,N_3425);
nor U5533 (N_5533,N_3518,N_4136);
nor U5534 (N_5534,N_3580,N_4489);
nor U5535 (N_5535,N_2905,N_3715);
nand U5536 (N_5536,N_3871,N_4699);
nor U5537 (N_5537,N_4837,N_4984);
xnor U5538 (N_5538,N_2522,N_4316);
and U5539 (N_5539,N_2512,N_2724);
or U5540 (N_5540,N_3779,N_4484);
nand U5541 (N_5541,N_3826,N_4309);
nor U5542 (N_5542,N_3219,N_4368);
nor U5543 (N_5543,N_3369,N_4611);
nand U5544 (N_5544,N_3494,N_4670);
nor U5545 (N_5545,N_3167,N_4589);
nor U5546 (N_5546,N_3548,N_4298);
or U5547 (N_5547,N_4194,N_4463);
nand U5548 (N_5548,N_3025,N_4680);
and U5549 (N_5549,N_4543,N_4769);
or U5550 (N_5550,N_3688,N_3542);
nand U5551 (N_5551,N_4584,N_3442);
nand U5552 (N_5552,N_4084,N_4950);
nor U5553 (N_5553,N_4743,N_4331);
nor U5554 (N_5554,N_4442,N_3661);
xnor U5555 (N_5555,N_3729,N_4218);
or U5556 (N_5556,N_3371,N_4694);
nand U5557 (N_5557,N_3506,N_4225);
nor U5558 (N_5558,N_2946,N_2887);
nor U5559 (N_5559,N_4517,N_3433);
xor U5560 (N_5560,N_3188,N_3644);
and U5561 (N_5561,N_4185,N_3129);
and U5562 (N_5562,N_4533,N_3628);
nor U5563 (N_5563,N_3460,N_4360);
nor U5564 (N_5564,N_4000,N_2773);
xor U5565 (N_5565,N_4775,N_3061);
nand U5566 (N_5566,N_4168,N_4125);
or U5567 (N_5567,N_3942,N_3237);
and U5568 (N_5568,N_3978,N_4118);
or U5569 (N_5569,N_4102,N_2701);
xor U5570 (N_5570,N_3435,N_4987);
nand U5571 (N_5571,N_4345,N_3546);
and U5572 (N_5572,N_3977,N_2586);
nand U5573 (N_5573,N_3155,N_4294);
nand U5574 (N_5574,N_4728,N_2794);
nor U5575 (N_5575,N_3680,N_4318);
nor U5576 (N_5576,N_3179,N_4754);
and U5577 (N_5577,N_3856,N_4054);
and U5578 (N_5578,N_4803,N_3375);
or U5579 (N_5579,N_3940,N_4953);
nor U5580 (N_5580,N_4493,N_3813);
nor U5581 (N_5581,N_3544,N_4907);
nor U5582 (N_5582,N_2552,N_4811);
or U5583 (N_5583,N_4173,N_2843);
and U5584 (N_5584,N_2615,N_3727);
or U5585 (N_5585,N_3170,N_3233);
or U5586 (N_5586,N_3805,N_4870);
xnor U5587 (N_5587,N_4030,N_4511);
xnor U5588 (N_5588,N_4571,N_4099);
nand U5589 (N_5589,N_3695,N_4557);
nor U5590 (N_5590,N_3549,N_3900);
nor U5591 (N_5591,N_3308,N_2696);
xor U5592 (N_5592,N_4550,N_4873);
xnor U5593 (N_5593,N_3594,N_2605);
and U5594 (N_5594,N_3762,N_4969);
and U5595 (N_5595,N_4486,N_4998);
xor U5596 (N_5596,N_4981,N_4304);
nand U5597 (N_5597,N_2950,N_3583);
nor U5598 (N_5598,N_4350,N_2967);
nor U5599 (N_5599,N_3324,N_4857);
xor U5600 (N_5600,N_3088,N_2802);
nand U5601 (N_5601,N_3158,N_4301);
nand U5602 (N_5602,N_4473,N_2728);
nand U5603 (N_5603,N_4414,N_3563);
xor U5604 (N_5604,N_4925,N_3863);
nor U5605 (N_5605,N_4238,N_3849);
xor U5606 (N_5606,N_3690,N_3556);
xor U5607 (N_5607,N_4217,N_3083);
nor U5608 (N_5608,N_4379,N_4305);
or U5609 (N_5609,N_4732,N_4332);
or U5610 (N_5610,N_3613,N_4166);
xnor U5611 (N_5611,N_2518,N_3513);
nand U5612 (N_5612,N_4620,N_3579);
nor U5613 (N_5613,N_4273,N_4330);
nor U5614 (N_5614,N_3795,N_3937);
nand U5615 (N_5615,N_3299,N_2503);
nor U5616 (N_5616,N_4449,N_3600);
or U5617 (N_5617,N_4333,N_4688);
and U5618 (N_5618,N_4383,N_3472);
xnor U5619 (N_5619,N_4652,N_4049);
nand U5620 (N_5620,N_3599,N_3981);
nand U5621 (N_5621,N_4827,N_4451);
and U5622 (N_5622,N_3504,N_4019);
nor U5623 (N_5623,N_4926,N_4229);
nor U5624 (N_5624,N_4660,N_2834);
or U5625 (N_5625,N_2592,N_3432);
nand U5626 (N_5626,N_4965,N_4406);
xnor U5627 (N_5627,N_3925,N_2721);
nand U5628 (N_5628,N_3275,N_3041);
nor U5629 (N_5629,N_3907,N_3436);
nor U5630 (N_5630,N_3756,N_4735);
nor U5631 (N_5631,N_4686,N_4407);
xor U5632 (N_5632,N_4849,N_3775);
and U5633 (N_5633,N_4056,N_4094);
and U5634 (N_5634,N_3809,N_4155);
nand U5635 (N_5635,N_4391,N_3948);
xor U5636 (N_5636,N_3020,N_3855);
nand U5637 (N_5637,N_3444,N_2601);
and U5638 (N_5638,N_4548,N_4936);
or U5639 (N_5639,N_2524,N_4905);
nand U5640 (N_5640,N_3136,N_4656);
and U5641 (N_5641,N_4748,N_4592);
nor U5642 (N_5642,N_3050,N_3707);
or U5643 (N_5643,N_3315,N_3227);
and U5644 (N_5644,N_4629,N_2952);
nor U5645 (N_5645,N_2725,N_3657);
or U5646 (N_5646,N_4068,N_3811);
nor U5647 (N_5647,N_3698,N_3322);
and U5648 (N_5648,N_3185,N_3768);
nor U5649 (N_5649,N_4828,N_3573);
xnor U5650 (N_5650,N_3422,N_4466);
nor U5651 (N_5651,N_4683,N_3663);
and U5652 (N_5652,N_4140,N_2555);
xnor U5653 (N_5653,N_3303,N_3499);
and U5654 (N_5654,N_4739,N_3493);
xnor U5655 (N_5655,N_3988,N_4035);
and U5656 (N_5656,N_4618,N_3685);
and U5657 (N_5657,N_4042,N_3959);
or U5658 (N_5658,N_4450,N_4556);
nor U5659 (N_5659,N_2945,N_2805);
nand U5660 (N_5660,N_3674,N_3082);
nand U5661 (N_5661,N_3547,N_3391);
xor U5662 (N_5662,N_3699,N_2927);
or U5663 (N_5663,N_4244,N_2587);
or U5664 (N_5664,N_4007,N_4180);
nand U5665 (N_5665,N_3866,N_3630);
nor U5666 (N_5666,N_3512,N_4904);
xnor U5667 (N_5667,N_2906,N_2878);
and U5668 (N_5668,N_4690,N_3810);
nand U5669 (N_5669,N_2690,N_2663);
xor U5670 (N_5670,N_4055,N_2533);
nand U5671 (N_5671,N_3689,N_2792);
nand U5672 (N_5672,N_3399,N_4445);
nor U5673 (N_5673,N_3807,N_2982);
and U5674 (N_5674,N_4650,N_4663);
xnor U5675 (N_5675,N_4416,N_3658);
xnor U5676 (N_5676,N_2528,N_4838);
and U5677 (N_5677,N_3002,N_3080);
nor U5678 (N_5678,N_3032,N_4558);
and U5679 (N_5679,N_3592,N_2674);
nand U5680 (N_5680,N_2556,N_2901);
and U5681 (N_5681,N_2816,N_3765);
and U5682 (N_5682,N_3420,N_3379);
nor U5683 (N_5683,N_4296,N_4995);
xnor U5684 (N_5684,N_4025,N_4271);
and U5685 (N_5685,N_4458,N_3491);
xor U5686 (N_5686,N_4946,N_2571);
xor U5687 (N_5687,N_3920,N_3545);
and U5688 (N_5688,N_2513,N_4131);
and U5689 (N_5689,N_3305,N_4328);
nor U5690 (N_5690,N_4952,N_3718);
xnor U5691 (N_5691,N_3394,N_4315);
nand U5692 (N_5692,N_3051,N_3205);
xnor U5693 (N_5693,N_4132,N_3409);
xor U5694 (N_5694,N_4409,N_4223);
xnor U5695 (N_5695,N_3086,N_2910);
nor U5696 (N_5696,N_2912,N_4447);
nand U5697 (N_5697,N_3189,N_3714);
nor U5698 (N_5698,N_4404,N_4257);
and U5699 (N_5699,N_3449,N_2966);
and U5700 (N_5700,N_4539,N_4597);
nand U5701 (N_5701,N_4801,N_3851);
and U5702 (N_5702,N_4248,N_4677);
nor U5703 (N_5703,N_3507,N_3049);
nand U5704 (N_5704,N_4288,N_4808);
or U5705 (N_5705,N_4721,N_2936);
xor U5706 (N_5706,N_3131,N_4745);
xnor U5707 (N_5707,N_4858,N_4544);
and U5708 (N_5708,N_3842,N_3744);
nor U5709 (N_5709,N_2902,N_2955);
xor U5710 (N_5710,N_2958,N_4141);
and U5711 (N_5711,N_3056,N_2781);
and U5712 (N_5712,N_4302,N_4337);
and U5713 (N_5713,N_4121,N_4116);
or U5714 (N_5714,N_4502,N_3717);
nand U5715 (N_5715,N_3958,N_4836);
nor U5716 (N_5716,N_2757,N_4742);
nand U5717 (N_5717,N_4945,N_3796);
xor U5718 (N_5718,N_2578,N_4982);
nand U5719 (N_5719,N_2657,N_3069);
and U5720 (N_5720,N_2741,N_2723);
nand U5721 (N_5721,N_3659,N_4362);
nand U5722 (N_5722,N_4559,N_3941);
nor U5723 (N_5723,N_4488,N_2951);
xnor U5724 (N_5724,N_4567,N_2869);
or U5725 (N_5725,N_2896,N_3323);
or U5726 (N_5726,N_4535,N_2785);
nor U5727 (N_5727,N_2542,N_4903);
xor U5728 (N_5728,N_4381,N_2807);
xor U5729 (N_5729,N_3327,N_4867);
xnor U5730 (N_5730,N_3278,N_4212);
xor U5731 (N_5731,N_4308,N_3385);
and U5732 (N_5732,N_2698,N_4195);
and U5733 (N_5733,N_2835,N_3576);
and U5734 (N_5734,N_4233,N_4037);
xnor U5735 (N_5735,N_2557,N_2983);
or U5736 (N_5736,N_2904,N_3225);
nor U5737 (N_5737,N_3144,N_4048);
nand U5738 (N_5738,N_2692,N_2682);
xor U5739 (N_5739,N_3214,N_2659);
nor U5740 (N_5740,N_4291,N_2964);
nor U5741 (N_5741,N_3609,N_4205);
nand U5742 (N_5742,N_2953,N_4812);
and U5743 (N_5743,N_4371,N_4524);
nor U5744 (N_5744,N_3326,N_2948);
nand U5745 (N_5745,N_3911,N_3636);
xnor U5746 (N_5746,N_4823,N_4191);
xor U5747 (N_5747,N_4284,N_4329);
and U5748 (N_5748,N_4580,N_4601);
nand U5749 (N_5749,N_3426,N_3401);
or U5750 (N_5750,N_2709,N_4851);
and U5751 (N_5751,N_4719,N_4610);
nand U5752 (N_5752,N_3828,N_3066);
xnor U5753 (N_5753,N_4272,N_2763);
nand U5754 (N_5754,N_4955,N_2770);
xnor U5755 (N_5755,N_3400,N_3016);
nor U5756 (N_5756,N_3833,N_3616);
nor U5757 (N_5757,N_2506,N_3622);
and U5758 (N_5758,N_2614,N_4105);
xnor U5759 (N_5759,N_2837,N_3538);
and U5760 (N_5760,N_2767,N_3417);
nand U5761 (N_5761,N_4576,N_3137);
xor U5762 (N_5762,N_2939,N_3953);
nor U5763 (N_5763,N_2716,N_3079);
and U5764 (N_5764,N_3655,N_4676);
and U5765 (N_5765,N_3908,N_3405);
or U5766 (N_5766,N_3192,N_3945);
xnor U5767 (N_5767,N_3165,N_3341);
xor U5768 (N_5768,N_2702,N_3438);
nand U5769 (N_5769,N_4135,N_3660);
or U5770 (N_5770,N_4453,N_3015);
and U5771 (N_5771,N_4786,N_4860);
xor U5772 (N_5772,N_4781,N_4464);
or U5773 (N_5773,N_4164,N_3142);
xnor U5774 (N_5774,N_3365,N_3153);
and U5775 (N_5775,N_4014,N_2553);
nand U5776 (N_5776,N_2707,N_4791);
or U5777 (N_5777,N_3822,N_4251);
and U5778 (N_5778,N_2788,N_2929);
nand U5779 (N_5779,N_2881,N_2749);
nor U5780 (N_5780,N_2639,N_3496);
nand U5781 (N_5781,N_4929,N_2677);
and U5782 (N_5782,N_4555,N_4813);
xor U5783 (N_5783,N_3224,N_3603);
or U5784 (N_5784,N_3581,N_3892);
xnor U5785 (N_5785,N_3620,N_4367);
and U5786 (N_5786,N_3993,N_3296);
or U5787 (N_5787,N_4268,N_3566);
or U5788 (N_5788,N_2620,N_3461);
and U5789 (N_5789,N_4796,N_4017);
nand U5790 (N_5790,N_3901,N_4046);
nor U5791 (N_5791,N_3473,N_4148);
nor U5792 (N_5792,N_3532,N_2697);
or U5793 (N_5793,N_3731,N_3593);
and U5794 (N_5794,N_3998,N_4593);
nand U5795 (N_5795,N_2548,N_3402);
and U5796 (N_5796,N_4990,N_4282);
or U5797 (N_5797,N_3589,N_4915);
or U5798 (N_5798,N_2711,N_3865);
or U5799 (N_5799,N_4231,N_2786);
or U5800 (N_5800,N_4342,N_3368);
and U5801 (N_5801,N_3210,N_3902);
nor U5802 (N_5802,N_4883,N_2916);
nor U5803 (N_5803,N_3463,N_3377);
xnor U5804 (N_5804,N_4630,N_4985);
nand U5805 (N_5805,N_4293,N_2981);
nand U5806 (N_5806,N_3075,N_2661);
and U5807 (N_5807,N_3274,N_3619);
nand U5808 (N_5808,N_4906,N_4138);
nand U5809 (N_5809,N_4182,N_3122);
nor U5810 (N_5810,N_2760,N_4659);
nand U5811 (N_5811,N_4770,N_4705);
or U5812 (N_5812,N_2850,N_3007);
or U5813 (N_5813,N_3396,N_4833);
nand U5814 (N_5814,N_4591,N_2703);
xor U5815 (N_5815,N_3625,N_3103);
nor U5816 (N_5816,N_3890,N_3154);
and U5817 (N_5817,N_2660,N_2907);
nand U5818 (N_5818,N_3711,N_4521);
xnor U5819 (N_5819,N_3360,N_3922);
nand U5820 (N_5820,N_3652,N_4758);
nand U5821 (N_5821,N_3186,N_3823);
or U5822 (N_5822,N_2510,N_4144);
nor U5823 (N_5823,N_3944,N_3147);
or U5824 (N_5824,N_3446,N_4078);
and U5825 (N_5825,N_3501,N_4174);
nor U5826 (N_5826,N_4418,N_3077);
nand U5827 (N_5827,N_3201,N_4712);
nor U5828 (N_5828,N_2531,N_4634);
nor U5829 (N_5829,N_3213,N_4079);
nor U5830 (N_5830,N_3386,N_4740);
and U5831 (N_5831,N_2938,N_3113);
nor U5832 (N_5832,N_3980,N_3839);
and U5833 (N_5833,N_4707,N_2566);
nor U5834 (N_5834,N_4335,N_4626);
and U5835 (N_5835,N_4983,N_2623);
nand U5836 (N_5836,N_2762,N_3927);
nor U5837 (N_5837,N_2818,N_3921);
xor U5838 (N_5838,N_2668,N_4112);
nor U5839 (N_5839,N_4766,N_3781);
nand U5840 (N_5840,N_3626,N_4184);
nand U5841 (N_5841,N_2954,N_3119);
xnor U5842 (N_5842,N_3006,N_2584);
xor U5843 (N_5843,N_3806,N_3074);
or U5844 (N_5844,N_3697,N_2591);
or U5845 (N_5845,N_3769,N_2516);
or U5846 (N_5846,N_3001,N_2526);
xnor U5847 (N_5847,N_3190,N_3372);
and U5848 (N_5848,N_4631,N_4043);
nor U5849 (N_5849,N_2886,N_4376);
nor U5850 (N_5850,N_2994,N_4541);
and U5851 (N_5851,N_3152,N_4841);
nor U5852 (N_5852,N_4785,N_3094);
nor U5853 (N_5853,N_3277,N_4887);
and U5854 (N_5854,N_3384,N_4087);
and U5855 (N_5855,N_2941,N_3704);
xnor U5856 (N_5856,N_3441,N_3759);
or U5857 (N_5857,N_2541,N_4888);
and U5858 (N_5858,N_3062,N_2689);
or U5859 (N_5859,N_4204,N_4989);
nand U5860 (N_5860,N_3182,N_4797);
nand U5861 (N_5861,N_4276,N_3469);
or U5862 (N_5862,N_3148,N_2935);
xor U5863 (N_5863,N_3725,N_4750);
and U5864 (N_5864,N_2722,N_4901);
or U5865 (N_5865,N_3198,N_3683);
and U5866 (N_5866,N_4151,N_4124);
nor U5867 (N_5867,N_4608,N_2891);
and U5868 (N_5868,N_4882,N_2699);
nand U5869 (N_5869,N_4896,N_2944);
xor U5870 (N_5870,N_3519,N_4523);
nor U5871 (N_5871,N_2629,N_4566);
nor U5872 (N_5872,N_4613,N_3554);
and U5873 (N_5873,N_4726,N_4958);
and U5874 (N_5874,N_4993,N_4850);
or U5875 (N_5875,N_3013,N_4072);
and U5876 (N_5876,N_4787,N_3346);
xor U5877 (N_5877,N_3964,N_4884);
or U5878 (N_5878,N_3099,N_4258);
nand U5879 (N_5879,N_3157,N_4457);
nand U5880 (N_5880,N_4587,N_4343);
xnor U5881 (N_5881,N_3848,N_3577);
xor U5882 (N_5882,N_4313,N_4574);
nor U5883 (N_5883,N_3132,N_3882);
xor U5884 (N_5884,N_4562,N_3009);
xnor U5885 (N_5885,N_4364,N_3335);
nand U5886 (N_5886,N_4267,N_4006);
nor U5887 (N_5887,N_4789,N_3868);
and U5888 (N_5888,N_3363,N_3700);
or U5889 (N_5889,N_3635,N_4263);
or U5890 (N_5890,N_3319,N_4369);
xor U5891 (N_5891,N_3361,N_2574);
nor U5892 (N_5892,N_4230,N_4960);
xnor U5893 (N_5893,N_3656,N_4848);
nand U5894 (N_5894,N_4643,N_3216);
xor U5895 (N_5895,N_2849,N_3380);
and U5896 (N_5896,N_4674,N_4162);
nand U5897 (N_5897,N_2570,N_3555);
nand U5898 (N_5898,N_2776,N_2979);
nor U5899 (N_5899,N_4126,N_2569);
xnor U5900 (N_5900,N_2745,N_4428);
xor U5901 (N_5901,N_3171,N_4914);
nor U5902 (N_5902,N_3138,N_4270);
xor U5903 (N_5903,N_4612,N_3076);
nor U5904 (N_5904,N_4899,N_2608);
nand U5905 (N_5905,N_3691,N_4249);
xor U5906 (N_5906,N_2809,N_4513);
nor U5907 (N_5907,N_4324,N_4648);
nand U5908 (N_5908,N_4855,N_3163);
nand U5909 (N_5909,N_4565,N_3357);
xnor U5910 (N_5910,N_4023,N_4004);
and U5911 (N_5911,N_3821,N_2796);
nor U5912 (N_5912,N_4115,N_3799);
nand U5913 (N_5913,N_3723,N_4795);
nor U5914 (N_5914,N_3162,N_3370);
nand U5915 (N_5915,N_3333,N_4510);
or U5916 (N_5916,N_2613,N_4246);
nor U5917 (N_5917,N_2685,N_4624);
and U5918 (N_5918,N_4977,N_3091);
xor U5919 (N_5919,N_3820,N_3968);
xnor U5920 (N_5920,N_4280,N_4235);
or U5921 (N_5921,N_4033,N_4700);
nor U5922 (N_5922,N_2523,N_3255);
nand U5923 (N_5923,N_4967,N_4875);
or U5924 (N_5924,N_4082,N_3903);
or U5925 (N_5925,N_3595,N_2590);
and U5926 (N_5926,N_3017,N_3533);
nand U5927 (N_5927,N_2700,N_2672);
xor U5928 (N_5928,N_3466,N_3916);
and U5929 (N_5929,N_4326,N_3489);
nor U5930 (N_5930,N_3430,N_4570);
nor U5931 (N_5931,N_4134,N_4255);
or U5932 (N_5932,N_3118,N_4657);
and U5933 (N_5933,N_3100,N_3312);
and U5934 (N_5934,N_3093,N_3053);
nand U5935 (N_5935,N_3708,N_3452);
nand U5936 (N_5936,N_4530,N_2821);
nor U5937 (N_5937,N_3633,N_3254);
xor U5938 (N_5938,N_4746,N_2600);
nand U5939 (N_5939,N_4625,N_4627);
xnor U5940 (N_5940,N_3304,N_2543);
nand U5941 (N_5941,N_2581,N_4088);
nand U5942 (N_5942,N_3352,N_4816);
nor U5943 (N_5943,N_4300,N_2836);
or U5944 (N_5944,N_3437,N_4150);
or U5945 (N_5945,N_3874,N_2942);
nand U5946 (N_5946,N_4996,N_4667);
xor U5947 (N_5947,N_3824,N_4375);
nand U5948 (N_5948,N_2922,N_4241);
xnor U5949 (N_5949,N_4192,N_3106);
or U5950 (N_5950,N_4202,N_4427);
or U5951 (N_5951,N_3414,N_3788);
xor U5952 (N_5952,N_4137,N_2892);
nor U5953 (N_5953,N_2934,N_3712);
nor U5954 (N_5954,N_3487,N_4265);
nand U5955 (N_5955,N_4572,N_3879);
and U5956 (N_5956,N_2857,N_3880);
and U5957 (N_5957,N_2873,N_2804);
and U5958 (N_5958,N_4232,N_4239);
xnor U5959 (N_5959,N_3843,N_2744);
or U5960 (N_5960,N_3585,N_3451);
or U5961 (N_5961,N_3087,N_2536);
and U5962 (N_5962,N_4871,N_4540);
and U5963 (N_5963,N_4253,N_4426);
xnor U5964 (N_5964,N_3270,N_2670);
or U5965 (N_5965,N_3877,N_4058);
nand U5966 (N_5966,N_4197,N_4590);
nor U5967 (N_5967,N_2758,N_4939);
xnor U5968 (N_5968,N_4696,N_2991);
xnor U5969 (N_5969,N_4607,N_3885);
or U5970 (N_5970,N_3367,N_3984);
and U5971 (N_5971,N_3485,N_2833);
nand U5972 (N_5972,N_2923,N_4312);
or U5973 (N_5973,N_3753,N_4800);
nor U5974 (N_5974,N_4057,N_2898);
and U5975 (N_5975,N_2987,N_3272);
and U5976 (N_5976,N_2628,N_3752);
or U5977 (N_5977,N_4546,N_2772);
and U5978 (N_5978,N_2735,N_4206);
nor U5979 (N_5979,N_2572,N_3837);
xor U5980 (N_5980,N_2787,N_4632);
nor U5981 (N_5981,N_3284,N_4188);
xnor U5982 (N_5982,N_2858,N_2631);
nand U5983 (N_5983,N_3281,N_4702);
or U5984 (N_5984,N_4736,N_4031);
nand U5985 (N_5985,N_4516,N_3300);
or U5986 (N_5986,N_4819,N_2978);
nand U5987 (N_5987,N_4160,N_4805);
and U5988 (N_5988,N_4895,N_4097);
nand U5989 (N_5989,N_3247,N_3072);
xnor U5990 (N_5990,N_4401,N_2980);
xor U5991 (N_5991,N_3672,N_2632);
nor U5992 (N_5992,N_4918,N_3735);
or U5993 (N_5993,N_3231,N_3939);
nor U5994 (N_5994,N_2861,N_3749);
xor U5995 (N_5995,N_4156,N_2998);
and U5996 (N_5996,N_3503,N_2997);
and U5997 (N_5997,N_4199,N_2790);
and U5998 (N_5998,N_2562,N_4462);
and U5999 (N_5999,N_3914,N_2619);
nand U6000 (N_6000,N_4306,N_3961);
or U6001 (N_6001,N_3209,N_3857);
or U6002 (N_6002,N_3354,N_2789);
nor U6003 (N_6003,N_3359,N_4520);
xor U6004 (N_6004,N_2995,N_2561);
xor U6005 (N_6005,N_3675,N_2598);
xor U6006 (N_6006,N_3411,N_3060);
nand U6007 (N_6007,N_2638,N_3390);
xor U6008 (N_6008,N_2580,N_4980);
and U6009 (N_6009,N_4415,N_2885);
nor U6010 (N_6010,N_3904,N_3101);
and U6011 (N_6011,N_3931,N_2919);
and U6012 (N_6012,N_4635,N_2717);
and U6013 (N_6013,N_3786,N_4976);
xor U6014 (N_6014,N_3802,N_3023);
or U6015 (N_6015,N_3867,N_4456);
nor U6016 (N_6016,N_4113,N_3389);
and U6017 (N_6017,N_2884,N_2784);
and U6018 (N_6018,N_3140,N_3747);
or U6019 (N_6019,N_3311,N_4003);
nor U6020 (N_6020,N_4961,N_3567);
and U6021 (N_6021,N_2797,N_2538);
nor U6022 (N_6022,N_3884,N_3611);
and U6023 (N_6023,N_3541,N_4149);
or U6024 (N_6024,N_4499,N_4356);
xnor U6025 (N_6025,N_4784,N_4454);
xnor U6026 (N_6026,N_3640,N_3126);
xnor U6027 (N_6027,N_4444,N_3845);
nand U6028 (N_6028,N_4954,N_4892);
nand U6029 (N_6029,N_3048,N_4890);
xnor U6030 (N_6030,N_3246,N_3395);
and U6031 (N_6031,N_2973,N_2612);
nor U6032 (N_6032,N_3760,N_2664);
and U6033 (N_6033,N_3288,N_2719);
and U6034 (N_6034,N_4994,N_3234);
and U6035 (N_6035,N_3037,N_3777);
nor U6036 (N_6036,N_4585,N_4474);
xnor U6037 (N_6037,N_3097,N_4090);
xnor U6038 (N_6038,N_4889,N_4254);
nor U6039 (N_6039,N_2635,N_3713);
nor U6040 (N_6040,N_2819,N_4411);
xor U6041 (N_6041,N_4908,N_3973);
and U6042 (N_6042,N_2737,N_3643);
nor U6043 (N_6043,N_3047,N_4637);
xor U6044 (N_6044,N_4423,N_4281);
or U6045 (N_6045,N_4881,N_3605);
and U6046 (N_6046,N_3528,N_4940);
and U6047 (N_6047,N_3650,N_3917);
nor U6048 (N_6048,N_3208,N_4211);
xor U6049 (N_6049,N_2899,N_3306);
or U6050 (N_6050,N_3754,N_3817);
and U6051 (N_6051,N_4130,N_2812);
xnor U6052 (N_6052,N_4038,N_4227);
nand U6053 (N_6053,N_4252,N_3151);
xnor U6054 (N_6054,N_4553,N_4083);
or U6055 (N_6055,N_3316,N_2730);
nor U6056 (N_6056,N_3134,N_2828);
and U6057 (N_6057,N_4478,N_3850);
or U6058 (N_6058,N_4798,N_2755);
or U6059 (N_6059,N_4956,N_3245);
nor U6060 (N_6060,N_3261,N_4214);
nor U6061 (N_6061,N_4807,N_4586);
nor U6062 (N_6062,N_4012,N_3292);
and U6063 (N_6063,N_4963,N_4928);
or U6064 (N_6064,N_4970,N_3745);
and U6065 (N_6065,N_4760,N_3338);
and U6066 (N_6066,N_4154,N_4026);
xor U6067 (N_6067,N_2779,N_4768);
nand U6068 (N_6068,N_3590,N_4846);
nand U6069 (N_6069,N_3095,N_3602);
nor U6070 (N_6070,N_3490,N_4642);
or U6071 (N_6071,N_3253,N_2791);
or U6072 (N_6072,N_2780,N_2890);
nand U6073 (N_6073,N_3364,N_3373);
xnor U6074 (N_6074,N_3258,N_4027);
nand U6075 (N_6075,N_3509,N_3036);
or U6076 (N_6076,N_4944,N_4602);
or U6077 (N_6077,N_2825,N_3693);
xor U6078 (N_6078,N_2913,N_4297);
nor U6079 (N_6079,N_2771,N_2863);
nor U6080 (N_6080,N_4485,N_4089);
and U6081 (N_6081,N_3282,N_4358);
and U6082 (N_6082,N_3345,N_2687);
nor U6083 (N_6083,N_3957,N_3651);
or U6084 (N_6084,N_4577,N_3318);
and U6085 (N_6085,N_3374,N_2567);
and U6086 (N_6086,N_3236,N_2975);
xor U6087 (N_6087,N_3740,N_3774);
or U6088 (N_6088,N_3588,N_2611);
xnor U6089 (N_6089,N_4186,N_3906);
nand U6090 (N_6090,N_2726,N_4603);
or U6091 (N_6091,N_4104,N_4438);
and U6092 (N_6092,N_4060,N_3869);
nor U6093 (N_6093,N_4310,N_3989);
or U6094 (N_6094,N_4283,N_3114);
nand U6095 (N_6095,N_3195,N_4716);
xnor U6096 (N_6096,N_4765,N_4598);
nand U6097 (N_6097,N_3150,N_4452);
and U6098 (N_6098,N_4886,N_4664);
nor U6099 (N_6099,N_3804,N_2962);
nand U6100 (N_6100,N_4704,N_3005);
nand U6101 (N_6101,N_4723,N_4560);
nand U6102 (N_6102,N_2748,N_4399);
or U6103 (N_6103,N_4009,N_4264);
and U6104 (N_6104,N_3615,N_4951);
nand U6105 (N_6105,N_3022,N_3477);
or U6106 (N_6106,N_4859,N_2521);
nand U6107 (N_6107,N_3068,N_2627);
nand U6108 (N_6108,N_4295,N_2643);
and U6109 (N_6109,N_3191,N_2879);
nand U6110 (N_6110,N_3447,N_4872);
or U6111 (N_6111,N_4853,N_4380);
or U6112 (N_6112,N_4734,N_4692);
or U6113 (N_6113,N_2596,N_4351);
nor U6114 (N_6114,N_2585,N_4044);
nor U6115 (N_6115,N_3766,N_4621);
nor U6116 (N_6116,N_4861,N_3476);
or U6117 (N_6117,N_3666,N_4568);
xnor U6118 (N_6118,N_4354,N_4941);
and U6119 (N_6119,N_2798,N_3954);
nor U6120 (N_6120,N_3608,N_4497);
nand U6121 (N_6121,N_4968,N_3889);
nor U6122 (N_6122,N_2554,N_4289);
and U6123 (N_6123,N_3991,N_3124);
and U6124 (N_6124,N_2937,N_3876);
nor U6125 (N_6125,N_3289,N_4737);
xnor U6126 (N_6126,N_2893,N_4299);
nand U6127 (N_6127,N_4999,N_2959);
or U6128 (N_6128,N_4290,N_3825);
nor U6129 (N_6129,N_4311,N_3468);
nor U6130 (N_6130,N_2733,N_3722);
xor U6131 (N_6131,N_2607,N_3896);
nand U6132 (N_6132,N_4831,N_3264);
and U6133 (N_6133,N_3701,N_3003);
or U6134 (N_6134,N_3480,N_3434);
nand U6135 (N_6135,N_4219,N_3358);
nor U6136 (N_6136,N_3290,N_2636);
and U6137 (N_6137,N_3293,N_4703);
xor U6138 (N_6138,N_3392,N_4064);
or U6139 (N_6139,N_3431,N_4661);
or U6140 (N_6140,N_2992,N_3669);
and U6141 (N_6141,N_4681,N_2695);
nor U6142 (N_6142,N_4261,N_3232);
xnor U6143 (N_6143,N_2866,N_4747);
xnor U6144 (N_6144,N_2795,N_3059);
xor U6145 (N_6145,N_4902,N_4378);
nor U6146 (N_6146,N_3974,N_4487);
nor U6147 (N_6147,N_3257,N_4815);
nand U6148 (N_6148,N_4834,N_2859);
nand U6149 (N_6149,N_4957,N_2583);
or U6150 (N_6150,N_2933,N_4843);
and U6151 (N_6151,N_4927,N_4480);
xnor U6152 (N_6152,N_2736,N_2565);
nand U6153 (N_6153,N_3832,N_3058);
nand U6154 (N_6154,N_4563,N_3791);
or U6155 (N_6155,N_2525,N_4988);
nand U6156 (N_6156,N_3027,N_3301);
nand U6157 (N_6157,N_2575,N_3928);
xnor U6158 (N_6158,N_4793,N_3249);
nand U6159 (N_6159,N_3737,N_2883);
or U6160 (N_6160,N_3110,N_2530);
nand U6161 (N_6161,N_3011,N_2947);
nand U6162 (N_6162,N_4685,N_4979);
or U6163 (N_6163,N_4594,N_4387);
or U6164 (N_6164,N_4413,N_2597);
or U6165 (N_6165,N_3878,N_4320);
and U6166 (N_6166,N_2710,N_2616);
xor U6167 (N_6167,N_4491,N_2704);
nor U6168 (N_6168,N_3570,N_4040);
nand U6169 (N_6169,N_3648,N_2509);
nor U6170 (N_6170,N_3862,N_3104);
nand U6171 (N_6171,N_3604,N_4198);
nor U6172 (N_6172,N_4525,N_4972);
nor U6173 (N_6173,N_4208,N_3475);
and U6174 (N_6174,N_4274,N_2517);
and U6175 (N_6175,N_4461,N_4774);
or U6176 (N_6176,N_4207,N_3317);
nand U6177 (N_6177,N_4440,N_3398);
nand U6178 (N_6178,N_3853,N_2957);
nand U6179 (N_6179,N_3523,N_4537);
and U6180 (N_6180,N_3562,N_4549);
nand U6181 (N_6181,N_4932,N_3706);
nand U6182 (N_6182,N_4477,N_4863);
nand U6183 (N_6183,N_3169,N_4938);
nand U6184 (N_6184,N_2599,N_2658);
nand U6185 (N_6185,N_3339,N_4804);
nand U6186 (N_6186,N_4325,N_2988);
and U6187 (N_6187,N_4605,N_4145);
or U6188 (N_6188,N_3797,N_3596);
or U6189 (N_6189,N_3355,N_4646);
xor U6190 (N_6190,N_2960,N_3019);
and U6191 (N_6191,N_2535,N_3778);
or U6192 (N_6192,N_3418,N_3645);
xor U6193 (N_6193,N_4002,N_4209);
xnor U6194 (N_6194,N_4923,N_3408);
xor U6195 (N_6195,N_4292,N_2595);
xnor U6196 (N_6196,N_3732,N_4794);
nand U6197 (N_6197,N_3458,N_2876);
nand U6198 (N_6198,N_3899,N_3298);
xor U6199 (N_6199,N_2505,N_4964);
nand U6200 (N_6200,N_3128,N_4614);
nor U6201 (N_6201,N_2826,N_4599);
or U6202 (N_6202,N_3415,N_2582);
and U6203 (N_6203,N_3387,N_4029);
nand U6204 (N_6204,N_4503,N_4353);
and U6205 (N_6205,N_2743,N_3913);
nor U6206 (N_6206,N_4096,N_3720);
xnor U6207 (N_6207,N_4847,N_3108);
or U6208 (N_6208,N_4538,N_3692);
xor U6209 (N_6209,N_3511,N_4101);
or U6210 (N_6210,N_4394,N_4243);
and U6211 (N_6211,N_4647,N_4679);
nand U6212 (N_6212,N_3337,N_4653);
or U6213 (N_6213,N_4879,N_3919);
or U6214 (N_6214,N_4744,N_4536);
and U6215 (N_6215,N_3505,N_4287);
nor U6216 (N_6216,N_3537,N_3342);
nor U6217 (N_6217,N_3883,N_4417);
xor U6218 (N_6218,N_3421,N_4405);
or U6219 (N_6219,N_4495,N_2633);
and U6220 (N_6220,N_4869,N_3343);
and U6221 (N_6221,N_3063,N_2801);
nand U6222 (N_6222,N_2673,N_4016);
or U6223 (N_6223,N_2688,N_4481);
nor U6224 (N_6224,N_4856,N_3291);
nor U6225 (N_6225,N_3196,N_3582);
and U6226 (N_6226,N_4697,N_4910);
xor U6227 (N_6227,N_2875,N_4658);
xor U6228 (N_6228,N_4771,N_3052);
nand U6229 (N_6229,N_3029,N_3222);
or U6230 (N_6230,N_2576,N_4852);
and U6231 (N_6231,N_3550,N_3428);
and U6232 (N_6232,N_3238,N_2642);
nor U6233 (N_6233,N_4256,N_2822);
and U6234 (N_6234,N_4398,N_4912);
xor U6235 (N_6235,N_3793,N_3330);
nor U6236 (N_6236,N_2648,N_3531);
nand U6237 (N_6237,N_4221,N_2769);
nand U6238 (N_6238,N_4388,N_3598);
xnor U6239 (N_6239,N_3574,N_3313);
and U6240 (N_6240,N_4269,N_4111);
nand U6241 (N_6241,N_4443,N_4015);
and U6242 (N_6242,N_3105,N_4344);
nand U6243 (N_6243,N_2646,N_2545);
xnor U6244 (N_6244,N_2588,N_4757);
and U6245 (N_6245,N_3256,N_3995);
nand U6246 (N_6246,N_4920,N_4429);
nor U6247 (N_6247,N_4402,N_3703);
or U6248 (N_6248,N_3212,N_4609);
nor U6249 (N_6249,N_4080,N_2559);
nor U6250 (N_6250,N_3259,N_4087);
and U6251 (N_6251,N_4859,N_2821);
nand U6252 (N_6252,N_3555,N_3248);
nand U6253 (N_6253,N_4305,N_4593);
nor U6254 (N_6254,N_3984,N_3049);
xnor U6255 (N_6255,N_2575,N_4877);
xnor U6256 (N_6256,N_3631,N_3938);
nor U6257 (N_6257,N_2976,N_3874);
and U6258 (N_6258,N_3716,N_3311);
and U6259 (N_6259,N_2737,N_2621);
nand U6260 (N_6260,N_3689,N_3534);
or U6261 (N_6261,N_2890,N_3221);
and U6262 (N_6262,N_3983,N_3846);
or U6263 (N_6263,N_2698,N_3491);
and U6264 (N_6264,N_3468,N_3881);
and U6265 (N_6265,N_3397,N_4830);
and U6266 (N_6266,N_2680,N_3049);
nor U6267 (N_6267,N_4751,N_3880);
xor U6268 (N_6268,N_3403,N_3800);
nand U6269 (N_6269,N_4312,N_4315);
or U6270 (N_6270,N_3285,N_4910);
and U6271 (N_6271,N_4272,N_2811);
and U6272 (N_6272,N_4263,N_2577);
nand U6273 (N_6273,N_3909,N_3730);
xnor U6274 (N_6274,N_4218,N_3902);
nand U6275 (N_6275,N_4425,N_2544);
or U6276 (N_6276,N_3118,N_4557);
xnor U6277 (N_6277,N_4942,N_4365);
and U6278 (N_6278,N_2778,N_4374);
nor U6279 (N_6279,N_4728,N_2538);
xor U6280 (N_6280,N_4914,N_2832);
nand U6281 (N_6281,N_3556,N_4504);
xnor U6282 (N_6282,N_3835,N_4845);
nor U6283 (N_6283,N_2959,N_4528);
nor U6284 (N_6284,N_4585,N_3034);
nand U6285 (N_6285,N_4053,N_3028);
nor U6286 (N_6286,N_4939,N_4289);
nand U6287 (N_6287,N_2574,N_4088);
or U6288 (N_6288,N_3381,N_3199);
xnor U6289 (N_6289,N_3037,N_4968);
nor U6290 (N_6290,N_4384,N_4435);
or U6291 (N_6291,N_2565,N_3549);
or U6292 (N_6292,N_3054,N_4645);
and U6293 (N_6293,N_2991,N_3870);
nand U6294 (N_6294,N_2831,N_4214);
and U6295 (N_6295,N_3378,N_4144);
xnor U6296 (N_6296,N_4765,N_4542);
and U6297 (N_6297,N_3523,N_4145);
or U6298 (N_6298,N_3181,N_2938);
or U6299 (N_6299,N_4696,N_2622);
nand U6300 (N_6300,N_2703,N_2554);
or U6301 (N_6301,N_4342,N_4808);
nand U6302 (N_6302,N_2706,N_2579);
or U6303 (N_6303,N_4146,N_3609);
xnor U6304 (N_6304,N_2746,N_4223);
xnor U6305 (N_6305,N_2513,N_3409);
and U6306 (N_6306,N_3492,N_4914);
nor U6307 (N_6307,N_4612,N_3994);
nand U6308 (N_6308,N_4970,N_2694);
nor U6309 (N_6309,N_4827,N_2653);
nor U6310 (N_6310,N_3929,N_4516);
xor U6311 (N_6311,N_2982,N_4014);
nor U6312 (N_6312,N_4315,N_3626);
nand U6313 (N_6313,N_4284,N_4159);
xor U6314 (N_6314,N_2940,N_3936);
xor U6315 (N_6315,N_4440,N_3986);
or U6316 (N_6316,N_4835,N_3189);
and U6317 (N_6317,N_4799,N_2967);
and U6318 (N_6318,N_4053,N_4856);
and U6319 (N_6319,N_3687,N_3888);
and U6320 (N_6320,N_3827,N_3595);
or U6321 (N_6321,N_4253,N_4689);
nor U6322 (N_6322,N_4451,N_4220);
nor U6323 (N_6323,N_3651,N_4461);
xnor U6324 (N_6324,N_3082,N_4481);
xnor U6325 (N_6325,N_4884,N_4961);
and U6326 (N_6326,N_2871,N_2644);
xor U6327 (N_6327,N_4122,N_2711);
xnor U6328 (N_6328,N_3693,N_3549);
xnor U6329 (N_6329,N_4960,N_4823);
xnor U6330 (N_6330,N_4148,N_4822);
nand U6331 (N_6331,N_2927,N_4966);
xor U6332 (N_6332,N_4124,N_3704);
and U6333 (N_6333,N_4792,N_4084);
xor U6334 (N_6334,N_4728,N_3601);
or U6335 (N_6335,N_2704,N_3270);
or U6336 (N_6336,N_3291,N_4356);
xor U6337 (N_6337,N_3102,N_3157);
nor U6338 (N_6338,N_3820,N_2737);
nor U6339 (N_6339,N_2871,N_4204);
and U6340 (N_6340,N_3134,N_2931);
nand U6341 (N_6341,N_3237,N_4390);
nand U6342 (N_6342,N_4253,N_4956);
or U6343 (N_6343,N_4079,N_3864);
nor U6344 (N_6344,N_4636,N_2756);
nor U6345 (N_6345,N_3870,N_4430);
nor U6346 (N_6346,N_3469,N_4218);
nand U6347 (N_6347,N_2992,N_4704);
xor U6348 (N_6348,N_2919,N_4799);
nand U6349 (N_6349,N_3771,N_3064);
nand U6350 (N_6350,N_4597,N_3386);
nor U6351 (N_6351,N_4251,N_2755);
and U6352 (N_6352,N_4863,N_3758);
nand U6353 (N_6353,N_3186,N_4415);
and U6354 (N_6354,N_4902,N_3115);
nor U6355 (N_6355,N_4686,N_4537);
nor U6356 (N_6356,N_4443,N_3829);
and U6357 (N_6357,N_4529,N_4563);
nor U6358 (N_6358,N_3243,N_3455);
nor U6359 (N_6359,N_3574,N_3532);
nand U6360 (N_6360,N_3474,N_4154);
and U6361 (N_6361,N_3364,N_3466);
nand U6362 (N_6362,N_2975,N_4218);
and U6363 (N_6363,N_4512,N_4456);
or U6364 (N_6364,N_2667,N_3166);
and U6365 (N_6365,N_4725,N_3855);
nand U6366 (N_6366,N_4951,N_3820);
nand U6367 (N_6367,N_4335,N_4323);
nor U6368 (N_6368,N_4650,N_2609);
nor U6369 (N_6369,N_2553,N_3140);
nand U6370 (N_6370,N_2886,N_3865);
nand U6371 (N_6371,N_4590,N_4029);
or U6372 (N_6372,N_2808,N_3798);
xnor U6373 (N_6373,N_4145,N_3505);
xor U6374 (N_6374,N_2799,N_4647);
xnor U6375 (N_6375,N_3924,N_4860);
xnor U6376 (N_6376,N_3100,N_3202);
nor U6377 (N_6377,N_3697,N_4848);
and U6378 (N_6378,N_3752,N_2879);
nor U6379 (N_6379,N_3602,N_3691);
nor U6380 (N_6380,N_2932,N_3211);
and U6381 (N_6381,N_3865,N_4844);
xnor U6382 (N_6382,N_2698,N_2502);
nor U6383 (N_6383,N_3658,N_3172);
nor U6384 (N_6384,N_4561,N_4016);
or U6385 (N_6385,N_3677,N_4267);
and U6386 (N_6386,N_3764,N_3967);
or U6387 (N_6387,N_4286,N_3277);
nor U6388 (N_6388,N_2984,N_4927);
and U6389 (N_6389,N_2799,N_3180);
nand U6390 (N_6390,N_4712,N_3817);
nor U6391 (N_6391,N_2950,N_3542);
xor U6392 (N_6392,N_4149,N_4062);
nor U6393 (N_6393,N_4268,N_2937);
nand U6394 (N_6394,N_2528,N_3612);
and U6395 (N_6395,N_2717,N_4433);
xnor U6396 (N_6396,N_3590,N_4450);
nand U6397 (N_6397,N_4155,N_3424);
or U6398 (N_6398,N_4284,N_3181);
and U6399 (N_6399,N_4663,N_4482);
nor U6400 (N_6400,N_4110,N_4828);
nor U6401 (N_6401,N_4220,N_2853);
nand U6402 (N_6402,N_3897,N_3271);
and U6403 (N_6403,N_4374,N_3144);
xnor U6404 (N_6404,N_4983,N_2829);
or U6405 (N_6405,N_3200,N_4304);
and U6406 (N_6406,N_4317,N_4246);
and U6407 (N_6407,N_4848,N_3587);
or U6408 (N_6408,N_4831,N_2870);
or U6409 (N_6409,N_3516,N_3920);
nand U6410 (N_6410,N_4052,N_2999);
and U6411 (N_6411,N_4322,N_4327);
or U6412 (N_6412,N_2552,N_4185);
and U6413 (N_6413,N_3864,N_4339);
nor U6414 (N_6414,N_2596,N_4056);
xor U6415 (N_6415,N_3867,N_3360);
nor U6416 (N_6416,N_4478,N_4991);
xor U6417 (N_6417,N_2963,N_3622);
or U6418 (N_6418,N_3921,N_3948);
nor U6419 (N_6419,N_4196,N_3865);
nor U6420 (N_6420,N_4865,N_3519);
nor U6421 (N_6421,N_4737,N_4874);
and U6422 (N_6422,N_2778,N_3605);
or U6423 (N_6423,N_4882,N_2705);
nand U6424 (N_6424,N_4302,N_3463);
nand U6425 (N_6425,N_4695,N_3690);
or U6426 (N_6426,N_3925,N_3857);
or U6427 (N_6427,N_3958,N_3328);
nor U6428 (N_6428,N_2786,N_4037);
nand U6429 (N_6429,N_3730,N_4510);
nand U6430 (N_6430,N_3721,N_3822);
or U6431 (N_6431,N_3159,N_2679);
or U6432 (N_6432,N_3821,N_3013);
nand U6433 (N_6433,N_2834,N_3183);
nand U6434 (N_6434,N_3986,N_4231);
nand U6435 (N_6435,N_3842,N_3228);
nor U6436 (N_6436,N_4687,N_3107);
or U6437 (N_6437,N_3247,N_3838);
nor U6438 (N_6438,N_3557,N_4673);
nor U6439 (N_6439,N_4901,N_3038);
and U6440 (N_6440,N_3317,N_3502);
nor U6441 (N_6441,N_4843,N_3607);
xor U6442 (N_6442,N_3671,N_4743);
or U6443 (N_6443,N_2674,N_2574);
nand U6444 (N_6444,N_2667,N_3026);
nor U6445 (N_6445,N_4711,N_4550);
xor U6446 (N_6446,N_3774,N_4514);
nor U6447 (N_6447,N_2881,N_4522);
nand U6448 (N_6448,N_3209,N_4725);
nand U6449 (N_6449,N_4845,N_2617);
nor U6450 (N_6450,N_4241,N_3382);
nor U6451 (N_6451,N_3539,N_2816);
nor U6452 (N_6452,N_3109,N_3814);
or U6453 (N_6453,N_4018,N_3807);
nand U6454 (N_6454,N_4196,N_4800);
xor U6455 (N_6455,N_4209,N_3145);
nand U6456 (N_6456,N_4386,N_4633);
or U6457 (N_6457,N_4415,N_4207);
nand U6458 (N_6458,N_3213,N_4243);
nor U6459 (N_6459,N_3984,N_2592);
or U6460 (N_6460,N_4400,N_4090);
nor U6461 (N_6461,N_4260,N_4483);
or U6462 (N_6462,N_2922,N_4118);
nand U6463 (N_6463,N_2544,N_3163);
xor U6464 (N_6464,N_3964,N_4012);
nor U6465 (N_6465,N_3528,N_4676);
xnor U6466 (N_6466,N_3005,N_4592);
xnor U6467 (N_6467,N_3557,N_2746);
nor U6468 (N_6468,N_3244,N_2571);
and U6469 (N_6469,N_3672,N_4112);
or U6470 (N_6470,N_4149,N_3335);
xor U6471 (N_6471,N_4824,N_4039);
xnor U6472 (N_6472,N_3031,N_4972);
nand U6473 (N_6473,N_4309,N_4282);
xnor U6474 (N_6474,N_3399,N_4030);
nor U6475 (N_6475,N_4729,N_3840);
nor U6476 (N_6476,N_4086,N_2668);
xor U6477 (N_6477,N_4825,N_4148);
or U6478 (N_6478,N_4363,N_3093);
nor U6479 (N_6479,N_4004,N_4618);
and U6480 (N_6480,N_3971,N_3737);
nand U6481 (N_6481,N_4375,N_3289);
nor U6482 (N_6482,N_4805,N_2561);
or U6483 (N_6483,N_4188,N_4148);
xor U6484 (N_6484,N_2651,N_3288);
xnor U6485 (N_6485,N_2629,N_3721);
and U6486 (N_6486,N_4152,N_4488);
nand U6487 (N_6487,N_3673,N_3454);
xor U6488 (N_6488,N_2852,N_3770);
and U6489 (N_6489,N_4535,N_3285);
xor U6490 (N_6490,N_3249,N_3230);
xnor U6491 (N_6491,N_3313,N_2936);
and U6492 (N_6492,N_3680,N_2951);
and U6493 (N_6493,N_3955,N_4833);
nand U6494 (N_6494,N_4669,N_4634);
nor U6495 (N_6495,N_4673,N_3763);
nor U6496 (N_6496,N_4644,N_2734);
xor U6497 (N_6497,N_4297,N_2518);
xnor U6498 (N_6498,N_4166,N_4155);
nand U6499 (N_6499,N_4346,N_3560);
nand U6500 (N_6500,N_3839,N_4964);
nor U6501 (N_6501,N_2937,N_3097);
nand U6502 (N_6502,N_4401,N_2667);
or U6503 (N_6503,N_2956,N_2634);
or U6504 (N_6504,N_2589,N_4055);
xnor U6505 (N_6505,N_2778,N_3498);
nand U6506 (N_6506,N_2879,N_3480);
or U6507 (N_6507,N_3230,N_2552);
nor U6508 (N_6508,N_4254,N_3681);
or U6509 (N_6509,N_2804,N_3779);
nor U6510 (N_6510,N_2555,N_4234);
xor U6511 (N_6511,N_3352,N_4699);
nor U6512 (N_6512,N_4811,N_3788);
xor U6513 (N_6513,N_4640,N_4537);
nor U6514 (N_6514,N_3244,N_3914);
and U6515 (N_6515,N_2530,N_4001);
nand U6516 (N_6516,N_4924,N_4609);
nand U6517 (N_6517,N_2658,N_4540);
nand U6518 (N_6518,N_3519,N_3428);
or U6519 (N_6519,N_2699,N_3541);
xnor U6520 (N_6520,N_3793,N_2858);
nor U6521 (N_6521,N_4306,N_3653);
and U6522 (N_6522,N_4133,N_4216);
xor U6523 (N_6523,N_3326,N_4037);
xnor U6524 (N_6524,N_3287,N_3146);
nor U6525 (N_6525,N_4880,N_3589);
xor U6526 (N_6526,N_3279,N_3104);
xnor U6527 (N_6527,N_4811,N_4502);
xnor U6528 (N_6528,N_4522,N_3806);
and U6529 (N_6529,N_3514,N_4639);
and U6530 (N_6530,N_2561,N_3674);
and U6531 (N_6531,N_4884,N_3883);
xor U6532 (N_6532,N_3684,N_3496);
and U6533 (N_6533,N_3033,N_3819);
and U6534 (N_6534,N_3789,N_2830);
or U6535 (N_6535,N_4450,N_3227);
nor U6536 (N_6536,N_3661,N_3202);
xor U6537 (N_6537,N_2963,N_2886);
nor U6538 (N_6538,N_3980,N_3646);
xnor U6539 (N_6539,N_4990,N_3921);
xnor U6540 (N_6540,N_3256,N_4606);
nand U6541 (N_6541,N_3031,N_4921);
xnor U6542 (N_6542,N_4377,N_4752);
nor U6543 (N_6543,N_2502,N_3450);
or U6544 (N_6544,N_3752,N_3479);
nor U6545 (N_6545,N_3354,N_2585);
xnor U6546 (N_6546,N_3820,N_3669);
and U6547 (N_6547,N_4785,N_3949);
or U6548 (N_6548,N_3714,N_4944);
or U6549 (N_6549,N_4490,N_3891);
or U6550 (N_6550,N_3345,N_4247);
xor U6551 (N_6551,N_4518,N_4392);
and U6552 (N_6552,N_3658,N_2896);
nand U6553 (N_6553,N_2848,N_4277);
nor U6554 (N_6554,N_4690,N_3234);
or U6555 (N_6555,N_2675,N_3194);
and U6556 (N_6556,N_4148,N_4208);
nor U6557 (N_6557,N_4412,N_3670);
xnor U6558 (N_6558,N_3060,N_2828);
and U6559 (N_6559,N_3585,N_3182);
xor U6560 (N_6560,N_3586,N_2878);
xnor U6561 (N_6561,N_4894,N_4281);
or U6562 (N_6562,N_3217,N_4008);
nor U6563 (N_6563,N_2711,N_3474);
and U6564 (N_6564,N_2547,N_3332);
xnor U6565 (N_6565,N_3067,N_4550);
and U6566 (N_6566,N_2873,N_3653);
nor U6567 (N_6567,N_3572,N_2737);
xnor U6568 (N_6568,N_4381,N_3196);
xnor U6569 (N_6569,N_2990,N_4235);
or U6570 (N_6570,N_4358,N_3601);
or U6571 (N_6571,N_3096,N_3058);
and U6572 (N_6572,N_2536,N_4515);
xnor U6573 (N_6573,N_3250,N_3193);
nor U6574 (N_6574,N_2502,N_4581);
nor U6575 (N_6575,N_4423,N_4597);
nor U6576 (N_6576,N_4457,N_2501);
xor U6577 (N_6577,N_4219,N_4461);
nand U6578 (N_6578,N_3408,N_2517);
or U6579 (N_6579,N_3362,N_2815);
and U6580 (N_6580,N_3500,N_2777);
xnor U6581 (N_6581,N_2529,N_4197);
nor U6582 (N_6582,N_2953,N_3082);
and U6583 (N_6583,N_3682,N_3358);
nor U6584 (N_6584,N_4775,N_4717);
nor U6585 (N_6585,N_4606,N_2882);
nand U6586 (N_6586,N_3584,N_4725);
xor U6587 (N_6587,N_2981,N_4321);
or U6588 (N_6588,N_4929,N_4282);
nand U6589 (N_6589,N_4273,N_4003);
nand U6590 (N_6590,N_3817,N_4156);
and U6591 (N_6591,N_3717,N_4230);
nor U6592 (N_6592,N_2963,N_3191);
and U6593 (N_6593,N_2685,N_4217);
nor U6594 (N_6594,N_4948,N_4226);
and U6595 (N_6595,N_3864,N_2830);
and U6596 (N_6596,N_3929,N_3986);
or U6597 (N_6597,N_2581,N_4596);
nand U6598 (N_6598,N_3622,N_3968);
and U6599 (N_6599,N_4502,N_3389);
nand U6600 (N_6600,N_2725,N_3451);
xnor U6601 (N_6601,N_3053,N_2774);
xnor U6602 (N_6602,N_4007,N_4288);
nor U6603 (N_6603,N_2987,N_3466);
or U6604 (N_6604,N_3490,N_2806);
and U6605 (N_6605,N_3815,N_4904);
or U6606 (N_6606,N_3642,N_4540);
nor U6607 (N_6607,N_3346,N_3248);
nand U6608 (N_6608,N_4483,N_3513);
nand U6609 (N_6609,N_3649,N_4574);
and U6610 (N_6610,N_4013,N_3271);
nor U6611 (N_6611,N_4197,N_2631);
xor U6612 (N_6612,N_3774,N_4322);
xnor U6613 (N_6613,N_2633,N_4363);
nand U6614 (N_6614,N_3883,N_2511);
nand U6615 (N_6615,N_4958,N_4868);
or U6616 (N_6616,N_2977,N_3834);
or U6617 (N_6617,N_3801,N_4345);
nor U6618 (N_6618,N_2736,N_4605);
and U6619 (N_6619,N_3936,N_3597);
and U6620 (N_6620,N_4656,N_3630);
or U6621 (N_6621,N_3369,N_4323);
and U6622 (N_6622,N_3574,N_3099);
or U6623 (N_6623,N_3998,N_3420);
or U6624 (N_6624,N_3790,N_3445);
and U6625 (N_6625,N_3246,N_3150);
and U6626 (N_6626,N_3264,N_4481);
nor U6627 (N_6627,N_4586,N_2970);
and U6628 (N_6628,N_3970,N_4288);
xor U6629 (N_6629,N_3380,N_4585);
xnor U6630 (N_6630,N_3461,N_3120);
nand U6631 (N_6631,N_4659,N_3808);
nor U6632 (N_6632,N_4095,N_4242);
nand U6633 (N_6633,N_4815,N_3665);
or U6634 (N_6634,N_3427,N_3802);
xnor U6635 (N_6635,N_4550,N_3571);
xor U6636 (N_6636,N_4997,N_4410);
xor U6637 (N_6637,N_4849,N_2523);
nor U6638 (N_6638,N_3927,N_2896);
nand U6639 (N_6639,N_4603,N_4495);
or U6640 (N_6640,N_4040,N_3292);
and U6641 (N_6641,N_3982,N_2862);
and U6642 (N_6642,N_2892,N_3466);
nor U6643 (N_6643,N_3570,N_4554);
xnor U6644 (N_6644,N_4890,N_3344);
and U6645 (N_6645,N_4852,N_3785);
nor U6646 (N_6646,N_3598,N_2616);
or U6647 (N_6647,N_2843,N_3323);
or U6648 (N_6648,N_4132,N_4119);
nor U6649 (N_6649,N_4570,N_3733);
or U6650 (N_6650,N_2718,N_4299);
and U6651 (N_6651,N_3710,N_3039);
xor U6652 (N_6652,N_2958,N_3436);
and U6653 (N_6653,N_4917,N_4883);
and U6654 (N_6654,N_3152,N_4394);
and U6655 (N_6655,N_4955,N_3087);
xnor U6656 (N_6656,N_3934,N_3898);
xor U6657 (N_6657,N_2829,N_2997);
or U6658 (N_6658,N_3517,N_3764);
xor U6659 (N_6659,N_3248,N_3850);
and U6660 (N_6660,N_2728,N_4320);
nand U6661 (N_6661,N_3171,N_4396);
nor U6662 (N_6662,N_3471,N_4731);
nand U6663 (N_6663,N_4593,N_4694);
and U6664 (N_6664,N_3911,N_2952);
and U6665 (N_6665,N_4913,N_2750);
nand U6666 (N_6666,N_3697,N_3298);
nand U6667 (N_6667,N_2952,N_2962);
or U6668 (N_6668,N_4753,N_4252);
nor U6669 (N_6669,N_4557,N_2627);
and U6670 (N_6670,N_3335,N_4899);
and U6671 (N_6671,N_4259,N_4343);
nand U6672 (N_6672,N_4331,N_3396);
nor U6673 (N_6673,N_3016,N_3574);
xnor U6674 (N_6674,N_4079,N_2526);
and U6675 (N_6675,N_3484,N_3765);
and U6676 (N_6676,N_2648,N_3449);
and U6677 (N_6677,N_4110,N_4694);
or U6678 (N_6678,N_3569,N_3739);
and U6679 (N_6679,N_4972,N_4590);
nand U6680 (N_6680,N_2784,N_4329);
and U6681 (N_6681,N_2969,N_3561);
or U6682 (N_6682,N_3638,N_2549);
nor U6683 (N_6683,N_3443,N_3942);
nand U6684 (N_6684,N_4944,N_4537);
nand U6685 (N_6685,N_4065,N_3526);
nand U6686 (N_6686,N_2918,N_4020);
nor U6687 (N_6687,N_3053,N_4181);
xor U6688 (N_6688,N_2518,N_3739);
nand U6689 (N_6689,N_4823,N_3666);
xor U6690 (N_6690,N_3586,N_4644);
nand U6691 (N_6691,N_4940,N_4422);
nand U6692 (N_6692,N_3020,N_3030);
nand U6693 (N_6693,N_4521,N_4905);
and U6694 (N_6694,N_4998,N_4665);
nor U6695 (N_6695,N_3631,N_3462);
or U6696 (N_6696,N_4961,N_4190);
and U6697 (N_6697,N_3639,N_4721);
and U6698 (N_6698,N_3170,N_3029);
xnor U6699 (N_6699,N_4739,N_2618);
or U6700 (N_6700,N_3192,N_3108);
nor U6701 (N_6701,N_4486,N_2568);
xnor U6702 (N_6702,N_3292,N_4418);
and U6703 (N_6703,N_3994,N_4260);
and U6704 (N_6704,N_4909,N_4609);
or U6705 (N_6705,N_2539,N_3153);
and U6706 (N_6706,N_4777,N_4530);
nor U6707 (N_6707,N_4961,N_3215);
nor U6708 (N_6708,N_4686,N_4209);
nor U6709 (N_6709,N_4412,N_2589);
or U6710 (N_6710,N_3972,N_2529);
nor U6711 (N_6711,N_3549,N_3114);
and U6712 (N_6712,N_3651,N_2939);
xnor U6713 (N_6713,N_4950,N_3429);
nand U6714 (N_6714,N_4109,N_4885);
or U6715 (N_6715,N_2937,N_4996);
and U6716 (N_6716,N_4160,N_4225);
or U6717 (N_6717,N_2939,N_4135);
and U6718 (N_6718,N_3696,N_2702);
and U6719 (N_6719,N_4095,N_3804);
or U6720 (N_6720,N_3580,N_4348);
and U6721 (N_6721,N_3159,N_2700);
nand U6722 (N_6722,N_3240,N_3457);
xnor U6723 (N_6723,N_2974,N_4882);
nor U6724 (N_6724,N_3713,N_2892);
nor U6725 (N_6725,N_3424,N_4824);
and U6726 (N_6726,N_2652,N_3353);
nand U6727 (N_6727,N_4971,N_3067);
xor U6728 (N_6728,N_3296,N_3502);
nor U6729 (N_6729,N_3849,N_4346);
or U6730 (N_6730,N_4019,N_3112);
nand U6731 (N_6731,N_3441,N_4408);
and U6732 (N_6732,N_4972,N_2711);
xor U6733 (N_6733,N_2999,N_4919);
xor U6734 (N_6734,N_4662,N_4230);
and U6735 (N_6735,N_3717,N_4217);
and U6736 (N_6736,N_3558,N_2976);
xnor U6737 (N_6737,N_3637,N_3923);
nor U6738 (N_6738,N_2504,N_2967);
nand U6739 (N_6739,N_4422,N_4741);
or U6740 (N_6740,N_3310,N_3392);
nor U6741 (N_6741,N_4499,N_3755);
nand U6742 (N_6742,N_4425,N_4687);
nand U6743 (N_6743,N_4171,N_4455);
xnor U6744 (N_6744,N_4578,N_3511);
nor U6745 (N_6745,N_4246,N_3794);
nand U6746 (N_6746,N_3949,N_3383);
nor U6747 (N_6747,N_2860,N_3627);
or U6748 (N_6748,N_3724,N_4894);
and U6749 (N_6749,N_4399,N_4206);
and U6750 (N_6750,N_4693,N_3204);
or U6751 (N_6751,N_4032,N_3715);
xnor U6752 (N_6752,N_3782,N_2736);
or U6753 (N_6753,N_4444,N_3529);
and U6754 (N_6754,N_4814,N_4382);
or U6755 (N_6755,N_3480,N_2581);
xnor U6756 (N_6756,N_3994,N_3397);
nor U6757 (N_6757,N_3184,N_2844);
nor U6758 (N_6758,N_3876,N_4688);
or U6759 (N_6759,N_4372,N_4616);
xor U6760 (N_6760,N_4890,N_2680);
or U6761 (N_6761,N_3108,N_4503);
xor U6762 (N_6762,N_4303,N_3705);
xor U6763 (N_6763,N_4619,N_2899);
nand U6764 (N_6764,N_4531,N_4885);
or U6765 (N_6765,N_4640,N_4869);
nand U6766 (N_6766,N_2524,N_3893);
nor U6767 (N_6767,N_3025,N_3492);
xor U6768 (N_6768,N_3167,N_2776);
nand U6769 (N_6769,N_2909,N_4424);
nand U6770 (N_6770,N_3031,N_4033);
nor U6771 (N_6771,N_4084,N_3375);
and U6772 (N_6772,N_4511,N_4521);
or U6773 (N_6773,N_4307,N_3234);
xor U6774 (N_6774,N_4681,N_4553);
nor U6775 (N_6775,N_3026,N_3332);
xnor U6776 (N_6776,N_4807,N_4805);
nand U6777 (N_6777,N_4368,N_2896);
or U6778 (N_6778,N_4158,N_4605);
nor U6779 (N_6779,N_4539,N_2747);
nor U6780 (N_6780,N_4700,N_4766);
xor U6781 (N_6781,N_2908,N_4737);
nor U6782 (N_6782,N_3363,N_4880);
nor U6783 (N_6783,N_3981,N_4441);
nor U6784 (N_6784,N_4743,N_4150);
nand U6785 (N_6785,N_3843,N_3870);
nand U6786 (N_6786,N_2617,N_3567);
xor U6787 (N_6787,N_2696,N_4311);
and U6788 (N_6788,N_2999,N_2852);
nor U6789 (N_6789,N_2605,N_4785);
or U6790 (N_6790,N_3049,N_4597);
or U6791 (N_6791,N_3999,N_2644);
and U6792 (N_6792,N_4824,N_3772);
nand U6793 (N_6793,N_2595,N_4866);
nand U6794 (N_6794,N_3951,N_4578);
and U6795 (N_6795,N_2853,N_4689);
nand U6796 (N_6796,N_4630,N_2746);
or U6797 (N_6797,N_3048,N_4909);
nand U6798 (N_6798,N_2849,N_3639);
xor U6799 (N_6799,N_3215,N_4076);
or U6800 (N_6800,N_4291,N_4889);
xnor U6801 (N_6801,N_2862,N_3718);
xnor U6802 (N_6802,N_4706,N_4512);
or U6803 (N_6803,N_2730,N_3576);
nand U6804 (N_6804,N_3276,N_3900);
nand U6805 (N_6805,N_4325,N_4984);
xor U6806 (N_6806,N_3652,N_4601);
nor U6807 (N_6807,N_4021,N_4094);
nor U6808 (N_6808,N_2628,N_3197);
or U6809 (N_6809,N_2552,N_3750);
nand U6810 (N_6810,N_3133,N_4861);
nor U6811 (N_6811,N_3805,N_2938);
nand U6812 (N_6812,N_4104,N_3609);
xnor U6813 (N_6813,N_4024,N_3555);
nor U6814 (N_6814,N_3490,N_3253);
xnor U6815 (N_6815,N_4516,N_3751);
and U6816 (N_6816,N_4283,N_4123);
or U6817 (N_6817,N_2792,N_4016);
nor U6818 (N_6818,N_3853,N_4057);
nor U6819 (N_6819,N_3118,N_3822);
nand U6820 (N_6820,N_3510,N_3860);
nor U6821 (N_6821,N_2739,N_3114);
nand U6822 (N_6822,N_4078,N_2517);
or U6823 (N_6823,N_4589,N_2654);
or U6824 (N_6824,N_3925,N_4416);
or U6825 (N_6825,N_3056,N_3332);
xnor U6826 (N_6826,N_4781,N_3936);
nand U6827 (N_6827,N_2761,N_2973);
and U6828 (N_6828,N_2560,N_3010);
nand U6829 (N_6829,N_4652,N_4051);
xor U6830 (N_6830,N_3994,N_3592);
and U6831 (N_6831,N_3224,N_4445);
and U6832 (N_6832,N_3458,N_2783);
and U6833 (N_6833,N_3631,N_3572);
or U6834 (N_6834,N_3599,N_4101);
xor U6835 (N_6835,N_4063,N_2734);
xnor U6836 (N_6836,N_4578,N_4646);
xor U6837 (N_6837,N_2861,N_3844);
xnor U6838 (N_6838,N_4916,N_4892);
and U6839 (N_6839,N_4261,N_3087);
or U6840 (N_6840,N_3972,N_3876);
xnor U6841 (N_6841,N_3698,N_4592);
nor U6842 (N_6842,N_3736,N_4001);
or U6843 (N_6843,N_4751,N_3977);
xnor U6844 (N_6844,N_3865,N_2792);
and U6845 (N_6845,N_3580,N_2551);
nand U6846 (N_6846,N_4138,N_3913);
xnor U6847 (N_6847,N_3658,N_3064);
or U6848 (N_6848,N_2669,N_3117);
nand U6849 (N_6849,N_3991,N_4754);
and U6850 (N_6850,N_3010,N_3836);
nor U6851 (N_6851,N_4222,N_2589);
or U6852 (N_6852,N_4326,N_2759);
nand U6853 (N_6853,N_4699,N_3001);
xnor U6854 (N_6854,N_2942,N_3549);
nand U6855 (N_6855,N_3069,N_3417);
xor U6856 (N_6856,N_2799,N_4492);
xor U6857 (N_6857,N_4795,N_3859);
nor U6858 (N_6858,N_2566,N_3037);
nand U6859 (N_6859,N_3706,N_2937);
nand U6860 (N_6860,N_3109,N_2692);
xnor U6861 (N_6861,N_2874,N_3053);
nand U6862 (N_6862,N_4877,N_3364);
or U6863 (N_6863,N_4191,N_3436);
nor U6864 (N_6864,N_3270,N_4514);
or U6865 (N_6865,N_4855,N_4153);
nand U6866 (N_6866,N_3799,N_4778);
nand U6867 (N_6867,N_3410,N_4004);
nand U6868 (N_6868,N_4645,N_3085);
nand U6869 (N_6869,N_2765,N_2635);
nor U6870 (N_6870,N_4926,N_3334);
and U6871 (N_6871,N_3072,N_4630);
and U6872 (N_6872,N_4348,N_3211);
nand U6873 (N_6873,N_4793,N_3461);
or U6874 (N_6874,N_4129,N_4524);
nor U6875 (N_6875,N_4815,N_3951);
xnor U6876 (N_6876,N_2897,N_2813);
nand U6877 (N_6877,N_4487,N_4390);
nor U6878 (N_6878,N_4680,N_3931);
and U6879 (N_6879,N_3836,N_3938);
nor U6880 (N_6880,N_4111,N_2804);
and U6881 (N_6881,N_3599,N_4974);
and U6882 (N_6882,N_4529,N_2960);
nand U6883 (N_6883,N_3393,N_4825);
nand U6884 (N_6884,N_3520,N_4092);
xor U6885 (N_6885,N_3252,N_3012);
xnor U6886 (N_6886,N_4357,N_4490);
or U6887 (N_6887,N_2988,N_4233);
nand U6888 (N_6888,N_2601,N_4158);
nand U6889 (N_6889,N_2746,N_3068);
nand U6890 (N_6890,N_4513,N_4587);
xnor U6891 (N_6891,N_3863,N_2648);
xnor U6892 (N_6892,N_3505,N_2909);
nor U6893 (N_6893,N_2574,N_3991);
or U6894 (N_6894,N_2535,N_4767);
xnor U6895 (N_6895,N_3015,N_3614);
nor U6896 (N_6896,N_3211,N_2570);
xnor U6897 (N_6897,N_2662,N_2845);
nand U6898 (N_6898,N_2867,N_4092);
or U6899 (N_6899,N_3964,N_2537);
or U6900 (N_6900,N_3654,N_3607);
xnor U6901 (N_6901,N_3612,N_4461);
nand U6902 (N_6902,N_3421,N_4988);
nor U6903 (N_6903,N_4835,N_4614);
xnor U6904 (N_6904,N_3739,N_4824);
xor U6905 (N_6905,N_2907,N_4921);
and U6906 (N_6906,N_2705,N_2557);
and U6907 (N_6907,N_3299,N_4991);
nand U6908 (N_6908,N_4467,N_2699);
xnor U6909 (N_6909,N_2626,N_3250);
nor U6910 (N_6910,N_2736,N_4226);
xnor U6911 (N_6911,N_4260,N_4071);
nor U6912 (N_6912,N_4294,N_4833);
xor U6913 (N_6913,N_3898,N_2555);
or U6914 (N_6914,N_4881,N_3888);
xor U6915 (N_6915,N_2955,N_3404);
nand U6916 (N_6916,N_4061,N_4210);
and U6917 (N_6917,N_3076,N_4169);
xor U6918 (N_6918,N_4922,N_2873);
nand U6919 (N_6919,N_4487,N_2768);
nor U6920 (N_6920,N_4057,N_4885);
and U6921 (N_6921,N_2868,N_3974);
xnor U6922 (N_6922,N_4437,N_3652);
nand U6923 (N_6923,N_2560,N_4929);
xnor U6924 (N_6924,N_2852,N_4777);
nand U6925 (N_6925,N_2840,N_3694);
nand U6926 (N_6926,N_2858,N_2676);
and U6927 (N_6927,N_2648,N_3068);
nand U6928 (N_6928,N_2620,N_3069);
and U6929 (N_6929,N_2868,N_4975);
and U6930 (N_6930,N_3432,N_4201);
and U6931 (N_6931,N_3869,N_3926);
nand U6932 (N_6932,N_3652,N_3834);
nor U6933 (N_6933,N_3808,N_3574);
nand U6934 (N_6934,N_3047,N_4795);
or U6935 (N_6935,N_2789,N_3725);
or U6936 (N_6936,N_4666,N_4229);
nand U6937 (N_6937,N_4588,N_4391);
or U6938 (N_6938,N_3548,N_3455);
and U6939 (N_6939,N_4057,N_4648);
nand U6940 (N_6940,N_4528,N_3928);
nand U6941 (N_6941,N_2986,N_4444);
xor U6942 (N_6942,N_2865,N_3727);
nor U6943 (N_6943,N_3138,N_4986);
nor U6944 (N_6944,N_4356,N_2565);
or U6945 (N_6945,N_3347,N_3129);
or U6946 (N_6946,N_4368,N_3853);
xnor U6947 (N_6947,N_2570,N_4062);
or U6948 (N_6948,N_4526,N_4754);
nand U6949 (N_6949,N_4424,N_3150);
or U6950 (N_6950,N_2984,N_3100);
xnor U6951 (N_6951,N_3802,N_3037);
xnor U6952 (N_6952,N_4982,N_3757);
and U6953 (N_6953,N_4259,N_4897);
and U6954 (N_6954,N_4725,N_4080);
xnor U6955 (N_6955,N_4881,N_3703);
nor U6956 (N_6956,N_3693,N_3157);
nand U6957 (N_6957,N_4445,N_4559);
nand U6958 (N_6958,N_2685,N_2701);
nand U6959 (N_6959,N_3639,N_4621);
or U6960 (N_6960,N_3594,N_2947);
nor U6961 (N_6961,N_2813,N_3312);
xnor U6962 (N_6962,N_3169,N_3578);
nor U6963 (N_6963,N_2831,N_4110);
and U6964 (N_6964,N_3407,N_3784);
xnor U6965 (N_6965,N_2707,N_3782);
and U6966 (N_6966,N_3080,N_2983);
or U6967 (N_6967,N_4951,N_4863);
xor U6968 (N_6968,N_3999,N_2605);
xor U6969 (N_6969,N_3184,N_4684);
xnor U6970 (N_6970,N_3337,N_3080);
nand U6971 (N_6971,N_3367,N_2828);
or U6972 (N_6972,N_2945,N_4607);
and U6973 (N_6973,N_3439,N_3307);
nand U6974 (N_6974,N_4471,N_3735);
nand U6975 (N_6975,N_2868,N_2770);
nand U6976 (N_6976,N_2934,N_4447);
and U6977 (N_6977,N_2854,N_4287);
nor U6978 (N_6978,N_4808,N_3333);
and U6979 (N_6979,N_4362,N_2811);
nor U6980 (N_6980,N_4648,N_2651);
nand U6981 (N_6981,N_4601,N_3103);
xnor U6982 (N_6982,N_4978,N_4294);
nand U6983 (N_6983,N_3637,N_4152);
and U6984 (N_6984,N_4863,N_4123);
xor U6985 (N_6985,N_2871,N_2806);
or U6986 (N_6986,N_2834,N_3762);
nand U6987 (N_6987,N_3837,N_2505);
nand U6988 (N_6988,N_4993,N_3519);
or U6989 (N_6989,N_4739,N_3192);
nand U6990 (N_6990,N_4540,N_2525);
xnor U6991 (N_6991,N_4129,N_4762);
nor U6992 (N_6992,N_4792,N_2914);
and U6993 (N_6993,N_2521,N_4597);
or U6994 (N_6994,N_3984,N_3482);
nand U6995 (N_6995,N_2655,N_2649);
nor U6996 (N_6996,N_3476,N_4567);
and U6997 (N_6997,N_4645,N_2510);
and U6998 (N_6998,N_3954,N_4867);
xor U6999 (N_6999,N_3705,N_3255);
or U7000 (N_7000,N_4259,N_4089);
nand U7001 (N_7001,N_3815,N_2502);
or U7002 (N_7002,N_3623,N_2803);
or U7003 (N_7003,N_3279,N_3790);
nor U7004 (N_7004,N_4844,N_2781);
nor U7005 (N_7005,N_4863,N_4987);
and U7006 (N_7006,N_3456,N_3294);
nand U7007 (N_7007,N_4618,N_3927);
xnor U7008 (N_7008,N_2878,N_3169);
nor U7009 (N_7009,N_3685,N_4186);
nor U7010 (N_7010,N_3749,N_4053);
nor U7011 (N_7011,N_4107,N_2551);
or U7012 (N_7012,N_3970,N_3725);
nand U7013 (N_7013,N_3107,N_2842);
or U7014 (N_7014,N_3423,N_4285);
or U7015 (N_7015,N_3284,N_3538);
and U7016 (N_7016,N_3831,N_2608);
nor U7017 (N_7017,N_4031,N_3808);
or U7018 (N_7018,N_4274,N_3225);
nor U7019 (N_7019,N_4757,N_3953);
nor U7020 (N_7020,N_3075,N_3444);
or U7021 (N_7021,N_4831,N_4948);
xnor U7022 (N_7022,N_3850,N_3707);
and U7023 (N_7023,N_3269,N_3198);
nand U7024 (N_7024,N_3768,N_2877);
nor U7025 (N_7025,N_4764,N_3606);
xnor U7026 (N_7026,N_3466,N_3473);
xor U7027 (N_7027,N_3424,N_2928);
xor U7028 (N_7028,N_2832,N_4835);
nor U7029 (N_7029,N_4837,N_4133);
nor U7030 (N_7030,N_4251,N_4741);
nor U7031 (N_7031,N_3866,N_4543);
nand U7032 (N_7032,N_4750,N_4754);
or U7033 (N_7033,N_4643,N_2763);
nand U7034 (N_7034,N_4153,N_4440);
or U7035 (N_7035,N_3969,N_4372);
xor U7036 (N_7036,N_3283,N_3120);
nor U7037 (N_7037,N_4755,N_4996);
or U7038 (N_7038,N_3003,N_4293);
nor U7039 (N_7039,N_3092,N_3472);
nand U7040 (N_7040,N_4258,N_2838);
nand U7041 (N_7041,N_3722,N_3430);
nand U7042 (N_7042,N_2786,N_4851);
nand U7043 (N_7043,N_3935,N_4368);
and U7044 (N_7044,N_4541,N_3126);
xnor U7045 (N_7045,N_3408,N_3503);
nor U7046 (N_7046,N_4430,N_4989);
xnor U7047 (N_7047,N_3164,N_3981);
or U7048 (N_7048,N_3570,N_3490);
nor U7049 (N_7049,N_3509,N_2776);
or U7050 (N_7050,N_2587,N_3491);
xor U7051 (N_7051,N_4053,N_4035);
nor U7052 (N_7052,N_3911,N_4546);
nand U7053 (N_7053,N_3445,N_3508);
or U7054 (N_7054,N_3382,N_3205);
nor U7055 (N_7055,N_4171,N_3682);
or U7056 (N_7056,N_4667,N_4161);
or U7057 (N_7057,N_2998,N_4871);
or U7058 (N_7058,N_4055,N_2742);
nor U7059 (N_7059,N_4836,N_4951);
xor U7060 (N_7060,N_4200,N_3752);
or U7061 (N_7061,N_3095,N_4750);
xnor U7062 (N_7062,N_3877,N_4013);
nand U7063 (N_7063,N_2766,N_3905);
xor U7064 (N_7064,N_4354,N_3735);
and U7065 (N_7065,N_3696,N_2868);
and U7066 (N_7066,N_3048,N_4096);
xnor U7067 (N_7067,N_4619,N_3097);
xor U7068 (N_7068,N_3883,N_2820);
or U7069 (N_7069,N_4393,N_4963);
xnor U7070 (N_7070,N_3219,N_2639);
and U7071 (N_7071,N_4863,N_3465);
nor U7072 (N_7072,N_4019,N_2877);
nand U7073 (N_7073,N_2947,N_3143);
nor U7074 (N_7074,N_4196,N_4927);
xor U7075 (N_7075,N_4146,N_2608);
and U7076 (N_7076,N_3169,N_3624);
or U7077 (N_7077,N_4364,N_4972);
and U7078 (N_7078,N_3324,N_3884);
xor U7079 (N_7079,N_3341,N_2940);
nand U7080 (N_7080,N_4627,N_3719);
and U7081 (N_7081,N_4183,N_4449);
xnor U7082 (N_7082,N_3222,N_3684);
nor U7083 (N_7083,N_3312,N_2730);
xnor U7084 (N_7084,N_4767,N_4273);
nor U7085 (N_7085,N_3196,N_4678);
nand U7086 (N_7086,N_3867,N_2550);
xor U7087 (N_7087,N_4962,N_4125);
nor U7088 (N_7088,N_4609,N_3728);
xnor U7089 (N_7089,N_4043,N_4374);
or U7090 (N_7090,N_4099,N_4634);
and U7091 (N_7091,N_3243,N_3522);
and U7092 (N_7092,N_3350,N_3818);
nor U7093 (N_7093,N_4979,N_3994);
and U7094 (N_7094,N_4597,N_4999);
or U7095 (N_7095,N_3362,N_3441);
xnor U7096 (N_7096,N_3015,N_4627);
or U7097 (N_7097,N_3021,N_4835);
nor U7098 (N_7098,N_4823,N_3615);
nand U7099 (N_7099,N_2593,N_3219);
and U7100 (N_7100,N_3422,N_4491);
nor U7101 (N_7101,N_3427,N_3254);
or U7102 (N_7102,N_4341,N_3089);
nand U7103 (N_7103,N_3011,N_3268);
xnor U7104 (N_7104,N_4089,N_4564);
or U7105 (N_7105,N_3329,N_3103);
or U7106 (N_7106,N_3531,N_3975);
or U7107 (N_7107,N_3941,N_2573);
and U7108 (N_7108,N_3603,N_4825);
xnor U7109 (N_7109,N_3367,N_2541);
or U7110 (N_7110,N_4244,N_4049);
or U7111 (N_7111,N_3371,N_2720);
xor U7112 (N_7112,N_3480,N_2629);
nand U7113 (N_7113,N_3865,N_4429);
or U7114 (N_7114,N_4900,N_4270);
nand U7115 (N_7115,N_4719,N_3990);
nand U7116 (N_7116,N_3856,N_4445);
and U7117 (N_7117,N_4065,N_2738);
nand U7118 (N_7118,N_2844,N_4565);
nand U7119 (N_7119,N_4653,N_3498);
or U7120 (N_7120,N_3749,N_2863);
nand U7121 (N_7121,N_3752,N_4018);
or U7122 (N_7122,N_3919,N_4047);
xnor U7123 (N_7123,N_4597,N_3217);
and U7124 (N_7124,N_3538,N_3483);
or U7125 (N_7125,N_3424,N_4736);
and U7126 (N_7126,N_3382,N_4455);
xor U7127 (N_7127,N_3752,N_3471);
or U7128 (N_7128,N_4243,N_3985);
or U7129 (N_7129,N_3280,N_3676);
xor U7130 (N_7130,N_2725,N_2722);
or U7131 (N_7131,N_2567,N_2583);
and U7132 (N_7132,N_4087,N_3028);
or U7133 (N_7133,N_4603,N_4829);
and U7134 (N_7134,N_2988,N_4157);
and U7135 (N_7135,N_2598,N_3550);
nand U7136 (N_7136,N_2834,N_3741);
nand U7137 (N_7137,N_3119,N_4868);
nor U7138 (N_7138,N_4170,N_2667);
or U7139 (N_7139,N_3312,N_3004);
or U7140 (N_7140,N_2873,N_2540);
xnor U7141 (N_7141,N_2621,N_4275);
nor U7142 (N_7142,N_2892,N_4575);
and U7143 (N_7143,N_4583,N_4031);
nor U7144 (N_7144,N_3270,N_4580);
nor U7145 (N_7145,N_2667,N_2754);
nor U7146 (N_7146,N_4729,N_2918);
xor U7147 (N_7147,N_2814,N_4452);
or U7148 (N_7148,N_4149,N_4165);
and U7149 (N_7149,N_3316,N_4995);
or U7150 (N_7150,N_3281,N_4645);
or U7151 (N_7151,N_4108,N_3249);
or U7152 (N_7152,N_4957,N_3273);
nand U7153 (N_7153,N_4307,N_3092);
xnor U7154 (N_7154,N_4656,N_3585);
xnor U7155 (N_7155,N_3648,N_2557);
or U7156 (N_7156,N_3992,N_3259);
nor U7157 (N_7157,N_3101,N_4961);
or U7158 (N_7158,N_4226,N_2584);
or U7159 (N_7159,N_3582,N_2831);
xnor U7160 (N_7160,N_3840,N_3982);
or U7161 (N_7161,N_3024,N_3279);
xnor U7162 (N_7162,N_2766,N_2575);
nand U7163 (N_7163,N_3938,N_2645);
nand U7164 (N_7164,N_3201,N_3367);
or U7165 (N_7165,N_4253,N_4606);
xor U7166 (N_7166,N_3050,N_3840);
nor U7167 (N_7167,N_2652,N_2895);
nor U7168 (N_7168,N_3697,N_4587);
and U7169 (N_7169,N_3611,N_2726);
nor U7170 (N_7170,N_2996,N_2705);
xor U7171 (N_7171,N_3115,N_2968);
nand U7172 (N_7172,N_3678,N_4212);
nand U7173 (N_7173,N_4649,N_3687);
nand U7174 (N_7174,N_3254,N_2766);
nand U7175 (N_7175,N_4158,N_3740);
xor U7176 (N_7176,N_2687,N_4843);
and U7177 (N_7177,N_3242,N_3675);
or U7178 (N_7178,N_2934,N_2572);
xor U7179 (N_7179,N_4959,N_2590);
or U7180 (N_7180,N_2718,N_3705);
nand U7181 (N_7181,N_4500,N_3141);
or U7182 (N_7182,N_4579,N_4239);
nor U7183 (N_7183,N_3202,N_2585);
or U7184 (N_7184,N_2604,N_2594);
nor U7185 (N_7185,N_2544,N_3806);
and U7186 (N_7186,N_3688,N_3910);
and U7187 (N_7187,N_3233,N_4129);
xnor U7188 (N_7188,N_3928,N_4634);
xnor U7189 (N_7189,N_3859,N_2833);
nor U7190 (N_7190,N_3625,N_2909);
nor U7191 (N_7191,N_4049,N_3138);
nor U7192 (N_7192,N_3629,N_4214);
nand U7193 (N_7193,N_2613,N_3311);
nand U7194 (N_7194,N_4666,N_4808);
or U7195 (N_7195,N_2642,N_4469);
or U7196 (N_7196,N_4661,N_4080);
nor U7197 (N_7197,N_4387,N_3776);
nor U7198 (N_7198,N_4773,N_3162);
and U7199 (N_7199,N_2621,N_2856);
nand U7200 (N_7200,N_2750,N_3798);
xnor U7201 (N_7201,N_3900,N_4521);
nand U7202 (N_7202,N_4181,N_3983);
or U7203 (N_7203,N_4405,N_3436);
xor U7204 (N_7204,N_4209,N_2580);
nor U7205 (N_7205,N_2529,N_4103);
nand U7206 (N_7206,N_4514,N_3502);
nor U7207 (N_7207,N_4439,N_2773);
nand U7208 (N_7208,N_3573,N_3504);
nor U7209 (N_7209,N_2567,N_3987);
xor U7210 (N_7210,N_3644,N_3126);
and U7211 (N_7211,N_2688,N_3152);
nor U7212 (N_7212,N_4386,N_2601);
and U7213 (N_7213,N_4765,N_2671);
and U7214 (N_7214,N_3018,N_4557);
xor U7215 (N_7215,N_4923,N_4074);
xor U7216 (N_7216,N_4599,N_3654);
xor U7217 (N_7217,N_3134,N_3697);
xnor U7218 (N_7218,N_3190,N_3217);
nor U7219 (N_7219,N_4929,N_2928);
xnor U7220 (N_7220,N_4659,N_3860);
or U7221 (N_7221,N_3013,N_4556);
nand U7222 (N_7222,N_3800,N_2966);
or U7223 (N_7223,N_3883,N_3130);
nor U7224 (N_7224,N_4913,N_2622);
nand U7225 (N_7225,N_3824,N_3565);
nand U7226 (N_7226,N_3414,N_2720);
nor U7227 (N_7227,N_4595,N_3266);
and U7228 (N_7228,N_4642,N_4598);
or U7229 (N_7229,N_4423,N_3215);
xnor U7230 (N_7230,N_3578,N_4804);
nor U7231 (N_7231,N_2773,N_2991);
and U7232 (N_7232,N_2573,N_4987);
nor U7233 (N_7233,N_4861,N_2658);
nor U7234 (N_7234,N_4362,N_3621);
xor U7235 (N_7235,N_3197,N_3590);
nor U7236 (N_7236,N_4110,N_2913);
and U7237 (N_7237,N_3749,N_2758);
or U7238 (N_7238,N_3237,N_3795);
and U7239 (N_7239,N_4503,N_2505);
and U7240 (N_7240,N_4239,N_3215);
and U7241 (N_7241,N_2737,N_3738);
nor U7242 (N_7242,N_2700,N_4773);
nand U7243 (N_7243,N_2596,N_2956);
or U7244 (N_7244,N_3660,N_3322);
nor U7245 (N_7245,N_3676,N_4194);
or U7246 (N_7246,N_4150,N_3505);
nor U7247 (N_7247,N_3442,N_3918);
xor U7248 (N_7248,N_4224,N_3597);
nor U7249 (N_7249,N_4392,N_4814);
and U7250 (N_7250,N_3591,N_4693);
and U7251 (N_7251,N_4235,N_4634);
or U7252 (N_7252,N_4794,N_4089);
nand U7253 (N_7253,N_4041,N_3800);
xor U7254 (N_7254,N_2560,N_3349);
nand U7255 (N_7255,N_4331,N_2800);
and U7256 (N_7256,N_2933,N_3155);
and U7257 (N_7257,N_4225,N_3524);
and U7258 (N_7258,N_2858,N_3613);
or U7259 (N_7259,N_3780,N_3785);
xnor U7260 (N_7260,N_3412,N_3415);
nand U7261 (N_7261,N_4850,N_3462);
xor U7262 (N_7262,N_4467,N_3937);
xnor U7263 (N_7263,N_2521,N_2570);
nand U7264 (N_7264,N_2568,N_4462);
or U7265 (N_7265,N_3871,N_3165);
xnor U7266 (N_7266,N_4061,N_2556);
nor U7267 (N_7267,N_4262,N_3388);
nor U7268 (N_7268,N_4832,N_3428);
nand U7269 (N_7269,N_2821,N_2725);
or U7270 (N_7270,N_3371,N_4061);
nand U7271 (N_7271,N_2777,N_4636);
nor U7272 (N_7272,N_4503,N_4549);
xnor U7273 (N_7273,N_4526,N_4260);
xor U7274 (N_7274,N_3314,N_3741);
nor U7275 (N_7275,N_3925,N_4818);
xnor U7276 (N_7276,N_4048,N_2784);
or U7277 (N_7277,N_4360,N_3582);
nor U7278 (N_7278,N_3104,N_4828);
xor U7279 (N_7279,N_2514,N_4342);
nand U7280 (N_7280,N_4758,N_3081);
nor U7281 (N_7281,N_4590,N_2820);
xnor U7282 (N_7282,N_4841,N_4005);
or U7283 (N_7283,N_4729,N_4478);
and U7284 (N_7284,N_2591,N_4369);
nor U7285 (N_7285,N_3594,N_3872);
and U7286 (N_7286,N_3915,N_2901);
xor U7287 (N_7287,N_3589,N_2841);
xnor U7288 (N_7288,N_3822,N_3959);
nor U7289 (N_7289,N_3847,N_4872);
or U7290 (N_7290,N_3203,N_3071);
xnor U7291 (N_7291,N_4301,N_3434);
nand U7292 (N_7292,N_3127,N_3919);
and U7293 (N_7293,N_4443,N_4376);
and U7294 (N_7294,N_4579,N_3687);
nand U7295 (N_7295,N_4683,N_4184);
or U7296 (N_7296,N_3097,N_3746);
and U7297 (N_7297,N_4017,N_3781);
xor U7298 (N_7298,N_4408,N_2732);
xnor U7299 (N_7299,N_2608,N_3013);
nor U7300 (N_7300,N_3925,N_3157);
xor U7301 (N_7301,N_4252,N_4690);
nand U7302 (N_7302,N_3289,N_3624);
or U7303 (N_7303,N_3604,N_3835);
or U7304 (N_7304,N_2569,N_4554);
or U7305 (N_7305,N_4269,N_3485);
or U7306 (N_7306,N_4777,N_4507);
and U7307 (N_7307,N_2882,N_4367);
nand U7308 (N_7308,N_4844,N_3713);
nor U7309 (N_7309,N_2560,N_3695);
and U7310 (N_7310,N_3259,N_4428);
nor U7311 (N_7311,N_3454,N_4727);
and U7312 (N_7312,N_3886,N_2944);
nand U7313 (N_7313,N_4199,N_3538);
nor U7314 (N_7314,N_2955,N_3394);
xor U7315 (N_7315,N_3168,N_3137);
xor U7316 (N_7316,N_4699,N_2555);
nand U7317 (N_7317,N_2695,N_3741);
or U7318 (N_7318,N_3513,N_3868);
nor U7319 (N_7319,N_4689,N_2646);
nor U7320 (N_7320,N_2595,N_3023);
or U7321 (N_7321,N_3162,N_3530);
and U7322 (N_7322,N_4405,N_4389);
or U7323 (N_7323,N_3836,N_4300);
nor U7324 (N_7324,N_3836,N_2846);
xor U7325 (N_7325,N_3469,N_2587);
or U7326 (N_7326,N_4759,N_4716);
or U7327 (N_7327,N_4808,N_3990);
xor U7328 (N_7328,N_3594,N_4858);
nor U7329 (N_7329,N_3319,N_4328);
nor U7330 (N_7330,N_3858,N_3050);
nand U7331 (N_7331,N_4011,N_4017);
or U7332 (N_7332,N_4148,N_3524);
xnor U7333 (N_7333,N_4323,N_3726);
or U7334 (N_7334,N_2851,N_3015);
or U7335 (N_7335,N_3301,N_3185);
xnor U7336 (N_7336,N_4696,N_4319);
nor U7337 (N_7337,N_3773,N_3162);
and U7338 (N_7338,N_4278,N_3959);
xor U7339 (N_7339,N_2862,N_2572);
and U7340 (N_7340,N_3113,N_3214);
or U7341 (N_7341,N_2954,N_3137);
and U7342 (N_7342,N_2982,N_4216);
nor U7343 (N_7343,N_3206,N_4301);
or U7344 (N_7344,N_4879,N_3096);
or U7345 (N_7345,N_3091,N_4701);
xnor U7346 (N_7346,N_4702,N_2592);
and U7347 (N_7347,N_4178,N_4182);
nand U7348 (N_7348,N_2912,N_3660);
or U7349 (N_7349,N_3197,N_3339);
nor U7350 (N_7350,N_3323,N_3260);
nand U7351 (N_7351,N_3485,N_4986);
or U7352 (N_7352,N_3491,N_3489);
nand U7353 (N_7353,N_4540,N_4477);
or U7354 (N_7354,N_4496,N_3560);
xor U7355 (N_7355,N_4965,N_2964);
or U7356 (N_7356,N_4805,N_4065);
nand U7357 (N_7357,N_3343,N_4347);
xor U7358 (N_7358,N_3088,N_3666);
nand U7359 (N_7359,N_4866,N_4734);
xnor U7360 (N_7360,N_3646,N_3882);
xnor U7361 (N_7361,N_4894,N_4490);
and U7362 (N_7362,N_3983,N_3156);
and U7363 (N_7363,N_3940,N_4267);
nor U7364 (N_7364,N_3456,N_4618);
and U7365 (N_7365,N_4873,N_3068);
and U7366 (N_7366,N_4290,N_3253);
and U7367 (N_7367,N_2864,N_3404);
nor U7368 (N_7368,N_4994,N_3608);
nor U7369 (N_7369,N_3239,N_3753);
nand U7370 (N_7370,N_4795,N_3779);
nand U7371 (N_7371,N_2952,N_3991);
and U7372 (N_7372,N_3547,N_2707);
nand U7373 (N_7373,N_4221,N_2835);
or U7374 (N_7374,N_3915,N_4464);
nor U7375 (N_7375,N_3583,N_2847);
xnor U7376 (N_7376,N_3249,N_3396);
or U7377 (N_7377,N_2981,N_3268);
and U7378 (N_7378,N_3236,N_3165);
and U7379 (N_7379,N_4281,N_3855);
and U7380 (N_7380,N_4489,N_3369);
nor U7381 (N_7381,N_3864,N_4337);
nor U7382 (N_7382,N_2550,N_3314);
or U7383 (N_7383,N_4671,N_4559);
and U7384 (N_7384,N_4578,N_4770);
xnor U7385 (N_7385,N_3074,N_4539);
xor U7386 (N_7386,N_2544,N_2849);
nor U7387 (N_7387,N_3885,N_4881);
or U7388 (N_7388,N_4725,N_3616);
nand U7389 (N_7389,N_3924,N_2803);
xnor U7390 (N_7390,N_4214,N_3730);
nor U7391 (N_7391,N_3676,N_3886);
xor U7392 (N_7392,N_4610,N_3901);
nor U7393 (N_7393,N_4930,N_3196);
or U7394 (N_7394,N_2985,N_2736);
xor U7395 (N_7395,N_2732,N_2858);
xnor U7396 (N_7396,N_4865,N_4104);
nor U7397 (N_7397,N_2876,N_4245);
and U7398 (N_7398,N_4579,N_4646);
nand U7399 (N_7399,N_4015,N_4710);
and U7400 (N_7400,N_4347,N_3893);
or U7401 (N_7401,N_4961,N_2609);
nor U7402 (N_7402,N_4206,N_3933);
nand U7403 (N_7403,N_3123,N_3296);
xnor U7404 (N_7404,N_4558,N_4666);
or U7405 (N_7405,N_2732,N_4498);
and U7406 (N_7406,N_3854,N_4998);
xor U7407 (N_7407,N_2619,N_2630);
and U7408 (N_7408,N_2753,N_4017);
xor U7409 (N_7409,N_4786,N_4327);
or U7410 (N_7410,N_2636,N_2717);
nand U7411 (N_7411,N_4596,N_4504);
nor U7412 (N_7412,N_4227,N_3229);
or U7413 (N_7413,N_4347,N_4927);
or U7414 (N_7414,N_3878,N_4519);
and U7415 (N_7415,N_4252,N_3567);
nand U7416 (N_7416,N_2922,N_4351);
or U7417 (N_7417,N_3091,N_4782);
or U7418 (N_7418,N_3119,N_3743);
xnor U7419 (N_7419,N_2805,N_4289);
nand U7420 (N_7420,N_3763,N_3514);
or U7421 (N_7421,N_3191,N_3477);
nand U7422 (N_7422,N_3398,N_3900);
nor U7423 (N_7423,N_2566,N_3391);
xnor U7424 (N_7424,N_3691,N_2899);
or U7425 (N_7425,N_4899,N_3831);
xnor U7426 (N_7426,N_4748,N_4822);
nor U7427 (N_7427,N_3364,N_2887);
xnor U7428 (N_7428,N_4242,N_4312);
or U7429 (N_7429,N_4648,N_4192);
nor U7430 (N_7430,N_2808,N_2800);
and U7431 (N_7431,N_3598,N_3412);
nor U7432 (N_7432,N_3677,N_4028);
or U7433 (N_7433,N_3319,N_4348);
or U7434 (N_7434,N_2598,N_3960);
or U7435 (N_7435,N_3179,N_3952);
xnor U7436 (N_7436,N_2550,N_3282);
or U7437 (N_7437,N_3573,N_3149);
or U7438 (N_7438,N_3508,N_3855);
nand U7439 (N_7439,N_2824,N_2574);
and U7440 (N_7440,N_2579,N_4669);
and U7441 (N_7441,N_3626,N_3533);
xnor U7442 (N_7442,N_4697,N_4482);
and U7443 (N_7443,N_4864,N_3383);
nor U7444 (N_7444,N_2630,N_4693);
or U7445 (N_7445,N_3181,N_4183);
or U7446 (N_7446,N_2613,N_4003);
nor U7447 (N_7447,N_4895,N_2759);
or U7448 (N_7448,N_4591,N_3382);
nor U7449 (N_7449,N_4231,N_4889);
xor U7450 (N_7450,N_2623,N_3598);
or U7451 (N_7451,N_2825,N_2883);
nor U7452 (N_7452,N_3851,N_2742);
nand U7453 (N_7453,N_4172,N_3706);
or U7454 (N_7454,N_4710,N_4464);
nand U7455 (N_7455,N_4756,N_3033);
nor U7456 (N_7456,N_2872,N_4100);
and U7457 (N_7457,N_3274,N_3174);
and U7458 (N_7458,N_3603,N_3862);
nand U7459 (N_7459,N_4155,N_2701);
and U7460 (N_7460,N_4487,N_4177);
and U7461 (N_7461,N_3390,N_3853);
and U7462 (N_7462,N_2644,N_3319);
or U7463 (N_7463,N_4874,N_4073);
and U7464 (N_7464,N_2758,N_3362);
or U7465 (N_7465,N_4357,N_2713);
and U7466 (N_7466,N_4717,N_3419);
nand U7467 (N_7467,N_3182,N_4015);
nor U7468 (N_7468,N_2807,N_4614);
or U7469 (N_7469,N_4524,N_4251);
nand U7470 (N_7470,N_2939,N_4027);
nor U7471 (N_7471,N_2527,N_4143);
or U7472 (N_7472,N_2596,N_4227);
and U7473 (N_7473,N_4897,N_2525);
xnor U7474 (N_7474,N_2681,N_3519);
nand U7475 (N_7475,N_3320,N_4333);
or U7476 (N_7476,N_3043,N_3762);
xnor U7477 (N_7477,N_4647,N_4244);
and U7478 (N_7478,N_4029,N_3513);
and U7479 (N_7479,N_3785,N_3103);
and U7480 (N_7480,N_3207,N_3005);
nor U7481 (N_7481,N_4955,N_2968);
and U7482 (N_7482,N_3159,N_2779);
and U7483 (N_7483,N_3901,N_2667);
or U7484 (N_7484,N_2898,N_4875);
nor U7485 (N_7485,N_4303,N_2996);
xor U7486 (N_7486,N_2684,N_2596);
or U7487 (N_7487,N_3538,N_4642);
nor U7488 (N_7488,N_4857,N_3793);
nor U7489 (N_7489,N_4047,N_4717);
nor U7490 (N_7490,N_3828,N_4930);
nand U7491 (N_7491,N_3757,N_4741);
and U7492 (N_7492,N_2757,N_4594);
or U7493 (N_7493,N_3726,N_3719);
or U7494 (N_7494,N_3298,N_2968);
or U7495 (N_7495,N_3583,N_2693);
or U7496 (N_7496,N_3950,N_3365);
and U7497 (N_7497,N_4745,N_2929);
or U7498 (N_7498,N_2704,N_4067);
and U7499 (N_7499,N_3923,N_4091);
xor U7500 (N_7500,N_6182,N_7082);
xnor U7501 (N_7501,N_6045,N_7481);
nand U7502 (N_7502,N_7342,N_5234);
nand U7503 (N_7503,N_7440,N_5746);
nand U7504 (N_7504,N_7244,N_6863);
nor U7505 (N_7505,N_6587,N_6386);
nand U7506 (N_7506,N_5687,N_5819);
nor U7507 (N_7507,N_7204,N_5487);
xor U7508 (N_7508,N_5760,N_6419);
nand U7509 (N_7509,N_6447,N_6212);
and U7510 (N_7510,N_5942,N_6731);
nor U7511 (N_7511,N_5464,N_6004);
nor U7512 (N_7512,N_6844,N_5765);
and U7513 (N_7513,N_6409,N_5008);
xnor U7514 (N_7514,N_6780,N_6924);
and U7515 (N_7515,N_6822,N_6125);
nor U7516 (N_7516,N_6883,N_6406);
nor U7517 (N_7517,N_5956,N_7181);
and U7518 (N_7518,N_7479,N_5501);
xor U7519 (N_7519,N_5770,N_5825);
xnor U7520 (N_7520,N_6410,N_5585);
or U7521 (N_7521,N_5118,N_7094);
or U7522 (N_7522,N_7049,N_7031);
nand U7523 (N_7523,N_5712,N_6626);
xor U7524 (N_7524,N_5223,N_6670);
or U7525 (N_7525,N_5399,N_6976);
nor U7526 (N_7526,N_5341,N_5104);
nand U7527 (N_7527,N_5214,N_5576);
or U7528 (N_7528,N_5451,N_5841);
nand U7529 (N_7529,N_5690,N_7421);
xor U7530 (N_7530,N_5333,N_6699);
or U7531 (N_7531,N_6355,N_6530);
nor U7532 (N_7532,N_7156,N_5862);
nor U7533 (N_7533,N_5930,N_6193);
and U7534 (N_7534,N_6224,N_5022);
or U7535 (N_7535,N_5338,N_6562);
nand U7536 (N_7536,N_6824,N_6818);
xnor U7537 (N_7537,N_6725,N_7086);
xnor U7538 (N_7538,N_6115,N_5351);
xnor U7539 (N_7539,N_6769,N_5416);
or U7540 (N_7540,N_6580,N_5482);
nor U7541 (N_7541,N_6717,N_6343);
nor U7542 (N_7542,N_5230,N_5850);
nor U7543 (N_7543,N_6013,N_6341);
nand U7544 (N_7544,N_6606,N_7363);
and U7545 (N_7545,N_5160,N_5443);
nor U7546 (N_7546,N_6990,N_6779);
xor U7547 (N_7547,N_6480,N_5721);
or U7548 (N_7548,N_7017,N_6254);
nor U7549 (N_7549,N_6302,N_7483);
or U7550 (N_7550,N_7229,N_7336);
xnor U7551 (N_7551,N_5190,N_5350);
and U7552 (N_7552,N_6886,N_5468);
or U7553 (N_7553,N_6711,N_5220);
xnor U7554 (N_7554,N_6881,N_7380);
nand U7555 (N_7555,N_6950,N_7476);
nor U7556 (N_7556,N_5218,N_5452);
nor U7557 (N_7557,N_6693,N_7404);
nand U7558 (N_7558,N_7489,N_6804);
xnor U7559 (N_7559,N_7217,N_6654);
nor U7560 (N_7560,N_6011,N_5096);
xnor U7561 (N_7561,N_6088,N_6984);
or U7562 (N_7562,N_7025,N_6887);
or U7563 (N_7563,N_6521,N_7293);
and U7564 (N_7564,N_6923,N_7304);
or U7565 (N_7565,N_6194,N_5724);
nand U7566 (N_7566,N_6590,N_6037);
and U7567 (N_7567,N_6897,N_6333);
and U7568 (N_7568,N_6032,N_6865);
nor U7569 (N_7569,N_7158,N_5592);
xor U7570 (N_7570,N_6700,N_5434);
xnor U7571 (N_7571,N_7376,N_7486);
or U7572 (N_7572,N_5682,N_5256);
nand U7573 (N_7573,N_5049,N_5442);
and U7574 (N_7574,N_6250,N_7493);
or U7575 (N_7575,N_6042,N_5678);
and U7576 (N_7576,N_5648,N_5984);
and U7577 (N_7577,N_5461,N_5433);
nand U7578 (N_7578,N_5507,N_7470);
and U7579 (N_7579,N_5463,N_6782);
or U7580 (N_7580,N_5853,N_6084);
and U7581 (N_7581,N_5974,N_6597);
xnor U7582 (N_7582,N_6891,N_5056);
or U7583 (N_7583,N_6370,N_7365);
nand U7584 (N_7584,N_6369,N_6953);
nor U7585 (N_7585,N_7182,N_5011);
and U7586 (N_7586,N_5559,N_6946);
nor U7587 (N_7587,N_6964,N_6970);
nand U7588 (N_7588,N_5939,N_6140);
and U7589 (N_7589,N_5345,N_6668);
nand U7590 (N_7590,N_6016,N_5334);
xnor U7591 (N_7591,N_7416,N_6272);
nand U7592 (N_7592,N_6335,N_5564);
xnor U7593 (N_7593,N_5880,N_7395);
nand U7594 (N_7594,N_5856,N_6726);
xor U7595 (N_7595,N_5315,N_7423);
xnor U7596 (N_7596,N_5567,N_6010);
nor U7597 (N_7597,N_6459,N_6526);
and U7598 (N_7598,N_5847,N_5739);
and U7599 (N_7599,N_5800,N_7409);
xor U7600 (N_7600,N_6702,N_7102);
and U7601 (N_7601,N_5221,N_7472);
xor U7602 (N_7602,N_7128,N_6623);
and U7603 (N_7603,N_5828,N_5549);
xor U7604 (N_7604,N_7157,N_6801);
or U7605 (N_7605,N_5167,N_6256);
or U7606 (N_7606,N_7055,N_6227);
xnor U7607 (N_7607,N_7253,N_7468);
and U7608 (N_7608,N_7324,N_6715);
nand U7609 (N_7609,N_6282,N_5976);
and U7610 (N_7610,N_5455,N_5275);
xor U7611 (N_7611,N_7311,N_7448);
nor U7612 (N_7612,N_6142,N_7482);
xnor U7613 (N_7613,N_5119,N_5578);
nor U7614 (N_7614,N_5055,N_6973);
nor U7615 (N_7615,N_6996,N_6301);
nand U7616 (N_7616,N_5405,N_6139);
xnor U7617 (N_7617,N_5863,N_7296);
nor U7618 (N_7618,N_7498,N_6729);
xnor U7619 (N_7619,N_7106,N_6705);
nand U7620 (N_7620,N_6443,N_5680);
xor U7621 (N_7621,N_7449,N_7381);
and U7622 (N_7622,N_6810,N_5077);
nand U7623 (N_7623,N_5208,N_7134);
nand U7624 (N_7624,N_5219,N_6709);
or U7625 (N_7625,N_6400,N_7133);
nand U7626 (N_7626,N_6754,N_6719);
xor U7627 (N_7627,N_7402,N_6251);
nand U7628 (N_7628,N_6422,N_5447);
or U7629 (N_7629,N_5868,N_5659);
and U7630 (N_7630,N_5824,N_6978);
or U7631 (N_7631,N_5728,N_7323);
nand U7632 (N_7632,N_5396,N_7183);
nand U7633 (N_7633,N_7178,N_7419);
or U7634 (N_7634,N_5618,N_7485);
nor U7635 (N_7635,N_5252,N_5432);
xor U7636 (N_7636,N_5222,N_7198);
xnor U7637 (N_7637,N_6491,N_5454);
or U7638 (N_7638,N_7054,N_6033);
xor U7639 (N_7639,N_6775,N_7499);
and U7640 (N_7640,N_6453,N_6299);
nor U7641 (N_7641,N_6330,N_5368);
and U7642 (N_7642,N_6920,N_5987);
or U7643 (N_7643,N_6947,N_6547);
nand U7644 (N_7644,N_7162,N_7463);
and U7645 (N_7645,N_5012,N_7043);
or U7646 (N_7646,N_5419,N_6306);
or U7647 (N_7647,N_6187,N_5854);
and U7648 (N_7648,N_6523,N_6470);
or U7649 (N_7649,N_7361,N_5748);
nor U7650 (N_7650,N_5059,N_7190);
nand U7651 (N_7651,N_5035,N_5000);
or U7652 (N_7652,N_5537,N_6936);
nor U7653 (N_7653,N_6956,N_7009);
and U7654 (N_7654,N_7452,N_6049);
or U7655 (N_7655,N_6092,N_6760);
or U7656 (N_7656,N_5099,N_5626);
nor U7657 (N_7657,N_6366,N_6701);
and U7658 (N_7658,N_6108,N_6211);
and U7659 (N_7659,N_6907,N_6872);
or U7660 (N_7660,N_5654,N_5964);
and U7661 (N_7661,N_7197,N_6681);
xor U7662 (N_7662,N_6979,N_5228);
xor U7663 (N_7663,N_5058,N_7491);
nor U7664 (N_7664,N_6359,N_7263);
nor U7665 (N_7665,N_6157,N_6235);
xnor U7666 (N_7666,N_6832,N_5371);
nor U7667 (N_7667,N_7005,N_5698);
nor U7668 (N_7668,N_5137,N_5028);
xnor U7669 (N_7669,N_5407,N_5440);
nor U7670 (N_7670,N_7427,N_6307);
and U7671 (N_7671,N_7152,N_5876);
xnor U7672 (N_7672,N_5356,N_5917);
nand U7673 (N_7673,N_6350,N_6089);
nand U7674 (N_7674,N_5362,N_5383);
or U7675 (N_7675,N_5882,N_6479);
and U7676 (N_7676,N_5753,N_5100);
nand U7677 (N_7677,N_6185,N_5267);
nand U7678 (N_7678,N_6908,N_6543);
nor U7679 (N_7679,N_6512,N_6389);
nand U7680 (N_7680,N_5354,N_7386);
xnor U7681 (N_7681,N_6146,N_6105);
or U7682 (N_7682,N_5312,N_5827);
xor U7683 (N_7683,N_7103,N_6721);
xnor U7684 (N_7684,N_5191,N_5823);
nor U7685 (N_7685,N_5706,N_7330);
nand U7686 (N_7686,N_7454,N_5936);
nor U7687 (N_7687,N_7292,N_6582);
xnor U7688 (N_7688,N_7131,N_6696);
or U7689 (N_7689,N_5384,N_5710);
xor U7690 (N_7690,N_6387,N_7033);
and U7691 (N_7691,N_6614,N_5397);
nand U7692 (N_7692,N_6348,N_5918);
nand U7693 (N_7693,N_6894,N_5558);
nand U7694 (N_7694,N_6163,N_5547);
and U7695 (N_7695,N_6794,N_6296);
and U7696 (N_7696,N_6091,N_6457);
nor U7697 (N_7697,N_5296,N_5241);
xor U7698 (N_7698,N_5750,N_6921);
or U7699 (N_7699,N_5701,N_6388);
nand U7700 (N_7700,N_5444,N_7159);
nor U7701 (N_7701,N_7412,N_5725);
xor U7702 (N_7702,N_6317,N_5877);
nor U7703 (N_7703,N_6879,N_6451);
and U7704 (N_7704,N_5611,N_7024);
and U7705 (N_7705,N_5971,N_7283);
nor U7706 (N_7706,N_5069,N_6893);
and U7707 (N_7707,N_6739,N_6075);
and U7708 (N_7708,N_7092,N_5121);
nand U7709 (N_7709,N_5061,N_6215);
nor U7710 (N_7710,N_5393,N_7126);
nand U7711 (N_7711,N_7313,N_5641);
xor U7712 (N_7712,N_5038,N_7431);
xor U7713 (N_7713,N_5184,N_5881);
xnor U7714 (N_7714,N_6464,N_5619);
and U7715 (N_7715,N_5144,N_6463);
nor U7716 (N_7716,N_6503,N_5587);
nand U7717 (N_7717,N_6809,N_6502);
and U7718 (N_7718,N_5217,N_5029);
nor U7719 (N_7719,N_5742,N_5289);
nand U7720 (N_7720,N_7069,N_6612);
nor U7721 (N_7721,N_5335,N_5584);
or U7722 (N_7722,N_7232,N_5838);
nor U7723 (N_7723,N_6339,N_5901);
xnor U7724 (N_7724,N_5538,N_5403);
nand U7725 (N_7725,N_6759,N_5183);
nor U7726 (N_7726,N_5782,N_5944);
xor U7727 (N_7727,N_5546,N_6213);
or U7728 (N_7728,N_7469,N_7127);
nor U7729 (N_7729,N_5635,N_5259);
xnor U7730 (N_7730,N_7037,N_5424);
nor U7731 (N_7731,N_6462,N_5488);
xor U7732 (N_7732,N_6855,N_7155);
or U7733 (N_7733,N_6876,N_6311);
xor U7734 (N_7734,N_5762,N_6154);
and U7735 (N_7735,N_6662,N_6461);
nor U7736 (N_7736,N_5814,N_6987);
and U7737 (N_7737,N_5166,N_5940);
or U7738 (N_7738,N_7279,N_7096);
nor U7739 (N_7739,N_6862,N_6636);
nor U7740 (N_7740,N_5398,N_6048);
xnor U7741 (N_7741,N_6177,N_6742);
xnor U7742 (N_7742,N_7369,N_5848);
and U7743 (N_7743,N_6203,N_7460);
or U7744 (N_7744,N_5629,N_6080);
nand U7745 (N_7745,N_6074,N_7374);
nor U7746 (N_7746,N_6003,N_5192);
nand U7747 (N_7747,N_7450,N_5965);
or U7748 (N_7748,N_5462,N_6267);
nand U7749 (N_7749,N_5209,N_5835);
xnor U7750 (N_7750,N_5647,N_5933);
nand U7751 (N_7751,N_5503,N_5543);
or U7752 (N_7752,N_7439,N_7325);
xnor U7753 (N_7753,N_5278,N_5291);
or U7754 (N_7754,N_6712,N_5873);
xor U7755 (N_7755,N_6516,N_6588);
and U7756 (N_7756,N_5821,N_6609);
nand U7757 (N_7757,N_5734,N_6860);
xor U7758 (N_7758,N_5411,N_5738);
nand U7759 (N_7759,N_6257,N_6489);
nand U7760 (N_7760,N_5589,N_5953);
and U7761 (N_7761,N_6234,N_6602);
nand U7762 (N_7762,N_5201,N_6637);
or U7763 (N_7763,N_7306,N_6196);
nor U7764 (N_7764,N_6038,N_5919);
nand U7765 (N_7765,N_5797,N_5309);
xor U7766 (N_7766,N_5804,N_5548);
nand U7767 (N_7767,N_5266,N_5229);
xor U7768 (N_7768,N_7383,N_5926);
nor U7769 (N_7769,N_6403,N_6585);
nand U7770 (N_7770,N_6751,N_5566);
and U7771 (N_7771,N_5126,N_5519);
and U7772 (N_7772,N_6214,N_5920);
xor U7773 (N_7773,N_7429,N_6795);
or U7774 (N_7774,N_7175,N_7091);
xnor U7775 (N_7775,N_7433,N_6188);
xor U7776 (N_7776,N_5740,N_5102);
and U7777 (N_7777,N_6361,N_7351);
or U7778 (N_7778,N_5524,N_5163);
nand U7779 (N_7779,N_5949,N_6732);
xor U7780 (N_7780,N_6675,N_7443);
and U7781 (N_7781,N_6054,N_6444);
nand U7782 (N_7782,N_7083,N_5955);
or U7783 (N_7783,N_6695,N_7435);
nand U7784 (N_7784,N_6315,N_7062);
and U7785 (N_7785,N_5176,N_5481);
nor U7786 (N_7786,N_6376,N_5046);
and U7787 (N_7787,N_5928,N_5977);
and U7788 (N_7788,N_6240,N_7068);
nand U7789 (N_7789,N_5401,N_5486);
and U7790 (N_7790,N_5431,N_7051);
or U7791 (N_7791,N_7099,N_5157);
nor U7792 (N_7792,N_5094,N_5255);
nor U7793 (N_7793,N_5895,N_7248);
and U7794 (N_7794,N_6815,N_6285);
nand U7795 (N_7795,N_6050,N_5025);
nor U7796 (N_7796,N_6399,N_6160);
xnor U7797 (N_7797,N_7337,N_6899);
or U7798 (N_7798,N_6773,N_7436);
nand U7799 (N_7799,N_7179,N_6689);
nand U7800 (N_7800,N_5237,N_5938);
nand U7801 (N_7801,N_6483,N_6991);
xor U7802 (N_7802,N_6407,N_5448);
nor U7803 (N_7803,N_6450,N_7393);
or U7804 (N_7804,N_6322,N_6039);
or U7805 (N_7805,N_5565,N_6498);
xnor U7806 (N_7806,N_6192,N_5131);
nand U7807 (N_7807,N_5831,N_6634);
nor U7808 (N_7808,N_5910,N_7187);
and U7809 (N_7809,N_5736,N_6232);
nor U7810 (N_7810,N_7312,N_5070);
nand U7811 (N_7811,N_6641,N_6857);
nor U7812 (N_7812,N_6639,N_7020);
and U7813 (N_7813,N_5013,N_5471);
xnor U7814 (N_7814,N_5653,N_7066);
xnor U7815 (N_7815,N_5437,N_7001);
nand U7816 (N_7816,N_6052,N_6768);
xnor U7817 (N_7817,N_7173,N_7455);
nand U7818 (N_7818,N_7141,N_6076);
nor U7819 (N_7819,N_7163,N_6245);
xnor U7820 (N_7820,N_7377,N_7041);
or U7821 (N_7821,N_6981,N_6613);
nor U7822 (N_7822,N_5865,N_6111);
nand U7823 (N_7823,N_6261,N_7471);
nor U7824 (N_7824,N_7274,N_5700);
or U7825 (N_7825,N_6026,N_5317);
xor U7826 (N_7826,N_6971,N_6536);
or U7827 (N_7827,N_6735,N_7390);
nand U7828 (N_7828,N_5210,N_7446);
xor U7829 (N_7829,N_7144,N_5914);
nand U7830 (N_7830,N_5427,N_6660);
or U7831 (N_7831,N_6798,N_6127);
or U7832 (N_7832,N_7359,N_6067);
and U7833 (N_7833,N_5662,N_5198);
nand U7834 (N_7834,N_5048,N_6869);
and U7835 (N_7835,N_6802,N_5394);
and U7836 (N_7836,N_5265,N_5834);
or U7837 (N_7837,N_5090,N_7310);
nand U7838 (N_7838,N_6698,N_6197);
nor U7839 (N_7839,N_6471,N_5604);
nand U7840 (N_7840,N_5189,N_5580);
and U7841 (N_7841,N_6481,N_5402);
and U7842 (N_7842,N_6218,N_5179);
xnor U7843 (N_7843,N_6746,N_6838);
xor U7844 (N_7844,N_5582,N_5084);
and U7845 (N_7845,N_5967,N_6053);
nor U7846 (N_7846,N_5044,N_6246);
xnor U7847 (N_7847,N_6046,N_5111);
nand U7848 (N_7848,N_6405,N_5385);
nor U7849 (N_7849,N_6066,N_5085);
nor U7850 (N_7850,N_5457,N_6647);
nand U7851 (N_7851,N_7466,N_5330);
or U7852 (N_7852,N_5340,N_6041);
nor U7853 (N_7853,N_5811,N_6594);
nand U7854 (N_7854,N_6610,N_6167);
nand U7855 (N_7855,N_6087,N_7050);
xnor U7856 (N_7856,N_5986,N_7494);
nand U7857 (N_7857,N_7277,N_7109);
and U7858 (N_7858,N_7286,N_5532);
or U7859 (N_7859,N_5705,N_6969);
and U7860 (N_7860,N_5624,N_5392);
nor U7861 (N_7861,N_5557,N_7453);
or U7862 (N_7862,N_6993,N_5115);
and U7863 (N_7863,N_6434,N_5140);
or U7864 (N_7864,N_6570,N_6002);
or U7865 (N_7865,N_5019,N_6685);
xnor U7866 (N_7866,N_6217,N_6925);
nor U7867 (N_7867,N_6520,N_7333);
and U7868 (N_7868,N_7490,N_6346);
xor U7869 (N_7869,N_5128,N_6043);
xor U7870 (N_7870,N_5318,N_6635);
xor U7871 (N_7871,N_6014,N_6786);
xnor U7872 (N_7872,N_7171,N_7213);
nand U7873 (N_7873,N_5134,N_7142);
or U7874 (N_7874,N_6166,N_6393);
xor U7875 (N_7875,N_6018,N_5861);
nand U7876 (N_7876,N_6210,N_7408);
and U7877 (N_7877,N_6247,N_6476);
nor U7878 (N_7878,N_5492,N_7172);
xor U7879 (N_7879,N_7139,N_7473);
or U7880 (N_7880,N_5525,N_6811);
nand U7881 (N_7881,N_7056,N_5952);
nor U7882 (N_7882,N_5321,N_5375);
and U7883 (N_7883,N_5129,N_6738);
or U7884 (N_7884,N_5522,N_6357);
nor U7885 (N_7885,N_6599,N_6354);
and U7886 (N_7886,N_5286,N_7065);
and U7887 (N_7887,N_5238,N_6394);
and U7888 (N_7888,N_5450,N_5946);
or U7889 (N_7889,N_7398,N_6659);
or U7890 (N_7890,N_6044,N_6770);
nor U7891 (N_7891,N_6961,N_5744);
xnor U7892 (N_7892,N_7006,N_5263);
xor U7893 (N_7893,N_6524,N_6509);
nor U7894 (N_7894,N_6029,N_7267);
or U7895 (N_7895,N_5718,N_7299);
or U7896 (N_7896,N_6432,N_5130);
nor U7897 (N_7897,N_6031,N_6648);
or U7898 (N_7898,N_5717,N_5032);
nor U7899 (N_7899,N_7437,N_6842);
or U7900 (N_7900,N_7147,N_6598);
xor U7901 (N_7901,N_6383,N_5535);
nand U7902 (N_7902,N_6501,N_7107);
or U7903 (N_7903,N_5670,N_7080);
xnor U7904 (N_7904,N_5631,N_5078);
nand U7905 (N_7905,N_5283,N_7215);
nor U7906 (N_7906,N_5526,N_5249);
nor U7907 (N_7907,N_5319,N_5388);
nand U7908 (N_7908,N_6007,N_5240);
nand U7909 (N_7909,N_6119,N_7093);
or U7910 (N_7910,N_5002,N_6324);
xor U7911 (N_7911,N_6922,N_5288);
xnor U7912 (N_7912,N_6102,N_5572);
xnor U7913 (N_7913,N_5591,N_6914);
nand U7914 (N_7914,N_5595,N_7237);
nand U7915 (N_7915,N_6850,N_6728);
xnor U7916 (N_7916,N_6423,N_5669);
nand U7917 (N_7917,N_7464,N_5818);
and U7918 (N_7918,N_6398,N_6847);
xnor U7919 (N_7919,N_5561,N_6927);
nor U7920 (N_7920,N_7276,N_5196);
or U7921 (N_7921,N_6047,N_6904);
and U7922 (N_7922,N_7095,N_5636);
nor U7923 (N_7923,N_7400,N_6116);
nand U7924 (N_7924,N_7251,N_6117);
xor U7925 (N_7925,N_5477,N_5139);
nor U7926 (N_7926,N_6421,N_6601);
or U7927 (N_7927,N_7184,N_5577);
nor U7928 (N_7928,N_5791,N_6334);
and U7929 (N_7929,N_5843,N_5328);
xor U7930 (N_7930,N_5248,N_6207);
nor U7931 (N_7931,N_6833,N_7321);
or U7932 (N_7932,N_6848,N_5363);
xnor U7933 (N_7933,N_5175,N_5520);
xnor U7934 (N_7934,N_5316,N_7034);
nor U7935 (N_7935,N_6082,N_5807);
nor U7936 (N_7936,N_5122,N_6999);
or U7937 (N_7937,N_7354,N_5232);
or U7938 (N_7938,N_6107,N_5245);
or U7939 (N_7939,N_6551,N_6475);
nand U7940 (N_7940,N_5658,N_7199);
or U7941 (N_7941,N_5787,N_6706);
xor U7942 (N_7942,N_6627,N_7018);
nand U7943 (N_7943,N_6237,N_5714);
nor U7944 (N_7944,N_5975,N_7048);
or U7945 (N_7945,N_5646,N_5999);
and U7946 (N_7946,N_7280,N_7222);
nor U7947 (N_7947,N_5478,N_6982);
and U7948 (N_7948,N_5713,N_7288);
nand U7949 (N_7949,N_5353,N_6063);
nor U7950 (N_7950,N_6487,N_6380);
or U7951 (N_7951,N_6112,N_6277);
xor U7952 (N_7952,N_6960,N_7252);
nand U7953 (N_7953,N_5555,N_5673);
nor U7954 (N_7954,N_5899,N_7261);
and U7955 (N_7955,N_6718,N_5845);
or U7956 (N_7956,N_6664,N_5904);
and U7957 (N_7957,N_7220,N_6439);
nor U7958 (N_7958,N_5366,N_5430);
or U7959 (N_7959,N_5164,N_6159);
xor U7960 (N_7960,N_6544,N_6426);
and U7961 (N_7961,N_5593,N_5988);
nand U7962 (N_7962,N_6424,N_6940);
nor U7963 (N_7963,N_6931,N_5389);
nor U7964 (N_7964,N_7451,N_6360);
and U7965 (N_7965,N_5685,N_7208);
and U7966 (N_7966,N_6226,N_7060);
nand U7967 (N_7967,N_5173,N_5943);
or U7968 (N_7968,N_6913,N_7211);
nor U7969 (N_7969,N_5103,N_5379);
and U7970 (N_7970,N_6778,N_5344);
xnor U7971 (N_7971,N_5387,N_6079);
nor U7972 (N_7972,N_5979,N_6945);
nor U7973 (N_7973,N_6870,N_7474);
and U7974 (N_7974,N_6515,N_5796);
xor U7975 (N_7975,N_5623,N_5530);
or U7976 (N_7976,N_6836,N_7297);
nand U7977 (N_7977,N_5124,N_6651);
nor U7978 (N_7978,N_5154,N_7239);
xnor U7979 (N_7979,N_5822,N_5866);
nand U7980 (N_7980,N_6320,N_7067);
and U7981 (N_7981,N_6929,N_6741);
and U7982 (N_7982,N_7216,N_6806);
xor U7983 (N_7983,N_6958,N_6325);
nor U7984 (N_7984,N_5799,N_7085);
nand U7985 (N_7985,N_7385,N_5798);
and U7986 (N_7986,N_7003,N_7212);
nand U7987 (N_7987,N_6259,N_5047);
or U7988 (N_7988,N_7344,N_5469);
or U7989 (N_7989,N_7161,N_5088);
and U7990 (N_7990,N_7338,N_7059);
xor U7991 (N_7991,N_6653,N_6534);
nor U7992 (N_7992,N_5305,N_6150);
xnor U7993 (N_7993,N_6578,N_7246);
or U7994 (N_7994,N_6596,N_5726);
xnor U7995 (N_7995,N_7477,N_5883);
and U7996 (N_7996,N_5622,N_7432);
and U7997 (N_7997,N_5470,N_6488);
or U7998 (N_7998,N_5844,N_5983);
nor U7999 (N_7999,N_5541,N_5258);
nor U8000 (N_8000,N_5380,N_5361);
or U8001 (N_8001,N_6104,N_5906);
or U8002 (N_8002,N_5982,N_7345);
nor U8003 (N_8003,N_6429,N_5364);
nor U8004 (N_8004,N_7078,N_6916);
nor U8005 (N_8005,N_5820,N_5846);
nor U8006 (N_8006,N_6716,N_5441);
nand U8007 (N_8007,N_6557,N_5573);
xor U8008 (N_8008,N_6934,N_5730);
nor U8009 (N_8009,N_5794,N_5274);
nand U8010 (N_8010,N_5276,N_5759);
nand U8011 (N_8011,N_7484,N_6500);
or U8012 (N_8012,N_6793,N_6015);
and U8013 (N_8013,N_6573,N_5420);
xor U8014 (N_8014,N_5802,N_5696);
or U8015 (N_8015,N_7240,N_7145);
nor U8016 (N_8016,N_6745,N_7036);
or U8017 (N_8017,N_5569,N_5185);
or U8018 (N_8018,N_6153,N_6055);
or U8019 (N_8019,N_6906,N_5023);
or U8020 (N_8020,N_7090,N_5540);
xor U8021 (N_8021,N_7135,N_6158);
or U8022 (N_8022,N_6508,N_6577);
and U8023 (N_8023,N_6310,N_6059);
or U8024 (N_8024,N_7011,N_7367);
xor U8025 (N_8025,N_6510,N_5298);
xor U8026 (N_8026,N_5417,N_6148);
or U8027 (N_8027,N_7070,N_6425);
nor U8028 (N_8028,N_5331,N_7290);
and U8029 (N_8029,N_6615,N_5072);
and U8030 (N_8030,N_5026,N_6085);
xor U8031 (N_8031,N_6995,N_7040);
nand U8032 (N_8032,N_6595,N_6518);
nand U8033 (N_8033,N_6060,N_6368);
and U8034 (N_8034,N_5150,N_5609);
nand U8035 (N_8035,N_7013,N_7072);
and U8036 (N_8036,N_6243,N_6710);
nand U8037 (N_8037,N_5141,N_6023);
or U8038 (N_8038,N_6083,N_7328);
or U8039 (N_8039,N_6808,N_7265);
or U8040 (N_8040,N_6145,N_6300);
and U8041 (N_8041,N_5499,N_5485);
xor U8042 (N_8042,N_5630,N_6284);
nor U8043 (N_8043,N_5043,N_6655);
xor U8044 (N_8044,N_5300,N_6415);
nand U8045 (N_8045,N_5500,N_6650);
xnor U8046 (N_8046,N_7285,N_6926);
xnor U8047 (N_8047,N_6430,N_5474);
nand U8048 (N_8048,N_6771,N_5842);
or U8049 (N_8049,N_7371,N_7241);
nor U8050 (N_8050,N_5512,N_7411);
nor U8051 (N_8051,N_6268,N_5033);
or U8052 (N_8052,N_6777,N_7264);
and U8053 (N_8053,N_6221,N_7257);
xor U8054 (N_8054,N_6807,N_6620);
nand U8055 (N_8055,N_5931,N_5172);
nand U8056 (N_8056,N_5517,N_5993);
and U8057 (N_8057,N_6704,N_5466);
nand U8058 (N_8058,N_6733,N_6090);
nand U8059 (N_8059,N_6165,N_6803);
nand U8060 (N_8060,N_6986,N_5060);
nor U8061 (N_8061,N_6629,N_6124);
or U8062 (N_8062,N_5251,N_6486);
xnor U8063 (N_8063,N_6199,N_6420);
xnor U8064 (N_8064,N_5628,N_7061);
and U8065 (N_8065,N_6448,N_7340);
nand U8066 (N_8066,N_5279,N_7287);
nand U8067 (N_8067,N_7235,N_5516);
nor U8068 (N_8068,N_6694,N_6255);
nor U8069 (N_8069,N_6499,N_5484);
nor U8070 (N_8070,N_6460,N_5064);
nand U8071 (N_8071,N_6347,N_6305);
or U8072 (N_8072,N_7326,N_5909);
nor U8073 (N_8073,N_7210,N_6445);
and U8074 (N_8074,N_6209,N_5686);
nor U8075 (N_8075,N_6624,N_5193);
and U8076 (N_8076,N_5142,N_5518);
or U8077 (N_8077,N_7100,N_6859);
and U8078 (N_8078,N_6068,N_6413);
xnor U8079 (N_8079,N_6723,N_7480);
xnor U8080 (N_8080,N_5887,N_6661);
nand U8081 (N_8081,N_5374,N_5858);
nand U8082 (N_8082,N_5915,N_5870);
nand U8083 (N_8083,N_6783,N_5376);
xor U8084 (N_8084,N_6740,N_7335);
nand U8085 (N_8085,N_5859,N_6169);
xor U8086 (N_8086,N_6431,N_6058);
nand U8087 (N_8087,N_6656,N_5065);
xnor U8088 (N_8088,N_7406,N_6414);
xnor U8089 (N_8089,N_5832,N_6586);
nand U8090 (N_8090,N_6545,N_6566);
and U8091 (N_8091,N_6841,N_5711);
xor U8092 (N_8092,N_6321,N_7028);
or U8093 (N_8093,N_6556,N_5400);
or U8094 (N_8094,N_6903,N_5284);
or U8095 (N_8095,N_6138,N_5852);
or U8096 (N_8096,N_7372,N_5600);
nand U8097 (N_8097,N_6938,N_5616);
and U8098 (N_8098,N_6939,N_7138);
nand U8099 (N_8099,N_7218,N_7167);
nor U8100 (N_8100,N_5067,N_5372);
nor U8101 (N_8101,N_7388,N_7149);
or U8102 (N_8102,N_5247,N_5197);
nor U8103 (N_8103,N_6223,N_6093);
xnor U8104 (N_8104,N_5735,N_6096);
nor U8105 (N_8105,N_6640,N_5194);
xor U8106 (N_8106,N_5213,N_6511);
and U8107 (N_8107,N_6281,N_5552);
and U8108 (N_8108,N_6184,N_6428);
nor U8109 (N_8109,N_5515,N_5073);
nor U8110 (N_8110,N_7415,N_6181);
and U8111 (N_8111,N_6309,N_5106);
nand U8112 (N_8112,N_6856,N_6064);
nand U8113 (N_8113,N_6895,N_5528);
or U8114 (N_8114,N_5539,N_6349);
xor U8115 (N_8115,N_7407,N_6677);
nand U8116 (N_8116,N_7064,N_5083);
or U8117 (N_8117,N_5849,N_6465);
or U8118 (N_8118,N_5490,N_6201);
or U8119 (N_8119,N_5644,N_5962);
and U8120 (N_8120,N_5575,N_7425);
nand U8121 (N_8121,N_7140,N_6937);
or U8122 (N_8122,N_6752,N_7194);
xor U8123 (N_8123,N_5171,N_5684);
nand U8124 (N_8124,N_6156,N_6094);
xnor U8125 (N_8125,N_5771,N_5709);
nand U8126 (N_8126,N_5349,N_7273);
xnor U8127 (N_8127,N_6417,N_5521);
or U8128 (N_8128,N_5370,N_5504);
nand U8129 (N_8129,N_6081,N_7193);
and U8130 (N_8130,N_5004,N_5836);
nand U8131 (N_8131,N_5010,N_6482);
xor U8132 (N_8132,N_7356,N_5148);
nand U8133 (N_8133,N_5970,N_6123);
nand U8134 (N_8134,N_6402,N_6069);
nor U8135 (N_8135,N_6630,N_6035);
or U8136 (N_8136,N_6478,N_5837);
xnor U8137 (N_8137,N_6130,N_5617);
nor U8138 (N_8138,N_5633,N_7255);
nand U8139 (N_8139,N_6671,N_6550);
and U8140 (N_8140,N_7262,N_5779);
and U8141 (N_8141,N_5950,N_6264);
or U8142 (N_8142,N_5749,N_5697);
nand U8143 (N_8143,N_5793,N_5667);
xor U8144 (N_8144,N_5649,N_7352);
and U8145 (N_8145,N_5720,N_6454);
or U8146 (N_8146,N_6581,N_7467);
or U8147 (N_8147,N_5311,N_5170);
nand U8148 (N_8148,N_5727,N_7174);
and U8149 (N_8149,N_5307,N_7116);
nand U8150 (N_8150,N_5708,N_7339);
nand U8151 (N_8151,N_7444,N_6252);
nand U8152 (N_8152,N_6030,N_5674);
and U8153 (N_8153,N_5603,N_5916);
or U8154 (N_8154,N_6538,N_5207);
nor U8155 (N_8155,N_7076,N_5151);
xnor U8156 (N_8156,N_6377,N_5108);
or U8157 (N_8157,N_5941,N_5123);
nor U8158 (N_8158,N_5270,N_5893);
xor U8159 (N_8159,N_6397,N_6051);
or U8160 (N_8160,N_5780,N_6800);
nand U8161 (N_8161,N_5888,N_5545);
and U8162 (N_8162,N_7089,N_6892);
and U8163 (N_8163,N_6722,N_5505);
nor U8164 (N_8164,N_6474,N_5467);
and U8165 (N_8165,N_6495,N_6957);
nor U8166 (N_8166,N_5874,N_6552);
and U8167 (N_8167,N_5007,N_5395);
and U8168 (N_8168,N_7188,N_5093);
xnor U8169 (N_8169,N_5923,N_6909);
nand U8170 (N_8170,N_5009,N_6469);
nand U8171 (N_8171,N_5781,N_5805);
or U8172 (N_8172,N_6834,N_7201);
nand U8173 (N_8173,N_5404,N_6944);
or U8174 (N_8174,N_6574,N_5018);
nor U8175 (N_8175,N_5105,N_6338);
and U8176 (N_8176,N_7035,N_7148);
and U8177 (N_8177,N_6097,N_5872);
xor U8178 (N_8178,N_6755,N_5343);
nand U8179 (N_8179,N_5097,N_5754);
nand U8180 (N_8180,N_6468,N_7387);
and U8181 (N_8181,N_5313,N_5337);
and U8182 (N_8182,N_6179,N_5116);
nand U8183 (N_8183,N_6707,N_6205);
xor U8184 (N_8184,N_5969,N_5594);
or U8185 (N_8185,N_5080,N_7382);
nand U8186 (N_8186,N_6323,N_6120);
nand U8187 (N_8187,N_6329,N_5006);
xnor U8188 (N_8188,N_7195,N_6382);
or U8189 (N_8189,N_7379,N_6446);
nand U8190 (N_8190,N_5891,N_7413);
xnor U8191 (N_8191,N_6571,N_6864);
or U8192 (N_8192,N_5257,N_7270);
nand U8193 (N_8193,N_5310,N_6270);
nor U8194 (N_8194,N_5365,N_6603);
nor U8195 (N_8195,N_5425,N_7146);
and U8196 (N_8196,N_6890,N_6827);
nand U8197 (N_8197,N_5810,N_5702);
nor U8198 (N_8198,N_5602,N_5803);
and U8199 (N_8199,N_6504,N_5068);
or U8200 (N_8200,N_6396,N_6875);
nand U8201 (N_8201,N_5775,N_6673);
nor U8202 (N_8202,N_5051,N_7219);
xnor U8203 (N_8203,N_6565,N_6766);
and U8204 (N_8204,N_5990,N_6072);
xnor U8205 (N_8205,N_6955,N_6458);
nand U8206 (N_8206,N_5693,N_5806);
or U8207 (N_8207,N_6493,N_6362);
or U8208 (N_8208,N_5066,N_5574);
nor U8209 (N_8209,N_6657,N_6787);
nand U8210 (N_8210,N_6390,N_6326);
nor U8211 (N_8211,N_7301,N_6918);
nor U8212 (N_8212,N_7320,N_5506);
xor U8213 (N_8213,N_6748,N_6812);
nor U8214 (N_8214,N_5612,N_7021);
nand U8215 (N_8215,N_7399,N_5063);
or U8216 (N_8216,N_6437,N_5159);
nand U8217 (N_8217,N_5260,N_5224);
nor U8218 (N_8218,N_6392,N_5980);
xor U8219 (N_8219,N_5005,N_7341);
nand U8220 (N_8220,N_6496,N_6379);
nor U8221 (N_8221,N_7104,N_5689);
nand U8222 (N_8222,N_5994,N_7308);
or U8223 (N_8223,N_7030,N_5905);
nand U8224 (N_8224,N_7166,N_5422);
and U8225 (N_8225,N_7180,N_6416);
nor U8226 (N_8226,N_5911,N_5973);
nand U8227 (N_8227,N_6293,N_5606);
or U8228 (N_8228,N_5015,N_6225);
nand U8229 (N_8229,N_7170,N_5155);
xor U8230 (N_8230,N_5830,N_6708);
xor U8231 (N_8231,N_6784,N_5086);
nand U8232 (N_8232,N_5491,N_6466);
and U8233 (N_8233,N_6744,N_7164);
or U8234 (N_8234,N_7110,N_6303);
nand U8235 (N_8235,N_6820,N_6776);
or U8236 (N_8236,N_6592,N_7132);
xor U8237 (N_8237,N_7426,N_6911);
nor U8238 (N_8238,N_7221,N_6762);
xnor U8239 (N_8239,N_6674,N_6149);
xor U8240 (N_8240,N_6724,N_5621);
nor U8241 (N_8241,N_5777,N_5180);
nand U8242 (N_8242,N_7442,N_6868);
xnor U8243 (N_8243,N_6008,N_6356);
and U8244 (N_8244,N_5985,N_5287);
nand U8245 (N_8245,N_5358,N_5867);
nor U8246 (N_8246,N_6858,N_7224);
nor U8247 (N_8247,N_6591,N_5929);
and U8248 (N_8248,N_5672,N_6128);
xor U8249 (N_8249,N_7016,N_5596);
nand U8250 (N_8250,N_6175,N_7403);
and U8251 (N_8251,N_6531,N_5570);
xnor U8252 (N_8252,N_5963,N_5182);
or U8253 (N_8253,N_6889,N_7000);
nand U8254 (N_8254,N_5186,N_7081);
nor U8255 (N_8255,N_6202,N_5741);
nor U8256 (N_8256,N_6375,N_5544);
xor U8257 (N_8257,N_6367,N_7275);
nor U8258 (N_8258,N_6691,N_5932);
or U8259 (N_8259,N_7410,N_7071);
or U8260 (N_8260,N_5774,N_6558);
xor U8261 (N_8261,N_5212,N_5381);
nor U8262 (N_8262,N_7137,N_6952);
xnor U8263 (N_8263,N_6684,N_7357);
xnor U8264 (N_8264,N_6514,N_5934);
or U8265 (N_8265,N_6646,N_5855);
or U8266 (N_8266,N_7366,N_6078);
nand U8267 (N_8267,N_7247,N_5996);
and U8268 (N_8268,N_5428,N_6915);
or U8269 (N_8269,N_5268,N_7260);
or U8270 (N_8270,N_6412,N_5768);
nand U8271 (N_8271,N_5095,N_6395);
nor U8272 (N_8272,N_7282,N_6371);
xnor U8273 (N_8273,N_6672,N_6583);
or U8274 (N_8274,N_6764,N_6204);
nand U8275 (N_8275,N_6477,N_5324);
nand U8276 (N_8276,N_5509,N_5699);
nand U8277 (N_8277,N_5579,N_6756);
and U8278 (N_8278,N_7254,N_7329);
or U8279 (N_8279,N_6319,N_7364);
and U8280 (N_8280,N_5523,N_5178);
and U8281 (N_8281,N_6024,N_6505);
and U8282 (N_8282,N_6455,N_5320);
and U8283 (N_8283,N_5897,N_6767);
xor U8284 (N_8284,N_5808,N_5113);
or U8285 (N_8285,N_5784,N_7014);
xnor U8286 (N_8286,N_6749,N_5666);
nand U8287 (N_8287,N_6830,N_5243);
or U8288 (N_8288,N_5688,N_5410);
xor U8289 (N_8289,N_6669,N_5813);
xor U8290 (N_8290,N_5704,N_7378);
nor U8291 (N_8291,N_5995,N_5945);
xor U8292 (N_8292,N_5205,N_6456);
and U8293 (N_8293,N_6180,N_5280);
or U8294 (N_8294,N_6242,N_6977);
and U8295 (N_8295,N_5342,N_7073);
or U8296 (N_8296,N_5125,N_6001);
nand U8297 (N_8297,N_6821,N_7039);
or U8298 (N_8298,N_5790,N_6019);
xnor U8299 (N_8299,N_6236,N_5840);
and U8300 (N_8300,N_6765,N_5082);
xnor U8301 (N_8301,N_7284,N_6992);
or U8302 (N_8302,N_7214,N_6172);
nor U8303 (N_8303,N_6276,N_6372);
nand U8304 (N_8304,N_6164,N_6962);
or U8305 (N_8305,N_5902,N_6294);
nand U8306 (N_8306,N_6440,N_5597);
xnor U8307 (N_8307,N_6230,N_6692);
or U8308 (N_8308,N_6758,N_5981);
xor U8309 (N_8309,N_6280,N_5878);
or U8310 (N_8310,N_7118,N_5511);
nor U8311 (N_8311,N_6028,N_6262);
and U8312 (N_8312,N_7042,N_6385);
nor U8313 (N_8313,N_6750,N_6073);
or U8314 (N_8314,N_7223,N_5293);
nand U8315 (N_8315,N_6611,N_6313);
nand U8316 (N_8316,N_6528,N_5513);
xor U8317 (N_8317,N_6697,N_6972);
nor U8318 (N_8318,N_5429,N_6625);
nand U8319 (N_8319,N_6077,N_6497);
nor U8320 (N_8320,N_7189,N_7101);
nand U8321 (N_8321,N_5826,N_5062);
xor U8322 (N_8322,N_6792,N_5306);
or U8323 (N_8323,N_5409,N_6265);
xor U8324 (N_8324,N_7309,N_5329);
nand U8325 (N_8325,N_5769,N_6433);
nand U8326 (N_8326,N_6122,N_7032);
and U8327 (N_8327,N_5638,N_5527);
and U8328 (N_8328,N_5227,N_5937);
or U8329 (N_8329,N_6679,N_6314);
or U8330 (N_8330,N_5998,N_5412);
or U8331 (N_8331,N_7302,N_5651);
xnor U8332 (N_8332,N_6555,N_6219);
nor U8333 (N_8333,N_5314,N_7114);
xor U8334 (N_8334,N_7046,N_6933);
xnor U8335 (N_8335,N_6747,N_6680);
and U8336 (N_8336,N_5339,N_5632);
and U8337 (N_8337,N_6831,N_6490);
nand U8338 (N_8338,N_5098,N_7058);
nand U8339 (N_8339,N_5894,N_6621);
and U8340 (N_8340,N_5277,N_5757);
xor U8341 (N_8341,N_7492,N_7084);
nor U8342 (N_8342,N_5677,N_6198);
and U8343 (N_8343,N_7269,N_7346);
nand U8344 (N_8344,N_6452,N_5801);
or U8345 (N_8345,N_6404,N_5560);
or U8346 (N_8346,N_5608,N_5960);
and U8347 (N_8347,N_5829,N_5533);
and U8348 (N_8348,N_7303,N_5352);
or U8349 (N_8349,N_7230,N_5377);
and U8350 (N_8350,N_5413,N_6100);
nand U8351 (N_8351,N_6753,N_6727);
nand U8352 (N_8352,N_7272,N_5132);
nand U8353 (N_8353,N_7459,N_7295);
or U8354 (N_8354,N_7242,N_5536);
xnor U8355 (N_8355,N_7488,N_7360);
or U8356 (N_8356,N_6649,N_7023);
xnor U8357 (N_8357,N_6954,N_7478);
xnor U8358 (N_8358,N_6572,N_7165);
nor U8359 (N_8359,N_6568,N_6825);
or U8360 (N_8360,N_6381,N_6983);
and U8361 (N_8361,N_5508,N_6260);
nor U8362 (N_8362,N_6567,N_6229);
or U8363 (N_8363,N_6101,N_5003);
nor U8364 (N_8364,N_7203,N_7079);
nand U8365 (N_8365,N_7315,N_6110);
and U8366 (N_8366,N_6126,N_6147);
nand U8367 (N_8367,N_5681,N_6563);
and U8368 (N_8368,N_7389,N_6682);
xnor U8369 (N_8369,N_7462,N_7154);
xnor U8370 (N_8370,N_5896,N_7186);
or U8371 (N_8371,N_5514,N_6607);
and U8372 (N_8372,N_5421,N_5112);
and U8373 (N_8373,N_5789,N_6846);
nand U8374 (N_8374,N_7305,N_7125);
or U8375 (N_8375,N_7112,N_5788);
and U8376 (N_8376,N_5851,N_5817);
xor U8377 (N_8377,N_5640,N_7129);
and U8378 (N_8378,N_6113,N_7294);
and U8379 (N_8379,N_6331,N_6155);
nand U8380 (N_8380,N_6533,N_6797);
xor U8381 (N_8381,N_6951,N_5639);
and U8382 (N_8382,N_5034,N_6560);
nor U8383 (N_8383,N_6837,N_6985);
and U8384 (N_8384,N_6579,N_6228);
and U8385 (N_8385,N_7153,N_5081);
nand U8386 (N_8386,N_5322,N_5074);
or U8387 (N_8387,N_6720,N_6902);
nand U8388 (N_8388,N_6829,N_5476);
nor U8389 (N_8389,N_7119,N_6291);
nand U8390 (N_8390,N_6327,N_5057);
nand U8391 (N_8391,N_7022,N_6884);
nor U8392 (N_8392,N_5426,N_5367);
or U8393 (N_8393,N_7445,N_6186);
nor U8394 (N_8394,N_7349,N_5169);
nand U8395 (N_8395,N_5764,N_5233);
or U8396 (N_8396,N_7348,N_6373);
or U8397 (N_8397,N_5109,N_5052);
nor U8398 (N_8398,N_6638,N_6195);
xor U8399 (N_8399,N_5386,N_7176);
xor U8400 (N_8400,N_5133,N_7414);
or U8401 (N_8401,N_6012,N_6619);
nand U8402 (N_8402,N_6663,N_6593);
nor U8403 (N_8403,N_6328,N_5763);
and U8404 (N_8404,N_6628,N_5913);
nor U8405 (N_8405,N_7394,N_5459);
nor U8406 (N_8406,N_5722,N_6312);
nor U8407 (N_8407,N_6438,N_7206);
and U8408 (N_8408,N_5326,N_7347);
or U8409 (N_8409,N_5152,N_6517);
nand U8410 (N_8410,N_5181,N_5449);
nand U8411 (N_8411,N_5966,N_5235);
xnor U8412 (N_8412,N_7447,N_5554);
or U8413 (N_8413,N_5348,N_5027);
nand U8414 (N_8414,N_7319,N_7192);
and U8415 (N_8415,N_5756,N_5303);
nor U8416 (N_8416,N_5271,N_5581);
nand U8417 (N_8417,N_7495,N_5202);
nor U8418 (N_8418,N_6342,N_5598);
xnor U8419 (N_8419,N_7461,N_7317);
nand U8420 (N_8420,N_6271,N_6963);
and U8421 (N_8421,N_5200,N_6888);
xnor U8422 (N_8422,N_5323,N_6542);
xnor U8423 (N_8423,N_7177,N_7057);
and U8424 (N_8424,N_6114,N_6279);
nor U8425 (N_8425,N_6882,N_6009);
xor U8426 (N_8426,N_6337,N_5737);
nor U8427 (N_8427,N_5809,N_5531);
or U8428 (N_8428,N_6548,N_6564);
nor U8429 (N_8429,N_7314,N_5613);
or U8430 (N_8430,N_6289,N_7291);
and U8431 (N_8431,N_6772,N_6345);
or U8432 (N_8432,N_7250,N_6930);
nor U8433 (N_8433,N_5325,N_7228);
or U8434 (N_8434,N_7298,N_6966);
nand U8435 (N_8435,N_6631,N_7289);
and U8436 (N_8436,N_5494,N_6546);
nand U8437 (N_8437,N_6849,N_7120);
xor U8438 (N_8438,N_5502,N_7150);
or U8439 (N_8439,N_6575,N_5188);
or U8440 (N_8440,N_7278,N_5703);
and U8441 (N_8441,N_6845,N_5458);
and U8442 (N_8442,N_7227,N_5605);
and U8443 (N_8443,N_5884,N_5959);
nor U8444 (N_8444,N_5301,N_6676);
xor U8445 (N_8445,N_7316,N_5489);
and U8446 (N_8446,N_6099,N_5295);
and U8447 (N_8447,N_6467,N_6248);
or U8448 (N_8448,N_7332,N_6384);
nand U8449 (N_8449,N_7258,N_6559);
nand U8450 (N_8450,N_6642,N_7151);
xor U8451 (N_8451,N_6788,N_5244);
xor U8452 (N_8452,N_5036,N_5795);
nor U8453 (N_8453,N_5715,N_7123);
xnor U8454 (N_8454,N_6132,N_5815);
xor U8455 (N_8455,N_7047,N_6170);
or U8456 (N_8456,N_6020,N_6569);
and U8457 (N_8457,N_5551,N_5290);
xnor U8458 (N_8458,N_6616,N_6442);
xor U8459 (N_8459,N_5497,N_6826);
and U8460 (N_8460,N_6898,N_7343);
nand U8461 (N_8461,N_5075,N_5907);
or U8462 (N_8462,N_5755,N_7111);
xor U8463 (N_8463,N_5542,N_6231);
nand U8464 (N_8464,N_6308,N_6994);
or U8465 (N_8465,N_5346,N_7397);
xor U8466 (N_8466,N_7350,N_5833);
nand U8467 (N_8467,N_6449,N_5908);
nor U8468 (N_8468,N_5695,N_6141);
or U8469 (N_8469,N_6290,N_6106);
xor U8470 (N_8470,N_6633,N_7233);
or U8471 (N_8471,N_5898,N_6644);
and U8472 (N_8472,N_5053,N_6877);
xnor U8473 (N_8473,N_5438,N_6241);
or U8474 (N_8474,N_7249,N_5174);
and U8475 (N_8475,N_5747,N_5890);
or U8476 (N_8476,N_7063,N_6000);
and U8477 (N_8477,N_6997,N_6363);
and U8478 (N_8478,N_5039,N_6686);
nand U8479 (N_8479,N_6866,N_5162);
or U8480 (N_8480,N_5892,N_7053);
or U8481 (N_8481,N_6391,N_7205);
and U8482 (N_8482,N_5045,N_5563);
xnor U8483 (N_8483,N_6851,N_6819);
or U8484 (N_8484,N_6297,N_6618);
nand U8485 (N_8485,N_7353,N_6736);
nand U8486 (N_8486,N_6688,N_6200);
xnor U8487 (N_8487,N_5889,N_7266);
nor U8488 (N_8488,N_5553,N_6604);
xnor U8489 (N_8489,N_5199,N_6418);
nor U8490 (N_8490,N_5031,N_5391);
xnor U8491 (N_8491,N_5206,N_6286);
and U8492 (N_8492,N_6988,N_5378);
xor U8493 (N_8493,N_5947,N_6304);
and U8494 (N_8494,N_6275,N_5707);
and U8495 (N_8495,N_6683,N_7026);
nor U8496 (N_8496,N_7207,N_6645);
xor U8497 (N_8497,N_6974,N_5101);
xor U8498 (N_8498,N_5510,N_6687);
or U8499 (N_8499,N_5357,N_7115);
or U8500 (N_8500,N_6441,N_7200);
nor U8501 (N_8501,N_6965,N_6086);
and U8502 (N_8502,N_5733,N_5439);
nor U8503 (N_8503,N_5239,N_5694);
nand U8504 (N_8504,N_6244,N_5772);
or U8505 (N_8505,N_5900,N_6358);
nor U8506 (N_8506,N_6513,N_5556);
nand U8507 (N_8507,N_6174,N_6492);
xnor U8508 (N_8508,N_6137,N_5871);
or U8509 (N_8509,N_5231,N_5042);
nand U8510 (N_8510,N_5496,N_6796);
xor U8511 (N_8511,N_7327,N_7196);
or U8512 (N_8512,N_7355,N_7375);
xnor U8513 (N_8513,N_5024,N_6103);
nor U8514 (N_8514,N_6351,N_6266);
nor U8515 (N_8515,N_6109,N_6900);
or U8516 (N_8516,N_7497,N_6529);
or U8517 (N_8517,N_5958,N_5885);
and U8518 (N_8518,N_7300,N_5187);
xor U8519 (N_8519,N_7334,N_6525);
xnor U8520 (N_8520,N_7281,N_6287);
nor U8521 (N_8521,N_6522,N_7420);
and U8522 (N_8522,N_6901,N_5590);
xor U8523 (N_8523,N_5117,N_6017);
nor U8524 (N_8524,N_6173,N_7038);
and U8525 (N_8525,N_5282,N_5273);
or U8526 (N_8526,N_6183,N_5498);
or U8527 (N_8527,N_5127,N_6133);
nand U8528 (N_8528,N_5614,N_6278);
nor U8529 (N_8529,N_6667,N_5886);
xor U8530 (N_8530,N_5143,N_5001);
xor U8531 (N_8531,N_5297,N_5691);
nand U8532 (N_8532,N_7045,N_5246);
xnor U8533 (N_8533,N_7430,N_5456);
xor U8534 (N_8534,N_5390,N_5761);
xor U8535 (N_8535,N_6880,N_6828);
nand U8536 (N_8536,N_5336,N_6919);
xnor U8537 (N_8537,N_6853,N_7384);
or U8538 (N_8538,N_5107,N_6189);
xnor U8539 (N_8539,N_5254,N_6854);
nand U8540 (N_8540,N_5583,N_6494);
or U8541 (N_8541,N_7097,N_7418);
or U8542 (N_8542,N_6161,N_5767);
nor U8543 (N_8543,N_6057,N_5758);
xnor U8544 (N_8544,N_6874,N_5479);
and U8545 (N_8545,N_6472,N_6835);
nor U8546 (N_8546,N_7434,N_5620);
xnor U8547 (N_8547,N_5729,N_6622);
xnor U8548 (N_8548,N_6485,N_5925);
and U8549 (N_8549,N_6171,N_7122);
nand U8550 (N_8550,N_5355,N_6168);
and U8551 (N_8551,N_6852,N_7010);
nor U8552 (N_8552,N_7428,N_5879);
nand U8553 (N_8553,N_5261,N_5211);
xor U8554 (N_8554,N_5302,N_7202);
nor U8555 (N_8555,N_5663,N_5954);
and U8556 (N_8556,N_5656,N_6233);
nand U8557 (N_8557,N_7121,N_5020);
nand U8558 (N_8558,N_5679,N_7236);
and U8559 (N_8559,N_5864,N_6666);
and U8560 (N_8560,N_7268,N_6118);
nand U8561 (N_8561,N_6005,N_7465);
nor U8562 (N_8562,N_7322,N_5327);
xnor U8563 (N_8563,N_6763,N_5610);
nand U8564 (N_8564,N_6813,N_5262);
nand U8565 (N_8565,N_7044,N_5972);
and U8566 (N_8566,N_6340,N_6617);
xor U8567 (N_8567,N_5869,N_7191);
xor U8568 (N_8568,N_6941,N_6036);
xnor U8569 (N_8569,N_5992,N_5079);
nand U8570 (N_8570,N_5961,N_5731);
and U8571 (N_8571,N_7002,N_6178);
or U8572 (N_8572,N_6968,N_6532);
nor U8573 (N_8573,N_6144,N_7331);
nand U8574 (N_8574,N_6539,N_7318);
nor U8575 (N_8575,N_6401,N_6998);
and U8576 (N_8576,N_7226,N_6949);
or U8577 (N_8577,N_6943,N_5415);
or U8578 (N_8578,N_6098,N_6152);
xnor U8579 (N_8579,N_5665,N_5601);
xnor U8580 (N_8580,N_5037,N_5465);
nor U8581 (N_8581,N_7087,N_5225);
or U8582 (N_8582,N_5136,N_7271);
or U8583 (N_8583,N_6799,N_5071);
xnor U8584 (N_8584,N_5216,N_7113);
and U8585 (N_8585,N_6411,N_6273);
nand U8586 (N_8586,N_6507,N_6823);
and U8587 (N_8587,N_6734,N_6408);
and U8588 (N_8588,N_7457,N_5661);
xor U8589 (N_8589,N_6730,N_5668);
or U8590 (N_8590,N_6643,N_5634);
xor U8591 (N_8591,N_6239,N_5017);
nand U8592 (N_8592,N_5957,N_6791);
nand U8593 (N_8593,N_7456,N_6352);
or U8594 (N_8594,N_5692,N_5483);
and U8595 (N_8595,N_6216,N_5607);
nand U8596 (N_8596,N_7075,N_6537);
nor U8597 (N_8597,N_5177,N_5588);
or U8598 (N_8598,N_6928,N_5660);
xnor U8599 (N_8599,N_5586,N_7362);
xor U8600 (N_8600,N_5016,N_6665);
nand U8601 (N_8601,N_7004,N_6632);
xor U8602 (N_8602,N_7029,N_5642);
nand U8603 (N_8603,N_6065,N_6344);
nor U8604 (N_8604,N_6910,N_5655);
nor U8605 (N_8605,N_6967,N_7143);
and U8606 (N_8606,N_6605,N_6790);
or U8607 (N_8607,N_6805,N_5671);
or U8608 (N_8608,N_5857,N_5168);
xor U8609 (N_8609,N_5991,N_5153);
and U8610 (N_8610,N_6162,N_5299);
nor U8611 (N_8611,N_7225,N_6027);
or U8612 (N_8612,N_5281,N_5091);
nand U8613 (N_8613,N_5453,N_5550);
xor U8614 (N_8614,N_6435,N_5968);
xor U8615 (N_8615,N_6151,N_5158);
or U8616 (N_8616,N_5114,N_6714);
xnor U8617 (N_8617,N_5285,N_5138);
xor U8618 (N_8618,N_6253,N_6713);
xor U8619 (N_8619,N_7117,N_6292);
xor U8620 (N_8620,N_5120,N_7124);
nand U8621 (N_8621,N_5423,N_6948);
and U8622 (N_8622,N_6817,N_7417);
and U8623 (N_8623,N_6316,N_5664);
or U8624 (N_8624,N_6743,N_5145);
and U8625 (N_8625,N_6378,N_7168);
nor U8626 (N_8626,N_5360,N_5408);
xnor U8627 (N_8627,N_7438,N_5050);
xor U8628 (N_8628,N_5812,N_6878);
nor U8629 (N_8629,N_6600,N_5161);
xor U8630 (N_8630,N_5792,N_6206);
nand U8631 (N_8631,N_5683,N_5373);
nor U8632 (N_8632,N_7185,N_7012);
nand U8633 (N_8633,N_6176,N_6220);
nand U8634 (N_8634,N_5816,N_6056);
and U8635 (N_8635,N_6989,N_5719);
nor U8636 (N_8636,N_6737,N_5446);
and U8637 (N_8637,N_7160,N_7008);
or U8638 (N_8638,N_6589,N_5204);
or U8639 (N_8639,N_7475,N_6473);
nor U8640 (N_8640,N_5460,N_5472);
and U8641 (N_8641,N_6873,N_5264);
and U8642 (N_8642,N_7368,N_5927);
nand U8643 (N_8643,N_5716,N_6364);
xor U8644 (N_8644,N_6288,N_7373);
nor U8645 (N_8645,N_7370,N_6561);
or U8646 (N_8646,N_5435,N_7007);
xnor U8647 (N_8647,N_6527,N_5625);
and U8648 (N_8648,N_7108,N_5480);
or U8649 (N_8649,N_5149,N_5087);
or U8650 (N_8650,N_6861,N_6191);
or U8651 (N_8651,N_6896,N_5743);
and U8652 (N_8652,N_5529,N_6336);
xor U8653 (N_8653,N_6365,N_5226);
xor U8654 (N_8654,N_7259,N_5308);
and U8655 (N_8655,N_6295,N_5369);
and U8656 (N_8656,N_7358,N_5165);
and U8657 (N_8657,N_6658,N_5250);
nor U8658 (N_8658,N_5921,N_5935);
xnor U8659 (N_8659,N_5040,N_5359);
or U8660 (N_8660,N_5599,N_6298);
nor U8661 (N_8661,N_7098,N_5236);
or U8662 (N_8662,N_6143,N_6980);
nor U8663 (N_8663,N_5135,N_5766);
xor U8664 (N_8664,N_5571,N_6208);
and U8665 (N_8665,N_7405,N_5776);
or U8666 (N_8666,N_7245,N_7169);
or U8667 (N_8667,N_7231,N_7209);
and U8668 (N_8668,N_6131,N_7396);
nand U8669 (N_8669,N_5030,N_6134);
xor U8670 (N_8670,N_6258,N_5272);
nor U8671 (N_8671,N_6374,N_5406);
and U8672 (N_8672,N_5110,N_5215);
nand U8673 (N_8673,N_5146,N_6519);
and U8674 (N_8674,N_5675,N_5875);
or U8675 (N_8675,N_7458,N_6789);
nand U8676 (N_8676,N_6576,N_6190);
nor U8677 (N_8677,N_5912,N_5041);
and U8678 (N_8678,N_5347,N_5948);
and U8679 (N_8679,N_7088,N_7487);
nand U8680 (N_8680,N_5054,N_5615);
and U8681 (N_8681,N_6070,N_6905);
nor U8682 (N_8682,N_6506,N_5723);
xnor U8683 (N_8683,N_6263,N_6584);
xor U8684 (N_8684,N_6703,N_5860);
nand U8685 (N_8685,N_5839,N_7074);
and U8686 (N_8686,N_5156,N_6814);
xnor U8687 (N_8687,N_6690,N_7496);
nand U8688 (N_8688,N_6269,N_5304);
and U8689 (N_8689,N_6062,N_5418);
nand U8690 (N_8690,N_6816,N_5147);
nor U8691 (N_8691,N_7105,N_7243);
and U8692 (N_8692,N_6006,N_5650);
nand U8693 (N_8693,N_5924,N_7422);
or U8694 (N_8694,N_5436,N_6975);
or U8695 (N_8695,N_6959,N_5778);
xor U8696 (N_8696,N_6761,N_5534);
xnor U8697 (N_8697,N_6840,N_5786);
or U8698 (N_8698,N_6871,N_6040);
and U8699 (N_8699,N_5568,N_6678);
and U8700 (N_8700,N_5473,N_5997);
nand U8701 (N_8701,N_5076,N_6867);
nor U8702 (N_8702,N_6484,N_6283);
nand U8703 (N_8703,N_6071,N_6652);
xnor U8704 (N_8704,N_5903,N_5195);
nor U8705 (N_8705,N_5773,N_5989);
nor U8706 (N_8706,N_7424,N_7307);
or U8707 (N_8707,N_5643,N_5292);
and U8708 (N_8708,N_6554,N_5021);
or U8709 (N_8709,N_6885,N_5253);
xor U8710 (N_8710,N_5562,N_6427);
nor U8711 (N_8711,N_6942,N_6757);
xnor U8712 (N_8712,N_6553,N_5978);
xor U8713 (N_8713,N_6781,N_7130);
or U8714 (N_8714,N_6022,N_5445);
or U8715 (N_8715,N_7401,N_6249);
nand U8716 (N_8716,N_5014,N_6912);
and U8717 (N_8717,N_6785,N_7238);
nor U8718 (N_8718,N_5951,N_7077);
nand U8719 (N_8719,N_7392,N_5652);
xnor U8720 (N_8720,N_5637,N_6332);
nand U8721 (N_8721,N_6932,N_6136);
nor U8722 (N_8722,N_5382,N_5203);
xor U8723 (N_8723,N_5785,N_5657);
and U8724 (N_8724,N_5294,N_5752);
or U8725 (N_8725,N_6353,N_5269);
and U8726 (N_8726,N_7234,N_5745);
or U8727 (N_8727,N_6535,N_5414);
or U8728 (N_8728,N_6839,N_6843);
xor U8729 (N_8729,N_5493,N_7256);
and U8730 (N_8730,N_6135,N_7015);
and U8731 (N_8731,N_6541,N_6025);
xnor U8732 (N_8732,N_6540,N_5922);
xor U8733 (N_8733,N_6034,N_5089);
nor U8734 (N_8734,N_6095,N_5495);
xnor U8735 (N_8735,N_6608,N_5645);
nor U8736 (N_8736,N_6318,N_5242);
and U8737 (N_8737,N_7027,N_6129);
nor U8738 (N_8738,N_5092,N_6935);
nand U8739 (N_8739,N_5475,N_5732);
and U8740 (N_8740,N_6238,N_7052);
nor U8741 (N_8741,N_6222,N_5627);
and U8742 (N_8742,N_5332,N_6061);
nand U8743 (N_8743,N_7136,N_5676);
nor U8744 (N_8744,N_6274,N_6774);
nand U8745 (N_8745,N_5783,N_6021);
and U8746 (N_8746,N_7391,N_6436);
nand U8747 (N_8747,N_6549,N_7019);
and U8748 (N_8748,N_5751,N_7441);
nand U8749 (N_8749,N_6121,N_6917);
or U8750 (N_8750,N_6375,N_5051);
and U8751 (N_8751,N_5890,N_5902);
or U8752 (N_8752,N_6494,N_7095);
xor U8753 (N_8753,N_7102,N_6789);
and U8754 (N_8754,N_7416,N_5939);
xnor U8755 (N_8755,N_6656,N_7329);
xor U8756 (N_8756,N_6128,N_5307);
nor U8757 (N_8757,N_5345,N_6062);
xnor U8758 (N_8758,N_7241,N_6651);
or U8759 (N_8759,N_5705,N_6190);
nor U8760 (N_8760,N_5578,N_6830);
nor U8761 (N_8761,N_5457,N_5490);
nand U8762 (N_8762,N_6979,N_7321);
nor U8763 (N_8763,N_7237,N_5674);
or U8764 (N_8764,N_5138,N_6881);
and U8765 (N_8765,N_5762,N_6719);
xor U8766 (N_8766,N_5673,N_5832);
nor U8767 (N_8767,N_6620,N_5024);
nor U8768 (N_8768,N_5314,N_6478);
nor U8769 (N_8769,N_5503,N_5009);
nor U8770 (N_8770,N_5780,N_5455);
nor U8771 (N_8771,N_6195,N_7276);
and U8772 (N_8772,N_6255,N_5854);
nor U8773 (N_8773,N_5979,N_7129);
nand U8774 (N_8774,N_6280,N_5552);
or U8775 (N_8775,N_7196,N_5078);
xor U8776 (N_8776,N_7242,N_5213);
and U8777 (N_8777,N_6880,N_5239);
and U8778 (N_8778,N_6588,N_7247);
nand U8779 (N_8779,N_6663,N_6038);
nor U8780 (N_8780,N_5896,N_6675);
and U8781 (N_8781,N_7378,N_7218);
nor U8782 (N_8782,N_6224,N_6952);
xor U8783 (N_8783,N_6939,N_6279);
xnor U8784 (N_8784,N_6946,N_7399);
and U8785 (N_8785,N_6849,N_5611);
nand U8786 (N_8786,N_5350,N_7119);
xor U8787 (N_8787,N_6559,N_6299);
nand U8788 (N_8788,N_6241,N_6685);
nand U8789 (N_8789,N_5531,N_5278);
nand U8790 (N_8790,N_5499,N_6035);
and U8791 (N_8791,N_5548,N_5056);
xnor U8792 (N_8792,N_5404,N_5190);
nand U8793 (N_8793,N_5759,N_7467);
nand U8794 (N_8794,N_5877,N_5518);
nor U8795 (N_8795,N_5487,N_6312);
and U8796 (N_8796,N_7423,N_7400);
and U8797 (N_8797,N_7248,N_6633);
nand U8798 (N_8798,N_5253,N_5912);
xor U8799 (N_8799,N_7010,N_5574);
nor U8800 (N_8800,N_5594,N_5478);
or U8801 (N_8801,N_6824,N_6219);
nor U8802 (N_8802,N_6508,N_6050);
xnor U8803 (N_8803,N_5898,N_5341);
or U8804 (N_8804,N_6859,N_7240);
xnor U8805 (N_8805,N_6863,N_7353);
and U8806 (N_8806,N_5142,N_7008);
xor U8807 (N_8807,N_5261,N_7259);
nand U8808 (N_8808,N_6976,N_7271);
and U8809 (N_8809,N_7431,N_5026);
nand U8810 (N_8810,N_5315,N_6088);
and U8811 (N_8811,N_5070,N_6217);
nand U8812 (N_8812,N_6000,N_6217);
xor U8813 (N_8813,N_6708,N_6033);
or U8814 (N_8814,N_7315,N_6787);
xnor U8815 (N_8815,N_5382,N_5747);
or U8816 (N_8816,N_6596,N_5228);
nand U8817 (N_8817,N_6000,N_5395);
nand U8818 (N_8818,N_7460,N_6344);
and U8819 (N_8819,N_6056,N_6747);
nor U8820 (N_8820,N_6619,N_6258);
nor U8821 (N_8821,N_5358,N_6581);
or U8822 (N_8822,N_7164,N_5738);
xnor U8823 (N_8823,N_5766,N_6649);
or U8824 (N_8824,N_5112,N_6115);
nand U8825 (N_8825,N_5986,N_5419);
nor U8826 (N_8826,N_7253,N_6049);
or U8827 (N_8827,N_7346,N_7055);
nand U8828 (N_8828,N_6449,N_6825);
nor U8829 (N_8829,N_5810,N_5388);
nand U8830 (N_8830,N_7239,N_6904);
nor U8831 (N_8831,N_5145,N_5682);
and U8832 (N_8832,N_6127,N_5816);
nor U8833 (N_8833,N_5103,N_6425);
xnor U8834 (N_8834,N_5778,N_6700);
nand U8835 (N_8835,N_6131,N_7156);
xor U8836 (N_8836,N_5103,N_5526);
and U8837 (N_8837,N_6894,N_6586);
nor U8838 (N_8838,N_6366,N_5472);
xnor U8839 (N_8839,N_7264,N_5946);
or U8840 (N_8840,N_7374,N_7474);
or U8841 (N_8841,N_7431,N_7430);
nor U8842 (N_8842,N_5324,N_6280);
or U8843 (N_8843,N_6205,N_6521);
nor U8844 (N_8844,N_6267,N_5260);
or U8845 (N_8845,N_7368,N_5595);
and U8846 (N_8846,N_5203,N_5742);
xnor U8847 (N_8847,N_7127,N_7185);
nand U8848 (N_8848,N_5971,N_6873);
and U8849 (N_8849,N_7456,N_6220);
nor U8850 (N_8850,N_7361,N_7019);
nand U8851 (N_8851,N_6066,N_5824);
or U8852 (N_8852,N_5635,N_6267);
nand U8853 (N_8853,N_6933,N_5872);
or U8854 (N_8854,N_5886,N_6537);
xnor U8855 (N_8855,N_5826,N_7389);
or U8856 (N_8856,N_6479,N_5881);
and U8857 (N_8857,N_5750,N_7498);
nand U8858 (N_8858,N_6901,N_6111);
and U8859 (N_8859,N_7475,N_6842);
and U8860 (N_8860,N_5286,N_7035);
and U8861 (N_8861,N_7285,N_6038);
nand U8862 (N_8862,N_5043,N_5746);
xnor U8863 (N_8863,N_6394,N_7470);
xor U8864 (N_8864,N_5264,N_5909);
and U8865 (N_8865,N_5255,N_5457);
nand U8866 (N_8866,N_6928,N_7433);
or U8867 (N_8867,N_6202,N_7480);
nand U8868 (N_8868,N_5079,N_5246);
nor U8869 (N_8869,N_5405,N_5935);
and U8870 (N_8870,N_6887,N_5785);
and U8871 (N_8871,N_5003,N_5826);
xnor U8872 (N_8872,N_6114,N_5460);
nor U8873 (N_8873,N_6759,N_5856);
nor U8874 (N_8874,N_6871,N_5043);
or U8875 (N_8875,N_6730,N_6996);
nand U8876 (N_8876,N_6753,N_5591);
or U8877 (N_8877,N_6577,N_6110);
nand U8878 (N_8878,N_6451,N_6472);
nand U8879 (N_8879,N_6739,N_7474);
nand U8880 (N_8880,N_7034,N_6760);
xor U8881 (N_8881,N_6485,N_5396);
or U8882 (N_8882,N_7087,N_5142);
nor U8883 (N_8883,N_7368,N_6118);
nor U8884 (N_8884,N_6504,N_5605);
nor U8885 (N_8885,N_5812,N_5886);
nor U8886 (N_8886,N_6704,N_6143);
xnor U8887 (N_8887,N_6940,N_6364);
or U8888 (N_8888,N_5523,N_6341);
nand U8889 (N_8889,N_5992,N_6368);
nor U8890 (N_8890,N_7001,N_5431);
xor U8891 (N_8891,N_5530,N_5341);
nand U8892 (N_8892,N_7380,N_6415);
nor U8893 (N_8893,N_5631,N_5039);
and U8894 (N_8894,N_6685,N_6938);
xor U8895 (N_8895,N_7402,N_6849);
xnor U8896 (N_8896,N_7477,N_5947);
xor U8897 (N_8897,N_7119,N_7494);
and U8898 (N_8898,N_6976,N_6360);
or U8899 (N_8899,N_5521,N_7368);
xor U8900 (N_8900,N_6932,N_5410);
and U8901 (N_8901,N_5520,N_5781);
xnor U8902 (N_8902,N_5449,N_7399);
or U8903 (N_8903,N_7002,N_6025);
xor U8904 (N_8904,N_5256,N_5884);
nand U8905 (N_8905,N_5827,N_7151);
nor U8906 (N_8906,N_6443,N_5417);
nor U8907 (N_8907,N_7461,N_6918);
nor U8908 (N_8908,N_7352,N_5730);
xnor U8909 (N_8909,N_5788,N_6085);
nor U8910 (N_8910,N_5297,N_5301);
and U8911 (N_8911,N_7143,N_5946);
nor U8912 (N_8912,N_5637,N_6239);
or U8913 (N_8913,N_6105,N_6912);
nand U8914 (N_8914,N_5636,N_6168);
and U8915 (N_8915,N_5650,N_6353);
and U8916 (N_8916,N_6622,N_6253);
nor U8917 (N_8917,N_5547,N_6562);
nand U8918 (N_8918,N_6297,N_7212);
xnor U8919 (N_8919,N_5967,N_5567);
and U8920 (N_8920,N_6560,N_6352);
nor U8921 (N_8921,N_5035,N_5376);
nand U8922 (N_8922,N_5615,N_6186);
nand U8923 (N_8923,N_6608,N_6336);
xnor U8924 (N_8924,N_5545,N_5325);
or U8925 (N_8925,N_5025,N_5187);
xor U8926 (N_8926,N_7389,N_5559);
and U8927 (N_8927,N_7055,N_7062);
nor U8928 (N_8928,N_7152,N_5678);
xor U8929 (N_8929,N_6704,N_6461);
nand U8930 (N_8930,N_6496,N_6167);
or U8931 (N_8931,N_7183,N_7424);
xor U8932 (N_8932,N_5027,N_6091);
nand U8933 (N_8933,N_6920,N_6462);
nor U8934 (N_8934,N_7327,N_6552);
or U8935 (N_8935,N_5265,N_5283);
or U8936 (N_8936,N_7240,N_7012);
or U8937 (N_8937,N_7430,N_5727);
nor U8938 (N_8938,N_7258,N_5534);
or U8939 (N_8939,N_6829,N_5632);
or U8940 (N_8940,N_7431,N_5959);
nor U8941 (N_8941,N_5190,N_7279);
and U8942 (N_8942,N_7438,N_5922);
nor U8943 (N_8943,N_6684,N_6325);
and U8944 (N_8944,N_6034,N_6261);
nand U8945 (N_8945,N_5203,N_6734);
or U8946 (N_8946,N_5243,N_5700);
or U8947 (N_8947,N_7247,N_6366);
nand U8948 (N_8948,N_7248,N_6333);
nor U8949 (N_8949,N_5991,N_6418);
nor U8950 (N_8950,N_7081,N_7470);
and U8951 (N_8951,N_5248,N_6606);
xnor U8952 (N_8952,N_5705,N_5332);
and U8953 (N_8953,N_7355,N_7149);
or U8954 (N_8954,N_5258,N_5380);
nand U8955 (N_8955,N_5718,N_7103);
or U8956 (N_8956,N_5519,N_5315);
xnor U8957 (N_8957,N_5064,N_6568);
and U8958 (N_8958,N_6643,N_6969);
or U8959 (N_8959,N_6486,N_5717);
nand U8960 (N_8960,N_6029,N_6216);
and U8961 (N_8961,N_6602,N_5220);
or U8962 (N_8962,N_6441,N_5899);
xor U8963 (N_8963,N_7040,N_6077);
or U8964 (N_8964,N_6884,N_7128);
nor U8965 (N_8965,N_5490,N_7215);
nand U8966 (N_8966,N_7069,N_6422);
nand U8967 (N_8967,N_5997,N_7307);
nand U8968 (N_8968,N_6034,N_5500);
nand U8969 (N_8969,N_5119,N_7118);
nor U8970 (N_8970,N_6319,N_7147);
nor U8971 (N_8971,N_5440,N_6004);
nand U8972 (N_8972,N_5669,N_7244);
xor U8973 (N_8973,N_5304,N_6863);
nor U8974 (N_8974,N_6246,N_5727);
xnor U8975 (N_8975,N_6712,N_5436);
nand U8976 (N_8976,N_6477,N_7209);
nor U8977 (N_8977,N_6187,N_6783);
and U8978 (N_8978,N_6033,N_5832);
and U8979 (N_8979,N_7314,N_5452);
nand U8980 (N_8980,N_6424,N_5293);
xor U8981 (N_8981,N_6875,N_6812);
and U8982 (N_8982,N_6340,N_6684);
and U8983 (N_8983,N_5758,N_5739);
nor U8984 (N_8984,N_6258,N_5301);
and U8985 (N_8985,N_5759,N_7114);
nand U8986 (N_8986,N_6116,N_7230);
and U8987 (N_8987,N_7075,N_5373);
xor U8988 (N_8988,N_5283,N_5028);
nor U8989 (N_8989,N_5323,N_6431);
nand U8990 (N_8990,N_7397,N_5765);
nor U8991 (N_8991,N_5465,N_7142);
nor U8992 (N_8992,N_6199,N_6699);
or U8993 (N_8993,N_7371,N_6717);
and U8994 (N_8994,N_7059,N_5683);
xor U8995 (N_8995,N_6010,N_7184);
nand U8996 (N_8996,N_6386,N_5710);
xor U8997 (N_8997,N_6745,N_5593);
nand U8998 (N_8998,N_5893,N_6069);
nand U8999 (N_8999,N_5885,N_6382);
or U9000 (N_9000,N_7457,N_6205);
nor U9001 (N_9001,N_5132,N_5944);
nand U9002 (N_9002,N_6199,N_5705);
or U9003 (N_9003,N_6665,N_7154);
xnor U9004 (N_9004,N_5040,N_6081);
nor U9005 (N_9005,N_6915,N_6253);
nand U9006 (N_9006,N_6886,N_5174);
nor U9007 (N_9007,N_6086,N_6108);
nand U9008 (N_9008,N_5930,N_5631);
nand U9009 (N_9009,N_7208,N_5936);
nand U9010 (N_9010,N_6494,N_6241);
and U9011 (N_9011,N_6379,N_6287);
nor U9012 (N_9012,N_7205,N_5829);
nor U9013 (N_9013,N_6657,N_6344);
nand U9014 (N_9014,N_5023,N_7065);
xor U9015 (N_9015,N_5132,N_5285);
nand U9016 (N_9016,N_6855,N_5075);
and U9017 (N_9017,N_6379,N_6047);
xnor U9018 (N_9018,N_7093,N_7379);
xor U9019 (N_9019,N_7134,N_6868);
or U9020 (N_9020,N_7148,N_6134);
xor U9021 (N_9021,N_6438,N_7284);
nor U9022 (N_9022,N_6850,N_5967);
xnor U9023 (N_9023,N_6282,N_7443);
or U9024 (N_9024,N_5038,N_6813);
or U9025 (N_9025,N_6425,N_6482);
xnor U9026 (N_9026,N_7363,N_7268);
nor U9027 (N_9027,N_5910,N_6586);
nand U9028 (N_9028,N_5251,N_6991);
nor U9029 (N_9029,N_7347,N_5545);
nor U9030 (N_9030,N_6861,N_5114);
and U9031 (N_9031,N_7324,N_7402);
nand U9032 (N_9032,N_6329,N_7017);
or U9033 (N_9033,N_5140,N_6029);
nor U9034 (N_9034,N_7297,N_6781);
or U9035 (N_9035,N_7269,N_7417);
or U9036 (N_9036,N_5048,N_5091);
xnor U9037 (N_9037,N_5308,N_5269);
nand U9038 (N_9038,N_7003,N_7138);
nor U9039 (N_9039,N_6124,N_6343);
xnor U9040 (N_9040,N_6442,N_5633);
nand U9041 (N_9041,N_5382,N_7059);
xnor U9042 (N_9042,N_6438,N_5259);
and U9043 (N_9043,N_7283,N_6717);
nand U9044 (N_9044,N_6905,N_5715);
nor U9045 (N_9045,N_5499,N_5018);
and U9046 (N_9046,N_6709,N_6881);
and U9047 (N_9047,N_7250,N_6297);
nor U9048 (N_9048,N_6655,N_6816);
nor U9049 (N_9049,N_7087,N_5067);
xnor U9050 (N_9050,N_6548,N_7462);
and U9051 (N_9051,N_7108,N_6777);
nor U9052 (N_9052,N_6796,N_6362);
nand U9053 (N_9053,N_5894,N_5304);
nand U9054 (N_9054,N_6340,N_5687);
nand U9055 (N_9055,N_5869,N_5202);
xnor U9056 (N_9056,N_5421,N_6848);
xnor U9057 (N_9057,N_6936,N_7224);
and U9058 (N_9058,N_5640,N_6469);
and U9059 (N_9059,N_6106,N_5465);
xor U9060 (N_9060,N_6819,N_6896);
nand U9061 (N_9061,N_5330,N_6025);
and U9062 (N_9062,N_6442,N_5920);
xnor U9063 (N_9063,N_6090,N_5163);
nand U9064 (N_9064,N_7151,N_6546);
nor U9065 (N_9065,N_5411,N_7366);
and U9066 (N_9066,N_6050,N_7009);
nor U9067 (N_9067,N_5725,N_6152);
nor U9068 (N_9068,N_6584,N_7123);
nand U9069 (N_9069,N_5742,N_7019);
and U9070 (N_9070,N_6093,N_6285);
or U9071 (N_9071,N_7113,N_7298);
nor U9072 (N_9072,N_6697,N_7409);
and U9073 (N_9073,N_5607,N_6250);
or U9074 (N_9074,N_7472,N_6607);
nand U9075 (N_9075,N_5130,N_5218);
nor U9076 (N_9076,N_5930,N_7007);
or U9077 (N_9077,N_7086,N_6147);
nor U9078 (N_9078,N_6262,N_7397);
xnor U9079 (N_9079,N_6356,N_5058);
or U9080 (N_9080,N_6476,N_6155);
nor U9081 (N_9081,N_5833,N_6688);
nor U9082 (N_9082,N_5205,N_5703);
xor U9083 (N_9083,N_6050,N_6046);
and U9084 (N_9084,N_5949,N_6408);
xor U9085 (N_9085,N_6691,N_6054);
or U9086 (N_9086,N_5215,N_6847);
and U9087 (N_9087,N_5855,N_6455);
and U9088 (N_9088,N_6968,N_7268);
or U9089 (N_9089,N_6382,N_6401);
and U9090 (N_9090,N_5333,N_5809);
or U9091 (N_9091,N_6455,N_5054);
or U9092 (N_9092,N_6706,N_6738);
xnor U9093 (N_9093,N_7214,N_6898);
or U9094 (N_9094,N_6902,N_6099);
nor U9095 (N_9095,N_5667,N_6812);
and U9096 (N_9096,N_6217,N_7164);
xor U9097 (N_9097,N_6526,N_6430);
nand U9098 (N_9098,N_5420,N_5363);
nor U9099 (N_9099,N_6334,N_5830);
nor U9100 (N_9100,N_6608,N_6883);
xnor U9101 (N_9101,N_5029,N_6503);
and U9102 (N_9102,N_5647,N_5843);
or U9103 (N_9103,N_5784,N_6583);
and U9104 (N_9104,N_7353,N_5069);
nand U9105 (N_9105,N_5106,N_6916);
xor U9106 (N_9106,N_6671,N_6458);
or U9107 (N_9107,N_6475,N_7411);
xor U9108 (N_9108,N_7118,N_5805);
xnor U9109 (N_9109,N_6245,N_6833);
and U9110 (N_9110,N_5443,N_5033);
xor U9111 (N_9111,N_6532,N_5080);
xnor U9112 (N_9112,N_5509,N_6054);
and U9113 (N_9113,N_6431,N_6434);
or U9114 (N_9114,N_5822,N_5493);
nor U9115 (N_9115,N_5229,N_6488);
nor U9116 (N_9116,N_5799,N_6318);
and U9117 (N_9117,N_5211,N_7230);
or U9118 (N_9118,N_7167,N_6009);
nor U9119 (N_9119,N_6387,N_6141);
xnor U9120 (N_9120,N_7042,N_5235);
and U9121 (N_9121,N_5506,N_7368);
and U9122 (N_9122,N_5206,N_5528);
nand U9123 (N_9123,N_5059,N_5451);
nand U9124 (N_9124,N_6273,N_6452);
and U9125 (N_9125,N_5268,N_7000);
xnor U9126 (N_9126,N_7223,N_6510);
nand U9127 (N_9127,N_5919,N_6905);
and U9128 (N_9128,N_6866,N_5527);
xor U9129 (N_9129,N_5039,N_6549);
and U9130 (N_9130,N_7034,N_5651);
nor U9131 (N_9131,N_7210,N_5309);
and U9132 (N_9132,N_5227,N_6563);
nor U9133 (N_9133,N_7351,N_7103);
nor U9134 (N_9134,N_5308,N_6695);
and U9135 (N_9135,N_5661,N_7370);
nand U9136 (N_9136,N_5354,N_5549);
and U9137 (N_9137,N_7224,N_7125);
xor U9138 (N_9138,N_5882,N_7427);
nand U9139 (N_9139,N_7189,N_6565);
and U9140 (N_9140,N_5932,N_5565);
nand U9141 (N_9141,N_6838,N_5270);
xor U9142 (N_9142,N_5461,N_5195);
nand U9143 (N_9143,N_7084,N_5844);
or U9144 (N_9144,N_5378,N_5848);
xor U9145 (N_9145,N_6669,N_6949);
and U9146 (N_9146,N_7078,N_7386);
nand U9147 (N_9147,N_7407,N_5960);
nor U9148 (N_9148,N_6946,N_7389);
or U9149 (N_9149,N_5933,N_5420);
xor U9150 (N_9150,N_6297,N_7040);
or U9151 (N_9151,N_6713,N_7026);
xnor U9152 (N_9152,N_6849,N_5158);
nand U9153 (N_9153,N_5566,N_5894);
or U9154 (N_9154,N_6745,N_6946);
nor U9155 (N_9155,N_5758,N_5744);
nand U9156 (N_9156,N_6071,N_6283);
nor U9157 (N_9157,N_5791,N_6462);
and U9158 (N_9158,N_6919,N_5026);
and U9159 (N_9159,N_5621,N_5980);
or U9160 (N_9160,N_6395,N_5875);
and U9161 (N_9161,N_7489,N_6995);
nor U9162 (N_9162,N_5477,N_7121);
and U9163 (N_9163,N_6762,N_5407);
xor U9164 (N_9164,N_5260,N_6357);
xnor U9165 (N_9165,N_5954,N_6950);
and U9166 (N_9166,N_6758,N_6918);
nand U9167 (N_9167,N_7430,N_6474);
nand U9168 (N_9168,N_6392,N_5788);
nand U9169 (N_9169,N_5161,N_7313);
xor U9170 (N_9170,N_5256,N_7362);
or U9171 (N_9171,N_6074,N_7265);
or U9172 (N_9172,N_6418,N_5339);
nand U9173 (N_9173,N_5850,N_5863);
and U9174 (N_9174,N_6703,N_5973);
xor U9175 (N_9175,N_6722,N_6441);
nand U9176 (N_9176,N_6779,N_5947);
nand U9177 (N_9177,N_5517,N_7109);
and U9178 (N_9178,N_7099,N_5824);
xor U9179 (N_9179,N_6305,N_7098);
or U9180 (N_9180,N_7318,N_6376);
nor U9181 (N_9181,N_5362,N_5947);
nand U9182 (N_9182,N_6726,N_6576);
xnor U9183 (N_9183,N_6258,N_7072);
and U9184 (N_9184,N_5972,N_5866);
nor U9185 (N_9185,N_6135,N_5736);
xor U9186 (N_9186,N_5860,N_5493);
xnor U9187 (N_9187,N_6123,N_6762);
nand U9188 (N_9188,N_7425,N_6781);
or U9189 (N_9189,N_7253,N_7190);
xnor U9190 (N_9190,N_5604,N_6175);
and U9191 (N_9191,N_5682,N_6949);
xor U9192 (N_9192,N_5531,N_6774);
nand U9193 (N_9193,N_5951,N_6029);
nor U9194 (N_9194,N_6497,N_5343);
nor U9195 (N_9195,N_7168,N_6249);
and U9196 (N_9196,N_6317,N_5435);
nand U9197 (N_9197,N_5087,N_5121);
xor U9198 (N_9198,N_5328,N_6228);
nand U9199 (N_9199,N_6328,N_6071);
nor U9200 (N_9200,N_6802,N_7207);
nand U9201 (N_9201,N_7091,N_5847);
nor U9202 (N_9202,N_6861,N_5662);
nand U9203 (N_9203,N_7071,N_5882);
or U9204 (N_9204,N_6882,N_5795);
xor U9205 (N_9205,N_6163,N_6463);
and U9206 (N_9206,N_5020,N_6871);
nor U9207 (N_9207,N_5796,N_5791);
xor U9208 (N_9208,N_6770,N_6581);
nand U9209 (N_9209,N_6390,N_6876);
and U9210 (N_9210,N_5379,N_6763);
nor U9211 (N_9211,N_7244,N_6235);
xor U9212 (N_9212,N_5024,N_5427);
nand U9213 (N_9213,N_6590,N_6021);
and U9214 (N_9214,N_5361,N_5252);
nor U9215 (N_9215,N_5175,N_5700);
nand U9216 (N_9216,N_6726,N_5073);
and U9217 (N_9217,N_6214,N_7274);
xor U9218 (N_9218,N_5404,N_6032);
xor U9219 (N_9219,N_5656,N_7170);
or U9220 (N_9220,N_7038,N_7234);
or U9221 (N_9221,N_6370,N_6432);
nand U9222 (N_9222,N_5816,N_6752);
nor U9223 (N_9223,N_7258,N_6241);
xor U9224 (N_9224,N_7010,N_5406);
xor U9225 (N_9225,N_6563,N_7063);
and U9226 (N_9226,N_6773,N_5768);
nand U9227 (N_9227,N_5649,N_5348);
xor U9228 (N_9228,N_5313,N_6862);
nor U9229 (N_9229,N_6841,N_5815);
and U9230 (N_9230,N_7339,N_6528);
and U9231 (N_9231,N_6547,N_5844);
xor U9232 (N_9232,N_6211,N_7422);
or U9233 (N_9233,N_7234,N_5129);
nand U9234 (N_9234,N_7345,N_5370);
nor U9235 (N_9235,N_6788,N_5641);
nor U9236 (N_9236,N_7274,N_6345);
nand U9237 (N_9237,N_7215,N_5945);
nand U9238 (N_9238,N_5374,N_7226);
nand U9239 (N_9239,N_5174,N_6927);
and U9240 (N_9240,N_6266,N_7407);
xnor U9241 (N_9241,N_6820,N_6466);
nor U9242 (N_9242,N_6443,N_5268);
xor U9243 (N_9243,N_5274,N_6059);
or U9244 (N_9244,N_5010,N_5279);
or U9245 (N_9245,N_6386,N_6879);
or U9246 (N_9246,N_5057,N_5889);
and U9247 (N_9247,N_5041,N_7343);
or U9248 (N_9248,N_5040,N_6922);
and U9249 (N_9249,N_5321,N_6488);
xnor U9250 (N_9250,N_5725,N_6386);
and U9251 (N_9251,N_7066,N_6737);
nand U9252 (N_9252,N_5131,N_5069);
xnor U9253 (N_9253,N_7071,N_7308);
nand U9254 (N_9254,N_6188,N_5340);
nand U9255 (N_9255,N_5821,N_6970);
xnor U9256 (N_9256,N_5721,N_7492);
or U9257 (N_9257,N_6184,N_5756);
and U9258 (N_9258,N_5303,N_5686);
nand U9259 (N_9259,N_7250,N_5879);
nor U9260 (N_9260,N_7083,N_6974);
xor U9261 (N_9261,N_6072,N_5581);
or U9262 (N_9262,N_6345,N_6025);
nand U9263 (N_9263,N_5543,N_5417);
nand U9264 (N_9264,N_7016,N_6547);
nor U9265 (N_9265,N_6190,N_6550);
xor U9266 (N_9266,N_6077,N_6388);
xor U9267 (N_9267,N_7466,N_7181);
nand U9268 (N_9268,N_6962,N_6752);
nand U9269 (N_9269,N_6845,N_7398);
or U9270 (N_9270,N_5512,N_6571);
and U9271 (N_9271,N_5017,N_7447);
and U9272 (N_9272,N_7402,N_6266);
xnor U9273 (N_9273,N_6218,N_6596);
or U9274 (N_9274,N_5917,N_7319);
or U9275 (N_9275,N_6533,N_6637);
and U9276 (N_9276,N_6544,N_6066);
nand U9277 (N_9277,N_5094,N_7308);
nand U9278 (N_9278,N_6533,N_5091);
nor U9279 (N_9279,N_5883,N_6226);
and U9280 (N_9280,N_5083,N_5294);
or U9281 (N_9281,N_6402,N_5142);
and U9282 (N_9282,N_5566,N_7276);
or U9283 (N_9283,N_7458,N_7298);
xor U9284 (N_9284,N_5052,N_7018);
and U9285 (N_9285,N_6248,N_6487);
and U9286 (N_9286,N_5873,N_5448);
xor U9287 (N_9287,N_6570,N_6057);
xor U9288 (N_9288,N_7341,N_5569);
nor U9289 (N_9289,N_6017,N_5413);
or U9290 (N_9290,N_6480,N_6175);
nand U9291 (N_9291,N_6388,N_6452);
nand U9292 (N_9292,N_7236,N_5077);
and U9293 (N_9293,N_5929,N_6228);
nor U9294 (N_9294,N_5767,N_5563);
and U9295 (N_9295,N_6199,N_5315);
xnor U9296 (N_9296,N_5466,N_7138);
and U9297 (N_9297,N_5145,N_5987);
and U9298 (N_9298,N_7476,N_6457);
and U9299 (N_9299,N_5559,N_6973);
and U9300 (N_9300,N_6950,N_7116);
or U9301 (N_9301,N_6082,N_6167);
and U9302 (N_9302,N_7253,N_5346);
nand U9303 (N_9303,N_5988,N_6578);
nor U9304 (N_9304,N_5037,N_7387);
and U9305 (N_9305,N_5853,N_6711);
or U9306 (N_9306,N_6481,N_5832);
xor U9307 (N_9307,N_6947,N_6920);
xor U9308 (N_9308,N_6133,N_7005);
or U9309 (N_9309,N_6268,N_7300);
xnor U9310 (N_9310,N_6948,N_6906);
or U9311 (N_9311,N_5906,N_6778);
nand U9312 (N_9312,N_7432,N_6900);
xor U9313 (N_9313,N_5283,N_7445);
nand U9314 (N_9314,N_6675,N_6692);
and U9315 (N_9315,N_5831,N_5867);
xnor U9316 (N_9316,N_5979,N_7338);
nor U9317 (N_9317,N_6300,N_6692);
nor U9318 (N_9318,N_6241,N_6509);
nand U9319 (N_9319,N_5628,N_5939);
and U9320 (N_9320,N_5163,N_5531);
xor U9321 (N_9321,N_6396,N_6658);
or U9322 (N_9322,N_6436,N_6950);
nand U9323 (N_9323,N_7487,N_7234);
or U9324 (N_9324,N_5233,N_7465);
and U9325 (N_9325,N_5005,N_6277);
or U9326 (N_9326,N_7028,N_5185);
xor U9327 (N_9327,N_6403,N_5673);
nor U9328 (N_9328,N_6711,N_7439);
nand U9329 (N_9329,N_5402,N_6753);
and U9330 (N_9330,N_6875,N_5068);
xnor U9331 (N_9331,N_5246,N_6478);
or U9332 (N_9332,N_5664,N_5966);
or U9333 (N_9333,N_5150,N_7346);
xnor U9334 (N_9334,N_5263,N_7446);
nor U9335 (N_9335,N_5589,N_5827);
or U9336 (N_9336,N_6204,N_6817);
xor U9337 (N_9337,N_5916,N_6451);
or U9338 (N_9338,N_7294,N_5423);
xor U9339 (N_9339,N_6547,N_6015);
xnor U9340 (N_9340,N_5660,N_5835);
or U9341 (N_9341,N_5775,N_5565);
or U9342 (N_9342,N_7180,N_5282);
and U9343 (N_9343,N_5755,N_5295);
nand U9344 (N_9344,N_5967,N_5986);
or U9345 (N_9345,N_5203,N_6783);
or U9346 (N_9346,N_6352,N_5458);
or U9347 (N_9347,N_5953,N_6913);
or U9348 (N_9348,N_5468,N_7139);
nor U9349 (N_9349,N_7154,N_6253);
and U9350 (N_9350,N_7396,N_6001);
or U9351 (N_9351,N_5012,N_6672);
nand U9352 (N_9352,N_6397,N_6673);
and U9353 (N_9353,N_5372,N_6020);
and U9354 (N_9354,N_5656,N_5205);
and U9355 (N_9355,N_6855,N_5201);
and U9356 (N_9356,N_5493,N_5845);
or U9357 (N_9357,N_5844,N_6154);
nor U9358 (N_9358,N_5832,N_5952);
or U9359 (N_9359,N_5080,N_7333);
nor U9360 (N_9360,N_7087,N_7221);
or U9361 (N_9361,N_5128,N_5850);
nand U9362 (N_9362,N_6201,N_6444);
nand U9363 (N_9363,N_7459,N_5884);
xnor U9364 (N_9364,N_5075,N_5929);
xor U9365 (N_9365,N_5388,N_7112);
and U9366 (N_9366,N_7076,N_7218);
nor U9367 (N_9367,N_5292,N_7335);
xor U9368 (N_9368,N_6445,N_5371);
or U9369 (N_9369,N_5952,N_5892);
nor U9370 (N_9370,N_6583,N_7304);
xor U9371 (N_9371,N_7431,N_6557);
nor U9372 (N_9372,N_6163,N_7452);
and U9373 (N_9373,N_6311,N_6487);
xor U9374 (N_9374,N_6569,N_5020);
and U9375 (N_9375,N_7234,N_5412);
and U9376 (N_9376,N_5765,N_6940);
xnor U9377 (N_9377,N_6926,N_6544);
or U9378 (N_9378,N_6406,N_5731);
xor U9379 (N_9379,N_5207,N_5443);
nand U9380 (N_9380,N_6783,N_5680);
or U9381 (N_9381,N_6047,N_5155);
or U9382 (N_9382,N_7392,N_6102);
or U9383 (N_9383,N_5937,N_5791);
and U9384 (N_9384,N_5596,N_5981);
and U9385 (N_9385,N_7239,N_6287);
and U9386 (N_9386,N_5471,N_7138);
or U9387 (N_9387,N_7161,N_5084);
nand U9388 (N_9388,N_6385,N_5915);
or U9389 (N_9389,N_5957,N_6722);
or U9390 (N_9390,N_5886,N_5583);
nor U9391 (N_9391,N_5177,N_7144);
nor U9392 (N_9392,N_6258,N_5648);
nand U9393 (N_9393,N_5220,N_6977);
nand U9394 (N_9394,N_5030,N_6677);
nor U9395 (N_9395,N_5318,N_5800);
or U9396 (N_9396,N_5550,N_7315);
xnor U9397 (N_9397,N_5617,N_5946);
xor U9398 (N_9398,N_5062,N_6352);
xnor U9399 (N_9399,N_7270,N_5564);
xnor U9400 (N_9400,N_6284,N_6359);
and U9401 (N_9401,N_6377,N_6872);
nor U9402 (N_9402,N_6694,N_7447);
nand U9403 (N_9403,N_6974,N_6062);
and U9404 (N_9404,N_5932,N_7267);
xnor U9405 (N_9405,N_6111,N_6221);
or U9406 (N_9406,N_7393,N_5499);
nand U9407 (N_9407,N_5238,N_5681);
xnor U9408 (N_9408,N_6726,N_5775);
xnor U9409 (N_9409,N_5188,N_6514);
nand U9410 (N_9410,N_6856,N_7486);
nand U9411 (N_9411,N_7146,N_7086);
nor U9412 (N_9412,N_7465,N_7422);
xnor U9413 (N_9413,N_5410,N_6403);
or U9414 (N_9414,N_5326,N_6649);
or U9415 (N_9415,N_6074,N_6992);
and U9416 (N_9416,N_6094,N_7439);
xor U9417 (N_9417,N_5904,N_6943);
nor U9418 (N_9418,N_5733,N_7359);
nor U9419 (N_9419,N_7071,N_6686);
nor U9420 (N_9420,N_6335,N_6400);
xor U9421 (N_9421,N_5075,N_5990);
xor U9422 (N_9422,N_7039,N_5887);
xor U9423 (N_9423,N_5741,N_7168);
nand U9424 (N_9424,N_6055,N_6609);
nand U9425 (N_9425,N_7119,N_5910);
nor U9426 (N_9426,N_5375,N_5608);
and U9427 (N_9427,N_6048,N_6902);
nor U9428 (N_9428,N_5539,N_5994);
and U9429 (N_9429,N_6429,N_5499);
or U9430 (N_9430,N_6023,N_5017);
and U9431 (N_9431,N_5528,N_7351);
and U9432 (N_9432,N_7499,N_6654);
or U9433 (N_9433,N_6914,N_5713);
nor U9434 (N_9434,N_5523,N_7003);
and U9435 (N_9435,N_6030,N_7190);
nor U9436 (N_9436,N_5568,N_6522);
nor U9437 (N_9437,N_5055,N_6863);
or U9438 (N_9438,N_5077,N_6477);
nor U9439 (N_9439,N_5869,N_5767);
or U9440 (N_9440,N_5349,N_6283);
and U9441 (N_9441,N_5299,N_6739);
nand U9442 (N_9442,N_5895,N_5910);
nand U9443 (N_9443,N_5199,N_5632);
or U9444 (N_9444,N_5836,N_6906);
nand U9445 (N_9445,N_6742,N_6221);
xnor U9446 (N_9446,N_6521,N_5200);
nor U9447 (N_9447,N_5006,N_6359);
and U9448 (N_9448,N_7431,N_6771);
or U9449 (N_9449,N_5000,N_5773);
and U9450 (N_9450,N_5176,N_6366);
nor U9451 (N_9451,N_7224,N_5816);
and U9452 (N_9452,N_7303,N_6697);
nand U9453 (N_9453,N_6978,N_7414);
and U9454 (N_9454,N_6935,N_7489);
nor U9455 (N_9455,N_5508,N_5452);
nor U9456 (N_9456,N_6374,N_5216);
xor U9457 (N_9457,N_5530,N_7161);
nor U9458 (N_9458,N_7343,N_6584);
nor U9459 (N_9459,N_7193,N_6891);
nand U9460 (N_9460,N_5217,N_6967);
nand U9461 (N_9461,N_5186,N_7353);
xnor U9462 (N_9462,N_7130,N_5028);
and U9463 (N_9463,N_6600,N_6828);
xnor U9464 (N_9464,N_5987,N_6457);
nor U9465 (N_9465,N_5216,N_7054);
or U9466 (N_9466,N_7314,N_6995);
and U9467 (N_9467,N_6463,N_5547);
and U9468 (N_9468,N_6359,N_6086);
nor U9469 (N_9469,N_6214,N_6277);
or U9470 (N_9470,N_7120,N_5290);
or U9471 (N_9471,N_5938,N_6828);
nor U9472 (N_9472,N_5805,N_5547);
nand U9473 (N_9473,N_5274,N_7393);
xnor U9474 (N_9474,N_5485,N_5650);
nor U9475 (N_9475,N_6619,N_7215);
nand U9476 (N_9476,N_6994,N_7434);
nor U9477 (N_9477,N_6952,N_5337);
xor U9478 (N_9478,N_5026,N_6699);
nor U9479 (N_9479,N_6243,N_6027);
xnor U9480 (N_9480,N_7410,N_7102);
nand U9481 (N_9481,N_7317,N_5114);
and U9482 (N_9482,N_7174,N_6184);
nor U9483 (N_9483,N_6228,N_5582);
or U9484 (N_9484,N_6429,N_5266);
and U9485 (N_9485,N_5610,N_6057);
xor U9486 (N_9486,N_7412,N_5555);
xnor U9487 (N_9487,N_5970,N_6404);
or U9488 (N_9488,N_7192,N_6352);
nor U9489 (N_9489,N_6703,N_6213);
xor U9490 (N_9490,N_6784,N_6807);
nand U9491 (N_9491,N_7047,N_6732);
xor U9492 (N_9492,N_7039,N_6473);
nand U9493 (N_9493,N_6380,N_5950);
and U9494 (N_9494,N_5787,N_6094);
xnor U9495 (N_9495,N_6599,N_7102);
or U9496 (N_9496,N_6952,N_5449);
nand U9497 (N_9497,N_6054,N_7101);
or U9498 (N_9498,N_7084,N_5055);
or U9499 (N_9499,N_7291,N_7104);
or U9500 (N_9500,N_6693,N_5909);
xnor U9501 (N_9501,N_6940,N_7085);
xnor U9502 (N_9502,N_5007,N_5599);
nand U9503 (N_9503,N_5990,N_6380);
xnor U9504 (N_9504,N_5008,N_7183);
nor U9505 (N_9505,N_5157,N_6120);
xor U9506 (N_9506,N_6150,N_5942);
nand U9507 (N_9507,N_7289,N_5839);
or U9508 (N_9508,N_5809,N_6313);
nand U9509 (N_9509,N_6150,N_7193);
or U9510 (N_9510,N_6609,N_6725);
xor U9511 (N_9511,N_6881,N_7109);
or U9512 (N_9512,N_6822,N_6154);
xor U9513 (N_9513,N_7166,N_7002);
nor U9514 (N_9514,N_5721,N_6756);
or U9515 (N_9515,N_6613,N_6931);
or U9516 (N_9516,N_6275,N_5319);
nor U9517 (N_9517,N_6345,N_6219);
nor U9518 (N_9518,N_6124,N_5633);
and U9519 (N_9519,N_6418,N_5547);
nand U9520 (N_9520,N_5600,N_7257);
xnor U9521 (N_9521,N_7016,N_5510);
nor U9522 (N_9522,N_7431,N_5018);
nor U9523 (N_9523,N_6371,N_6657);
or U9524 (N_9524,N_7437,N_6541);
or U9525 (N_9525,N_5244,N_7479);
nand U9526 (N_9526,N_6631,N_6366);
xnor U9527 (N_9527,N_6054,N_6004);
and U9528 (N_9528,N_7078,N_6374);
nand U9529 (N_9529,N_7443,N_5631);
nand U9530 (N_9530,N_5542,N_6700);
nor U9531 (N_9531,N_5202,N_6145);
nor U9532 (N_9532,N_6325,N_6209);
xor U9533 (N_9533,N_5025,N_5440);
xor U9534 (N_9534,N_6700,N_5925);
nor U9535 (N_9535,N_6994,N_5032);
nand U9536 (N_9536,N_6069,N_7274);
and U9537 (N_9537,N_6832,N_6720);
xor U9538 (N_9538,N_6680,N_5499);
xnor U9539 (N_9539,N_7166,N_6796);
and U9540 (N_9540,N_6512,N_7385);
nand U9541 (N_9541,N_5839,N_5978);
and U9542 (N_9542,N_7174,N_6501);
nor U9543 (N_9543,N_6908,N_7473);
and U9544 (N_9544,N_6916,N_6056);
and U9545 (N_9545,N_6314,N_6644);
nand U9546 (N_9546,N_5302,N_5403);
nor U9547 (N_9547,N_6809,N_5878);
and U9548 (N_9548,N_6746,N_5407);
and U9549 (N_9549,N_6426,N_7120);
nand U9550 (N_9550,N_5647,N_5359);
nand U9551 (N_9551,N_6508,N_7305);
nor U9552 (N_9552,N_6985,N_6153);
and U9553 (N_9553,N_5895,N_5869);
xor U9554 (N_9554,N_6415,N_6867);
nand U9555 (N_9555,N_5614,N_7285);
xnor U9556 (N_9556,N_6046,N_6117);
or U9557 (N_9557,N_7075,N_7045);
or U9558 (N_9558,N_7167,N_6319);
and U9559 (N_9559,N_5718,N_5775);
nand U9560 (N_9560,N_5568,N_5073);
xnor U9561 (N_9561,N_7370,N_5861);
nor U9562 (N_9562,N_5044,N_5846);
xnor U9563 (N_9563,N_5572,N_5485);
xnor U9564 (N_9564,N_7459,N_5410);
and U9565 (N_9565,N_5088,N_5521);
or U9566 (N_9566,N_5762,N_6297);
or U9567 (N_9567,N_6509,N_6233);
xnor U9568 (N_9568,N_6405,N_5402);
and U9569 (N_9569,N_6377,N_6839);
or U9570 (N_9570,N_6782,N_6475);
nand U9571 (N_9571,N_6921,N_5401);
or U9572 (N_9572,N_6010,N_6431);
nand U9573 (N_9573,N_6548,N_6855);
nor U9574 (N_9574,N_6554,N_5283);
nand U9575 (N_9575,N_6511,N_5055);
nor U9576 (N_9576,N_5438,N_6061);
xnor U9577 (N_9577,N_6769,N_6531);
nor U9578 (N_9578,N_5824,N_6855);
and U9579 (N_9579,N_5802,N_5495);
and U9580 (N_9580,N_7469,N_7032);
nand U9581 (N_9581,N_6169,N_6974);
nand U9582 (N_9582,N_5689,N_5366);
nor U9583 (N_9583,N_5760,N_5365);
nor U9584 (N_9584,N_5191,N_6117);
or U9585 (N_9585,N_7064,N_6340);
xor U9586 (N_9586,N_5657,N_6148);
nand U9587 (N_9587,N_6397,N_7439);
and U9588 (N_9588,N_5882,N_6980);
or U9589 (N_9589,N_6663,N_7355);
or U9590 (N_9590,N_7384,N_5194);
or U9591 (N_9591,N_5638,N_5328);
xnor U9592 (N_9592,N_7035,N_5307);
nand U9593 (N_9593,N_6744,N_7247);
or U9594 (N_9594,N_5971,N_5684);
nor U9595 (N_9595,N_5721,N_6479);
and U9596 (N_9596,N_5825,N_6770);
or U9597 (N_9597,N_6630,N_6783);
xor U9598 (N_9598,N_5872,N_6990);
nor U9599 (N_9599,N_6683,N_6179);
and U9600 (N_9600,N_6143,N_6472);
xnor U9601 (N_9601,N_7434,N_5645);
or U9602 (N_9602,N_7218,N_6890);
nor U9603 (N_9603,N_5051,N_5226);
nand U9604 (N_9604,N_7061,N_7417);
xnor U9605 (N_9605,N_5561,N_5082);
or U9606 (N_9606,N_6239,N_7126);
xnor U9607 (N_9607,N_6118,N_5488);
nand U9608 (N_9608,N_5219,N_6605);
xor U9609 (N_9609,N_6383,N_5842);
xnor U9610 (N_9610,N_5382,N_7068);
nor U9611 (N_9611,N_5812,N_6857);
or U9612 (N_9612,N_5144,N_5845);
nand U9613 (N_9613,N_5847,N_7077);
or U9614 (N_9614,N_5891,N_5188);
xor U9615 (N_9615,N_5944,N_6552);
xnor U9616 (N_9616,N_5379,N_7341);
and U9617 (N_9617,N_6463,N_6254);
or U9618 (N_9618,N_5377,N_5170);
nor U9619 (N_9619,N_5870,N_5767);
or U9620 (N_9620,N_6103,N_5841);
nand U9621 (N_9621,N_5754,N_5212);
xor U9622 (N_9622,N_6966,N_6543);
nand U9623 (N_9623,N_6894,N_5540);
or U9624 (N_9624,N_7304,N_6017);
xor U9625 (N_9625,N_6254,N_5996);
nand U9626 (N_9626,N_6890,N_6208);
or U9627 (N_9627,N_5725,N_6943);
or U9628 (N_9628,N_7026,N_5172);
nand U9629 (N_9629,N_7333,N_5494);
and U9630 (N_9630,N_7361,N_5676);
xnor U9631 (N_9631,N_5871,N_5492);
nand U9632 (N_9632,N_5899,N_6730);
or U9633 (N_9633,N_5763,N_6005);
nand U9634 (N_9634,N_5507,N_6046);
and U9635 (N_9635,N_6116,N_5909);
xor U9636 (N_9636,N_6333,N_7495);
nor U9637 (N_9637,N_7375,N_7177);
or U9638 (N_9638,N_6220,N_6389);
nand U9639 (N_9639,N_7493,N_5685);
nor U9640 (N_9640,N_6415,N_6732);
and U9641 (N_9641,N_6283,N_5795);
nand U9642 (N_9642,N_7405,N_6143);
nand U9643 (N_9643,N_6226,N_5490);
xor U9644 (N_9644,N_6006,N_5832);
nor U9645 (N_9645,N_7424,N_5830);
and U9646 (N_9646,N_6201,N_7235);
nor U9647 (N_9647,N_5377,N_7084);
xor U9648 (N_9648,N_6110,N_7075);
xor U9649 (N_9649,N_5811,N_6451);
nand U9650 (N_9650,N_5814,N_6052);
xnor U9651 (N_9651,N_6525,N_7442);
or U9652 (N_9652,N_7071,N_7022);
nor U9653 (N_9653,N_6030,N_6674);
or U9654 (N_9654,N_7391,N_6306);
nor U9655 (N_9655,N_6907,N_5553);
nor U9656 (N_9656,N_5406,N_5239);
or U9657 (N_9657,N_5147,N_7130);
or U9658 (N_9658,N_6327,N_7344);
or U9659 (N_9659,N_5543,N_7219);
or U9660 (N_9660,N_5621,N_6333);
xor U9661 (N_9661,N_5735,N_6332);
xnor U9662 (N_9662,N_7302,N_7208);
nand U9663 (N_9663,N_6326,N_5789);
and U9664 (N_9664,N_5848,N_5883);
xnor U9665 (N_9665,N_6590,N_7313);
nor U9666 (N_9666,N_7209,N_5622);
nand U9667 (N_9667,N_5848,N_7387);
and U9668 (N_9668,N_5023,N_5450);
nand U9669 (N_9669,N_6179,N_7086);
or U9670 (N_9670,N_5879,N_6059);
xor U9671 (N_9671,N_6897,N_6272);
and U9672 (N_9672,N_5452,N_6425);
nor U9673 (N_9673,N_5507,N_6890);
nor U9674 (N_9674,N_6982,N_7471);
and U9675 (N_9675,N_7153,N_7465);
or U9676 (N_9676,N_6855,N_6767);
and U9677 (N_9677,N_5548,N_6150);
xor U9678 (N_9678,N_5872,N_6709);
xor U9679 (N_9679,N_5320,N_5611);
nor U9680 (N_9680,N_5701,N_7125);
nor U9681 (N_9681,N_6910,N_6211);
or U9682 (N_9682,N_6176,N_5968);
and U9683 (N_9683,N_5255,N_5883);
and U9684 (N_9684,N_6786,N_5577);
and U9685 (N_9685,N_5739,N_6545);
and U9686 (N_9686,N_7212,N_6041);
nor U9687 (N_9687,N_6368,N_6344);
and U9688 (N_9688,N_5570,N_7010);
nand U9689 (N_9689,N_5891,N_7442);
and U9690 (N_9690,N_5771,N_6609);
and U9691 (N_9691,N_5196,N_5744);
nor U9692 (N_9692,N_5466,N_6192);
nor U9693 (N_9693,N_6213,N_6910);
or U9694 (N_9694,N_6360,N_6908);
and U9695 (N_9695,N_5086,N_5278);
nand U9696 (N_9696,N_6302,N_6597);
and U9697 (N_9697,N_7283,N_5376);
or U9698 (N_9698,N_6089,N_5411);
nand U9699 (N_9699,N_5406,N_6983);
nand U9700 (N_9700,N_6031,N_6941);
nor U9701 (N_9701,N_5223,N_5693);
or U9702 (N_9702,N_5251,N_7139);
and U9703 (N_9703,N_5088,N_6803);
nor U9704 (N_9704,N_5275,N_5296);
or U9705 (N_9705,N_6973,N_5188);
and U9706 (N_9706,N_5032,N_5243);
and U9707 (N_9707,N_7129,N_6811);
xor U9708 (N_9708,N_6270,N_6950);
and U9709 (N_9709,N_5529,N_7381);
or U9710 (N_9710,N_6816,N_6659);
nor U9711 (N_9711,N_6388,N_6755);
nor U9712 (N_9712,N_7364,N_5205);
and U9713 (N_9713,N_5992,N_7075);
nor U9714 (N_9714,N_6644,N_6366);
nand U9715 (N_9715,N_5607,N_5488);
nor U9716 (N_9716,N_6482,N_7166);
or U9717 (N_9717,N_6290,N_7282);
nor U9718 (N_9718,N_7007,N_7000);
nor U9719 (N_9719,N_7127,N_6074);
xor U9720 (N_9720,N_5844,N_5965);
and U9721 (N_9721,N_5006,N_6121);
nand U9722 (N_9722,N_6167,N_7267);
nor U9723 (N_9723,N_5021,N_7358);
nand U9724 (N_9724,N_6050,N_6470);
xor U9725 (N_9725,N_6465,N_5527);
nand U9726 (N_9726,N_5936,N_5870);
nand U9727 (N_9727,N_6501,N_5839);
xnor U9728 (N_9728,N_5001,N_6228);
nand U9729 (N_9729,N_6942,N_7053);
or U9730 (N_9730,N_6490,N_6895);
nor U9731 (N_9731,N_5642,N_5339);
xnor U9732 (N_9732,N_5771,N_5328);
and U9733 (N_9733,N_5743,N_7040);
and U9734 (N_9734,N_7039,N_5843);
nand U9735 (N_9735,N_7334,N_7066);
xor U9736 (N_9736,N_6628,N_7247);
and U9737 (N_9737,N_6207,N_6462);
nand U9738 (N_9738,N_5742,N_5982);
nor U9739 (N_9739,N_7494,N_7422);
and U9740 (N_9740,N_5387,N_5212);
or U9741 (N_9741,N_5707,N_5423);
nor U9742 (N_9742,N_6341,N_5219);
nand U9743 (N_9743,N_5443,N_7187);
or U9744 (N_9744,N_6181,N_6557);
and U9745 (N_9745,N_7110,N_5386);
xor U9746 (N_9746,N_6074,N_6295);
nor U9747 (N_9747,N_5815,N_6802);
and U9748 (N_9748,N_6986,N_5890);
nor U9749 (N_9749,N_6589,N_5272);
nand U9750 (N_9750,N_5113,N_7305);
nor U9751 (N_9751,N_5072,N_5748);
xnor U9752 (N_9752,N_7265,N_5849);
nor U9753 (N_9753,N_5385,N_5140);
and U9754 (N_9754,N_7075,N_6524);
and U9755 (N_9755,N_5333,N_5920);
and U9756 (N_9756,N_6249,N_7237);
nor U9757 (N_9757,N_5553,N_5996);
or U9758 (N_9758,N_6753,N_6601);
xor U9759 (N_9759,N_7037,N_6210);
or U9760 (N_9760,N_6138,N_6720);
or U9761 (N_9761,N_5525,N_6942);
nor U9762 (N_9762,N_5389,N_5072);
nor U9763 (N_9763,N_6730,N_5760);
xor U9764 (N_9764,N_6806,N_7420);
nand U9765 (N_9765,N_5435,N_7421);
nand U9766 (N_9766,N_6184,N_5394);
nand U9767 (N_9767,N_5416,N_7320);
xor U9768 (N_9768,N_6270,N_7357);
nor U9769 (N_9769,N_6367,N_5009);
and U9770 (N_9770,N_5609,N_6119);
and U9771 (N_9771,N_7379,N_5859);
xnor U9772 (N_9772,N_6807,N_5094);
or U9773 (N_9773,N_5669,N_6445);
nor U9774 (N_9774,N_6058,N_7209);
xnor U9775 (N_9775,N_5725,N_5888);
and U9776 (N_9776,N_6767,N_5045);
xnor U9777 (N_9777,N_5197,N_5598);
nor U9778 (N_9778,N_6296,N_7383);
nor U9779 (N_9779,N_7022,N_7375);
nand U9780 (N_9780,N_6159,N_7093);
or U9781 (N_9781,N_6415,N_7434);
nor U9782 (N_9782,N_5545,N_6853);
nand U9783 (N_9783,N_5529,N_5081);
and U9784 (N_9784,N_5091,N_6766);
nor U9785 (N_9785,N_7118,N_6558);
xnor U9786 (N_9786,N_6536,N_5937);
xnor U9787 (N_9787,N_6248,N_6087);
xnor U9788 (N_9788,N_6694,N_7369);
xnor U9789 (N_9789,N_6059,N_5185);
and U9790 (N_9790,N_5205,N_7491);
xor U9791 (N_9791,N_5385,N_5079);
or U9792 (N_9792,N_7087,N_5015);
xor U9793 (N_9793,N_7289,N_6106);
nor U9794 (N_9794,N_5370,N_5277);
nand U9795 (N_9795,N_5425,N_6277);
or U9796 (N_9796,N_7190,N_5988);
nor U9797 (N_9797,N_5470,N_7125);
and U9798 (N_9798,N_5493,N_6108);
nor U9799 (N_9799,N_5552,N_5466);
nand U9800 (N_9800,N_6574,N_6907);
and U9801 (N_9801,N_5014,N_6395);
xnor U9802 (N_9802,N_7380,N_6746);
nor U9803 (N_9803,N_5481,N_6411);
nand U9804 (N_9804,N_5963,N_5916);
and U9805 (N_9805,N_5043,N_6380);
nor U9806 (N_9806,N_5329,N_6623);
and U9807 (N_9807,N_6053,N_5038);
nand U9808 (N_9808,N_6724,N_7203);
or U9809 (N_9809,N_5765,N_5576);
xor U9810 (N_9810,N_5075,N_5876);
xnor U9811 (N_9811,N_5048,N_5556);
and U9812 (N_9812,N_6647,N_7265);
and U9813 (N_9813,N_6902,N_6685);
and U9814 (N_9814,N_5072,N_5959);
nand U9815 (N_9815,N_7484,N_5607);
or U9816 (N_9816,N_6472,N_5552);
or U9817 (N_9817,N_5751,N_5392);
nor U9818 (N_9818,N_7281,N_6703);
nand U9819 (N_9819,N_5106,N_7006);
nor U9820 (N_9820,N_5273,N_6024);
nor U9821 (N_9821,N_5982,N_5899);
nand U9822 (N_9822,N_7306,N_6760);
nor U9823 (N_9823,N_6006,N_6118);
and U9824 (N_9824,N_5368,N_5078);
nand U9825 (N_9825,N_7060,N_5306);
and U9826 (N_9826,N_6292,N_5437);
nor U9827 (N_9827,N_5105,N_5044);
and U9828 (N_9828,N_5556,N_7269);
nand U9829 (N_9829,N_6455,N_5777);
xor U9830 (N_9830,N_7028,N_5413);
or U9831 (N_9831,N_6585,N_7135);
or U9832 (N_9832,N_5824,N_6696);
xnor U9833 (N_9833,N_7095,N_6243);
xor U9834 (N_9834,N_6928,N_5110);
nand U9835 (N_9835,N_5348,N_6925);
or U9836 (N_9836,N_5340,N_5558);
or U9837 (N_9837,N_7365,N_5782);
nor U9838 (N_9838,N_7421,N_7400);
nor U9839 (N_9839,N_6502,N_5957);
nand U9840 (N_9840,N_5359,N_7474);
nor U9841 (N_9841,N_7114,N_7390);
and U9842 (N_9842,N_7001,N_5629);
nor U9843 (N_9843,N_7365,N_6592);
and U9844 (N_9844,N_5182,N_6129);
xor U9845 (N_9845,N_6827,N_6809);
xor U9846 (N_9846,N_6772,N_6607);
nand U9847 (N_9847,N_7333,N_5517);
xnor U9848 (N_9848,N_7440,N_7332);
or U9849 (N_9849,N_5376,N_6392);
and U9850 (N_9850,N_7324,N_7070);
xor U9851 (N_9851,N_5855,N_6620);
nor U9852 (N_9852,N_6411,N_6587);
xor U9853 (N_9853,N_5825,N_5852);
nor U9854 (N_9854,N_6383,N_7016);
or U9855 (N_9855,N_7437,N_5737);
xnor U9856 (N_9856,N_7277,N_5063);
nand U9857 (N_9857,N_5673,N_5350);
nor U9858 (N_9858,N_5428,N_6326);
nor U9859 (N_9859,N_7043,N_6532);
and U9860 (N_9860,N_6417,N_5198);
and U9861 (N_9861,N_7232,N_7183);
or U9862 (N_9862,N_6660,N_5998);
and U9863 (N_9863,N_7379,N_5789);
and U9864 (N_9864,N_7206,N_6656);
xor U9865 (N_9865,N_5231,N_5290);
xnor U9866 (N_9866,N_5266,N_5104);
or U9867 (N_9867,N_7259,N_6857);
xnor U9868 (N_9868,N_6954,N_5596);
nand U9869 (N_9869,N_5897,N_7039);
and U9870 (N_9870,N_5469,N_7329);
nand U9871 (N_9871,N_5287,N_5731);
and U9872 (N_9872,N_6773,N_5764);
xnor U9873 (N_9873,N_5031,N_5706);
nand U9874 (N_9874,N_5080,N_5970);
and U9875 (N_9875,N_5872,N_6437);
and U9876 (N_9876,N_5320,N_5983);
xor U9877 (N_9877,N_5339,N_6465);
nor U9878 (N_9878,N_5160,N_5395);
and U9879 (N_9879,N_7003,N_5943);
or U9880 (N_9880,N_6784,N_5560);
or U9881 (N_9881,N_6633,N_5934);
xnor U9882 (N_9882,N_5977,N_7392);
xor U9883 (N_9883,N_6113,N_5656);
and U9884 (N_9884,N_6141,N_7392);
nor U9885 (N_9885,N_5128,N_6864);
or U9886 (N_9886,N_6709,N_5660);
or U9887 (N_9887,N_7275,N_7101);
nor U9888 (N_9888,N_7085,N_7283);
and U9889 (N_9889,N_6051,N_5356);
or U9890 (N_9890,N_6998,N_7368);
and U9891 (N_9891,N_5179,N_6153);
xnor U9892 (N_9892,N_7150,N_7224);
nor U9893 (N_9893,N_6421,N_6559);
xor U9894 (N_9894,N_5997,N_6367);
nor U9895 (N_9895,N_6377,N_6860);
nor U9896 (N_9896,N_5522,N_5998);
nand U9897 (N_9897,N_5095,N_7424);
nor U9898 (N_9898,N_7175,N_5663);
and U9899 (N_9899,N_6856,N_5463);
xor U9900 (N_9900,N_6559,N_7355);
nor U9901 (N_9901,N_7392,N_6634);
nand U9902 (N_9902,N_7165,N_6046);
nand U9903 (N_9903,N_5881,N_5170);
or U9904 (N_9904,N_7347,N_6264);
nand U9905 (N_9905,N_6434,N_6911);
nor U9906 (N_9906,N_6858,N_5517);
and U9907 (N_9907,N_6461,N_5667);
and U9908 (N_9908,N_5851,N_7057);
or U9909 (N_9909,N_7306,N_7066);
or U9910 (N_9910,N_7232,N_7053);
nand U9911 (N_9911,N_6423,N_6314);
and U9912 (N_9912,N_6086,N_5228);
nor U9913 (N_9913,N_6046,N_5808);
xnor U9914 (N_9914,N_5173,N_6118);
xnor U9915 (N_9915,N_5709,N_5213);
or U9916 (N_9916,N_7227,N_7368);
and U9917 (N_9917,N_5487,N_6369);
nor U9918 (N_9918,N_7465,N_6170);
or U9919 (N_9919,N_5309,N_5874);
and U9920 (N_9920,N_7405,N_5421);
nand U9921 (N_9921,N_6106,N_5438);
nor U9922 (N_9922,N_6227,N_5728);
nor U9923 (N_9923,N_5038,N_7085);
and U9924 (N_9924,N_6101,N_7413);
nor U9925 (N_9925,N_5807,N_5206);
nor U9926 (N_9926,N_7306,N_6914);
nand U9927 (N_9927,N_6707,N_6602);
or U9928 (N_9928,N_6033,N_6577);
nand U9929 (N_9929,N_5176,N_5192);
or U9930 (N_9930,N_5312,N_6413);
or U9931 (N_9931,N_7415,N_5462);
or U9932 (N_9932,N_5835,N_5376);
nand U9933 (N_9933,N_7152,N_5736);
and U9934 (N_9934,N_6887,N_7034);
or U9935 (N_9935,N_6866,N_6895);
nor U9936 (N_9936,N_7257,N_6532);
and U9937 (N_9937,N_5335,N_7008);
and U9938 (N_9938,N_6300,N_6141);
or U9939 (N_9939,N_6521,N_7104);
and U9940 (N_9940,N_5457,N_7264);
or U9941 (N_9941,N_5479,N_6897);
or U9942 (N_9942,N_6304,N_6184);
xnor U9943 (N_9943,N_5179,N_5858);
and U9944 (N_9944,N_6677,N_5423);
nor U9945 (N_9945,N_6593,N_5213);
and U9946 (N_9946,N_5567,N_5159);
nor U9947 (N_9947,N_7280,N_6002);
xnor U9948 (N_9948,N_5634,N_5747);
nand U9949 (N_9949,N_5412,N_6185);
nor U9950 (N_9950,N_6046,N_7048);
xor U9951 (N_9951,N_5442,N_5554);
or U9952 (N_9952,N_5053,N_7156);
and U9953 (N_9953,N_5751,N_7155);
nand U9954 (N_9954,N_6207,N_6682);
nor U9955 (N_9955,N_7459,N_6413);
xnor U9956 (N_9956,N_5360,N_5801);
nor U9957 (N_9957,N_6769,N_5829);
nor U9958 (N_9958,N_5553,N_7014);
nand U9959 (N_9959,N_5100,N_7089);
or U9960 (N_9960,N_6436,N_7245);
nand U9961 (N_9961,N_6733,N_6322);
nor U9962 (N_9962,N_5202,N_6251);
nor U9963 (N_9963,N_6458,N_6228);
xor U9964 (N_9964,N_6357,N_5900);
and U9965 (N_9965,N_6252,N_5105);
nor U9966 (N_9966,N_6099,N_6293);
or U9967 (N_9967,N_6285,N_6237);
or U9968 (N_9968,N_6375,N_7394);
nor U9969 (N_9969,N_6525,N_5667);
or U9970 (N_9970,N_7062,N_7156);
and U9971 (N_9971,N_6483,N_7359);
and U9972 (N_9972,N_5581,N_5075);
or U9973 (N_9973,N_6558,N_7012);
or U9974 (N_9974,N_6377,N_6402);
or U9975 (N_9975,N_6735,N_7479);
or U9976 (N_9976,N_5532,N_6045);
nand U9977 (N_9977,N_7499,N_5639);
or U9978 (N_9978,N_6624,N_5266);
and U9979 (N_9979,N_7495,N_6544);
nand U9980 (N_9980,N_6448,N_5258);
or U9981 (N_9981,N_5032,N_6080);
xor U9982 (N_9982,N_6617,N_7355);
nand U9983 (N_9983,N_6894,N_5377);
and U9984 (N_9984,N_6651,N_6598);
and U9985 (N_9985,N_7428,N_6357);
nand U9986 (N_9986,N_6221,N_5472);
and U9987 (N_9987,N_6685,N_5472);
or U9988 (N_9988,N_6802,N_5359);
nor U9989 (N_9989,N_6286,N_6790);
or U9990 (N_9990,N_5150,N_7014);
nor U9991 (N_9991,N_6087,N_7298);
nor U9992 (N_9992,N_5009,N_5105);
nor U9993 (N_9993,N_6677,N_6777);
nor U9994 (N_9994,N_5334,N_5860);
nor U9995 (N_9995,N_5332,N_6224);
and U9996 (N_9996,N_5666,N_6854);
xor U9997 (N_9997,N_6508,N_6298);
nor U9998 (N_9998,N_5662,N_6214);
or U9999 (N_9999,N_6263,N_6256);
nor U10000 (N_10000,N_8471,N_9805);
or U10001 (N_10001,N_8986,N_8666);
nor U10002 (N_10002,N_8037,N_9249);
and U10003 (N_10003,N_8810,N_8224);
nor U10004 (N_10004,N_9827,N_9722);
xor U10005 (N_10005,N_9442,N_8347);
or U10006 (N_10006,N_8166,N_9558);
xnor U10007 (N_10007,N_9374,N_9617);
or U10008 (N_10008,N_8739,N_8923);
xnor U10009 (N_10009,N_8256,N_9107);
and U10010 (N_10010,N_9269,N_9109);
nor U10011 (N_10011,N_9653,N_9673);
nor U10012 (N_10012,N_8747,N_7966);
or U10013 (N_10013,N_9809,N_8641);
xor U10014 (N_10014,N_9942,N_7613);
nor U10015 (N_10015,N_7668,N_8989);
and U10016 (N_10016,N_7573,N_9169);
nand U10017 (N_10017,N_8764,N_8834);
nand U10018 (N_10018,N_7770,N_8964);
nand U10019 (N_10019,N_7689,N_8795);
or U10020 (N_10020,N_7672,N_8302);
or U10021 (N_10021,N_9990,N_9583);
or U10022 (N_10022,N_8853,N_8353);
and U10023 (N_10023,N_9529,N_7790);
nor U10024 (N_10024,N_8000,N_9449);
and U10025 (N_10025,N_8540,N_9039);
and U10026 (N_10026,N_9407,N_8813);
nor U10027 (N_10027,N_8112,N_8275);
and U10028 (N_10028,N_7891,N_8741);
nand U10029 (N_10029,N_7878,N_8549);
and U10030 (N_10030,N_8143,N_9776);
and U10031 (N_10031,N_7918,N_9871);
nand U10032 (N_10032,N_9175,N_8245);
nand U10033 (N_10033,N_7522,N_9058);
nand U10034 (N_10034,N_8953,N_8064);
and U10035 (N_10035,N_8421,N_9493);
nand U10036 (N_10036,N_7859,N_7812);
or U10037 (N_10037,N_8100,N_8161);
nor U10038 (N_10038,N_9873,N_8823);
and U10039 (N_10039,N_8790,N_8287);
xor U10040 (N_10040,N_8393,N_9959);
nor U10041 (N_10041,N_8910,N_9286);
xor U10042 (N_10042,N_8822,N_8878);
nor U10043 (N_10043,N_8581,N_9657);
xor U10044 (N_10044,N_8090,N_9489);
nor U10045 (N_10045,N_8400,N_7657);
xor U10046 (N_10046,N_9250,N_9160);
xor U10047 (N_10047,N_8525,N_9447);
nor U10048 (N_10048,N_9495,N_7775);
and U10049 (N_10049,N_8313,N_8365);
nand U10050 (N_10050,N_9606,N_9114);
or U10051 (N_10051,N_8983,N_8176);
nand U10052 (N_10052,N_9779,N_9123);
and U10053 (N_10053,N_9046,N_7777);
nand U10054 (N_10054,N_7888,N_8005);
xnor U10055 (N_10055,N_8455,N_9317);
and U10056 (N_10056,N_9865,N_7528);
or U10057 (N_10057,N_9567,N_7693);
and U10058 (N_10058,N_8887,N_9263);
nor U10059 (N_10059,N_9518,N_8402);
nor U10060 (N_10060,N_9751,N_9487);
nor U10061 (N_10061,N_8031,N_7665);
or U10062 (N_10062,N_9773,N_9678);
and U10063 (N_10063,N_8268,N_8093);
nor U10064 (N_10064,N_8837,N_9026);
nand U10065 (N_10065,N_7509,N_8065);
nor U10066 (N_10066,N_7887,N_8059);
nor U10067 (N_10067,N_9542,N_8618);
xnor U10068 (N_10068,N_8619,N_7929);
xnor U10069 (N_10069,N_7728,N_9488);
xnor U10070 (N_10070,N_9130,N_9102);
or U10071 (N_10071,N_7815,N_8382);
xor U10072 (N_10072,N_9986,N_7588);
or U10073 (N_10073,N_7861,N_9354);
nor U10074 (N_10074,N_9611,N_9648);
or U10075 (N_10075,N_7541,N_7510);
or U10076 (N_10076,N_9584,N_9173);
xor U10077 (N_10077,N_7963,N_9635);
nor U10078 (N_10078,N_8477,N_9017);
nor U10079 (N_10079,N_9920,N_9804);
or U10080 (N_10080,N_8684,N_9812);
nand U10081 (N_10081,N_9117,N_9034);
and U10082 (N_10082,N_7726,N_7952);
xnor U10083 (N_10083,N_7897,N_9690);
xor U10084 (N_10084,N_8572,N_7596);
nand U10085 (N_10085,N_7618,N_8013);
or U10086 (N_10086,N_8979,N_8791);
nand U10087 (N_10087,N_7710,N_9701);
nor U10088 (N_10088,N_8009,N_9721);
nor U10089 (N_10089,N_9861,N_9378);
or U10090 (N_10090,N_8939,N_9900);
or U10091 (N_10091,N_9131,N_8945);
xnor U10092 (N_10092,N_9180,N_7727);
or U10093 (N_10093,N_8295,N_7637);
nand U10094 (N_10094,N_7896,N_8766);
nand U10095 (N_10095,N_8575,N_8431);
or U10096 (N_10096,N_9353,N_9057);
and U10097 (N_10097,N_8179,N_8902);
nor U10098 (N_10098,N_8976,N_8818);
nand U10099 (N_10099,N_9260,N_8794);
nand U10100 (N_10100,N_7526,N_7636);
xnor U10101 (N_10101,N_8772,N_7702);
nor U10102 (N_10102,N_8218,N_9790);
nand U10103 (N_10103,N_9326,N_7956);
nand U10104 (N_10104,N_7539,N_8323);
or U10105 (N_10105,N_9282,N_8025);
xnor U10106 (N_10106,N_9283,N_9170);
nor U10107 (N_10107,N_7764,N_9957);
nand U10108 (N_10108,N_8120,N_8631);
xor U10109 (N_10109,N_8066,N_9868);
nand U10110 (N_10110,N_8929,N_8523);
nor U10111 (N_10111,N_9824,N_9348);
xor U10112 (N_10112,N_9535,N_8962);
and U10113 (N_10113,N_8160,N_9491);
or U10114 (N_10114,N_8630,N_9032);
xor U10115 (N_10115,N_8776,N_8909);
nand U10116 (N_10116,N_7698,N_8901);
nand U10117 (N_10117,N_9415,N_9705);
nand U10118 (N_10118,N_9176,N_7638);
nor U10119 (N_10119,N_8088,N_9884);
and U10120 (N_10120,N_9695,N_8940);
and U10121 (N_10121,N_8960,N_9025);
xor U10122 (N_10122,N_9023,N_7611);
nand U10123 (N_10123,N_9465,N_8977);
xnor U10124 (N_10124,N_7543,N_8310);
and U10125 (N_10125,N_8105,N_8634);
nand U10126 (N_10126,N_9745,N_8532);
and U10127 (N_10127,N_9016,N_8286);
nor U10128 (N_10128,N_8384,N_9171);
and U10129 (N_10129,N_7898,N_8513);
nor U10130 (N_10130,N_7562,N_9055);
nor U10131 (N_10131,N_8686,N_8459);
and U10132 (N_10132,N_9662,N_8846);
or U10133 (N_10133,N_8872,N_9620);
xnor U10134 (N_10134,N_9943,N_9853);
xnor U10135 (N_10135,N_9687,N_7792);
xor U10136 (N_10136,N_7754,N_8707);
nor U10137 (N_10137,N_9640,N_9060);
nand U10138 (N_10138,N_9400,N_9811);
and U10139 (N_10139,N_7523,N_7752);
and U10140 (N_10140,N_7818,N_7984);
nand U10141 (N_10141,N_9852,N_8080);
nand U10142 (N_10142,N_9191,N_9343);
xor U10143 (N_10143,N_7604,N_8348);
xor U10144 (N_10144,N_7530,N_9710);
and U10145 (N_10145,N_7940,N_7660);
nor U10146 (N_10146,N_8524,N_8679);
nand U10147 (N_10147,N_7756,N_7524);
and U10148 (N_10148,N_9295,N_7848);
or U10149 (N_10149,N_8079,N_7701);
and U10150 (N_10150,N_7648,N_9364);
nand U10151 (N_10151,N_8915,N_8985);
and U10152 (N_10152,N_9737,N_9480);
or U10153 (N_10153,N_9674,N_9887);
xor U10154 (N_10154,N_7595,N_9818);
xnor U10155 (N_10155,N_8495,N_9053);
or U10156 (N_10156,N_9228,N_8174);
or U10157 (N_10157,N_9822,N_9429);
nor U10158 (N_10158,N_8370,N_8696);
nor U10159 (N_10159,N_7691,N_7890);
nand U10160 (N_10160,N_9328,N_7977);
or U10161 (N_10161,N_8324,N_7631);
or U10162 (N_10162,N_9076,N_9788);
and U10163 (N_10163,N_9557,N_8635);
and U10164 (N_10164,N_7570,N_8547);
nor U10165 (N_10165,N_8596,N_8607);
and U10166 (N_10166,N_7685,N_8531);
nand U10167 (N_10167,N_8774,N_8767);
nor U10168 (N_10168,N_8705,N_8423);
and U10169 (N_10169,N_7627,N_8492);
xnor U10170 (N_10170,N_9450,N_8297);
or U10171 (N_10171,N_9508,N_8210);
xnor U10172 (N_10172,N_9154,N_8724);
or U10173 (N_10173,N_8994,N_9443);
or U10174 (N_10174,N_7656,N_8487);
xor U10175 (N_10175,N_9038,N_7797);
nand U10176 (N_10176,N_8553,N_8116);
xnor U10177 (N_10177,N_8717,N_9708);
or U10178 (N_10178,N_7617,N_7823);
nor U10179 (N_10179,N_9009,N_8197);
nand U10180 (N_10180,N_8503,N_9251);
xnor U10181 (N_10181,N_8900,N_8828);
and U10182 (N_10182,N_9668,N_9659);
xor U10183 (N_10183,N_7577,N_8738);
and U10184 (N_10184,N_9514,N_9292);
and U10185 (N_10185,N_7587,N_9490);
and U10186 (N_10186,N_9340,N_8711);
nand U10187 (N_10187,N_9670,N_8558);
or U10188 (N_10188,N_8498,N_8778);
xor U10189 (N_10189,N_8072,N_8293);
xor U10190 (N_10190,N_8918,N_8329);
xor U10191 (N_10191,N_9172,N_9071);
xor U10192 (N_10192,N_9424,N_9219);
nand U10193 (N_10193,N_8950,N_8163);
xnor U10194 (N_10194,N_9882,N_8202);
nand U10195 (N_10195,N_8022,N_9952);
and U10196 (N_10196,N_8017,N_8792);
nand U10197 (N_10197,N_8113,N_7941);
or U10198 (N_10198,N_9540,N_7585);
nand U10199 (N_10199,N_8139,N_8627);
or U10200 (N_10200,N_9164,N_7873);
xor U10201 (N_10201,N_9122,N_8255);
nor U10202 (N_10202,N_7601,N_8427);
nand U10203 (N_10203,N_9444,N_9379);
nand U10204 (N_10204,N_9096,N_9578);
nor U10205 (N_10205,N_9004,N_8869);
and U10206 (N_10206,N_8941,N_8083);
nand U10207 (N_10207,N_8095,N_9763);
or U10208 (N_10208,N_7690,N_8959);
xnor U10209 (N_10209,N_7748,N_9619);
nor U10210 (N_10210,N_9483,N_8451);
nand U10211 (N_10211,N_7678,N_7742);
or U10212 (N_10212,N_7817,N_7615);
nand U10213 (N_10213,N_9361,N_9598);
xnor U10214 (N_10214,N_8593,N_9561);
nand U10215 (N_10215,N_9864,N_8861);
nand U10216 (N_10216,N_7767,N_9696);
and U10217 (N_10217,N_8155,N_9387);
or U10218 (N_10218,N_7677,N_9116);
xnor U10219 (N_10219,N_8538,N_8749);
nor U10220 (N_10220,N_9319,N_7659);
nand U10221 (N_10221,N_9182,N_9280);
nand U10222 (N_10222,N_9137,N_8483);
nand U10223 (N_10223,N_8533,N_9586);
xor U10224 (N_10224,N_8067,N_8735);
xnor U10225 (N_10225,N_8335,N_7582);
xor U10226 (N_10226,N_9995,N_9065);
nand U10227 (N_10227,N_9371,N_8107);
nand U10228 (N_10228,N_9425,N_9199);
nand U10229 (N_10229,N_8290,N_8673);
nand U10230 (N_10230,N_8482,N_8512);
xnor U10231 (N_10231,N_8658,N_8264);
and U10232 (N_10232,N_7948,N_8809);
xor U10233 (N_10233,N_7856,N_8308);
nand U10234 (N_10234,N_9515,N_8562);
and U10235 (N_10235,N_8737,N_8074);
nor U10236 (N_10236,N_8611,N_8559);
or U10237 (N_10237,N_7839,N_9869);
nor U10238 (N_10238,N_9746,N_9481);
nand U10239 (N_10239,N_7899,N_8052);
xor U10240 (N_10240,N_7924,N_7938);
xnor U10241 (N_10241,N_7734,N_9936);
or U10242 (N_10242,N_8889,N_9974);
or U10243 (N_10243,N_9024,N_8015);
and U10244 (N_10244,N_8567,N_9607);
and U10245 (N_10245,N_8151,N_8118);
nor U10246 (N_10246,N_9841,N_8949);
nand U10247 (N_10247,N_9667,N_9468);
or U10248 (N_10248,N_7546,N_8243);
nand U10249 (N_10249,N_7560,N_7982);
xnor U10250 (N_10250,N_9625,N_8781);
nor U10251 (N_10251,N_7789,N_9200);
and U10252 (N_10252,N_9433,N_7833);
or U10253 (N_10253,N_8289,N_9842);
or U10254 (N_10254,N_8729,N_9834);
xor U10255 (N_10255,N_8319,N_8371);
and U10256 (N_10256,N_7713,N_7592);
nand U10257 (N_10257,N_7569,N_7894);
xor U10258 (N_10258,N_9077,N_8510);
nand U10259 (N_10259,N_9523,N_8699);
nand U10260 (N_10260,N_7766,N_7739);
xor U10261 (N_10261,N_8053,N_8680);
and U10262 (N_10262,N_8515,N_9599);
nand U10263 (N_10263,N_9042,N_9927);
nor U10264 (N_10264,N_9413,N_9639);
nand U10265 (N_10265,N_9944,N_9338);
and U10266 (N_10266,N_9820,N_8903);
nand U10267 (N_10267,N_9215,N_8479);
nand U10268 (N_10268,N_7531,N_8480);
or U10269 (N_10269,N_8316,N_7574);
or U10270 (N_10270,N_9289,N_8320);
and U10271 (N_10271,N_9382,N_9422);
or U10272 (N_10272,N_7553,N_8473);
nor U10273 (N_10273,N_9671,N_8615);
xnor U10274 (N_10274,N_8842,N_8396);
nand U10275 (N_10275,N_8338,N_8725);
and U10276 (N_10276,N_7863,N_7557);
nand U10277 (N_10277,N_9187,N_9547);
or U10278 (N_10278,N_8674,N_8250);
and U10279 (N_10279,N_7658,N_8401);
and U10280 (N_10280,N_8154,N_9496);
xnor U10281 (N_10281,N_9126,N_9110);
or U10282 (N_10282,N_9898,N_8660);
nor U10283 (N_10283,N_8168,N_8638);
xnor U10284 (N_10284,N_7709,N_8858);
or U10285 (N_10285,N_8392,N_9632);
xnor U10286 (N_10286,N_9596,N_9795);
nor U10287 (N_10287,N_9531,N_8980);
nor U10288 (N_10288,N_9571,N_8582);
or U10289 (N_10289,N_9955,N_8586);
nor U10290 (N_10290,N_7719,N_8351);
and U10291 (N_10291,N_9087,N_9152);
and U10292 (N_10292,N_8123,N_8847);
and U10293 (N_10293,N_9150,N_7651);
nor U10294 (N_10294,N_7556,N_8133);
nor U10295 (N_10295,N_7842,N_9717);
nand U10296 (N_10296,N_9587,N_9305);
and U10297 (N_10297,N_7808,N_7852);
nand U10298 (N_10298,N_8667,N_8456);
or U10299 (N_10299,N_9513,N_7537);
nor U10300 (N_10300,N_9127,N_9556);
nand U10301 (N_10301,N_9778,N_9120);
nor U10302 (N_10302,N_9405,N_7786);
nor U10303 (N_10303,N_9235,N_8311);
nand U10304 (N_10304,N_9147,N_9297);
xor U10305 (N_10305,N_8178,N_9649);
xnor U10306 (N_10306,N_9789,N_8598);
nor U10307 (N_10307,N_7681,N_8405);
xnor U10308 (N_10308,N_8502,N_8075);
and U10309 (N_10309,N_7921,N_9651);
and U10310 (N_10310,N_8691,N_9086);
xnor U10311 (N_10311,N_8734,N_8010);
nor U10312 (N_10312,N_9091,N_9933);
nor U10313 (N_10313,N_9461,N_9962);
nor U10314 (N_10314,N_7821,N_9186);
xor U10315 (N_10315,N_7518,N_7608);
nor U10316 (N_10316,N_9580,N_8981);
nor U10317 (N_10317,N_9498,N_8942);
nand U10318 (N_10318,N_9234,N_9181);
nand U10319 (N_10319,N_9934,N_7935);
nor U10320 (N_10320,N_7960,N_8821);
xnor U10321 (N_10321,N_9321,N_9534);
or U10322 (N_10322,N_9497,N_8127);
or U10323 (N_10323,N_8998,N_7559);
nand U10324 (N_10324,N_9434,N_8325);
and U10325 (N_10325,N_8879,N_8955);
nand U10326 (N_10326,N_9526,N_7731);
nand U10327 (N_10327,N_8991,N_9828);
xnor U10328 (N_10328,N_9904,N_8805);
nand U10329 (N_10329,N_7741,N_9672);
or U10330 (N_10330,N_7825,N_8261);
nor U10331 (N_10331,N_8211,N_8346);
and U10332 (N_10332,N_9350,N_7561);
xor U10333 (N_10333,N_9681,N_8406);
or U10334 (N_10334,N_8181,N_9241);
or U10335 (N_10335,N_7540,N_8466);
or U10336 (N_10336,N_9978,N_8369);
or U10337 (N_10337,N_9101,N_8521);
and U10338 (N_10338,N_7504,N_9665);
and U10339 (N_10339,N_9727,N_8399);
nor U10340 (N_10340,N_8101,N_9248);
nand U10341 (N_10341,N_8831,N_9363);
nand U10342 (N_10342,N_7914,N_9499);
and U10343 (N_10343,N_7536,N_8445);
nand U10344 (N_10344,N_7923,N_8645);
xor U10345 (N_10345,N_8356,N_8233);
and U10346 (N_10346,N_9312,N_9610);
xnor U10347 (N_10347,N_9192,N_9268);
nand U10348 (N_10348,N_7605,N_8432);
nor U10349 (N_10349,N_8084,N_8156);
and U10350 (N_10350,N_9766,N_9764);
and U10351 (N_10351,N_9119,N_9485);
xor U10352 (N_10352,N_7760,N_7999);
or U10353 (N_10353,N_9698,N_9726);
and U10354 (N_10354,N_9486,N_9738);
and U10355 (N_10355,N_9728,N_7901);
nand U10356 (N_10356,N_9896,N_8897);
nor U10357 (N_10357,N_8868,N_8060);
xor U10358 (N_10358,N_9781,N_8771);
nand U10359 (N_10359,N_9198,N_7942);
xor U10360 (N_10360,N_7933,N_7674);
or U10361 (N_10361,N_9644,N_9206);
and U10362 (N_10362,N_7931,N_9801);
nor U10363 (N_10363,N_7550,N_9229);
and U10364 (N_10364,N_8337,N_8036);
or U10365 (N_10365,N_8601,N_8653);
nand U10366 (N_10366,N_8336,N_8561);
nor U10367 (N_10367,N_9167,N_7620);
nor U10368 (N_10368,N_8603,N_9782);
nor U10369 (N_10369,N_9356,N_7866);
and U10370 (N_10370,N_8448,N_9381);
or U10371 (N_10371,N_9362,N_8284);
or U10372 (N_10372,N_8722,N_9702);
and U10373 (N_10373,N_8258,N_8770);
xnor U10374 (N_10374,N_8437,N_8625);
nand U10375 (N_10375,N_8508,N_8605);
xor U10376 (N_10376,N_9807,N_9970);
or U10377 (N_10377,N_8675,N_9089);
xnor U10378 (N_10378,N_8806,N_9437);
or U10379 (N_10379,N_7567,N_9941);
and U10380 (N_10380,N_8071,N_8937);
and U10381 (N_10381,N_8591,N_8049);
and U10382 (N_10382,N_9050,N_9504);
xor U10383 (N_10383,N_9637,N_8125);
nor U10384 (N_10384,N_9857,N_9118);
and U10385 (N_10385,N_8623,N_9045);
nor U10386 (N_10386,N_8140,N_8409);
or U10387 (N_10387,N_8249,N_9293);
xor U10388 (N_10388,N_7973,N_7972);
nor U10389 (N_10389,N_8424,N_7841);
and U10390 (N_10390,N_9479,N_7794);
and U10391 (N_10391,N_9783,N_9720);
or U10392 (N_10392,N_8494,N_9047);
nand U10393 (N_10393,N_8038,N_9153);
xor U10394 (N_10394,N_8137,N_9616);
nor U10395 (N_10395,N_9652,N_8470);
or U10396 (N_10396,N_7505,N_8914);
or U10397 (N_10397,N_7769,N_8085);
nand U10398 (N_10398,N_9262,N_8142);
and U10399 (N_10399,N_7597,N_8159);
xor U10400 (N_10400,N_8871,N_9072);
and U10401 (N_10401,N_8438,N_9345);
or U10402 (N_10402,N_8291,N_8807);
or U10403 (N_10403,N_9858,N_9037);
or U10404 (N_10404,N_9965,N_8906);
nor U10405 (N_10405,N_9151,N_9628);
or U10406 (N_10406,N_8373,N_9684);
or U10407 (N_10407,N_8930,N_9184);
and U10408 (N_10408,N_9860,N_8762);
and U10409 (N_10409,N_8236,N_9360);
and U10410 (N_10410,N_9462,N_9877);
xnor U10411 (N_10411,N_8435,N_8965);
or U10412 (N_10412,N_8162,N_7967);
nand U10413 (N_10413,N_7759,N_9418);
nor U10414 (N_10414,N_8463,N_9816);
xor U10415 (N_10415,N_8732,N_8069);
xor U10416 (N_10416,N_9837,N_7813);
xnor U10417 (N_10417,N_7809,N_8870);
nand U10418 (N_10418,N_8700,N_9592);
xor U10419 (N_10419,N_8543,N_8309);
nand U10420 (N_10420,N_9281,N_8678);
xor U10421 (N_10421,N_7544,N_8779);
nand U10422 (N_10422,N_8460,N_9654);
nand U10423 (N_10423,N_8086,N_9802);
nand U10424 (N_10424,N_8514,N_8226);
nand U10425 (N_10425,N_9569,N_9439);
or U10426 (N_10426,N_9718,N_9862);
and U10427 (N_10427,N_9749,N_9600);
or U10428 (N_10428,N_7774,N_7520);
nand U10429 (N_10429,N_8604,N_8121);
nor U10430 (N_10430,N_7936,N_7555);
or U10431 (N_10431,N_7954,N_9675);
or U10432 (N_10432,N_8895,N_8177);
nand U10433 (N_10433,N_8345,N_7614);
nand U10434 (N_10434,N_7882,N_9484);
nand U10435 (N_10435,N_8661,N_8447);
xor U10436 (N_10436,N_7986,N_7598);
nand U10437 (N_10437,N_8327,N_8759);
xor U10438 (N_10438,N_8988,N_8442);
or U10439 (N_10439,N_9724,N_9035);
and U10440 (N_10440,N_8589,N_9257);
xor U10441 (N_10441,N_8963,N_8136);
xnor U10442 (N_10442,N_9703,N_7634);
xnor U10443 (N_10443,N_9845,N_9922);
and U10444 (N_10444,N_8755,N_7684);
or U10445 (N_10445,N_9608,N_7642);
and U10446 (N_10446,N_8306,N_9815);
and U10447 (N_10447,N_7905,N_8650);
nor U10448 (N_10448,N_8124,N_9935);
nand U10449 (N_10449,N_8683,N_9377);
nor U10450 (N_10450,N_8788,N_8129);
or U10451 (N_10451,N_7744,N_9950);
xnor U10452 (N_10452,N_8785,N_8288);
nor U10453 (N_10453,N_8551,N_9448);
and U10454 (N_10454,N_8225,N_7575);
nor U10455 (N_10455,N_9430,N_8318);
xor U10456 (N_10456,N_7893,N_8223);
nand U10457 (N_10457,N_9658,N_7793);
nor U10458 (N_10458,N_8583,N_8070);
nor U10459 (N_10459,N_8272,N_9201);
or U10460 (N_10460,N_8404,N_9386);
nor U10461 (N_10461,N_9097,N_9840);
xor U10462 (N_10462,N_9367,N_8726);
and U10463 (N_10463,N_8746,N_8023);
nor U10464 (N_10464,N_9892,N_9022);
or U10465 (N_10465,N_9748,N_8153);
and U10466 (N_10466,N_8709,N_9300);
nand U10467 (N_10467,N_7732,N_9758);
or U10468 (N_10468,N_7886,N_8600);
and U10469 (N_10469,N_8135,N_7837);
or U10470 (N_10470,N_7937,N_9762);
and U10471 (N_10471,N_7953,N_9881);
nor U10472 (N_10472,N_9049,N_9976);
or U10473 (N_10473,N_9015,N_8195);
nor U10474 (N_10474,N_9279,N_9225);
xnor U10475 (N_10475,N_8920,N_9156);
or U10476 (N_10476,N_9564,N_8784);
and U10477 (N_10477,N_9438,N_9709);
nand U10478 (N_10478,N_9209,N_7699);
nor U10479 (N_10479,N_8633,N_7950);
xor U10480 (N_10480,N_8966,N_9355);
nor U10481 (N_10481,N_8260,N_9264);
nand U10482 (N_10482,N_8481,N_8548);
nand U10483 (N_10483,N_7889,N_8342);
xnor U10484 (N_10484,N_8706,N_7811);
nand U10485 (N_10485,N_8854,N_8899);
and U10486 (N_10486,N_7600,N_9919);
or U10487 (N_10487,N_9937,N_9453);
and U10488 (N_10488,N_8816,N_8167);
nor U10489 (N_10489,N_9886,N_8349);
nor U10490 (N_10490,N_9211,N_9551);
xnor U10491 (N_10491,N_8907,N_7581);
xor U10492 (N_10492,N_8954,N_8413);
nor U10493 (N_10493,N_8916,N_9189);
nand U10494 (N_10494,N_8656,N_8580);
and U10495 (N_10495,N_7957,N_9786);
nand U10496 (N_10496,N_7927,N_9274);
and U10497 (N_10497,N_8362,N_7644);
nand U10498 (N_10498,N_7694,N_8281);
xnor U10499 (N_10499,N_9638,N_7500);
xnor U10500 (N_10500,N_9288,N_7643);
xor U10501 (N_10501,N_7535,N_8058);
or U10502 (N_10502,N_9666,N_8912);
and U10503 (N_10503,N_9174,N_7737);
nor U10504 (N_10504,N_9823,N_8728);
xor U10505 (N_10505,N_9525,N_8554);
or U10506 (N_10506,N_9104,N_9793);
xnor U10507 (N_10507,N_9792,N_8511);
nor U10508 (N_10508,N_9613,N_9646);
or U10509 (N_10509,N_9591,N_8134);
or U10510 (N_10510,N_8990,N_8882);
and U10511 (N_10511,N_8363,N_8537);
and U10512 (N_10512,N_9716,N_7983);
xor U10513 (N_10513,N_8092,N_7705);
and U10514 (N_10514,N_8044,N_7554);
nor U10515 (N_10515,N_8305,N_8993);
or U10516 (N_10516,N_9875,N_8698);
nand U10517 (N_10517,N_8130,N_8609);
nor U10518 (N_10518,N_8585,N_7566);
or U10519 (N_10519,N_7572,N_8693);
xnor U10520 (N_10520,N_7565,N_8866);
nand U10521 (N_10521,N_8317,N_9622);
nor U10522 (N_10522,N_7853,N_9020);
xor U10523 (N_10523,N_7563,N_8565);
nand U10524 (N_10524,N_8014,N_7867);
or U10525 (N_10525,N_9302,N_9915);
nor U10526 (N_10526,N_9366,N_8782);
and U10527 (N_10527,N_9278,N_7773);
nor U10528 (N_10528,N_9222,N_9237);
xnor U10529 (N_10529,N_8849,N_9954);
or U10530 (N_10530,N_8995,N_7511);
nor U10531 (N_10531,N_7768,N_9029);
xnor U10532 (N_10532,N_9601,N_7916);
xnor U10533 (N_10533,N_9383,N_9230);
nor U10534 (N_10534,N_8799,N_8283);
nand U10535 (N_10535,N_8266,N_9033);
and U10536 (N_10536,N_8681,N_9204);
and U10537 (N_10537,N_7804,N_8588);
nand U10538 (N_10538,N_8383,N_7549);
xor U10539 (N_10539,N_8886,N_9146);
nor U10540 (N_10540,N_8221,N_8885);
nor U10541 (N_10541,N_8668,N_9165);
nor U10542 (N_10542,N_8632,N_9000);
and U10543 (N_10543,N_8274,N_9577);
and U10544 (N_10544,N_9063,N_7751);
and U10545 (N_10545,N_9105,N_9346);
nand U10546 (N_10546,N_8997,N_7949);
and U10547 (N_10547,N_7951,N_9918);
nor U10548 (N_10548,N_8682,N_9958);
nand U10549 (N_10549,N_8235,N_8220);
nand U10550 (N_10550,N_9889,N_8826);
xnor U10551 (N_10551,N_8815,N_8676);
nand U10552 (N_10552,N_8372,N_9233);
xnor U10553 (N_10553,N_8057,N_8944);
nor U10554 (N_10554,N_8186,N_8131);
nand U10555 (N_10555,N_9290,N_7579);
nor U10556 (N_10556,N_9589,N_9414);
nor U10557 (N_10557,N_7796,N_9081);
nand U10558 (N_10558,N_9419,N_7532);
nand U10559 (N_10559,N_7992,N_8951);
xor U10560 (N_10560,N_8663,N_7917);
nand U10561 (N_10561,N_8180,N_8417);
and U10562 (N_10562,N_9276,N_9643);
nor U10563 (N_10563,N_9991,N_9618);
xnor U10564 (N_10564,N_8394,N_8242);
or U10565 (N_10565,N_8122,N_9798);
xnor U10566 (N_10566,N_9981,N_9421);
nand U10567 (N_10567,N_9012,N_8462);
and U10568 (N_10568,N_9519,N_7667);
nand U10569 (N_10569,N_8672,N_7947);
nor U10570 (N_10570,N_8573,N_9203);
nor U10571 (N_10571,N_8214,N_8205);
nand U10572 (N_10572,N_8269,N_8689);
xnor U10573 (N_10573,N_9909,N_9707);
nor U10574 (N_10574,N_9100,N_8303);
and U10575 (N_10575,N_9409,N_9902);
or U10576 (N_10576,N_8946,N_7755);
or U10577 (N_10577,N_9917,N_8412);
nand U10578 (N_10578,N_7663,N_9907);
nand U10579 (N_10579,N_8814,N_8050);
xor U10580 (N_10580,N_8203,N_9759);
and U10581 (N_10581,N_8570,N_9817);
and U10582 (N_10582,N_8545,N_8355);
nand U10583 (N_10583,N_9085,N_7753);
nand U10584 (N_10584,N_8578,N_7787);
nand U10585 (N_10585,N_8924,N_8298);
nor U10586 (N_10586,N_8873,N_8852);
or U10587 (N_10587,N_7788,N_9923);
and U10588 (N_10588,N_7883,N_9030);
nand U10589 (N_10589,N_9541,N_8144);
nor U10590 (N_10590,N_9469,N_8103);
nor U10591 (N_10591,N_7703,N_8138);
and U10592 (N_10592,N_8388,N_7623);
nand U10593 (N_10593,N_8217,N_9401);
nand U10594 (N_10594,N_9412,N_8563);
or U10595 (N_10595,N_7589,N_9926);
xor U10596 (N_10596,N_8428,N_7962);
or U10597 (N_10597,N_9370,N_9634);
and U10598 (N_10598,N_8877,N_9124);
and U10599 (N_10599,N_9966,N_8671);
or U10600 (N_10600,N_8434,N_9683);
xnor U10601 (N_10601,N_8259,N_7835);
or U10602 (N_10602,N_8204,N_7610);
xnor U10603 (N_10603,N_7871,N_8522);
xnor U10604 (N_10604,N_7987,N_9254);
and U10605 (N_10605,N_8271,N_7622);
or U10606 (N_10606,N_8062,N_8368);
nor U10607 (N_10607,N_9121,N_7609);
nand U10608 (N_10608,N_8566,N_8378);
xnor U10609 (N_10609,N_9924,N_7879);
and U10610 (N_10610,N_8097,N_9477);
xor U10611 (N_10611,N_9575,N_9036);
xor U10612 (N_10612,N_9832,N_9520);
or U10613 (N_10613,N_7991,N_9190);
and U10614 (N_10614,N_9604,N_9427);
xnor U10615 (N_10615,N_7746,N_9850);
and U10616 (N_10616,N_8840,N_7649);
or U10617 (N_10617,N_9975,N_8334);
xnor U10618 (N_10618,N_7692,N_8708);
or U10619 (N_10619,N_7519,N_8652);
nand U10620 (N_10620,N_9179,N_9048);
nor U10621 (N_10621,N_9092,N_8051);
nand U10622 (N_10622,N_9744,N_9775);
nand U10623 (N_10623,N_9207,N_7514);
nand U10624 (N_10624,N_9890,N_8263);
xor U10625 (N_10625,N_9851,N_8340);
nand U10626 (N_10626,N_9028,N_9844);
xor U10627 (N_10627,N_8126,N_9391);
or U10628 (N_10628,N_8606,N_9780);
nor U10629 (N_10629,N_8517,N_9715);
nand U10630 (N_10630,N_7645,N_8257);
xor U10631 (N_10631,N_7740,N_8301);
xnor U10632 (N_10632,N_9277,N_9500);
and U10633 (N_10633,N_8331,N_8328);
xnor U10634 (N_10634,N_7978,N_7624);
nand U10635 (N_10635,N_8248,N_8364);
and U10636 (N_10636,N_9691,N_8703);
and U10637 (N_10637,N_8757,N_8485);
xnor U10638 (N_10638,N_9385,N_8253);
xnor U10639 (N_10639,N_8232,N_9987);
or U10640 (N_10640,N_8552,N_9971);
nor U10641 (N_10641,N_8931,N_8616);
xor U10642 (N_10642,N_8354,N_8820);
or U10643 (N_10643,N_7822,N_8662);
or U10644 (N_10644,N_8875,N_7971);
xnor U10645 (N_10645,N_9743,N_9392);
or U10646 (N_10646,N_7968,N_8824);
xnor U10647 (N_10647,N_9772,N_8386);
or U10648 (N_10648,N_7607,N_9602);
nor U10649 (N_10649,N_8106,N_8262);
and U10650 (N_10650,N_9399,N_9428);
xor U10651 (N_10651,N_9594,N_9258);
and U10652 (N_10652,N_9993,N_7771);
nor U10653 (N_10653,N_9471,N_7830);
xor U10654 (N_10654,N_8801,N_7862);
nor U10655 (N_10655,N_8252,N_7881);
nand U10656 (N_10656,N_8265,N_7745);
nand U10657 (N_10657,N_7646,N_8802);
nand U10658 (N_10658,N_9568,N_9894);
nand U10659 (N_10659,N_7718,N_7641);
xor U10660 (N_10660,N_9532,N_9455);
and U10661 (N_10661,N_8157,N_9947);
and U10662 (N_10662,N_9051,N_8829);
nand U10663 (N_10663,N_7847,N_8825);
and U10664 (N_10664,N_7819,N_9380);
nand U10665 (N_10665,N_8622,N_9474);
nand U10666 (N_10666,N_7591,N_9309);
or U10667 (N_10667,N_7860,N_7725);
or U10668 (N_10668,N_9870,N_9576);
or U10669 (N_10669,N_8564,N_9888);
and U10670 (N_10670,N_9784,N_7568);
nand U10671 (N_10671,N_9090,N_9210);
and U10672 (N_10672,N_7946,N_8380);
and U10673 (N_10673,N_9339,N_7993);
xor U10674 (N_10674,N_8381,N_8061);
nand U10675 (N_10675,N_7803,N_9059);
xor U10676 (N_10676,N_9636,N_8307);
xor U10677 (N_10677,N_9612,N_8206);
or U10678 (N_10678,N_8296,N_8836);
or U10679 (N_10679,N_8390,N_7529);
nor U10680 (N_10680,N_8246,N_8748);
and U10681 (N_10681,N_7981,N_9372);
and U10682 (N_10682,N_9559,N_8172);
or U10683 (N_10683,N_8509,N_7594);
or U10684 (N_10684,N_8943,N_9298);
nor U10685 (N_10685,N_9908,N_8377);
nand U10686 (N_10686,N_9574,N_7723);
xor U10687 (N_10687,N_7855,N_7621);
or U10688 (N_10688,N_7876,N_8867);
or U10689 (N_10689,N_8475,N_8500);
nand U10690 (N_10690,N_9061,N_8183);
or U10691 (N_10691,N_7508,N_9733);
or U10692 (N_10692,N_8196,N_8612);
nand U10693 (N_10693,N_9661,N_8029);
xor U10694 (N_10694,N_9501,N_8001);
nand U10695 (N_10695,N_8695,N_9195);
nand U10696 (N_10696,N_8207,N_7998);
and U10697 (N_10697,N_7629,N_9482);
xor U10698 (N_10698,N_7943,N_7516);
xor U10699 (N_10699,N_8933,N_7828);
and U10700 (N_10700,N_8714,N_8769);
and U10701 (N_10701,N_9375,N_8191);
or U10702 (N_10702,N_8114,N_9626);
nand U10703 (N_10703,N_9757,N_8111);
and U10704 (N_10704,N_9344,N_9040);
and U10705 (N_10705,N_9337,N_8045);
nor U10706 (N_10706,N_9982,N_9863);
and U10707 (N_10707,N_8375,N_8629);
or U10708 (N_10708,N_8568,N_9318);
xor U10709 (N_10709,N_9799,N_8670);
or U10710 (N_10710,N_8198,N_9313);
and U10711 (N_10711,N_9218,N_7655);
nor U10712 (N_10712,N_9062,N_9940);
xor U10713 (N_10713,N_8892,N_7653);
and U10714 (N_10714,N_9143,N_9369);
nand U10715 (N_10715,N_9068,N_8189);
nor U10716 (N_10716,N_7980,N_9645);
xnor U10717 (N_10717,N_8397,N_9614);
or U10718 (N_10718,N_7959,N_9895);
and U10719 (N_10719,N_8190,N_8636);
nand U10720 (N_10720,N_9291,N_9951);
and U10721 (N_10721,N_9492,N_9441);
and U10722 (N_10722,N_7955,N_8359);
xor U10723 (N_10723,N_9194,N_9013);
xnor U10724 (N_10724,N_8947,N_7743);
nor U10725 (N_10725,N_8241,N_8464);
or U10726 (N_10726,N_7716,N_8008);
nand U10727 (N_10727,N_7909,N_8043);
nor U10728 (N_10728,N_8247,N_8528);
and U10729 (N_10729,N_8796,N_7884);
or U10730 (N_10730,N_9641,N_7895);
and U10731 (N_10731,N_7548,N_9755);
xor U10732 (N_10732,N_7507,N_8228);
nor U10733 (N_10733,N_7715,N_8379);
nor U10734 (N_10734,N_8890,N_7782);
nor U10735 (N_10735,N_8832,N_9074);
nand U10736 (N_10736,N_9906,N_7925);
xor U10737 (N_10737,N_8555,N_8506);
nor U10738 (N_10738,N_7571,N_9159);
nand U10739 (N_10739,N_9785,N_8389);
xnor U10740 (N_10740,N_8024,N_9466);
nor U10741 (N_10741,N_9390,N_7934);
and U10742 (N_10742,N_9977,N_9185);
nor U10743 (N_10743,N_9243,N_8620);
nand U10744 (N_10744,N_8222,N_8999);
and U10745 (N_10745,N_9082,N_9740);
and U10746 (N_10746,N_8486,N_8326);
xnor U10747 (N_10747,N_9752,N_9572);
nor U10748 (N_10748,N_9463,N_9760);
and U10749 (N_10749,N_9803,N_9676);
nor U10750 (N_10750,N_8934,N_9544);
and U10751 (N_10751,N_9141,N_7688);
or U10752 (N_10752,N_9098,N_9158);
xnor U10753 (N_10753,N_7877,N_9879);
and U10754 (N_10754,N_8830,N_8975);
and U10755 (N_10755,N_7708,N_9731);
nand U10756 (N_10756,N_8476,N_9005);
nor U10757 (N_10757,N_8628,N_8002);
nand U10758 (N_10758,N_7919,N_8970);
nor U10759 (N_10759,N_7910,N_7749);
xor U10760 (N_10760,N_9964,N_9573);
nand U10761 (N_10761,N_9265,N_8637);
nand U10762 (N_10762,N_8694,N_8584);
and U10763 (N_10763,N_8430,N_9682);
nand U10764 (N_10764,N_9913,N_8702);
and U10765 (N_10765,N_8571,N_9213);
nand U10766 (N_10766,N_9872,N_8439);
nand U10767 (N_10767,N_8874,N_9548);
or U10768 (N_10768,N_7997,N_8690);
nand U10769 (N_10769,N_9010,N_8797);
nor U10770 (N_10770,N_9664,N_9358);
nand U10771 (N_10771,N_8688,N_9403);
xor U10772 (N_10772,N_9953,N_7625);
and U10773 (N_10773,N_8018,N_9070);
nor U10774 (N_10774,N_9079,N_7633);
xor U10775 (N_10775,N_7995,N_8465);
and U10776 (N_10776,N_7806,N_9960);
nand U10777 (N_10777,N_7904,N_8039);
nand U10778 (N_10778,N_7836,N_7829);
nor U10779 (N_10779,N_9761,N_9899);
xnor U10780 (N_10780,N_8147,N_7932);
or U10781 (N_10781,N_8646,N_8279);
xnor U10782 (N_10782,N_8712,N_9212);
nor U10783 (N_10783,N_8416,N_8992);
nor U10784 (N_10784,N_7851,N_8789);
nand U10785 (N_10785,N_9064,N_8519);
nand U10786 (N_10786,N_9825,N_9730);
xnor U10787 (N_10787,N_7586,N_9627);
or U10788 (N_10788,N_9725,N_8736);
or U10789 (N_10789,N_8030,N_9697);
and U10790 (N_10790,N_9729,N_7920);
and U10791 (N_10791,N_9562,N_9256);
and U10792 (N_10792,N_9445,N_8560);
xnor U10793 (N_10793,N_8750,N_8200);
or U10794 (N_10794,N_7845,N_7945);
nor U10795 (N_10795,N_9679,N_9402);
nand U10796 (N_10796,N_7673,N_9304);
and U10797 (N_10797,N_9244,N_8420);
or U10798 (N_10798,N_8913,N_8542);
nand U10799 (N_10799,N_9259,N_9996);
nor U10800 (N_10800,N_9972,N_8894);
nor U10801 (N_10801,N_8841,N_8893);
xnor U10802 (N_10802,N_9945,N_8648);
and U10803 (N_10803,N_9436,N_9831);
or U10804 (N_10804,N_7680,N_7724);
and U10805 (N_10805,N_7584,N_8507);
nand U10806 (N_10806,N_9472,N_7647);
or U10807 (N_10807,N_8642,N_7762);
xnor U10808 (N_10808,N_7857,N_8657);
or U10809 (N_10809,N_9836,N_8016);
and U10810 (N_10810,N_7784,N_8928);
or U10811 (N_10811,N_8744,N_9867);
or U10812 (N_10812,N_9352,N_9912);
nor U10813 (N_10813,N_8880,N_9685);
and U10814 (N_10814,N_7545,N_9075);
xor U10815 (N_10815,N_8956,N_9088);
and U10816 (N_10816,N_7780,N_9570);
nand U10817 (N_10817,N_8104,N_8032);
nand U10818 (N_10818,N_8273,N_8425);
xor U10819 (N_10819,N_9538,N_8721);
nand U10820 (N_10820,N_8610,N_9723);
or U10821 (N_10821,N_9750,N_7552);
nand U10822 (N_10822,N_7730,N_9099);
or U10823 (N_10823,N_8613,N_7912);
and U10824 (N_10824,N_9460,N_8285);
or U10825 (N_10825,N_8033,N_9330);
or U10826 (N_10826,N_9008,N_9142);
or U10827 (N_10827,N_9188,N_7911);
and U10828 (N_10828,N_8787,N_8501);
and U10829 (N_10829,N_8027,N_7930);
or U10830 (N_10830,N_9267,N_9224);
nand U10831 (N_10831,N_8777,N_8704);
nand U10832 (N_10832,N_8827,N_9303);
or U10833 (N_10833,N_9739,N_9989);
xnor U10834 (N_10834,N_8932,N_8530);
nand U10835 (N_10835,N_7885,N_8426);
and U10836 (N_10836,N_8185,N_8786);
nand U10837 (N_10837,N_9406,N_9713);
nor U10838 (N_10838,N_7534,N_8716);
nand U10839 (N_10839,N_8597,N_9359);
or U10840 (N_10840,N_9843,N_8278);
nand U10841 (N_10841,N_9517,N_9163);
nor U10842 (N_10842,N_9826,N_9595);
xor U10843 (N_10843,N_8237,N_8398);
or U10844 (N_10844,N_8469,N_8768);
nand U10845 (N_10845,N_8864,N_8967);
nor U10846 (N_10846,N_8978,N_8165);
xnor U10847 (N_10847,N_9044,N_9133);
nand U10848 (N_10848,N_9226,N_8550);
and U10849 (N_10849,N_9315,N_8957);
and U10850 (N_10850,N_8440,N_7781);
or U10851 (N_10851,N_9113,N_9408);
nand U10852 (N_10852,N_8367,N_8727);
nand U10853 (N_10853,N_8839,N_9311);
nor U10854 (N_10854,N_9554,N_9411);
nor U10855 (N_10855,N_7906,N_9939);
nor U10856 (N_10856,N_9553,N_9656);
nor U10857 (N_10857,N_9261,N_8187);
xor U10858 (N_10858,N_7765,N_9994);
and U10859 (N_10859,N_8798,N_9901);
xor U10860 (N_10860,N_9157,N_9903);
nand U10861 (N_10861,N_9320,N_9694);
xnor U10862 (N_10862,N_8280,N_9080);
nand U10863 (N_10863,N_7619,N_8452);
or U10864 (N_10864,N_8299,N_9533);
nand U10865 (N_10865,N_7757,N_9208);
xor U10866 (N_10866,N_8478,N_8193);
or U10867 (N_10867,N_8450,N_8819);
and U10868 (N_10868,N_8715,N_9813);
and U10869 (N_10869,N_7961,N_7512);
nand U10870 (N_10870,N_8982,N_8692);
xnor U10871 (N_10871,N_9819,N_9323);
nand U10872 (N_10872,N_9395,N_8361);
nor U10873 (N_10873,N_8387,N_7626);
and U10874 (N_10874,N_9988,N_9855);
nor U10875 (N_10875,N_9754,N_9066);
nand U10876 (N_10876,N_7580,N_8188);
or U10877 (N_10877,N_7988,N_8422);
and U10878 (N_10878,N_9459,N_7671);
xnor U10879 (N_10879,N_7844,N_9910);
nor U10880 (N_10880,N_9770,N_7722);
nor U10881 (N_10881,N_9054,N_9916);
nand U10882 (N_10882,N_8904,N_9997);
nand U10883 (N_10883,N_9041,N_8227);
nor U10884 (N_10884,N_8835,N_8411);
and U10885 (N_10885,N_8783,N_9078);
and U10886 (N_10886,N_9177,N_8516);
nand U10887 (N_10887,N_9835,N_7686);
nor U10888 (N_10888,N_9686,N_9605);
nand U10889 (N_10889,N_9810,N_9007);
and U10890 (N_10890,N_8576,N_8294);
xor U10891 (N_10891,N_8539,N_8742);
nand U10892 (N_10892,N_8863,N_9247);
xor U10893 (N_10893,N_9921,N_8056);
xnor U10894 (N_10894,N_9467,N_9322);
nor U10895 (N_10895,N_9094,N_8034);
nor U10896 (N_10896,N_8357,N_9555);
nor U10897 (N_10897,N_8454,N_8865);
nor U10898 (N_10898,N_8626,N_9394);
nand U10899 (N_10899,N_9239,N_9753);
and U10900 (N_10900,N_9973,N_9543);
and U10901 (N_10901,N_8152,N_7738);
or U10902 (N_10902,N_8011,N_7503);
or U10903 (N_10903,N_9106,N_8883);
and U10904 (N_10904,N_9767,N_9162);
xor U10905 (N_10905,N_9949,N_8925);
and U10906 (N_10906,N_9384,N_8004);
or U10907 (N_10907,N_9948,N_8763);
nor U10908 (N_10908,N_9756,N_9506);
nor U10909 (N_10909,N_9223,N_8491);
nand U10910 (N_10910,N_9306,N_9452);
xor U10911 (N_10911,N_8199,N_9502);
or U10912 (N_10912,N_8208,N_8215);
nand U10913 (N_10913,N_7779,N_9866);
xnor U10914 (N_10914,N_8414,N_7652);
or U10915 (N_10915,N_7975,N_7542);
xnor U10916 (N_10916,N_9324,N_8624);
and U10917 (N_10917,N_8640,N_7670);
and U10918 (N_10918,N_9388,N_9522);
and U10919 (N_10919,N_8891,N_9549);
nand U10920 (N_10920,N_8330,N_9351);
or U10921 (N_10921,N_7778,N_8594);
or U10922 (N_10922,N_9516,N_8775);
xor U10923 (N_10923,N_7603,N_9205);
or U10924 (N_10924,N_9967,N_8665);
xnor U10925 (N_10925,N_8527,N_9911);
nand U10926 (N_10926,N_7639,N_8429);
nor U10927 (N_10927,N_7802,N_9563);
and U10928 (N_10928,N_8751,N_9112);
and U10929 (N_10929,N_8898,N_8687);
nand U10930 (N_10930,N_9704,N_9928);
nand U10931 (N_10931,N_8251,N_9769);
and U10932 (N_10932,N_9566,N_8194);
nor U10933 (N_10933,N_9998,N_9511);
or U10934 (N_10934,N_9938,N_9168);
xnor U10935 (N_10935,N_7974,N_9593);
nor U10936 (N_10936,N_9647,N_8240);
nand U10937 (N_10937,N_7902,N_7717);
nor U10938 (N_10938,N_9027,N_7846);
nor U10939 (N_10939,N_9132,N_8132);
xor U10940 (N_10940,N_9314,N_9376);
and U10941 (N_10941,N_8756,N_9932);
and U10942 (N_10942,N_9002,N_7606);
xor U10943 (N_10943,N_9446,N_8800);
nand U10944 (N_10944,N_8012,N_8664);
and U10945 (N_10945,N_9527,N_9979);
xnor U10946 (N_10946,N_8149,N_9420);
and U10947 (N_10947,N_7831,N_9883);
and U10948 (N_10948,N_8958,N_9478);
xor U10949 (N_10949,N_8128,N_8444);
nor U10950 (N_10950,N_9680,N_9255);
and U10951 (N_10951,N_8119,N_8109);
xor U10952 (N_10952,N_8843,N_8649);
and U10953 (N_10953,N_9677,N_8219);
nor U10954 (N_10954,N_8856,N_8489);
or U10955 (N_10955,N_8449,N_7747);
xor U10956 (N_10956,N_8322,N_9706);
nand U10957 (N_10957,N_9270,N_9404);
and U10958 (N_10958,N_7772,N_8518);
nand U10959 (N_10959,N_8720,N_8209);
and U10960 (N_10960,N_9285,N_7515);
nand U10961 (N_10961,N_9615,N_9397);
nand U10962 (N_10962,N_7664,N_8192);
nor U10963 (N_10963,N_9253,N_8851);
nor U10964 (N_10964,N_9155,N_8765);
or U10965 (N_10965,N_9093,N_8608);
nand U10966 (N_10966,N_8433,N_8150);
and U10967 (N_10967,N_7864,N_8110);
or U10968 (N_10968,N_8146,N_9011);
xor U10969 (N_10969,N_9914,N_9633);
xnor U10970 (N_10970,N_8723,N_7669);
or U10971 (N_10971,N_8761,N_9545);
xnor U10972 (N_10972,N_8254,N_8753);
or U10973 (N_10973,N_8076,N_8366);
nor U10974 (N_10974,N_8651,N_8639);
nor U10975 (N_10975,N_9398,N_9202);
nor U10976 (N_10976,N_8046,N_8973);
nor U10977 (N_10977,N_9747,N_7679);
xnor U10978 (N_10978,N_9510,N_8896);
and U10979 (N_10979,N_8148,N_8876);
and U10980 (N_10980,N_7697,N_8556);
and U10981 (N_10981,N_7869,N_7810);
or U10982 (N_10982,N_7826,N_8350);
nor U10983 (N_10983,N_9125,N_9876);
nor U10984 (N_10984,N_9216,N_9014);
nor U10985 (N_10985,N_7989,N_7976);
and U10986 (N_10986,N_7870,N_8655);
nand U10987 (N_10987,N_8041,N_8312);
xnor U10988 (N_10988,N_9521,N_8927);
nand U10989 (N_10989,N_7735,N_8419);
nor U10990 (N_10990,N_9536,N_8115);
or U10991 (N_10991,N_8457,N_9590);
or U10992 (N_10992,N_8905,N_9507);
or U10993 (N_10993,N_8850,N_8754);
or U10994 (N_10994,N_8230,N_7907);
nor U10995 (N_10995,N_9968,N_8926);
xor U10996 (N_10996,N_8496,N_7599);
and U10997 (N_10997,N_8793,N_8082);
xor U10998 (N_10998,N_7517,N_9494);
nor U10999 (N_10999,N_7750,N_9742);
and U11000 (N_11000,N_8804,N_9473);
nand U11001 (N_11001,N_8042,N_9961);
and U11002 (N_11002,N_9985,N_9144);
xnor U11003 (N_11003,N_8647,N_7564);
nand U11004 (N_11004,N_9806,N_8087);
nor U11005 (N_11005,N_9585,N_9885);
xor U11006 (N_11006,N_9537,N_8376);
nor U11007 (N_11007,N_9505,N_9245);
and U11008 (N_11008,N_8654,N_8169);
or U11009 (N_11009,N_8595,N_8535);
nand U11010 (N_11010,N_9830,N_7583);
xor U11011 (N_11011,N_8969,N_8812);
or U11012 (N_11012,N_7640,N_9714);
xor U11013 (N_11013,N_9693,N_7729);
and U11014 (N_11014,N_8752,N_9546);
nand U11015 (N_11015,N_7834,N_8003);
nand U11016 (N_11016,N_7628,N_8234);
and U11017 (N_11017,N_9067,N_9509);
xor U11018 (N_11018,N_7994,N_9458);
and U11019 (N_11019,N_9539,N_8536);
or U11020 (N_11020,N_9797,N_8713);
or U11021 (N_11021,N_9475,N_8569);
nand U11022 (N_11022,N_9930,N_8773);
nor U11023 (N_11023,N_7650,N_7616);
and U11024 (N_11024,N_7558,N_8833);
and U11025 (N_11025,N_8332,N_9240);
and U11026 (N_11026,N_9417,N_8935);
and U11027 (N_11027,N_9847,N_8987);
xnor U11028 (N_11028,N_8078,N_9272);
nand U11029 (N_11029,N_8685,N_7922);
nand U11030 (N_11030,N_9006,N_9095);
and U11031 (N_11031,N_8182,N_9084);
nor U11032 (N_11032,N_7843,N_7915);
xnor U11033 (N_11033,N_9284,N_9984);
and U11034 (N_11034,N_9246,N_8213);
or U11035 (N_11035,N_8961,N_7763);
or U11036 (N_11036,N_7513,N_8231);
nor U11037 (N_11037,N_9771,N_9307);
nor U11038 (N_11038,N_9581,N_9115);
or U11039 (N_11039,N_9992,N_7630);
nor U11040 (N_11040,N_8731,N_7687);
xor U11041 (N_11041,N_9621,N_7824);
nand U11042 (N_11042,N_7602,N_8020);
and U11043 (N_11043,N_9878,N_8141);
and U11044 (N_11044,N_7695,N_7892);
nor U11045 (N_11045,N_8395,N_9333);
and U11046 (N_11046,N_9193,N_9476);
nor U11047 (N_11047,N_9021,N_8936);
and U11048 (N_11048,N_9464,N_9349);
and U11049 (N_11049,N_8526,N_8077);
xor U11050 (N_11050,N_9560,N_8488);
nand U11051 (N_11051,N_7865,N_9252);
nor U11052 (N_11052,N_7880,N_9629);
nor U11053 (N_11053,N_8292,N_9396);
or U11054 (N_11054,N_7533,N_7521);
nor U11055 (N_11055,N_7527,N_7593);
nor U11056 (N_11056,N_9287,N_8474);
xor U11057 (N_11057,N_9301,N_8229);
nor U11058 (N_11058,N_9849,N_9221);
xnor U11059 (N_11059,N_7985,N_9631);
and U11060 (N_11060,N_8599,N_8845);
and U11061 (N_11061,N_9719,N_8803);
or U11062 (N_11062,N_9018,N_8592);
nor U11063 (N_11063,N_8019,N_8344);
nor U11064 (N_11064,N_8838,N_9838);
or U11065 (N_11065,N_9456,N_9454);
or U11066 (N_11066,N_9905,N_9897);
nand U11067 (N_11067,N_8096,N_9524);
nor U11068 (N_11068,N_7872,N_9166);
and U11069 (N_11069,N_7578,N_8701);
or U11070 (N_11070,N_8621,N_8164);
or U11071 (N_11071,N_9839,N_8574);
xnor U11072 (N_11072,N_7799,N_9712);
nand U11073 (N_11073,N_9138,N_8175);
and U11074 (N_11074,N_9134,N_9765);
and U11075 (N_11075,N_8238,N_8467);
nand U11076 (N_11076,N_7783,N_9451);
xnor U11077 (N_11077,N_8021,N_8458);
nand U11078 (N_11078,N_9236,N_8099);
and U11079 (N_11079,N_9108,N_9859);
nor U11080 (N_11080,N_8971,N_7662);
nor U11081 (N_11081,N_7551,N_9741);
nand U11082 (N_11082,N_9470,N_8276);
or U11083 (N_11083,N_9736,N_8472);
or U11084 (N_11084,N_9083,N_9196);
nor U11085 (N_11085,N_8277,N_7979);
and U11086 (N_11086,N_7996,N_9052);
and U11087 (N_11087,N_9768,N_8602);
or U11088 (N_11088,N_8358,N_9660);
nor U11089 (N_11089,N_9735,N_9946);
nand U11090 (N_11090,N_9699,N_7832);
nand U11091 (N_11091,N_9800,N_9214);
nor U11092 (N_11092,N_7908,N_9431);
xor U11093 (N_11093,N_7547,N_8418);
nor U11094 (N_11094,N_8996,N_8468);
nand U11095 (N_11095,N_8117,N_8441);
or U11096 (N_11096,N_9325,N_9848);
and U11097 (N_11097,N_7807,N_8055);
and U11098 (N_11098,N_7721,N_8808);
nor U11099 (N_11099,N_8073,N_7675);
and U11100 (N_11100,N_9161,N_9777);
xor U11101 (N_11101,N_8529,N_9149);
nand U11102 (N_11102,N_8760,N_8089);
nor U11103 (N_11103,N_9787,N_7875);
or U11104 (N_11104,N_8857,N_8811);
or U11105 (N_11105,N_8710,N_9980);
or U11106 (N_11106,N_8577,N_8081);
or U11107 (N_11107,N_8659,N_9854);
and U11108 (N_11108,N_9550,N_9069);
xor U11109 (N_11109,N_9136,N_9669);
nor U11110 (N_11110,N_9178,N_7590);
xnor U11111 (N_11111,N_9874,N_9273);
nand U11112 (N_11112,N_7858,N_7733);
nand U11113 (N_11113,N_9588,N_7501);
nand U11114 (N_11114,N_8173,N_9073);
and U11115 (N_11115,N_7612,N_7939);
and U11116 (N_11116,N_8267,N_9796);
or U11117 (N_11117,N_7712,N_8719);
or U11118 (N_11118,N_7903,N_8848);
xor U11119 (N_11119,N_8743,N_7958);
xnor U11120 (N_11120,N_9373,N_8048);
nor U11121 (N_11121,N_8490,N_7761);
and U11122 (N_11122,N_7800,N_9530);
or U11123 (N_11123,N_8314,N_9791);
nand U11124 (N_11124,N_8888,N_9393);
and U11125 (N_11125,N_8968,N_7758);
or U11126 (N_11126,N_8446,N_8158);
xor U11127 (N_11127,N_8171,N_9347);
xnor U11128 (N_11128,N_9336,N_7840);
xnor U11129 (N_11129,N_9833,N_8860);
or U11130 (N_11130,N_9732,N_8403);
or U11131 (N_11131,N_8415,N_9642);
nor U11132 (N_11132,N_7795,N_9700);
and U11133 (N_11133,N_7798,N_9410);
xor U11134 (N_11134,N_9334,N_8579);
and U11135 (N_11135,N_8557,N_9624);
xnor U11136 (N_11136,N_7538,N_9821);
nor U11137 (N_11137,N_9145,N_8339);
nor U11138 (N_11138,N_9931,N_9426);
xnor U11139 (N_11139,N_9296,N_8028);
nand U11140 (N_11140,N_7816,N_8938);
xnor U11141 (N_11141,N_8733,N_9692);
xnor U11142 (N_11142,N_9929,N_9880);
nor U11143 (N_11143,N_9689,N_9332);
nor U11144 (N_11144,N_7964,N_9688);
and U11145 (N_11145,N_9663,N_8035);
and U11146 (N_11146,N_7900,N_7776);
and U11147 (N_11147,N_7736,N_9435);
or U11148 (N_11148,N_9582,N_7654);
xor U11149 (N_11149,N_7965,N_7525);
or U11150 (N_11150,N_7676,N_7714);
nand U11151 (N_11151,N_9139,N_8974);
nand U11152 (N_11152,N_9103,N_8391);
or U11153 (N_11153,N_8407,N_7801);
nand U11154 (N_11154,N_7838,N_9650);
and U11155 (N_11155,N_8453,N_8244);
nand U11156 (N_11156,N_9294,N_8352);
xor U11157 (N_11157,N_8972,N_8544);
and U11158 (N_11158,N_8216,N_9111);
nand U11159 (N_11159,N_8617,N_9711);
xor U11160 (N_11160,N_9774,N_8270);
or U11161 (N_11161,N_7576,N_7944);
nand U11162 (N_11162,N_8505,N_9579);
and U11163 (N_11163,N_8911,N_9969);
nor U11164 (N_11164,N_9457,N_9316);
xor U11165 (N_11165,N_8917,N_9275);
and U11166 (N_11166,N_8497,N_7635);
and U11167 (N_11167,N_8730,N_8541);
or U11168 (N_11168,N_9963,N_8170);
nor U11169 (N_11169,N_8758,N_8341);
or U11170 (N_11170,N_8102,N_8780);
xor U11171 (N_11171,N_8304,N_9001);
and U11172 (N_11172,N_8493,N_9503);
or U11173 (N_11173,N_8862,N_9440);
nor U11174 (N_11174,N_9983,N_9423);
xor U11175 (N_11175,N_9956,N_7820);
or U11176 (N_11176,N_8201,N_8817);
and U11177 (N_11177,N_8006,N_9999);
nand U11178 (N_11178,N_7868,N_8921);
and U11179 (N_11179,N_9043,N_9220);
xor U11180 (N_11180,N_9227,N_9003);
or U11181 (N_11181,N_9331,N_9893);
nor U11182 (N_11182,N_7700,N_8408);
and U11183 (N_11183,N_8855,N_8859);
nand U11184 (N_11184,N_8063,N_7928);
nor U11185 (N_11185,N_8908,N_8047);
and U11186 (N_11186,N_8108,N_8587);
or U11187 (N_11187,N_8360,N_8844);
xnor U11188 (N_11188,N_9597,N_9528);
and U11189 (N_11189,N_8745,N_8922);
xnor U11190 (N_11190,N_8534,N_7854);
xor U11191 (N_11191,N_9512,N_8952);
nand U11192 (N_11192,N_8677,N_9183);
and U11193 (N_11193,N_7682,N_7850);
and U11194 (N_11194,N_8054,N_8504);
or U11195 (N_11195,N_9357,N_9432);
nand U11196 (N_11196,N_8520,N_7720);
nor U11197 (N_11197,N_7913,N_8461);
xor U11198 (N_11198,N_7502,N_7706);
or U11199 (N_11199,N_8614,N_9630);
nor U11200 (N_11200,N_9368,N_9329);
and U11201 (N_11201,N_7849,N_8374);
xnor U11202 (N_11202,N_9242,N_9135);
nand U11203 (N_11203,N_8881,N_7827);
and U11204 (N_11204,N_7814,N_8410);
nand U11205 (N_11205,N_9299,N_8919);
nand U11206 (N_11206,N_9814,N_7506);
nand U11207 (N_11207,N_8212,N_8884);
nor U11208 (N_11208,N_8026,N_8948);
and U11209 (N_11209,N_9623,N_7666);
nand U11210 (N_11210,N_8546,N_8644);
nand U11211 (N_11211,N_8385,N_8984);
and U11212 (N_11212,N_9310,N_9891);
nor U11213 (N_11213,N_9416,N_9808);
xnor U11214 (N_11214,N_9365,N_7683);
nor U11215 (N_11215,N_7791,N_7874);
nand U11216 (N_11216,N_9389,N_8007);
nand U11217 (N_11217,N_8094,N_7696);
or U11218 (N_11218,N_8321,N_7970);
or U11219 (N_11219,N_9197,N_8697);
nand U11220 (N_11220,N_9056,N_7990);
or U11221 (N_11221,N_7632,N_8091);
xor U11222 (N_11222,N_9217,N_9829);
and U11223 (N_11223,N_8590,N_9341);
nand U11224 (N_11224,N_8239,N_9552);
nor U11225 (N_11225,N_8098,N_8343);
nor U11226 (N_11226,N_8040,N_7969);
and U11227 (N_11227,N_9609,N_9846);
and U11228 (N_11228,N_9342,N_9327);
nor U11229 (N_11229,N_9129,N_7785);
or U11230 (N_11230,N_7805,N_9603);
nand U11231 (N_11231,N_8315,N_7704);
or U11232 (N_11232,N_9655,N_8333);
nor U11233 (N_11233,N_8145,N_8740);
or U11234 (N_11234,N_9231,N_8436);
or U11235 (N_11235,N_8669,N_9128);
and U11236 (N_11236,N_9734,N_8643);
and U11237 (N_11237,N_8443,N_8499);
nand U11238 (N_11238,N_9148,N_9565);
or U11239 (N_11239,N_9238,N_9308);
nand U11240 (N_11240,N_8300,N_8484);
nand U11241 (N_11241,N_9794,N_9925);
nor U11242 (N_11242,N_9856,N_7661);
nor U11243 (N_11243,N_9271,N_8184);
and U11244 (N_11244,N_8282,N_7711);
xor U11245 (N_11245,N_9232,N_7707);
and U11246 (N_11246,N_9019,N_9031);
xor U11247 (N_11247,N_9266,N_8068);
and U11248 (N_11248,N_7926,N_9335);
nand U11249 (N_11249,N_9140,N_8718);
xor U11250 (N_11250,N_7541,N_8776);
nor U11251 (N_11251,N_8728,N_9569);
or U11252 (N_11252,N_8857,N_8039);
xnor U11253 (N_11253,N_7786,N_8153);
or U11254 (N_11254,N_8488,N_8087);
nand U11255 (N_11255,N_7836,N_9907);
and U11256 (N_11256,N_9004,N_9525);
nand U11257 (N_11257,N_8763,N_9711);
and U11258 (N_11258,N_8628,N_9635);
xor U11259 (N_11259,N_8468,N_8571);
nand U11260 (N_11260,N_7781,N_9838);
and U11261 (N_11261,N_9124,N_9487);
nor U11262 (N_11262,N_8311,N_7780);
nor U11263 (N_11263,N_9878,N_8731);
and U11264 (N_11264,N_9794,N_8485);
and U11265 (N_11265,N_8478,N_8609);
nor U11266 (N_11266,N_9819,N_9032);
nor U11267 (N_11267,N_8607,N_9050);
nor U11268 (N_11268,N_9534,N_9949);
nor U11269 (N_11269,N_8076,N_8866);
nor U11270 (N_11270,N_7982,N_8904);
nand U11271 (N_11271,N_7887,N_9934);
nor U11272 (N_11272,N_8854,N_9688);
xor U11273 (N_11273,N_8967,N_8243);
and U11274 (N_11274,N_9609,N_9496);
xnor U11275 (N_11275,N_9502,N_9861);
and U11276 (N_11276,N_7520,N_8290);
nand U11277 (N_11277,N_9017,N_8224);
xor U11278 (N_11278,N_8755,N_8238);
or U11279 (N_11279,N_9928,N_7677);
nand U11280 (N_11280,N_8183,N_9370);
or U11281 (N_11281,N_8606,N_7586);
or U11282 (N_11282,N_7593,N_9577);
xor U11283 (N_11283,N_8958,N_9275);
xor U11284 (N_11284,N_8330,N_8295);
or U11285 (N_11285,N_8943,N_8227);
xnor U11286 (N_11286,N_8589,N_8310);
xor U11287 (N_11287,N_8350,N_9310);
or U11288 (N_11288,N_9861,N_9977);
xor U11289 (N_11289,N_9982,N_9533);
xnor U11290 (N_11290,N_9494,N_7946);
xnor U11291 (N_11291,N_8058,N_8340);
xor U11292 (N_11292,N_8017,N_8993);
nor U11293 (N_11293,N_7645,N_9201);
nor U11294 (N_11294,N_9631,N_8043);
or U11295 (N_11295,N_8057,N_8741);
nor U11296 (N_11296,N_8341,N_7995);
or U11297 (N_11297,N_8341,N_7970);
nand U11298 (N_11298,N_9402,N_9032);
or U11299 (N_11299,N_8035,N_9982);
xnor U11300 (N_11300,N_8592,N_9493);
and U11301 (N_11301,N_9737,N_8461);
xnor U11302 (N_11302,N_9057,N_9959);
nor U11303 (N_11303,N_8437,N_8073);
or U11304 (N_11304,N_7950,N_7600);
nor U11305 (N_11305,N_7596,N_9765);
and U11306 (N_11306,N_9615,N_8584);
nor U11307 (N_11307,N_7810,N_7607);
nor U11308 (N_11308,N_8958,N_8369);
or U11309 (N_11309,N_8013,N_8208);
nand U11310 (N_11310,N_8295,N_9699);
or U11311 (N_11311,N_9517,N_9308);
nor U11312 (N_11312,N_7826,N_9729);
or U11313 (N_11313,N_8042,N_7873);
and U11314 (N_11314,N_8581,N_8941);
nand U11315 (N_11315,N_8061,N_9325);
nand U11316 (N_11316,N_7877,N_9873);
and U11317 (N_11317,N_8325,N_7584);
and U11318 (N_11318,N_9357,N_9878);
or U11319 (N_11319,N_9516,N_8268);
nor U11320 (N_11320,N_8173,N_8860);
nor U11321 (N_11321,N_7931,N_9749);
and U11322 (N_11322,N_9168,N_9349);
or U11323 (N_11323,N_7688,N_9060);
nand U11324 (N_11324,N_8068,N_9200);
xor U11325 (N_11325,N_8477,N_8583);
xor U11326 (N_11326,N_9041,N_8700);
nor U11327 (N_11327,N_9207,N_8632);
nand U11328 (N_11328,N_9579,N_8390);
nand U11329 (N_11329,N_9952,N_9729);
nand U11330 (N_11330,N_8291,N_8758);
or U11331 (N_11331,N_8250,N_8246);
or U11332 (N_11332,N_9501,N_7605);
or U11333 (N_11333,N_8057,N_9841);
xor U11334 (N_11334,N_7929,N_9075);
and U11335 (N_11335,N_8311,N_8105);
xnor U11336 (N_11336,N_7763,N_9806);
nor U11337 (N_11337,N_8965,N_9667);
nor U11338 (N_11338,N_9426,N_8368);
and U11339 (N_11339,N_7751,N_7894);
or U11340 (N_11340,N_9249,N_8651);
nand U11341 (N_11341,N_9602,N_7922);
nor U11342 (N_11342,N_9311,N_9839);
nor U11343 (N_11343,N_7511,N_8132);
xnor U11344 (N_11344,N_9418,N_9880);
nand U11345 (N_11345,N_9778,N_9723);
and U11346 (N_11346,N_9230,N_8427);
nand U11347 (N_11347,N_7583,N_7700);
nand U11348 (N_11348,N_9211,N_9060);
nand U11349 (N_11349,N_8928,N_9031);
and U11350 (N_11350,N_9327,N_7788);
nand U11351 (N_11351,N_8102,N_8802);
and U11352 (N_11352,N_9915,N_9881);
nand U11353 (N_11353,N_8186,N_7615);
or U11354 (N_11354,N_8219,N_8662);
xor U11355 (N_11355,N_9883,N_9915);
nand U11356 (N_11356,N_7739,N_8198);
nor U11357 (N_11357,N_8774,N_8908);
xor U11358 (N_11358,N_7536,N_7646);
or U11359 (N_11359,N_8510,N_9260);
xor U11360 (N_11360,N_8069,N_9578);
xor U11361 (N_11361,N_9296,N_7945);
xnor U11362 (N_11362,N_8750,N_7576);
and U11363 (N_11363,N_9053,N_8492);
nand U11364 (N_11364,N_7686,N_8902);
nand U11365 (N_11365,N_8737,N_9209);
or U11366 (N_11366,N_9665,N_8569);
nor U11367 (N_11367,N_8383,N_9061);
and U11368 (N_11368,N_8503,N_9407);
or U11369 (N_11369,N_8455,N_9708);
or U11370 (N_11370,N_9166,N_7946);
or U11371 (N_11371,N_8494,N_8626);
and U11372 (N_11372,N_9340,N_7706);
xor U11373 (N_11373,N_9704,N_9468);
xnor U11374 (N_11374,N_7840,N_8235);
and U11375 (N_11375,N_9777,N_9542);
nor U11376 (N_11376,N_8567,N_8143);
or U11377 (N_11377,N_9698,N_7625);
or U11378 (N_11378,N_9246,N_9542);
nand U11379 (N_11379,N_9552,N_8723);
or U11380 (N_11380,N_7580,N_7610);
xnor U11381 (N_11381,N_8181,N_9516);
and U11382 (N_11382,N_7961,N_9459);
or U11383 (N_11383,N_8993,N_9896);
xnor U11384 (N_11384,N_7671,N_9500);
and U11385 (N_11385,N_9414,N_7868);
nor U11386 (N_11386,N_7789,N_7855);
xnor U11387 (N_11387,N_9291,N_9755);
xor U11388 (N_11388,N_8601,N_8392);
and U11389 (N_11389,N_8553,N_9884);
nor U11390 (N_11390,N_7529,N_9873);
xor U11391 (N_11391,N_9274,N_9053);
or U11392 (N_11392,N_8135,N_7836);
xor U11393 (N_11393,N_9467,N_9303);
nand U11394 (N_11394,N_8498,N_8851);
or U11395 (N_11395,N_8235,N_8253);
xor U11396 (N_11396,N_8067,N_8288);
or U11397 (N_11397,N_8174,N_9673);
and U11398 (N_11398,N_9833,N_9717);
xnor U11399 (N_11399,N_9416,N_8030);
xnor U11400 (N_11400,N_9256,N_8480);
or U11401 (N_11401,N_9728,N_7720);
nor U11402 (N_11402,N_8733,N_8224);
or U11403 (N_11403,N_9815,N_7692);
and U11404 (N_11404,N_9326,N_7761);
or U11405 (N_11405,N_8220,N_7837);
nor U11406 (N_11406,N_9361,N_9660);
and U11407 (N_11407,N_7724,N_9692);
xor U11408 (N_11408,N_7777,N_7562);
xor U11409 (N_11409,N_8793,N_9317);
nor U11410 (N_11410,N_8848,N_9969);
nand U11411 (N_11411,N_8569,N_9388);
or U11412 (N_11412,N_7880,N_8527);
xnor U11413 (N_11413,N_9890,N_9376);
xor U11414 (N_11414,N_9524,N_8699);
nand U11415 (N_11415,N_7670,N_8236);
nor U11416 (N_11416,N_8454,N_7879);
nand U11417 (N_11417,N_8039,N_9719);
or U11418 (N_11418,N_8115,N_7871);
nand U11419 (N_11419,N_9412,N_7556);
or U11420 (N_11420,N_8814,N_8287);
xor U11421 (N_11421,N_9307,N_8552);
xnor U11422 (N_11422,N_9679,N_8483);
or U11423 (N_11423,N_8312,N_9908);
and U11424 (N_11424,N_8125,N_7612);
or U11425 (N_11425,N_7747,N_7741);
nand U11426 (N_11426,N_7936,N_8981);
nand U11427 (N_11427,N_9197,N_9365);
and U11428 (N_11428,N_7673,N_9743);
nor U11429 (N_11429,N_9398,N_7951);
nand U11430 (N_11430,N_7686,N_8434);
xor U11431 (N_11431,N_8763,N_7623);
or U11432 (N_11432,N_8331,N_8378);
nand U11433 (N_11433,N_9667,N_9763);
and U11434 (N_11434,N_7647,N_8354);
nor U11435 (N_11435,N_8773,N_9429);
and U11436 (N_11436,N_8380,N_9987);
nor U11437 (N_11437,N_9006,N_9784);
and U11438 (N_11438,N_8481,N_9936);
and U11439 (N_11439,N_8893,N_8757);
xnor U11440 (N_11440,N_9229,N_7714);
nor U11441 (N_11441,N_7607,N_8429);
xnor U11442 (N_11442,N_7606,N_8589);
xnor U11443 (N_11443,N_8756,N_8941);
nor U11444 (N_11444,N_7529,N_7713);
nand U11445 (N_11445,N_9188,N_8773);
or U11446 (N_11446,N_9011,N_9454);
nor U11447 (N_11447,N_7699,N_8091);
nor U11448 (N_11448,N_8973,N_9860);
or U11449 (N_11449,N_8247,N_7830);
nand U11450 (N_11450,N_7805,N_8086);
nand U11451 (N_11451,N_7932,N_8963);
and U11452 (N_11452,N_8294,N_8652);
nor U11453 (N_11453,N_8068,N_9711);
and U11454 (N_11454,N_8834,N_7867);
nand U11455 (N_11455,N_9889,N_9585);
nand U11456 (N_11456,N_8673,N_7743);
and U11457 (N_11457,N_7912,N_8710);
nand U11458 (N_11458,N_9015,N_9882);
or U11459 (N_11459,N_8301,N_8304);
nand U11460 (N_11460,N_9952,N_8508);
nand U11461 (N_11461,N_7655,N_8021);
or U11462 (N_11462,N_9410,N_9452);
and U11463 (N_11463,N_9733,N_8672);
nand U11464 (N_11464,N_7741,N_8437);
or U11465 (N_11465,N_8447,N_8967);
and U11466 (N_11466,N_8811,N_9961);
nor U11467 (N_11467,N_8316,N_9884);
nor U11468 (N_11468,N_8942,N_9635);
nand U11469 (N_11469,N_8543,N_7725);
nor U11470 (N_11470,N_9958,N_9496);
nand U11471 (N_11471,N_7919,N_9193);
or U11472 (N_11472,N_7889,N_8940);
xnor U11473 (N_11473,N_8156,N_7614);
nor U11474 (N_11474,N_7621,N_8763);
nand U11475 (N_11475,N_9588,N_9431);
nor U11476 (N_11476,N_7627,N_9549);
nand U11477 (N_11477,N_9007,N_8321);
and U11478 (N_11478,N_8231,N_7943);
and U11479 (N_11479,N_9388,N_9804);
xor U11480 (N_11480,N_8535,N_8214);
xor U11481 (N_11481,N_9028,N_8394);
nor U11482 (N_11482,N_7959,N_7960);
nor U11483 (N_11483,N_7873,N_9646);
xnor U11484 (N_11484,N_8548,N_8059);
nor U11485 (N_11485,N_9841,N_9853);
or U11486 (N_11486,N_9819,N_7501);
xnor U11487 (N_11487,N_9502,N_9138);
xnor U11488 (N_11488,N_9331,N_7907);
or U11489 (N_11489,N_9560,N_8901);
xnor U11490 (N_11490,N_8844,N_8700);
nor U11491 (N_11491,N_8155,N_9057);
nand U11492 (N_11492,N_7790,N_8604);
nor U11493 (N_11493,N_9461,N_7764);
xnor U11494 (N_11494,N_9999,N_9722);
xnor U11495 (N_11495,N_9551,N_9164);
xor U11496 (N_11496,N_7635,N_8966);
nand U11497 (N_11497,N_8279,N_9813);
and U11498 (N_11498,N_7547,N_9658);
and U11499 (N_11499,N_8378,N_9341);
nand U11500 (N_11500,N_9151,N_9050);
xor U11501 (N_11501,N_8312,N_8506);
nand U11502 (N_11502,N_9947,N_7619);
nor U11503 (N_11503,N_8284,N_9154);
or U11504 (N_11504,N_7522,N_9294);
or U11505 (N_11505,N_7599,N_8812);
xor U11506 (N_11506,N_9784,N_9255);
nor U11507 (N_11507,N_9932,N_8719);
or U11508 (N_11508,N_7718,N_9667);
nor U11509 (N_11509,N_8058,N_9555);
xor U11510 (N_11510,N_9405,N_8294);
and U11511 (N_11511,N_8062,N_8264);
and U11512 (N_11512,N_8779,N_9367);
nand U11513 (N_11513,N_7729,N_8263);
xnor U11514 (N_11514,N_7998,N_9902);
and U11515 (N_11515,N_8384,N_8235);
and U11516 (N_11516,N_8085,N_9671);
nor U11517 (N_11517,N_7543,N_9686);
xnor U11518 (N_11518,N_8310,N_9520);
and U11519 (N_11519,N_9239,N_9156);
xor U11520 (N_11520,N_7592,N_8056);
and U11521 (N_11521,N_9237,N_8780);
xnor U11522 (N_11522,N_7910,N_8011);
or U11523 (N_11523,N_9291,N_8193);
xor U11524 (N_11524,N_9674,N_9380);
and U11525 (N_11525,N_9312,N_7650);
nor U11526 (N_11526,N_8674,N_9680);
xor U11527 (N_11527,N_7567,N_9408);
xor U11528 (N_11528,N_8974,N_8945);
nand U11529 (N_11529,N_8396,N_8082);
or U11530 (N_11530,N_9786,N_8307);
or U11531 (N_11531,N_9115,N_7860);
nor U11532 (N_11532,N_8962,N_8334);
and U11533 (N_11533,N_9029,N_9008);
and U11534 (N_11534,N_9885,N_8812);
xor U11535 (N_11535,N_8270,N_9639);
nand U11536 (N_11536,N_9158,N_7788);
or U11537 (N_11537,N_8963,N_9364);
nand U11538 (N_11538,N_9811,N_7720);
and U11539 (N_11539,N_8113,N_9793);
and U11540 (N_11540,N_8562,N_8645);
and U11541 (N_11541,N_9652,N_7601);
nor U11542 (N_11542,N_9482,N_9664);
and U11543 (N_11543,N_9034,N_9504);
xor U11544 (N_11544,N_7872,N_8267);
xnor U11545 (N_11545,N_8697,N_8264);
and U11546 (N_11546,N_8046,N_9832);
or U11547 (N_11547,N_8867,N_8648);
nand U11548 (N_11548,N_8325,N_8712);
nor U11549 (N_11549,N_9648,N_8383);
nor U11550 (N_11550,N_8096,N_9359);
xnor U11551 (N_11551,N_8288,N_9872);
and U11552 (N_11552,N_9378,N_7653);
xor U11553 (N_11553,N_9475,N_7885);
xnor U11554 (N_11554,N_7616,N_9866);
and U11555 (N_11555,N_9189,N_8018);
nor U11556 (N_11556,N_9218,N_8020);
nand U11557 (N_11557,N_9682,N_8023);
nand U11558 (N_11558,N_9735,N_9189);
and U11559 (N_11559,N_9856,N_7873);
nor U11560 (N_11560,N_8253,N_7978);
nor U11561 (N_11561,N_8107,N_8233);
or U11562 (N_11562,N_9129,N_9561);
nor U11563 (N_11563,N_8194,N_7903);
and U11564 (N_11564,N_9049,N_7827);
nor U11565 (N_11565,N_8241,N_8918);
and U11566 (N_11566,N_9075,N_8419);
nor U11567 (N_11567,N_8164,N_8332);
nand U11568 (N_11568,N_9274,N_9817);
xor U11569 (N_11569,N_9213,N_7828);
xnor U11570 (N_11570,N_9255,N_8413);
xnor U11571 (N_11571,N_9841,N_8155);
nand U11572 (N_11572,N_7528,N_8858);
nor U11573 (N_11573,N_9250,N_9563);
nor U11574 (N_11574,N_9611,N_9208);
or U11575 (N_11575,N_7762,N_8982);
and U11576 (N_11576,N_9670,N_9000);
nand U11577 (N_11577,N_7882,N_9178);
xor U11578 (N_11578,N_8525,N_8676);
xnor U11579 (N_11579,N_8244,N_8128);
nor U11580 (N_11580,N_8366,N_9883);
xnor U11581 (N_11581,N_7999,N_8851);
xor U11582 (N_11582,N_8804,N_9209);
nand U11583 (N_11583,N_8973,N_9757);
xor U11584 (N_11584,N_8505,N_9378);
nand U11585 (N_11585,N_7781,N_7500);
nand U11586 (N_11586,N_8347,N_9446);
nand U11587 (N_11587,N_9345,N_9084);
or U11588 (N_11588,N_8765,N_9402);
nand U11589 (N_11589,N_9766,N_7972);
nor U11590 (N_11590,N_7934,N_8392);
and U11591 (N_11591,N_8443,N_9312);
nand U11592 (N_11592,N_8482,N_8659);
xor U11593 (N_11593,N_9999,N_8421);
nand U11594 (N_11594,N_9677,N_9929);
or U11595 (N_11595,N_8709,N_8018);
nor U11596 (N_11596,N_8463,N_9448);
nand U11597 (N_11597,N_7725,N_9044);
nor U11598 (N_11598,N_9962,N_8829);
or U11599 (N_11599,N_9108,N_8627);
nor U11600 (N_11600,N_7527,N_9787);
or U11601 (N_11601,N_9682,N_9300);
xnor U11602 (N_11602,N_9756,N_8441);
or U11603 (N_11603,N_9773,N_9752);
nand U11604 (N_11604,N_9349,N_7817);
and U11605 (N_11605,N_8560,N_9723);
nand U11606 (N_11606,N_8504,N_9936);
and U11607 (N_11607,N_8335,N_9735);
nand U11608 (N_11608,N_8369,N_7696);
nor U11609 (N_11609,N_8358,N_7813);
nor U11610 (N_11610,N_8553,N_9054);
xnor U11611 (N_11611,N_7750,N_9524);
xor U11612 (N_11612,N_9259,N_9823);
and U11613 (N_11613,N_8462,N_8314);
xnor U11614 (N_11614,N_9874,N_9779);
or U11615 (N_11615,N_9966,N_7886);
nand U11616 (N_11616,N_9366,N_7593);
nor U11617 (N_11617,N_8127,N_9939);
and U11618 (N_11618,N_9432,N_9813);
xnor U11619 (N_11619,N_9541,N_8796);
xor U11620 (N_11620,N_9823,N_9917);
xor U11621 (N_11621,N_9482,N_8112);
nor U11622 (N_11622,N_9758,N_9721);
nand U11623 (N_11623,N_8183,N_8283);
xnor U11624 (N_11624,N_9730,N_9611);
nand U11625 (N_11625,N_9143,N_8343);
or U11626 (N_11626,N_9632,N_9305);
nor U11627 (N_11627,N_9550,N_8902);
xnor U11628 (N_11628,N_9532,N_9887);
nand U11629 (N_11629,N_7705,N_9687);
nor U11630 (N_11630,N_9844,N_9184);
and U11631 (N_11631,N_9231,N_7975);
or U11632 (N_11632,N_9396,N_7906);
and U11633 (N_11633,N_8831,N_8397);
and U11634 (N_11634,N_7511,N_9070);
nor U11635 (N_11635,N_7865,N_8400);
nor U11636 (N_11636,N_9835,N_8105);
nand U11637 (N_11637,N_7604,N_8296);
xor U11638 (N_11638,N_8926,N_8575);
or U11639 (N_11639,N_8072,N_9998);
or U11640 (N_11640,N_7639,N_8362);
or U11641 (N_11641,N_7884,N_9850);
or U11642 (N_11642,N_9803,N_8247);
and U11643 (N_11643,N_7716,N_9781);
nand U11644 (N_11644,N_9605,N_8389);
nor U11645 (N_11645,N_8409,N_9573);
xnor U11646 (N_11646,N_7524,N_9087);
xnor U11647 (N_11647,N_7723,N_8521);
xor U11648 (N_11648,N_7954,N_9927);
nand U11649 (N_11649,N_7855,N_9124);
and U11650 (N_11650,N_9564,N_8259);
and U11651 (N_11651,N_8206,N_7713);
or U11652 (N_11652,N_8260,N_7795);
xnor U11653 (N_11653,N_8229,N_9824);
nand U11654 (N_11654,N_9272,N_9369);
or U11655 (N_11655,N_9619,N_9894);
xor U11656 (N_11656,N_9460,N_9837);
xor U11657 (N_11657,N_7600,N_8498);
xor U11658 (N_11658,N_8051,N_9499);
and U11659 (N_11659,N_8719,N_8977);
nor U11660 (N_11660,N_9312,N_7865);
and U11661 (N_11661,N_9240,N_7889);
and U11662 (N_11662,N_8137,N_9892);
nor U11663 (N_11663,N_8028,N_7817);
or U11664 (N_11664,N_9257,N_8126);
or U11665 (N_11665,N_9605,N_8605);
nor U11666 (N_11666,N_8983,N_7839);
nand U11667 (N_11667,N_8391,N_9560);
xor U11668 (N_11668,N_8335,N_9116);
nor U11669 (N_11669,N_9914,N_7502);
nand U11670 (N_11670,N_9628,N_9701);
nor U11671 (N_11671,N_8020,N_9358);
nor U11672 (N_11672,N_9757,N_7515);
nor U11673 (N_11673,N_9387,N_8540);
and U11674 (N_11674,N_7715,N_8542);
nor U11675 (N_11675,N_8444,N_7895);
nor U11676 (N_11676,N_9134,N_9737);
and U11677 (N_11677,N_8191,N_8867);
xor U11678 (N_11678,N_9581,N_7824);
nor U11679 (N_11679,N_9040,N_9411);
nand U11680 (N_11680,N_8725,N_8495);
or U11681 (N_11681,N_8995,N_7728);
and U11682 (N_11682,N_8077,N_9210);
or U11683 (N_11683,N_9884,N_8122);
nand U11684 (N_11684,N_7789,N_7614);
nand U11685 (N_11685,N_9732,N_9143);
or U11686 (N_11686,N_8312,N_9988);
and U11687 (N_11687,N_9825,N_8613);
nor U11688 (N_11688,N_8400,N_8850);
nor U11689 (N_11689,N_9856,N_8145);
xor U11690 (N_11690,N_8196,N_7825);
nor U11691 (N_11691,N_7660,N_8143);
and U11692 (N_11692,N_8784,N_9169);
nor U11693 (N_11693,N_9700,N_8363);
xor U11694 (N_11694,N_7620,N_8939);
or U11695 (N_11695,N_8812,N_9895);
or U11696 (N_11696,N_8193,N_8741);
or U11697 (N_11697,N_7646,N_8974);
and U11698 (N_11698,N_8454,N_7605);
nor U11699 (N_11699,N_9300,N_9375);
nor U11700 (N_11700,N_7699,N_8329);
and U11701 (N_11701,N_9659,N_8604);
nor U11702 (N_11702,N_9716,N_9888);
nor U11703 (N_11703,N_9971,N_9710);
nand U11704 (N_11704,N_9551,N_8003);
or U11705 (N_11705,N_9105,N_9925);
nor U11706 (N_11706,N_9898,N_8329);
nor U11707 (N_11707,N_9644,N_7544);
xor U11708 (N_11708,N_9922,N_7865);
or U11709 (N_11709,N_8349,N_9982);
nand U11710 (N_11710,N_9415,N_9031);
and U11711 (N_11711,N_9131,N_9115);
or U11712 (N_11712,N_7829,N_9512);
or U11713 (N_11713,N_9291,N_7501);
or U11714 (N_11714,N_8007,N_8612);
and U11715 (N_11715,N_8783,N_8994);
or U11716 (N_11716,N_8116,N_9519);
xnor U11717 (N_11717,N_8044,N_8633);
or U11718 (N_11718,N_8906,N_8937);
nor U11719 (N_11719,N_8783,N_7555);
nand U11720 (N_11720,N_7974,N_8212);
and U11721 (N_11721,N_9668,N_8705);
or U11722 (N_11722,N_8376,N_8168);
nand U11723 (N_11723,N_9462,N_7904);
or U11724 (N_11724,N_7707,N_8753);
or U11725 (N_11725,N_9846,N_8125);
xor U11726 (N_11726,N_9789,N_9961);
or U11727 (N_11727,N_7563,N_8498);
xor U11728 (N_11728,N_8370,N_9657);
or U11729 (N_11729,N_9073,N_9072);
xnor U11730 (N_11730,N_8688,N_8327);
nor U11731 (N_11731,N_8605,N_9187);
nand U11732 (N_11732,N_7903,N_9765);
xnor U11733 (N_11733,N_8861,N_9397);
and U11734 (N_11734,N_9772,N_9562);
and U11735 (N_11735,N_9789,N_7653);
and U11736 (N_11736,N_8561,N_9298);
or U11737 (N_11737,N_9673,N_7693);
or U11738 (N_11738,N_9082,N_8103);
and U11739 (N_11739,N_8449,N_7651);
or U11740 (N_11740,N_7845,N_7545);
nand U11741 (N_11741,N_8614,N_8210);
or U11742 (N_11742,N_9044,N_9527);
or U11743 (N_11743,N_8141,N_8292);
nand U11744 (N_11744,N_8722,N_9686);
nand U11745 (N_11745,N_8214,N_8926);
and U11746 (N_11746,N_8847,N_9474);
or U11747 (N_11747,N_7512,N_7700);
or U11748 (N_11748,N_7969,N_8548);
xor U11749 (N_11749,N_7737,N_8293);
and U11750 (N_11750,N_8147,N_8907);
xnor U11751 (N_11751,N_9393,N_8919);
nand U11752 (N_11752,N_8087,N_9637);
or U11753 (N_11753,N_8045,N_9894);
or U11754 (N_11754,N_8198,N_8990);
nand U11755 (N_11755,N_9787,N_9509);
xnor U11756 (N_11756,N_8352,N_8537);
xor U11757 (N_11757,N_8161,N_9714);
and U11758 (N_11758,N_7823,N_9306);
xor U11759 (N_11759,N_8319,N_9696);
nor U11760 (N_11760,N_7796,N_9713);
and U11761 (N_11761,N_9303,N_8013);
and U11762 (N_11762,N_8124,N_8477);
and U11763 (N_11763,N_8296,N_7915);
nor U11764 (N_11764,N_9932,N_9811);
nand U11765 (N_11765,N_8638,N_8840);
nor U11766 (N_11766,N_8178,N_9430);
xor U11767 (N_11767,N_7811,N_8551);
nand U11768 (N_11768,N_8508,N_8330);
nand U11769 (N_11769,N_9408,N_9303);
nand U11770 (N_11770,N_9687,N_8596);
nor U11771 (N_11771,N_9362,N_9935);
and U11772 (N_11772,N_8266,N_8987);
and U11773 (N_11773,N_8099,N_9581);
or U11774 (N_11774,N_9882,N_7534);
or U11775 (N_11775,N_9938,N_8950);
xnor U11776 (N_11776,N_8937,N_7946);
nand U11777 (N_11777,N_8284,N_9198);
xnor U11778 (N_11778,N_9419,N_8263);
nor U11779 (N_11779,N_7549,N_8703);
nand U11780 (N_11780,N_8459,N_8629);
nor U11781 (N_11781,N_8003,N_7942);
or U11782 (N_11782,N_9945,N_9444);
nor U11783 (N_11783,N_9886,N_8322);
or U11784 (N_11784,N_9967,N_8201);
or U11785 (N_11785,N_8644,N_8188);
or U11786 (N_11786,N_9800,N_9683);
and U11787 (N_11787,N_9449,N_8740);
or U11788 (N_11788,N_8993,N_7796);
xor U11789 (N_11789,N_8639,N_7924);
and U11790 (N_11790,N_9613,N_9853);
nand U11791 (N_11791,N_8334,N_9425);
nand U11792 (N_11792,N_9519,N_9688);
or U11793 (N_11793,N_7786,N_9790);
nand U11794 (N_11794,N_8455,N_9196);
and U11795 (N_11795,N_9087,N_9438);
and U11796 (N_11796,N_8669,N_9728);
nor U11797 (N_11797,N_7700,N_8784);
or U11798 (N_11798,N_8482,N_9200);
or U11799 (N_11799,N_7608,N_8774);
nor U11800 (N_11800,N_8963,N_8716);
and U11801 (N_11801,N_7768,N_9184);
xnor U11802 (N_11802,N_9100,N_9764);
xnor U11803 (N_11803,N_8053,N_7836);
and U11804 (N_11804,N_9542,N_9184);
xnor U11805 (N_11805,N_8484,N_7512);
xor U11806 (N_11806,N_8308,N_9251);
nor U11807 (N_11807,N_7610,N_8416);
xnor U11808 (N_11808,N_7918,N_8359);
or U11809 (N_11809,N_9860,N_9571);
or U11810 (N_11810,N_9258,N_7893);
and U11811 (N_11811,N_9294,N_8913);
nor U11812 (N_11812,N_8840,N_8523);
and U11813 (N_11813,N_8874,N_9566);
or U11814 (N_11814,N_8778,N_8924);
nor U11815 (N_11815,N_8542,N_9533);
nor U11816 (N_11816,N_7650,N_8975);
nor U11817 (N_11817,N_9150,N_7683);
and U11818 (N_11818,N_8744,N_9261);
nor U11819 (N_11819,N_7596,N_8306);
nor U11820 (N_11820,N_9226,N_9081);
nor U11821 (N_11821,N_9796,N_7544);
and U11822 (N_11822,N_8634,N_8491);
and U11823 (N_11823,N_8452,N_8649);
or U11824 (N_11824,N_9316,N_8019);
nand U11825 (N_11825,N_8503,N_8515);
nand U11826 (N_11826,N_7821,N_8767);
nor U11827 (N_11827,N_7788,N_9866);
and U11828 (N_11828,N_9828,N_9990);
nand U11829 (N_11829,N_9693,N_9450);
or U11830 (N_11830,N_8729,N_8457);
or U11831 (N_11831,N_8344,N_9543);
xnor U11832 (N_11832,N_8196,N_8962);
and U11833 (N_11833,N_8977,N_9237);
or U11834 (N_11834,N_9405,N_8124);
nor U11835 (N_11835,N_9949,N_9974);
nand U11836 (N_11836,N_9988,N_8204);
and U11837 (N_11837,N_9425,N_9948);
nor U11838 (N_11838,N_7889,N_9511);
or U11839 (N_11839,N_9043,N_9931);
nor U11840 (N_11840,N_9264,N_7936);
nor U11841 (N_11841,N_9167,N_7675);
and U11842 (N_11842,N_7690,N_9583);
or U11843 (N_11843,N_8490,N_9983);
nand U11844 (N_11844,N_9374,N_8995);
or U11845 (N_11845,N_8161,N_8747);
nor U11846 (N_11846,N_9472,N_8900);
nor U11847 (N_11847,N_8077,N_8730);
xor U11848 (N_11848,N_7918,N_7569);
and U11849 (N_11849,N_8233,N_9143);
nor U11850 (N_11850,N_7641,N_7984);
nand U11851 (N_11851,N_8625,N_7794);
nand U11852 (N_11852,N_9647,N_7885);
nand U11853 (N_11853,N_8513,N_8130);
or U11854 (N_11854,N_9385,N_8331);
nand U11855 (N_11855,N_7666,N_8155);
nor U11856 (N_11856,N_9433,N_7831);
and U11857 (N_11857,N_7987,N_7533);
nand U11858 (N_11858,N_7506,N_7972);
and U11859 (N_11859,N_9241,N_8904);
or U11860 (N_11860,N_8513,N_7581);
or U11861 (N_11861,N_9191,N_8604);
and U11862 (N_11862,N_9654,N_8246);
and U11863 (N_11863,N_8993,N_8333);
nor U11864 (N_11864,N_9830,N_9911);
or U11865 (N_11865,N_8715,N_8197);
nor U11866 (N_11866,N_9528,N_7987);
xnor U11867 (N_11867,N_9161,N_9030);
and U11868 (N_11868,N_7563,N_9186);
xor U11869 (N_11869,N_8829,N_7763);
or U11870 (N_11870,N_9119,N_8664);
nor U11871 (N_11871,N_9841,N_9479);
and U11872 (N_11872,N_7691,N_7578);
nand U11873 (N_11873,N_8966,N_9185);
or U11874 (N_11874,N_8762,N_9558);
nand U11875 (N_11875,N_9468,N_7559);
nand U11876 (N_11876,N_7923,N_7665);
and U11877 (N_11877,N_9373,N_8027);
nand U11878 (N_11878,N_9338,N_8627);
and U11879 (N_11879,N_8669,N_7880);
and U11880 (N_11880,N_9712,N_9954);
xor U11881 (N_11881,N_9443,N_9033);
and U11882 (N_11882,N_8120,N_8129);
nand U11883 (N_11883,N_8175,N_8832);
and U11884 (N_11884,N_7622,N_9853);
xor U11885 (N_11885,N_9051,N_9201);
or U11886 (N_11886,N_7889,N_7899);
nor U11887 (N_11887,N_8360,N_9276);
xor U11888 (N_11888,N_9683,N_8949);
or U11889 (N_11889,N_8764,N_8863);
or U11890 (N_11890,N_8165,N_9122);
and U11891 (N_11891,N_8675,N_9395);
and U11892 (N_11892,N_9618,N_9751);
nor U11893 (N_11893,N_7973,N_8892);
nor U11894 (N_11894,N_9854,N_8889);
nand U11895 (N_11895,N_9805,N_9621);
or U11896 (N_11896,N_8540,N_8067);
xnor U11897 (N_11897,N_9490,N_9730);
xnor U11898 (N_11898,N_9707,N_9574);
xnor U11899 (N_11899,N_9876,N_8044);
and U11900 (N_11900,N_8865,N_9197);
or U11901 (N_11901,N_9356,N_9152);
and U11902 (N_11902,N_7647,N_9329);
or U11903 (N_11903,N_9396,N_7912);
or U11904 (N_11904,N_9060,N_9704);
xnor U11905 (N_11905,N_8222,N_8274);
or U11906 (N_11906,N_7878,N_7865);
nand U11907 (N_11907,N_7689,N_7562);
nor U11908 (N_11908,N_9877,N_7739);
nand U11909 (N_11909,N_7940,N_8183);
nand U11910 (N_11910,N_8342,N_9608);
nor U11911 (N_11911,N_9551,N_7618);
nor U11912 (N_11912,N_9460,N_7964);
nand U11913 (N_11913,N_9774,N_9846);
xnor U11914 (N_11914,N_8539,N_8713);
and U11915 (N_11915,N_8402,N_9933);
xnor U11916 (N_11916,N_7578,N_7721);
nand U11917 (N_11917,N_9779,N_9889);
xnor U11918 (N_11918,N_8443,N_9923);
nor U11919 (N_11919,N_8007,N_8199);
nand U11920 (N_11920,N_7965,N_9314);
xnor U11921 (N_11921,N_8098,N_8596);
nor U11922 (N_11922,N_8472,N_9169);
nor U11923 (N_11923,N_9259,N_7875);
and U11924 (N_11924,N_9853,N_9013);
and U11925 (N_11925,N_7533,N_8711);
nor U11926 (N_11926,N_8318,N_8018);
nand U11927 (N_11927,N_9739,N_7712);
nor U11928 (N_11928,N_7958,N_8111);
and U11929 (N_11929,N_8294,N_8772);
nor U11930 (N_11930,N_8857,N_9768);
or U11931 (N_11931,N_8075,N_9811);
xor U11932 (N_11932,N_9898,N_8856);
xor U11933 (N_11933,N_8203,N_8451);
and U11934 (N_11934,N_8572,N_7552);
nor U11935 (N_11935,N_7607,N_9412);
nor U11936 (N_11936,N_9935,N_7776);
nor U11937 (N_11937,N_8356,N_9151);
xor U11938 (N_11938,N_8791,N_9924);
and U11939 (N_11939,N_8975,N_7963);
and U11940 (N_11940,N_8327,N_8964);
nand U11941 (N_11941,N_7664,N_9391);
xnor U11942 (N_11942,N_9570,N_9066);
nand U11943 (N_11943,N_9461,N_8028);
nor U11944 (N_11944,N_7794,N_8220);
and U11945 (N_11945,N_9373,N_7511);
or U11946 (N_11946,N_7898,N_9028);
or U11947 (N_11947,N_9095,N_9818);
nand U11948 (N_11948,N_7952,N_9314);
xor U11949 (N_11949,N_8755,N_7988);
or U11950 (N_11950,N_9718,N_7846);
nand U11951 (N_11951,N_8530,N_9511);
nor U11952 (N_11952,N_7675,N_8710);
or U11953 (N_11953,N_9891,N_9000);
nand U11954 (N_11954,N_9413,N_9241);
nor U11955 (N_11955,N_8737,N_8061);
xnor U11956 (N_11956,N_8673,N_8788);
nor U11957 (N_11957,N_9125,N_9406);
xor U11958 (N_11958,N_8930,N_9861);
or U11959 (N_11959,N_9950,N_8780);
nor U11960 (N_11960,N_8308,N_8964);
xor U11961 (N_11961,N_8861,N_9298);
nor U11962 (N_11962,N_9548,N_8321);
and U11963 (N_11963,N_7579,N_9333);
xor U11964 (N_11964,N_9617,N_8962);
nand U11965 (N_11965,N_7672,N_9520);
or U11966 (N_11966,N_9014,N_9632);
and U11967 (N_11967,N_8741,N_7771);
nand U11968 (N_11968,N_9016,N_9081);
and U11969 (N_11969,N_8253,N_9369);
and U11970 (N_11970,N_8140,N_9077);
nand U11971 (N_11971,N_8686,N_8716);
and U11972 (N_11972,N_7979,N_9261);
nor U11973 (N_11973,N_8453,N_9281);
nand U11974 (N_11974,N_9420,N_7970);
nor U11975 (N_11975,N_8486,N_8229);
and U11976 (N_11976,N_9896,N_9413);
xnor U11977 (N_11977,N_9918,N_9099);
nand U11978 (N_11978,N_9017,N_7692);
nor U11979 (N_11979,N_8868,N_9768);
or U11980 (N_11980,N_8438,N_8504);
nor U11981 (N_11981,N_9856,N_9280);
and U11982 (N_11982,N_9851,N_8399);
xor U11983 (N_11983,N_9511,N_7778);
and U11984 (N_11984,N_9141,N_9240);
nor U11985 (N_11985,N_8860,N_9992);
nand U11986 (N_11986,N_9414,N_8090);
nand U11987 (N_11987,N_8700,N_9832);
or U11988 (N_11988,N_9106,N_8065);
nand U11989 (N_11989,N_8622,N_9947);
and U11990 (N_11990,N_9524,N_9161);
nand U11991 (N_11991,N_7865,N_8863);
or U11992 (N_11992,N_8781,N_8951);
nor U11993 (N_11993,N_8734,N_9933);
and U11994 (N_11994,N_7547,N_9596);
nand U11995 (N_11995,N_7582,N_9062);
nand U11996 (N_11996,N_9054,N_9446);
or U11997 (N_11997,N_8446,N_7518);
and U11998 (N_11998,N_8929,N_9833);
and U11999 (N_11999,N_8506,N_7889);
nand U12000 (N_12000,N_8808,N_7882);
nor U12001 (N_12001,N_9277,N_8957);
nand U12002 (N_12002,N_8827,N_9241);
xnor U12003 (N_12003,N_8359,N_7596);
and U12004 (N_12004,N_9009,N_7759);
nand U12005 (N_12005,N_8602,N_9777);
nor U12006 (N_12006,N_8610,N_9783);
or U12007 (N_12007,N_7631,N_9041);
and U12008 (N_12008,N_9878,N_9072);
and U12009 (N_12009,N_9827,N_9805);
and U12010 (N_12010,N_9288,N_8757);
xnor U12011 (N_12011,N_8726,N_8810);
xor U12012 (N_12012,N_9056,N_8564);
nand U12013 (N_12013,N_9881,N_8535);
or U12014 (N_12014,N_8745,N_8102);
or U12015 (N_12015,N_8013,N_9908);
xnor U12016 (N_12016,N_7617,N_8661);
or U12017 (N_12017,N_7515,N_8397);
nor U12018 (N_12018,N_8964,N_7659);
nor U12019 (N_12019,N_9572,N_9716);
nor U12020 (N_12020,N_9934,N_9358);
xnor U12021 (N_12021,N_8453,N_8868);
nand U12022 (N_12022,N_8457,N_8295);
and U12023 (N_12023,N_9865,N_9248);
xor U12024 (N_12024,N_8505,N_9769);
nor U12025 (N_12025,N_7815,N_7945);
nand U12026 (N_12026,N_7832,N_8699);
and U12027 (N_12027,N_8712,N_7998);
or U12028 (N_12028,N_8811,N_8630);
nor U12029 (N_12029,N_8726,N_8020);
nand U12030 (N_12030,N_8412,N_9693);
nor U12031 (N_12031,N_9430,N_8156);
xor U12032 (N_12032,N_9161,N_8667);
or U12033 (N_12033,N_8251,N_7698);
or U12034 (N_12034,N_8424,N_8671);
xor U12035 (N_12035,N_8764,N_7663);
or U12036 (N_12036,N_9722,N_8508);
and U12037 (N_12037,N_9661,N_8037);
nor U12038 (N_12038,N_8045,N_7522);
nor U12039 (N_12039,N_8518,N_8519);
and U12040 (N_12040,N_9775,N_8883);
nor U12041 (N_12041,N_8549,N_9868);
nor U12042 (N_12042,N_7785,N_9365);
xor U12043 (N_12043,N_7811,N_8175);
or U12044 (N_12044,N_9586,N_7579);
nor U12045 (N_12045,N_9942,N_8749);
nand U12046 (N_12046,N_8744,N_8500);
nor U12047 (N_12047,N_9884,N_8882);
nor U12048 (N_12048,N_9256,N_7593);
nand U12049 (N_12049,N_9114,N_9276);
or U12050 (N_12050,N_8889,N_8240);
nand U12051 (N_12051,N_9456,N_9397);
xnor U12052 (N_12052,N_8977,N_7649);
xor U12053 (N_12053,N_8519,N_8284);
or U12054 (N_12054,N_8958,N_7509);
nand U12055 (N_12055,N_8655,N_8665);
or U12056 (N_12056,N_9064,N_8661);
xor U12057 (N_12057,N_9037,N_8104);
and U12058 (N_12058,N_7569,N_8469);
or U12059 (N_12059,N_9261,N_8593);
nor U12060 (N_12060,N_8828,N_8246);
or U12061 (N_12061,N_7706,N_7511);
or U12062 (N_12062,N_8236,N_7773);
or U12063 (N_12063,N_9660,N_9916);
nor U12064 (N_12064,N_8241,N_8984);
or U12065 (N_12065,N_8244,N_8394);
and U12066 (N_12066,N_9068,N_8063);
or U12067 (N_12067,N_7556,N_7585);
nor U12068 (N_12068,N_9443,N_8823);
xor U12069 (N_12069,N_8453,N_7566);
xnor U12070 (N_12070,N_7671,N_7807);
and U12071 (N_12071,N_7943,N_9408);
and U12072 (N_12072,N_8768,N_9778);
or U12073 (N_12073,N_9375,N_9892);
or U12074 (N_12074,N_7706,N_8991);
and U12075 (N_12075,N_8770,N_8036);
or U12076 (N_12076,N_8544,N_9877);
xor U12077 (N_12077,N_9737,N_9662);
xor U12078 (N_12078,N_9634,N_9317);
or U12079 (N_12079,N_8615,N_9242);
xor U12080 (N_12080,N_9058,N_8428);
nand U12081 (N_12081,N_7962,N_9198);
and U12082 (N_12082,N_8661,N_9079);
and U12083 (N_12083,N_7798,N_9698);
or U12084 (N_12084,N_9515,N_9629);
xor U12085 (N_12085,N_8575,N_9655);
xor U12086 (N_12086,N_9424,N_8852);
xor U12087 (N_12087,N_9520,N_7735);
xnor U12088 (N_12088,N_9504,N_9253);
or U12089 (N_12089,N_8081,N_8901);
nor U12090 (N_12090,N_7987,N_9162);
nand U12091 (N_12091,N_9934,N_9687);
nand U12092 (N_12092,N_8848,N_9070);
nor U12093 (N_12093,N_7558,N_8605);
xnor U12094 (N_12094,N_9630,N_8056);
and U12095 (N_12095,N_8671,N_8704);
nor U12096 (N_12096,N_8388,N_9473);
or U12097 (N_12097,N_9419,N_7625);
and U12098 (N_12098,N_7812,N_8238);
and U12099 (N_12099,N_9026,N_9617);
and U12100 (N_12100,N_8231,N_9285);
xor U12101 (N_12101,N_7738,N_8864);
nand U12102 (N_12102,N_8848,N_9826);
or U12103 (N_12103,N_9638,N_8164);
or U12104 (N_12104,N_8175,N_9296);
and U12105 (N_12105,N_7767,N_8161);
nor U12106 (N_12106,N_8214,N_8956);
and U12107 (N_12107,N_9926,N_8093);
nor U12108 (N_12108,N_9318,N_8135);
nand U12109 (N_12109,N_8821,N_7982);
nor U12110 (N_12110,N_8558,N_8100);
nor U12111 (N_12111,N_8096,N_8015);
or U12112 (N_12112,N_7664,N_9626);
nand U12113 (N_12113,N_8311,N_8020);
nand U12114 (N_12114,N_8943,N_9597);
xnor U12115 (N_12115,N_9521,N_8553);
nor U12116 (N_12116,N_8766,N_7557);
xnor U12117 (N_12117,N_8246,N_9076);
and U12118 (N_12118,N_9832,N_7997);
nor U12119 (N_12119,N_9921,N_9528);
and U12120 (N_12120,N_8917,N_8257);
nor U12121 (N_12121,N_8453,N_9179);
xor U12122 (N_12122,N_9122,N_7595);
or U12123 (N_12123,N_9685,N_9624);
nor U12124 (N_12124,N_8243,N_9772);
xor U12125 (N_12125,N_8808,N_9676);
nor U12126 (N_12126,N_9859,N_9069);
nor U12127 (N_12127,N_7579,N_7750);
nor U12128 (N_12128,N_8789,N_9672);
and U12129 (N_12129,N_9454,N_7847);
nor U12130 (N_12130,N_8869,N_9172);
nor U12131 (N_12131,N_8163,N_8078);
nor U12132 (N_12132,N_9716,N_9072);
or U12133 (N_12133,N_7931,N_8796);
nand U12134 (N_12134,N_7614,N_9705);
and U12135 (N_12135,N_8919,N_8516);
xor U12136 (N_12136,N_9186,N_8461);
and U12137 (N_12137,N_9969,N_8196);
and U12138 (N_12138,N_9569,N_9773);
nor U12139 (N_12139,N_7650,N_8077);
and U12140 (N_12140,N_8408,N_9453);
nor U12141 (N_12141,N_9642,N_8188);
or U12142 (N_12142,N_8859,N_9700);
nor U12143 (N_12143,N_7994,N_8692);
nand U12144 (N_12144,N_9784,N_9350);
nand U12145 (N_12145,N_8459,N_8718);
or U12146 (N_12146,N_7980,N_7990);
xor U12147 (N_12147,N_9736,N_8692);
xnor U12148 (N_12148,N_7934,N_7708);
nand U12149 (N_12149,N_7641,N_7543);
and U12150 (N_12150,N_8766,N_9294);
or U12151 (N_12151,N_9141,N_9400);
xnor U12152 (N_12152,N_8820,N_8428);
nor U12153 (N_12153,N_8365,N_8175);
xor U12154 (N_12154,N_7575,N_9393);
or U12155 (N_12155,N_8889,N_9219);
and U12156 (N_12156,N_8505,N_7830);
and U12157 (N_12157,N_8635,N_8334);
nor U12158 (N_12158,N_8619,N_8423);
or U12159 (N_12159,N_7782,N_9670);
nor U12160 (N_12160,N_9050,N_9377);
and U12161 (N_12161,N_9180,N_8729);
or U12162 (N_12162,N_7815,N_9784);
and U12163 (N_12163,N_9677,N_8776);
and U12164 (N_12164,N_9594,N_7767);
xor U12165 (N_12165,N_7858,N_8573);
xor U12166 (N_12166,N_9159,N_8880);
nor U12167 (N_12167,N_9137,N_7500);
xor U12168 (N_12168,N_8924,N_8705);
nor U12169 (N_12169,N_8982,N_8859);
nand U12170 (N_12170,N_8473,N_9880);
nand U12171 (N_12171,N_8983,N_9997);
xnor U12172 (N_12172,N_9462,N_8021);
or U12173 (N_12173,N_9492,N_9853);
nand U12174 (N_12174,N_8092,N_8122);
nand U12175 (N_12175,N_9372,N_8758);
or U12176 (N_12176,N_9013,N_8687);
or U12177 (N_12177,N_8666,N_9065);
or U12178 (N_12178,N_8620,N_8959);
nand U12179 (N_12179,N_9910,N_8466);
or U12180 (N_12180,N_8386,N_8426);
and U12181 (N_12181,N_7730,N_8867);
xnor U12182 (N_12182,N_8891,N_9573);
nand U12183 (N_12183,N_9879,N_9070);
and U12184 (N_12184,N_9233,N_8661);
or U12185 (N_12185,N_8020,N_8727);
xor U12186 (N_12186,N_7571,N_9343);
or U12187 (N_12187,N_7963,N_8752);
nor U12188 (N_12188,N_8795,N_8100);
or U12189 (N_12189,N_9721,N_8937);
nand U12190 (N_12190,N_8837,N_9914);
or U12191 (N_12191,N_7810,N_9355);
nand U12192 (N_12192,N_9049,N_8891);
or U12193 (N_12193,N_9534,N_8808);
nor U12194 (N_12194,N_8483,N_8941);
nor U12195 (N_12195,N_7622,N_9715);
or U12196 (N_12196,N_8593,N_8916);
nor U12197 (N_12197,N_9652,N_8173);
nand U12198 (N_12198,N_8910,N_7649);
nand U12199 (N_12199,N_8472,N_8747);
xor U12200 (N_12200,N_8507,N_7985);
xnor U12201 (N_12201,N_9110,N_8507);
and U12202 (N_12202,N_8015,N_8855);
nand U12203 (N_12203,N_9717,N_7667);
or U12204 (N_12204,N_9907,N_8156);
or U12205 (N_12205,N_7610,N_9159);
xnor U12206 (N_12206,N_8345,N_8713);
and U12207 (N_12207,N_8776,N_8853);
and U12208 (N_12208,N_9843,N_9054);
nand U12209 (N_12209,N_9064,N_9224);
and U12210 (N_12210,N_7654,N_7998);
nand U12211 (N_12211,N_7804,N_8505);
and U12212 (N_12212,N_7815,N_9415);
nand U12213 (N_12213,N_7658,N_9242);
nor U12214 (N_12214,N_7934,N_8015);
nand U12215 (N_12215,N_7558,N_8255);
xnor U12216 (N_12216,N_9262,N_9352);
nand U12217 (N_12217,N_7770,N_9909);
and U12218 (N_12218,N_8582,N_8649);
nand U12219 (N_12219,N_9559,N_9662);
or U12220 (N_12220,N_7578,N_9667);
xnor U12221 (N_12221,N_9142,N_8967);
and U12222 (N_12222,N_8891,N_8471);
or U12223 (N_12223,N_8978,N_8670);
and U12224 (N_12224,N_8858,N_7903);
nand U12225 (N_12225,N_8319,N_9245);
and U12226 (N_12226,N_9394,N_7570);
or U12227 (N_12227,N_9920,N_8730);
nand U12228 (N_12228,N_8568,N_9778);
and U12229 (N_12229,N_9177,N_8086);
xnor U12230 (N_12230,N_9522,N_9905);
xor U12231 (N_12231,N_8917,N_9553);
nand U12232 (N_12232,N_7614,N_7940);
nand U12233 (N_12233,N_8962,N_8036);
or U12234 (N_12234,N_9222,N_8127);
and U12235 (N_12235,N_8097,N_9009);
nor U12236 (N_12236,N_9616,N_8332);
nor U12237 (N_12237,N_9874,N_8381);
nand U12238 (N_12238,N_9619,N_8696);
and U12239 (N_12239,N_9127,N_8481);
or U12240 (N_12240,N_8822,N_8419);
nand U12241 (N_12241,N_9862,N_8078);
or U12242 (N_12242,N_8303,N_8887);
or U12243 (N_12243,N_8219,N_7748);
or U12244 (N_12244,N_8226,N_7631);
nand U12245 (N_12245,N_8964,N_9070);
nand U12246 (N_12246,N_9834,N_7689);
and U12247 (N_12247,N_8349,N_9960);
xor U12248 (N_12248,N_7982,N_8472);
xnor U12249 (N_12249,N_9604,N_8978);
nor U12250 (N_12250,N_9451,N_7726);
nor U12251 (N_12251,N_9151,N_9842);
or U12252 (N_12252,N_8975,N_7975);
or U12253 (N_12253,N_8772,N_9963);
nand U12254 (N_12254,N_9304,N_7953);
or U12255 (N_12255,N_7718,N_8328);
xnor U12256 (N_12256,N_9625,N_9218);
xnor U12257 (N_12257,N_7994,N_7526);
nand U12258 (N_12258,N_9484,N_8046);
and U12259 (N_12259,N_7678,N_8811);
nand U12260 (N_12260,N_8981,N_8765);
nor U12261 (N_12261,N_9551,N_8071);
or U12262 (N_12262,N_8347,N_9059);
xor U12263 (N_12263,N_9054,N_9857);
xor U12264 (N_12264,N_9228,N_8491);
or U12265 (N_12265,N_9851,N_8355);
or U12266 (N_12266,N_8526,N_9509);
nor U12267 (N_12267,N_8772,N_7706);
and U12268 (N_12268,N_8447,N_9141);
xor U12269 (N_12269,N_7999,N_9267);
or U12270 (N_12270,N_9394,N_8893);
nor U12271 (N_12271,N_9608,N_7899);
nor U12272 (N_12272,N_9249,N_7786);
nand U12273 (N_12273,N_8286,N_7966);
nand U12274 (N_12274,N_8286,N_8936);
and U12275 (N_12275,N_9433,N_7677);
nor U12276 (N_12276,N_8854,N_7804);
and U12277 (N_12277,N_9547,N_9084);
and U12278 (N_12278,N_7597,N_9227);
nor U12279 (N_12279,N_8938,N_8349);
and U12280 (N_12280,N_8016,N_7687);
and U12281 (N_12281,N_8317,N_8041);
nand U12282 (N_12282,N_7976,N_8560);
or U12283 (N_12283,N_8866,N_7617);
or U12284 (N_12284,N_7548,N_7541);
xor U12285 (N_12285,N_9954,N_9614);
nor U12286 (N_12286,N_8797,N_9409);
xnor U12287 (N_12287,N_7639,N_9098);
and U12288 (N_12288,N_9829,N_9576);
nand U12289 (N_12289,N_8325,N_8043);
or U12290 (N_12290,N_8215,N_7880);
nor U12291 (N_12291,N_8635,N_7560);
nand U12292 (N_12292,N_9121,N_9252);
xnor U12293 (N_12293,N_7698,N_8997);
nand U12294 (N_12294,N_8379,N_8955);
nor U12295 (N_12295,N_8731,N_8381);
or U12296 (N_12296,N_9735,N_8378);
and U12297 (N_12297,N_9555,N_9050);
and U12298 (N_12298,N_7622,N_8558);
or U12299 (N_12299,N_9842,N_9945);
and U12300 (N_12300,N_7803,N_9491);
nand U12301 (N_12301,N_7704,N_9592);
or U12302 (N_12302,N_8636,N_9636);
nand U12303 (N_12303,N_8532,N_8671);
nor U12304 (N_12304,N_9580,N_7988);
or U12305 (N_12305,N_9323,N_8241);
or U12306 (N_12306,N_9495,N_8168);
and U12307 (N_12307,N_7917,N_7846);
nor U12308 (N_12308,N_7592,N_9703);
xor U12309 (N_12309,N_8121,N_8506);
xnor U12310 (N_12310,N_9745,N_8445);
or U12311 (N_12311,N_8334,N_9364);
nor U12312 (N_12312,N_9486,N_8183);
or U12313 (N_12313,N_9670,N_9427);
or U12314 (N_12314,N_8276,N_9244);
xnor U12315 (N_12315,N_9208,N_7954);
or U12316 (N_12316,N_8935,N_8976);
and U12317 (N_12317,N_8500,N_8980);
and U12318 (N_12318,N_9242,N_7626);
and U12319 (N_12319,N_9660,N_9169);
or U12320 (N_12320,N_9522,N_8798);
xor U12321 (N_12321,N_8719,N_7999);
and U12322 (N_12322,N_8148,N_8746);
and U12323 (N_12323,N_8768,N_9744);
or U12324 (N_12324,N_7959,N_9843);
nor U12325 (N_12325,N_8497,N_8852);
nor U12326 (N_12326,N_9778,N_8006);
or U12327 (N_12327,N_8201,N_8819);
xnor U12328 (N_12328,N_8844,N_9845);
nand U12329 (N_12329,N_7548,N_7544);
and U12330 (N_12330,N_8869,N_8358);
and U12331 (N_12331,N_7751,N_9161);
xor U12332 (N_12332,N_8162,N_7640);
or U12333 (N_12333,N_7603,N_9053);
nand U12334 (N_12334,N_8990,N_8308);
nand U12335 (N_12335,N_8449,N_9453);
and U12336 (N_12336,N_7647,N_9867);
nor U12337 (N_12337,N_8815,N_8276);
and U12338 (N_12338,N_7795,N_8000);
or U12339 (N_12339,N_7689,N_9959);
and U12340 (N_12340,N_9560,N_8861);
and U12341 (N_12341,N_9248,N_9672);
nand U12342 (N_12342,N_9079,N_9894);
xnor U12343 (N_12343,N_8733,N_7582);
xor U12344 (N_12344,N_8340,N_7846);
or U12345 (N_12345,N_9124,N_8394);
xor U12346 (N_12346,N_7622,N_9731);
and U12347 (N_12347,N_8557,N_7655);
or U12348 (N_12348,N_9683,N_8955);
nor U12349 (N_12349,N_8454,N_7551);
or U12350 (N_12350,N_9922,N_8921);
xnor U12351 (N_12351,N_9667,N_9901);
nor U12352 (N_12352,N_7932,N_9076);
xor U12353 (N_12353,N_7536,N_9433);
nor U12354 (N_12354,N_7565,N_8399);
xor U12355 (N_12355,N_8148,N_9788);
or U12356 (N_12356,N_8230,N_8722);
or U12357 (N_12357,N_7853,N_9800);
and U12358 (N_12358,N_9805,N_8683);
and U12359 (N_12359,N_9058,N_8591);
and U12360 (N_12360,N_8656,N_8416);
nor U12361 (N_12361,N_9832,N_8018);
and U12362 (N_12362,N_8108,N_7834);
xnor U12363 (N_12363,N_7713,N_8411);
or U12364 (N_12364,N_9136,N_9515);
nor U12365 (N_12365,N_9268,N_8826);
nand U12366 (N_12366,N_8950,N_9866);
nand U12367 (N_12367,N_8259,N_8150);
or U12368 (N_12368,N_9785,N_7970);
xor U12369 (N_12369,N_8339,N_8748);
and U12370 (N_12370,N_9301,N_9797);
nor U12371 (N_12371,N_7522,N_7621);
nand U12372 (N_12372,N_7882,N_8225);
or U12373 (N_12373,N_8847,N_9630);
and U12374 (N_12374,N_9038,N_9293);
and U12375 (N_12375,N_9727,N_8190);
xor U12376 (N_12376,N_7889,N_8858);
xnor U12377 (N_12377,N_9778,N_7638);
nand U12378 (N_12378,N_9314,N_7724);
xnor U12379 (N_12379,N_8355,N_8761);
xnor U12380 (N_12380,N_8439,N_7606);
nand U12381 (N_12381,N_9927,N_8652);
nand U12382 (N_12382,N_9629,N_7512);
xor U12383 (N_12383,N_7997,N_9803);
or U12384 (N_12384,N_9975,N_8085);
and U12385 (N_12385,N_9974,N_7822);
xnor U12386 (N_12386,N_8628,N_8844);
and U12387 (N_12387,N_8248,N_9230);
or U12388 (N_12388,N_9514,N_9492);
and U12389 (N_12389,N_7810,N_7564);
xor U12390 (N_12390,N_7551,N_7594);
and U12391 (N_12391,N_9789,N_8460);
or U12392 (N_12392,N_8097,N_7658);
or U12393 (N_12393,N_9979,N_9453);
nor U12394 (N_12394,N_7857,N_9280);
and U12395 (N_12395,N_9693,N_8529);
or U12396 (N_12396,N_9593,N_9952);
nor U12397 (N_12397,N_8654,N_9733);
or U12398 (N_12398,N_8102,N_8958);
nand U12399 (N_12399,N_8192,N_8315);
nand U12400 (N_12400,N_8409,N_9452);
nand U12401 (N_12401,N_8335,N_9740);
and U12402 (N_12402,N_7694,N_8634);
nor U12403 (N_12403,N_9388,N_8605);
xor U12404 (N_12404,N_9731,N_7682);
nand U12405 (N_12405,N_9313,N_7703);
or U12406 (N_12406,N_9225,N_9659);
nand U12407 (N_12407,N_7639,N_9113);
and U12408 (N_12408,N_8365,N_9986);
or U12409 (N_12409,N_9741,N_7950);
nor U12410 (N_12410,N_8403,N_7764);
xnor U12411 (N_12411,N_8973,N_7501);
nand U12412 (N_12412,N_7946,N_9305);
nand U12413 (N_12413,N_7712,N_9870);
xnor U12414 (N_12414,N_9221,N_9655);
and U12415 (N_12415,N_9367,N_9492);
and U12416 (N_12416,N_7960,N_7629);
nand U12417 (N_12417,N_7614,N_8528);
nand U12418 (N_12418,N_7565,N_9845);
or U12419 (N_12419,N_9542,N_8947);
nand U12420 (N_12420,N_8555,N_9854);
xnor U12421 (N_12421,N_9571,N_9993);
nor U12422 (N_12422,N_9125,N_7652);
nand U12423 (N_12423,N_7661,N_7582);
nand U12424 (N_12424,N_8167,N_7928);
nand U12425 (N_12425,N_8500,N_8724);
xor U12426 (N_12426,N_7739,N_8847);
and U12427 (N_12427,N_8455,N_8405);
or U12428 (N_12428,N_9591,N_8465);
or U12429 (N_12429,N_7923,N_7852);
xor U12430 (N_12430,N_9533,N_9212);
nor U12431 (N_12431,N_8807,N_9343);
nand U12432 (N_12432,N_8887,N_8270);
xor U12433 (N_12433,N_9750,N_9130);
or U12434 (N_12434,N_7825,N_7542);
and U12435 (N_12435,N_8796,N_8780);
and U12436 (N_12436,N_9685,N_9840);
or U12437 (N_12437,N_8473,N_9158);
or U12438 (N_12438,N_8499,N_9787);
nand U12439 (N_12439,N_9041,N_8324);
nor U12440 (N_12440,N_7762,N_8530);
xor U12441 (N_12441,N_9152,N_7566);
nor U12442 (N_12442,N_8222,N_8929);
nor U12443 (N_12443,N_9830,N_9276);
nor U12444 (N_12444,N_8300,N_8789);
or U12445 (N_12445,N_8059,N_7593);
and U12446 (N_12446,N_8219,N_8628);
and U12447 (N_12447,N_7589,N_9663);
nand U12448 (N_12448,N_9934,N_9824);
nand U12449 (N_12449,N_8609,N_9946);
nand U12450 (N_12450,N_9781,N_9731);
nand U12451 (N_12451,N_8083,N_7689);
xnor U12452 (N_12452,N_7734,N_8840);
xor U12453 (N_12453,N_9992,N_7620);
nand U12454 (N_12454,N_9918,N_9874);
nor U12455 (N_12455,N_8448,N_7855);
nand U12456 (N_12456,N_8648,N_9021);
or U12457 (N_12457,N_9886,N_9497);
or U12458 (N_12458,N_8008,N_8258);
nor U12459 (N_12459,N_7560,N_8257);
and U12460 (N_12460,N_9294,N_9573);
or U12461 (N_12461,N_7879,N_9604);
xor U12462 (N_12462,N_9772,N_8342);
or U12463 (N_12463,N_8276,N_9045);
xnor U12464 (N_12464,N_8005,N_8019);
nand U12465 (N_12465,N_7731,N_8803);
nand U12466 (N_12466,N_8812,N_8792);
xor U12467 (N_12467,N_9153,N_8429);
xnor U12468 (N_12468,N_7896,N_9796);
xnor U12469 (N_12469,N_8756,N_8603);
nor U12470 (N_12470,N_8885,N_8098);
xnor U12471 (N_12471,N_8187,N_9785);
and U12472 (N_12472,N_8543,N_9105);
and U12473 (N_12473,N_8197,N_9275);
xnor U12474 (N_12474,N_7592,N_9533);
xnor U12475 (N_12475,N_8812,N_9615);
or U12476 (N_12476,N_9162,N_7925);
or U12477 (N_12477,N_8268,N_9715);
and U12478 (N_12478,N_8898,N_8571);
xnor U12479 (N_12479,N_8154,N_8409);
or U12480 (N_12480,N_9355,N_9717);
nand U12481 (N_12481,N_9504,N_8564);
and U12482 (N_12482,N_9618,N_7524);
and U12483 (N_12483,N_7960,N_7648);
nand U12484 (N_12484,N_7629,N_8012);
nand U12485 (N_12485,N_9421,N_9070);
nor U12486 (N_12486,N_9322,N_7971);
xnor U12487 (N_12487,N_9826,N_8092);
or U12488 (N_12488,N_9401,N_9322);
and U12489 (N_12489,N_8520,N_9523);
or U12490 (N_12490,N_8417,N_9455);
nand U12491 (N_12491,N_9942,N_7865);
nand U12492 (N_12492,N_8297,N_9884);
or U12493 (N_12493,N_8512,N_8814);
and U12494 (N_12494,N_9600,N_7886);
and U12495 (N_12495,N_8373,N_8831);
or U12496 (N_12496,N_7700,N_8499);
or U12497 (N_12497,N_8360,N_9425);
xnor U12498 (N_12498,N_7643,N_8210);
xor U12499 (N_12499,N_9028,N_8417);
xnor U12500 (N_12500,N_10274,N_10360);
nor U12501 (N_12501,N_10868,N_11224);
nor U12502 (N_12502,N_12044,N_11027);
xor U12503 (N_12503,N_10689,N_10064);
nand U12504 (N_12504,N_11421,N_11418);
nand U12505 (N_12505,N_11452,N_10690);
and U12506 (N_12506,N_12489,N_11200);
or U12507 (N_12507,N_10912,N_12485);
xnor U12508 (N_12508,N_10907,N_10219);
and U12509 (N_12509,N_11708,N_11087);
nand U12510 (N_12510,N_12120,N_10968);
nand U12511 (N_12511,N_11943,N_11619);
nor U12512 (N_12512,N_11600,N_10032);
xnor U12513 (N_12513,N_12170,N_10528);
or U12514 (N_12514,N_10386,N_11387);
xor U12515 (N_12515,N_10674,N_11383);
xnor U12516 (N_12516,N_12481,N_12220);
nor U12517 (N_12517,N_10910,N_11401);
nand U12518 (N_12518,N_10278,N_11522);
or U12519 (N_12519,N_10477,N_10415);
nand U12520 (N_12520,N_11426,N_12098);
and U12521 (N_12521,N_10444,N_11833);
and U12522 (N_12522,N_10359,N_11235);
nand U12523 (N_12523,N_11834,N_11288);
or U12524 (N_12524,N_12115,N_10916);
or U12525 (N_12525,N_12331,N_10704);
nor U12526 (N_12526,N_10580,N_10022);
nand U12527 (N_12527,N_11502,N_12209);
or U12528 (N_12528,N_10930,N_11237);
nand U12529 (N_12529,N_10093,N_11225);
nand U12530 (N_12530,N_11613,N_11503);
or U12531 (N_12531,N_10756,N_10697);
xnor U12532 (N_12532,N_12433,N_11272);
nand U12533 (N_12533,N_10098,N_12017);
xnor U12534 (N_12534,N_10561,N_11403);
or U12535 (N_12535,N_12211,N_11763);
nor U12536 (N_12536,N_10285,N_11591);
nor U12537 (N_12537,N_12392,N_11628);
xor U12538 (N_12538,N_10110,N_10221);
or U12539 (N_12539,N_11805,N_10152);
or U12540 (N_12540,N_10198,N_10836);
or U12541 (N_12541,N_12424,N_10288);
nand U12542 (N_12542,N_10725,N_11466);
and U12543 (N_12543,N_10914,N_11956);
xnor U12544 (N_12544,N_12068,N_10891);
or U12545 (N_12545,N_11411,N_11438);
nand U12546 (N_12546,N_11923,N_11340);
or U12547 (N_12547,N_12451,N_10331);
nor U12548 (N_12548,N_11663,N_10333);
nor U12549 (N_12549,N_12284,N_10672);
nor U12550 (N_12550,N_11084,N_11378);
nand U12551 (N_12551,N_10352,N_12383);
nand U12552 (N_12552,N_10925,N_10183);
nand U12553 (N_12553,N_12131,N_12029);
nand U12554 (N_12554,N_10945,N_11526);
or U12555 (N_12555,N_11456,N_10962);
nand U12556 (N_12556,N_10675,N_11262);
xor U12557 (N_12557,N_10727,N_11658);
and U12558 (N_12558,N_11268,N_11880);
nor U12559 (N_12559,N_11062,N_11020);
nand U12560 (N_12560,N_11915,N_10099);
nor U12561 (N_12561,N_12113,N_10133);
nor U12562 (N_12562,N_10519,N_11656);
or U12563 (N_12563,N_10170,N_12348);
xnor U12564 (N_12564,N_10542,N_10699);
or U12565 (N_12565,N_10624,N_11960);
xor U12566 (N_12566,N_11926,N_11415);
nand U12567 (N_12567,N_10403,N_11698);
xor U12568 (N_12568,N_10065,N_12292);
and U12569 (N_12569,N_10339,N_11890);
or U12570 (N_12570,N_10536,N_11207);
nor U12571 (N_12571,N_10223,N_10114);
nand U12572 (N_12572,N_10370,N_12180);
and U12573 (N_12573,N_12327,N_11443);
xnor U12574 (N_12574,N_10668,N_10490);
and U12575 (N_12575,N_12403,N_12206);
nand U12576 (N_12576,N_12215,N_10841);
nor U12577 (N_12577,N_11579,N_10751);
nand U12578 (N_12578,N_11813,N_10642);
nor U12579 (N_12579,N_11105,N_10545);
or U12580 (N_12580,N_12336,N_11530);
nand U12581 (N_12581,N_10900,N_10382);
nor U12582 (N_12582,N_12116,N_11718);
xnor U12583 (N_12583,N_10397,N_10984);
xnor U12584 (N_12584,N_10892,N_10760);
and U12585 (N_12585,N_10829,N_12085);
nor U12586 (N_12586,N_11148,N_11147);
nand U12587 (N_12587,N_12151,N_10436);
and U12588 (N_12588,N_12338,N_12373);
and U12589 (N_12589,N_10995,N_11390);
and U12590 (N_12590,N_12160,N_10908);
xnor U12591 (N_12591,N_11719,N_10940);
nand U12592 (N_12592,N_12013,N_10532);
xor U12593 (N_12593,N_10412,N_11817);
xnor U12594 (N_12594,N_10304,N_12107);
or U12595 (N_12595,N_10389,N_11664);
or U12596 (N_12596,N_10346,N_10050);
xor U12597 (N_12597,N_10119,N_11536);
nor U12598 (N_12598,N_10613,N_12465);
xor U12599 (N_12599,N_10802,N_11382);
nor U12600 (N_12600,N_10465,N_10427);
and U12601 (N_12601,N_11811,N_11531);
nand U12602 (N_12602,N_12357,N_11463);
nand U12603 (N_12603,N_12397,N_12100);
or U12604 (N_12604,N_11073,N_10696);
nand U12605 (N_12605,N_11238,N_12388);
nand U12606 (N_12606,N_12036,N_10160);
xor U12607 (N_12607,N_11815,N_10564);
xor U12608 (N_12608,N_10862,N_11611);
and U12609 (N_12609,N_11374,N_11747);
nand U12610 (N_12610,N_10002,N_10623);
nand U12611 (N_12611,N_12181,N_10101);
and U12612 (N_12612,N_10358,N_11824);
nand U12613 (N_12613,N_11046,N_12124);
nand U12614 (N_12614,N_12095,N_11540);
or U12615 (N_12615,N_11699,N_11353);
and U12616 (N_12616,N_11313,N_11596);
and U12617 (N_12617,N_12256,N_11341);
nor U12618 (N_12618,N_10373,N_12468);
and U12619 (N_12619,N_12239,N_10821);
xor U12620 (N_12620,N_10144,N_11895);
nand U12621 (N_12621,N_10020,N_10535);
nand U12622 (N_12622,N_12214,N_11850);
or U12623 (N_12623,N_11585,N_11686);
nand U12624 (N_12624,N_11129,N_11928);
or U12625 (N_12625,N_11060,N_10383);
or U12626 (N_12626,N_11731,N_11292);
nor U12627 (N_12627,N_12138,N_11840);
or U12628 (N_12628,N_11762,N_12409);
or U12629 (N_12629,N_10431,N_11480);
or U12630 (N_12630,N_11655,N_11196);
nand U12631 (N_12631,N_10733,N_10377);
nor U12632 (N_12632,N_11819,N_10941);
and U12633 (N_12633,N_12461,N_10424);
nand U12634 (N_12634,N_11888,N_11214);
or U12635 (N_12635,N_11727,N_10217);
and U12636 (N_12636,N_10454,N_10628);
xnor U12637 (N_12637,N_10812,N_10216);
xnor U12638 (N_12638,N_12079,N_11528);
or U12639 (N_12639,N_12266,N_11583);
nor U12640 (N_12640,N_12447,N_11462);
nor U12641 (N_12641,N_12456,N_12423);
xor U12642 (N_12642,N_11539,N_10834);
and U12643 (N_12643,N_11761,N_11575);
xnor U12644 (N_12644,N_11209,N_12498);
nand U12645 (N_12645,N_10316,N_12493);
nand U12646 (N_12646,N_11158,N_11465);
nor U12647 (N_12647,N_10630,N_11553);
nor U12648 (N_12648,N_11991,N_10512);
nor U12649 (N_12649,N_10635,N_12166);
nor U12650 (N_12650,N_12006,N_11038);
nor U12651 (N_12651,N_10385,N_11995);
nand U12652 (N_12652,N_10860,N_10882);
nor U12653 (N_12653,N_12484,N_10839);
nor U12654 (N_12654,N_12159,N_12222);
and U12655 (N_12655,N_10446,N_11851);
and U12656 (N_12656,N_11395,N_10023);
and U12657 (N_12657,N_11801,N_11001);
nor U12658 (N_12658,N_11793,N_11612);
nand U12659 (N_12659,N_11831,N_12398);
xor U12660 (N_12660,N_10788,N_11344);
xor U12661 (N_12661,N_10418,N_11832);
or U12662 (N_12662,N_10703,N_11461);
xor U12663 (N_12663,N_11634,N_11822);
or U12664 (N_12664,N_11681,N_11752);
or U12665 (N_12665,N_10572,N_10779);
and U12666 (N_12666,N_11270,N_11018);
xnor U12667 (N_12667,N_12261,N_12466);
nor U12668 (N_12668,N_11396,N_11644);
or U12669 (N_12669,N_10885,N_12470);
or U12670 (N_12670,N_12007,N_10737);
nor U12671 (N_12671,N_11798,N_11356);
nand U12672 (N_12672,N_10429,N_12272);
xor U12673 (N_12673,N_11343,N_10033);
or U12674 (N_12674,N_10665,N_10344);
or U12675 (N_12675,N_11232,N_11180);
or U12676 (N_12676,N_11803,N_10749);
nand U12677 (N_12677,N_11035,N_12232);
and U12678 (N_12678,N_10207,N_11970);
or U12679 (N_12679,N_10190,N_10939);
nand U12680 (N_12680,N_10103,N_11735);
nor U12681 (N_12681,N_12449,N_12428);
and U12682 (N_12682,N_11215,N_11513);
nor U12683 (N_12683,N_11052,N_11725);
xor U12684 (N_12684,N_10709,N_11173);
xnor U12685 (N_12685,N_10606,N_11988);
xor U12686 (N_12686,N_10565,N_11379);
or U12687 (N_12687,N_10075,N_11726);
xor U12688 (N_12688,N_12018,N_10148);
nand U12689 (N_12689,N_11629,N_11555);
and U12690 (N_12690,N_11687,N_12027);
and U12691 (N_12691,N_10247,N_11181);
and U12692 (N_12692,N_11568,N_10987);
and U12693 (N_12693,N_10809,N_10482);
nand U12694 (N_12694,N_10248,N_10125);
or U12695 (N_12695,N_11707,N_12390);
or U12696 (N_12696,N_11742,N_12434);
nand U12697 (N_12697,N_11593,N_10327);
and U12698 (N_12698,N_11077,N_11566);
nand U12699 (N_12699,N_11032,N_11512);
or U12700 (N_12700,N_10085,N_12250);
or U12701 (N_12701,N_11859,N_10250);
or U12702 (N_12702,N_12490,N_11041);
nor U12703 (N_12703,N_12235,N_11448);
nor U12704 (N_12704,N_12418,N_11716);
xnor U12705 (N_12705,N_10426,N_10899);
and U12706 (N_12706,N_12395,N_10234);
and U12707 (N_12707,N_12311,N_12453);
and U12708 (N_12708,N_11584,N_12060);
xor U12709 (N_12709,N_11508,N_10789);
or U12710 (N_12710,N_12426,N_10971);
and U12711 (N_12711,N_11008,N_10157);
nor U12712 (N_12712,N_10557,N_11095);
nand U12713 (N_12713,N_10341,N_11184);
nor U12714 (N_12714,N_11906,N_12057);
nand U12715 (N_12715,N_10781,N_11141);
xor U12716 (N_12716,N_11767,N_10854);
or U12717 (N_12717,N_11236,N_11240);
or U12718 (N_12718,N_11051,N_11867);
and U12719 (N_12719,N_10330,N_10244);
xor U12720 (N_12720,N_11352,N_12469);
and U12721 (N_12721,N_10662,N_11549);
nor U12722 (N_12722,N_10670,N_10633);
nand U12723 (N_12723,N_10437,N_10086);
nand U12724 (N_12724,N_10451,N_12431);
nor U12725 (N_12725,N_12023,N_11693);
or U12726 (N_12726,N_11674,N_11004);
and U12727 (N_12727,N_10182,N_11304);
or U12728 (N_12728,N_11932,N_12302);
nor U12729 (N_12729,N_12346,N_10209);
nor U12730 (N_12730,N_10222,N_11376);
or U12731 (N_12731,N_10993,N_11857);
or U12732 (N_12732,N_10793,N_10413);
or U12733 (N_12733,N_10156,N_10736);
nor U12734 (N_12734,N_12408,N_10745);
nand U12735 (N_12735,N_11063,N_12016);
nand U12736 (N_12736,N_10878,N_10752);
nand U12737 (N_12737,N_11080,N_10440);
nor U12738 (N_12738,N_11252,N_11517);
or U12739 (N_12739,N_12251,N_10608);
nor U12740 (N_12740,N_11564,N_11778);
xor U12741 (N_12741,N_11099,N_12003);
nand U12742 (N_12742,N_11162,N_10425);
nor U12743 (N_12743,N_11800,N_10100);
nor U12744 (N_12744,N_10473,N_12201);
xnor U12745 (N_12745,N_10634,N_10459);
and U12746 (N_12746,N_10599,N_12416);
nor U12747 (N_12747,N_12177,N_11921);
or U12748 (N_12748,N_12146,N_12330);
and U12749 (N_12749,N_11437,N_11524);
nor U12750 (N_12750,N_10422,N_10602);
xor U12751 (N_12751,N_12129,N_11188);
and U12752 (N_12752,N_11602,N_11739);
nand U12753 (N_12753,N_10231,N_11460);
and U12754 (N_12754,N_11828,N_10072);
nand U12755 (N_12755,N_12110,N_11706);
xor U12756 (N_12756,N_11552,N_12143);
or U12757 (N_12757,N_10291,N_12169);
and U12758 (N_12758,N_11160,N_11829);
nor U12759 (N_12759,N_10428,N_11122);
nand U12760 (N_12760,N_11820,N_11996);
nand U12761 (N_12761,N_11729,N_11975);
nor U12762 (N_12762,N_12178,N_10953);
and U12763 (N_12763,N_11050,N_10353);
nand U12764 (N_12764,N_10011,N_11082);
or U12765 (N_12765,N_10158,N_11042);
nand U12766 (N_12766,N_12460,N_11717);
or U12767 (N_12767,N_11254,N_10872);
or U12768 (N_12768,N_11696,N_11359);
nand U12769 (N_12769,N_10070,N_10457);
or U12770 (N_12770,N_10518,N_11590);
and U12771 (N_12771,N_11806,N_11483);
and U12772 (N_12772,N_10584,N_11759);
or U12773 (N_12773,N_11000,N_12478);
nor U12774 (N_12774,N_11302,N_12070);
and U12775 (N_12775,N_10325,N_11896);
or U12776 (N_12776,N_10343,N_10306);
or U12777 (N_12777,N_12422,N_10254);
nor U12778 (N_12778,N_11887,N_10006);
nor U12779 (N_12779,N_10111,N_12174);
nor U12780 (N_12780,N_10673,N_11825);
and U12781 (N_12781,N_10766,N_12358);
nor U12782 (N_12782,N_12226,N_12241);
nor U12783 (N_12783,N_11788,N_12375);
nor U12784 (N_12784,N_12074,N_11106);
nand U12785 (N_12785,N_10363,N_11659);
nand U12786 (N_12786,N_11457,N_10530);
xnor U12787 (N_12787,N_12237,N_10494);
nor U12788 (N_12788,N_11058,N_12233);
xor U12789 (N_12789,N_10671,N_11787);
and U12790 (N_12790,N_11711,N_12076);
or U12791 (N_12791,N_10263,N_10989);
and U12792 (N_12792,N_11569,N_10270);
and U12793 (N_12793,N_12114,N_10186);
nand U12794 (N_12794,N_11219,N_10113);
nor U12795 (N_12795,N_10267,N_10816);
nand U12796 (N_12796,N_12259,N_11627);
xor U12797 (N_12797,N_12406,N_10702);
nand U12798 (N_12798,N_11357,N_12312);
nand U12799 (N_12799,N_10558,N_11433);
nand U12800 (N_12800,N_10786,N_11349);
nand U12801 (N_12801,N_10400,N_10596);
nor U12802 (N_12802,N_11449,N_10901);
nand U12803 (N_12803,N_11835,N_10271);
nor U12804 (N_12804,N_10355,N_10488);
xor U12805 (N_12805,N_11734,N_11497);
or U12806 (N_12806,N_10852,N_10479);
nand U12807 (N_12807,N_10825,N_10563);
nand U12808 (N_12808,N_11957,N_11355);
nor U12809 (N_12809,N_12377,N_12260);
nand U12810 (N_12810,N_10265,N_11201);
and U12811 (N_12811,N_12126,N_11470);
xnor U12812 (N_12812,N_10594,N_11936);
xor U12813 (N_12813,N_11757,N_10879);
nor U12814 (N_12814,N_12366,N_11227);
or U12815 (N_12815,N_12341,N_10287);
xor U12816 (N_12816,N_11478,N_11998);
nor U12817 (N_12817,N_10835,N_10959);
nor U12818 (N_12818,N_10143,N_11958);
xnor U12819 (N_12819,N_12046,N_11535);
xnor U12820 (N_12820,N_11640,N_12372);
or U12821 (N_12821,N_10305,N_10047);
nor U12822 (N_12822,N_10129,N_11431);
nor U12823 (N_12823,N_11327,N_11258);
nor U12824 (N_12824,N_10362,N_12244);
and U12825 (N_12825,N_10475,N_10711);
xnor U12826 (N_12826,N_10094,N_10461);
nor U12827 (N_12827,N_11159,N_12202);
nand U12828 (N_12828,N_10754,N_10474);
nor U12829 (N_12829,N_10057,N_10338);
nor U12830 (N_12830,N_10522,N_11588);
nand U12831 (N_12831,N_10615,N_10458);
or U12832 (N_12832,N_10693,N_10650);
nand U12833 (N_12833,N_11559,N_10089);
xnor U12834 (N_12834,N_11940,N_11786);
and U12835 (N_12835,N_11984,N_11871);
xnor U12836 (N_12836,N_10128,N_10738);
xor U12837 (N_12837,N_11518,N_10447);
nand U12838 (N_12838,N_10975,N_12005);
nor U12839 (N_12839,N_10617,N_12118);
nand U12840 (N_12840,N_11864,N_12314);
and U12841 (N_12841,N_11618,N_11033);
or U12842 (N_12842,N_11978,N_10847);
nand U12843 (N_12843,N_11673,N_11900);
nor U12844 (N_12844,N_10205,N_12248);
nand U12845 (N_12845,N_11654,N_11295);
nor U12846 (N_12846,N_10357,N_12228);
xor U12847 (N_12847,N_10664,N_10501);
xnor U12848 (N_12848,N_10753,N_11405);
xor U12849 (N_12849,N_10813,N_11102);
and U12850 (N_12850,N_11467,N_10603);
and U12851 (N_12851,N_11135,N_11323);
nand U12852 (N_12852,N_10515,N_12389);
xor U12853 (N_12853,N_11837,N_11101);
nor U12854 (N_12854,N_11140,N_11675);
and U12855 (N_12855,N_11551,N_10846);
or U12856 (N_12856,N_11784,N_10493);
xor U12857 (N_12857,N_12323,N_11565);
or U12858 (N_12858,N_11691,N_10298);
or U12859 (N_12859,N_10108,N_10645);
nor U12860 (N_12860,N_11769,N_10356);
nor U12861 (N_12861,N_10589,N_10349);
nor U12862 (N_12862,N_10394,N_11679);
xnor U12863 (N_12863,N_11592,N_11257);
nand U12864 (N_12864,N_11486,N_12197);
and U12865 (N_12865,N_11648,N_12148);
xor U12866 (N_12866,N_12163,N_11743);
and U12867 (N_12867,N_10629,N_10188);
xnor U12868 (N_12868,N_11878,N_10611);
xor U12869 (N_12869,N_11218,N_12385);
and U12870 (N_12870,N_11324,N_11556);
xnor U12871 (N_12871,N_11119,N_10388);
or U12872 (N_12872,N_12452,N_11002);
xor U12873 (N_12873,N_11375,N_12391);
nand U12874 (N_12874,N_12119,N_11479);
and U12875 (N_12875,N_12263,N_10131);
or U12876 (N_12876,N_11208,N_12142);
nand U12877 (N_12877,N_12299,N_10658);
or U12878 (N_12878,N_12035,N_10233);
nand U12879 (N_12879,N_11416,N_11003);
and U12880 (N_12880,N_10230,N_11578);
nor U12881 (N_12881,N_11816,N_10007);
and U12882 (N_12882,N_11931,N_12155);
and U12883 (N_12883,N_12295,N_11741);
or U12884 (N_12884,N_11774,N_10199);
nor U12885 (N_12885,N_11315,N_10295);
nand U12886 (N_12886,N_12473,N_10000);
nor U12887 (N_12887,N_12328,N_11514);
and U12888 (N_12888,N_11715,N_10019);
nor U12889 (N_12889,N_10238,N_11336);
and U12890 (N_12890,N_10215,N_11910);
and U12891 (N_12891,N_11425,N_10317);
and U12892 (N_12892,N_10951,N_11891);
and U12893 (N_12893,N_11977,N_11746);
nand U12894 (N_12894,N_11190,N_10071);
xnor U12895 (N_12895,N_11969,N_11283);
xor U12896 (N_12896,N_10520,N_10124);
or U12897 (N_12897,N_11849,N_10965);
and U12898 (N_12898,N_11049,N_10652);
nor U12899 (N_12899,N_11519,N_11233);
or U12900 (N_12900,N_10053,N_12072);
nand U12901 (N_12901,N_10336,N_11814);
and U12902 (N_12902,N_11484,N_10112);
or U12903 (N_12903,N_11226,N_12450);
or U12904 (N_12904,N_10919,N_12363);
and U12905 (N_12905,N_11439,N_11862);
nand U12906 (N_12906,N_12313,N_11221);
and U12907 (N_12907,N_10942,N_11332);
and U12908 (N_12908,N_11557,N_10396);
nor U12909 (N_12909,N_10342,N_10442);
and U12910 (N_12910,N_12227,N_10008);
or U12911 (N_12911,N_12084,N_10136);
xnor U12912 (N_12912,N_12015,N_10243);
nor U12913 (N_12913,N_11948,N_11869);
xnor U12914 (N_12914,N_10078,N_11874);
and U12915 (N_12915,N_10402,N_10299);
xnor U12916 (N_12916,N_11916,N_10149);
nand U12917 (N_12917,N_10875,N_11770);
xnor U12918 (N_12918,N_10607,N_10682);
xor U12919 (N_12919,N_11019,N_12047);
and U12920 (N_12920,N_12264,N_10311);
nand U12921 (N_12921,N_11176,N_10393);
xor U12922 (N_12922,N_11964,N_10547);
or U12923 (N_12923,N_11368,N_12186);
nand U12924 (N_12924,N_11599,N_11532);
nor U12925 (N_12925,N_12188,N_10294);
nand U12926 (N_12926,N_10903,N_11229);
xor U12927 (N_12927,N_12185,N_10641);
xnor U12928 (N_12928,N_11143,N_12402);
xnor U12929 (N_12929,N_12002,N_10277);
nand U12930 (N_12930,N_11377,N_10768);
nand U12931 (N_12931,N_10313,N_11317);
xnor U12932 (N_12932,N_11400,N_11447);
or U12933 (N_12933,N_10573,N_12109);
xnor U12934 (N_12934,N_11281,N_12189);
xor U12935 (N_12935,N_11054,N_12171);
nor U12936 (N_12936,N_10102,N_11848);
xor U12937 (N_12937,N_10934,N_11444);
and U12938 (N_12938,N_11182,N_10997);
nor U12939 (N_12939,N_10978,N_11495);
or U12940 (N_12940,N_10782,N_11510);
nand U12941 (N_12941,N_11607,N_12200);
nand U12942 (N_12942,N_10368,N_11412);
or U12943 (N_12943,N_10687,N_10445);
nand U12944 (N_12944,N_11782,N_12464);
nand U12945 (N_12945,N_10977,N_12135);
or U12946 (N_12946,N_10419,N_10562);
nor U12947 (N_12947,N_11677,N_11130);
nand U12948 (N_12948,N_12471,N_10184);
or U12949 (N_12949,N_11284,N_11321);
and U12950 (N_12950,N_10139,N_10449);
or U12951 (N_12951,N_10241,N_10856);
or U12952 (N_12952,N_11212,N_11821);
or U12953 (N_12953,N_10175,N_12400);
nor U12954 (N_12954,N_12356,N_11308);
and U12955 (N_12955,N_10491,N_11464);
or U12956 (N_12956,N_12309,N_10492);
nor U12957 (N_12957,N_10224,N_10864);
nand U12958 (N_12958,N_12304,N_11955);
and U12959 (N_12959,N_11914,N_12307);
nor U12960 (N_12960,N_10721,N_10191);
and U12961 (N_12961,N_10843,N_11090);
and U12962 (N_12962,N_12288,N_11987);
or U12963 (N_12963,N_10472,N_11543);
and U12964 (N_12964,N_10016,N_11203);
nand U12965 (N_12965,N_11951,N_11429);
nor U12966 (N_12966,N_11328,N_10320);
and U12967 (N_12967,N_10038,N_12308);
xnor U12968 (N_12968,N_11633,N_10718);
or U12969 (N_12969,N_10496,N_12128);
nor U12970 (N_12970,N_10500,N_11785);
xor U12971 (N_12971,N_11710,N_10116);
nand U12972 (N_12972,N_11131,N_11604);
or U12973 (N_12973,N_12369,N_12194);
nor U12974 (N_12974,N_12103,N_11685);
nand U12975 (N_12975,N_11172,N_10544);
xor U12976 (N_12976,N_10130,N_12430);
or U12977 (N_12977,N_10297,N_10218);
nand U12978 (N_12978,N_10042,N_11239);
xnor U12979 (N_12979,N_10917,N_11736);
or U12980 (N_12980,N_10525,N_10783);
nand U12981 (N_12981,N_11015,N_11053);
and U12982 (N_12982,N_11608,N_10135);
and U12983 (N_12983,N_10163,N_11507);
or U12984 (N_12984,N_11198,N_10894);
and U12985 (N_12985,N_11312,N_12296);
xnor U12986 (N_12986,N_11610,N_10514);
nand U12987 (N_12987,N_11927,N_10443);
and U12988 (N_12988,N_12218,N_11337);
or U12989 (N_12989,N_10967,N_11234);
nor U12990 (N_12990,N_10329,N_12495);
or U12991 (N_12991,N_11504,N_10541);
nor U12992 (N_12992,N_11256,N_11597);
nor U12993 (N_12993,N_10722,N_10036);
xor U12994 (N_12994,N_11149,N_11653);
nand U12995 (N_12995,N_12083,N_12168);
and U12996 (N_12996,N_11802,N_11075);
xor U12997 (N_12997,N_12405,N_11723);
and U12998 (N_12998,N_11609,N_11515);
or U12999 (N_12999,N_11758,N_11365);
xor U13000 (N_13000,N_10761,N_12153);
or U13001 (N_13001,N_10734,N_11986);
and U13002 (N_13002,N_12184,N_12253);
and U13003 (N_13003,N_12410,N_10591);
and U13004 (N_13004,N_10531,N_10744);
xnor U13005 (N_13005,N_11812,N_10137);
or U13006 (N_13006,N_11213,N_12380);
xnor U13007 (N_13007,N_11886,N_11025);
xor U13008 (N_13008,N_11720,N_10235);
nand U13009 (N_13009,N_10414,N_10268);
xnor U13010 (N_13010,N_10080,N_11605);
xor U13011 (N_13011,N_11563,N_12243);
or U13012 (N_13012,N_10765,N_10374);
xor U13013 (N_13013,N_11547,N_10621);
or U13014 (N_13014,N_10076,N_10620);
or U13015 (N_13015,N_12443,N_11897);
xor U13016 (N_13016,N_11917,N_11827);
or U13017 (N_13017,N_10716,N_11039);
and U13018 (N_13018,N_10730,N_10166);
nand U13019 (N_13019,N_10932,N_10289);
nand U13020 (N_13020,N_11309,N_10555);
or U13021 (N_13021,N_11870,N_12090);
or U13022 (N_13022,N_12167,N_10326);
xnor U13023 (N_13023,N_10986,N_11351);
xnor U13024 (N_13024,N_12032,N_10147);
nand U13025 (N_13025,N_11210,N_11841);
or U13026 (N_13026,N_11126,N_12454);
nor U13027 (N_13027,N_11624,N_10253);
nand U13028 (N_13028,N_11363,N_12351);
xnor U13029 (N_13029,N_10487,N_10969);
and U13030 (N_13030,N_10605,N_12140);
xnor U13031 (N_13031,N_10947,N_10842);
and U13032 (N_13032,N_10588,N_11721);
nor U13033 (N_13033,N_12359,N_12091);
or U13034 (N_13034,N_11866,N_11133);
nor U13035 (N_13035,N_11189,N_10484);
xor U13036 (N_13036,N_10808,N_11169);
and U13037 (N_13037,N_10938,N_11523);
nor U13038 (N_13038,N_10804,N_10087);
nor U13039 (N_13039,N_12286,N_12279);
and U13040 (N_13040,N_10746,N_11354);
xor U13041 (N_13041,N_10398,N_10954);
nand U13042 (N_13042,N_11294,N_10666);
nor U13043 (N_13043,N_10778,N_10764);
and U13044 (N_13044,N_10340,N_10551);
or U13045 (N_13045,N_11930,N_11322);
or U13046 (N_13046,N_11282,N_10164);
nor U13047 (N_13047,N_10911,N_10031);
or U13048 (N_13048,N_10062,N_12082);
or U13049 (N_13049,N_11473,N_12097);
nor U13050 (N_13050,N_11586,N_12001);
nor U13051 (N_13051,N_10796,N_12472);
and U13052 (N_13052,N_12483,N_11279);
xnor U13053 (N_13053,N_10082,N_10961);
nand U13054 (N_13054,N_12413,N_12317);
nor U13055 (N_13055,N_11748,N_11333);
or U13056 (N_13056,N_10240,N_11098);
nor U13057 (N_13057,N_11124,N_10909);
xnor U13058 (N_13058,N_12127,N_11451);
nor U13059 (N_13059,N_11974,N_11253);
and U13060 (N_13060,N_11638,N_11952);
xor U13061 (N_13061,N_10194,N_12049);
nor U13062 (N_13062,N_10172,N_11070);
nand U13063 (N_13063,N_10044,N_10348);
xnor U13064 (N_13064,N_10873,N_11538);
xor U13065 (N_13065,N_11858,N_12217);
or U13066 (N_13066,N_10537,N_11083);
xor U13067 (N_13067,N_10467,N_11022);
and U13068 (N_13068,N_10228,N_11167);
and U13069 (N_13069,N_11132,N_10318);
nand U13070 (N_13070,N_10324,N_10210);
or U13071 (N_13071,N_10861,N_10345);
and U13072 (N_13072,N_12300,N_10534);
and U13073 (N_13073,N_11485,N_11847);
nand U13074 (N_13074,N_10884,N_12052);
xnor U13075 (N_13075,N_10970,N_11965);
and U13076 (N_13076,N_12139,N_10074);
nand U13077 (N_13077,N_11286,N_11211);
nor U13078 (N_13078,N_11005,N_10090);
nor U13079 (N_13079,N_12078,N_10701);
or U13080 (N_13080,N_10798,N_10260);
nand U13081 (N_13081,N_12306,N_11263);
xnor U13082 (N_13082,N_12077,N_11408);
and U13083 (N_13083,N_12234,N_10855);
nor U13084 (N_13084,N_10871,N_11902);
and U13085 (N_13085,N_10404,N_10740);
and U13086 (N_13086,N_11391,N_11245);
xor U13087 (N_13087,N_12303,N_12064);
nor U13088 (N_13088,N_12378,N_11668);
nor U13089 (N_13089,N_12051,N_10275);
xnor U13090 (N_13090,N_11064,N_12324);
and U13091 (N_13091,N_12316,N_10550);
and U13092 (N_13092,N_11280,N_12164);
xnor U13093 (N_13093,N_11966,N_10463);
or U13094 (N_13094,N_10375,N_11385);
and U13095 (N_13095,N_12394,N_11919);
and U13096 (N_13096,N_11667,N_10197);
xnor U13097 (N_13097,N_10631,N_12496);
and U13098 (N_13098,N_10416,N_10169);
nand U13099 (N_13099,N_11863,N_10805);
or U13100 (N_13100,N_10392,N_10632);
or U13101 (N_13101,N_11067,N_10845);
and U13102 (N_13102,N_11562,N_12474);
or U13103 (N_13103,N_10549,N_11392);
nand U13104 (N_13104,N_11487,N_12195);
and U13105 (N_13105,N_12179,N_11093);
nor U13106 (N_13106,N_10937,N_11220);
xnor U13107 (N_13107,N_11577,N_10933);
nand U13108 (N_13108,N_11950,N_11047);
nand U13109 (N_13109,N_10548,N_10239);
nor U13110 (N_13110,N_11259,N_11750);
xor U13111 (N_13111,N_10755,N_12354);
xnor U13112 (N_13112,N_10853,N_10800);
nor U13113 (N_13113,N_10213,N_10378);
nand U13114 (N_13114,N_12105,N_10647);
or U13115 (N_13115,N_11703,N_11029);
nand U13116 (N_13116,N_10141,N_10104);
nand U13117 (N_13117,N_11620,N_12048);
xor U13118 (N_13118,N_10742,N_10840);
and U13119 (N_13119,N_10739,N_11889);
nand U13120 (N_13120,N_10464,N_10012);
nor U13121 (N_13121,N_11048,N_10772);
nor U13122 (N_13122,N_12058,N_11990);
xor U13123 (N_13123,N_10117,N_10045);
nand U13124 (N_13124,N_12310,N_11981);
xnor U13125 (N_13125,N_11476,N_10923);
xor U13126 (N_13126,N_12355,N_11136);
nor U13127 (N_13127,N_11968,N_10068);
or U13128 (N_13128,N_12420,N_11657);
or U13129 (N_13129,N_10203,N_12026);
nor U13130 (N_13130,N_10988,N_11366);
nor U13131 (N_13131,N_11737,N_10708);
or U13132 (N_13132,N_12347,N_12238);
or U13133 (N_13133,N_11044,N_10059);
xnor U13134 (N_13134,N_11178,N_12287);
nand U13135 (N_13135,N_12277,N_12106);
or U13136 (N_13136,N_10717,N_11034);
nand U13137 (N_13137,N_12339,N_12183);
or U13138 (N_13138,N_11338,N_11676);
nand U13139 (N_13139,N_10120,N_10092);
and U13140 (N_13140,N_10035,N_10171);
or U13141 (N_13141,N_11231,N_10025);
and U13142 (N_13142,N_12122,N_10826);
nor U13143 (N_13143,N_11271,N_10657);
nand U13144 (N_13144,N_10180,N_12320);
nor U13145 (N_13145,N_11794,N_10096);
and U13146 (N_13146,N_12432,N_11490);
xnor U13147 (N_13147,N_10767,N_11548);
or U13148 (N_13148,N_12298,N_10540);
or U13149 (N_13149,N_11527,N_10161);
nor U13150 (N_13150,N_11846,N_12353);
nand U13151 (N_13151,N_12069,N_10552);
or U13152 (N_13152,N_12425,N_11339);
xor U13153 (N_13153,N_10817,N_10890);
nor U13154 (N_13154,N_10159,N_11300);
or U13155 (N_13155,N_10931,N_11855);
nor U13156 (N_13156,N_10983,N_10524);
or U13157 (N_13157,N_12137,N_11055);
xnor U13158 (N_13158,N_10401,N_11079);
xnor U13159 (N_13159,N_11617,N_10126);
and U13160 (N_13160,N_12089,N_10323);
xor U13161 (N_13161,N_11799,N_11645);
or U13162 (N_13162,N_10529,N_10134);
xnor U13163 (N_13163,N_12204,N_12219);
nand U13164 (N_13164,N_12192,N_11089);
xor U13165 (N_13165,N_10994,N_10801);
nor U13166 (N_13166,N_11740,N_12096);
or U13167 (N_13167,N_11195,N_12230);
and U13168 (N_13168,N_12290,N_10502);
nor U13169 (N_13169,N_12283,N_11768);
or U13170 (N_13170,N_11939,N_10799);
nor U13171 (N_13171,N_11689,N_11334);
nand U13172 (N_13172,N_10151,N_11838);
nor U13173 (N_13173,N_10819,N_11468);
or U13174 (N_13174,N_10677,N_10204);
nor U13175 (N_13175,N_12480,N_12059);
and U13176 (N_13176,N_12368,N_11206);
xor U13177 (N_13177,N_10880,N_10284);
xor U13178 (N_13178,N_11753,N_10844);
or U13179 (N_13179,N_10063,N_10455);
nand U13180 (N_13180,N_10735,N_10556);
or U13181 (N_13181,N_12056,N_11844);
nand U13182 (N_13182,N_10731,N_11573);
nand U13183 (N_13183,N_10948,N_11545);
nor U13184 (N_13184,N_11795,N_11804);
xnor U13185 (N_13185,N_10200,N_11771);
and U13186 (N_13186,N_12268,N_10167);
nand U13187 (N_13187,N_10705,N_10384);
and U13188 (N_13188,N_10037,N_11472);
nand U13189 (N_13189,N_12071,N_12319);
nor U13190 (N_13190,N_11296,N_10379);
nand U13191 (N_13191,N_12132,N_10214);
nand U13192 (N_13192,N_11371,N_11407);
or U13193 (N_13193,N_10784,N_11276);
nand U13194 (N_13194,N_12344,N_11285);
nand U13195 (N_13195,N_11009,N_11386);
or U13196 (N_13196,N_11694,N_12086);
nor U13197 (N_13197,N_11040,N_10262);
xor U13198 (N_13198,N_10504,N_12289);
nand U13199 (N_13199,N_11908,N_11247);
xor U13200 (N_13200,N_10229,N_11491);
nor U13201 (N_13201,N_10820,N_11925);
nand U13202 (N_13202,N_10546,N_12455);
or U13203 (N_13203,N_11021,N_11037);
xnor U13204 (N_13204,N_11157,N_10319);
xor U13205 (N_13205,N_10831,N_11695);
or U13206 (N_13206,N_10091,N_11320);
nor U13207 (N_13207,N_11185,N_11255);
nor U13208 (N_13208,N_10405,N_11881);
xor U13209 (N_13209,N_11142,N_12335);
nor U13210 (N_13210,N_12145,N_11192);
xnor U13211 (N_13211,N_11013,N_10471);
nor U13212 (N_13212,N_10902,N_10526);
xnor U13213 (N_13213,N_10220,N_11116);
nand U13214 (N_13214,N_11097,N_10009);
or U13215 (N_13215,N_10990,N_10771);
nor U13216 (N_13216,N_11883,N_12325);
and U13217 (N_13217,N_12343,N_11861);
nand U13218 (N_13218,N_12370,N_11078);
xnor U13219 (N_13219,N_11670,N_10433);
xor U13220 (N_13220,N_11455,N_10806);
xnor U13221 (N_13221,N_11170,N_11128);
and U13222 (N_13222,N_11301,N_11250);
and U13223 (N_13223,N_12067,N_11641);
and U13224 (N_13224,N_10048,N_10073);
nor U13225 (N_13225,N_11419,N_11790);
and U13226 (N_13226,N_12442,N_10123);
nor U13227 (N_13227,N_11650,N_10476);
or U13228 (N_13228,N_12212,N_11024);
or U13229 (N_13229,N_12438,N_11537);
nand U13230 (N_13230,N_10310,N_10371);
and U13231 (N_13231,N_10700,N_12280);
nand U13232 (N_13232,N_10350,N_12240);
and U13233 (N_13233,N_10577,N_10655);
nor U13234 (N_13234,N_10688,N_12121);
and U13235 (N_13235,N_12275,N_11108);
or U13236 (N_13236,N_12224,N_11318);
and U13237 (N_13237,N_11775,N_11007);
nor U13238 (N_13238,N_10980,N_10193);
nand U13239 (N_13239,N_11030,N_11297);
and U13240 (N_13240,N_10337,N_11469);
or U13241 (N_13241,N_10478,N_12458);
nand U13242 (N_13242,N_10365,N_11091);
xor U13243 (N_13243,N_11779,N_11652);
and U13244 (N_13244,N_11683,N_11151);
and U13245 (N_13245,N_10935,N_12419);
and U13246 (N_13246,N_11348,N_10669);
nand U13247 (N_13247,N_11223,N_12075);
and U13248 (N_13248,N_10127,N_12254);
nor U13249 (N_13249,N_10849,N_12342);
nand U13250 (N_13250,N_12246,N_11241);
or U13251 (N_13251,N_10005,N_11477);
and U13252 (N_13252,N_10162,N_11230);
xor U13253 (N_13253,N_10266,N_11516);
or U13254 (N_13254,N_10757,N_10636);
nand U13255 (N_13255,N_11642,N_11595);
nor U13256 (N_13256,N_10279,N_12322);
xor U13257 (N_13257,N_10583,N_10122);
nor U13258 (N_13258,N_10575,N_11631);
or U13259 (N_13259,N_11496,N_10301);
and U13260 (N_13260,N_11427,N_12033);
and U13261 (N_13261,N_12411,N_10196);
nand U13262 (N_13262,N_10028,N_10889);
nor U13263 (N_13263,N_10077,N_10354);
and U13264 (N_13264,N_12271,N_10960);
xor U13265 (N_13265,N_10280,N_10395);
or U13266 (N_13266,N_10334,N_10017);
xor U13267 (N_13267,N_12223,N_10347);
nand U13268 (N_13268,N_11440,N_11587);
nor U13269 (N_13269,N_11766,N_11912);
xnor U13270 (N_13270,N_12198,N_11894);
nand U13271 (N_13271,N_12326,N_11409);
or U13272 (N_13272,N_12273,N_11066);
nor U13273 (N_13273,N_10619,N_10081);
nand U13274 (N_13274,N_11012,N_11306);
nand U13275 (N_13275,N_11603,N_12479);
nor U13276 (N_13276,N_10420,N_12414);
xnor U13277 (N_13277,N_11789,N_10982);
nor U13278 (N_13278,N_11350,N_10795);
xor U13279 (N_13279,N_11414,N_10877);
nand U13280 (N_13280,N_10649,N_11704);
and U13281 (N_13281,N_10810,N_11705);
nand U13282 (N_13282,N_10283,N_12231);
nand U13283 (N_13283,N_11432,N_12364);
and U13284 (N_13284,N_12281,N_10920);
nor U13285 (N_13285,N_10773,N_10896);
or U13286 (N_13286,N_10707,N_10264);
or U13287 (N_13287,N_10469,N_11892);
and U13288 (N_13288,N_12332,N_12088);
or U13289 (N_13289,N_11017,N_12073);
or U13290 (N_13290,N_12467,N_11164);
and U13291 (N_13291,N_10595,N_11922);
nand U13292 (N_13292,N_11406,N_11319);
nor U13293 (N_13293,N_10435,N_11287);
and U13294 (N_13294,N_10539,N_10787);
and U13295 (N_13295,N_10527,N_11567);
nor U13296 (N_13296,N_12014,N_11305);
nor U13297 (N_13297,N_10448,N_11985);
xnor U13298 (N_13298,N_12221,N_10276);
nor U13299 (N_13299,N_10390,N_10296);
xor U13300 (N_13300,N_11949,N_10888);
nor U13301 (N_13301,N_10638,N_11872);
nand U13302 (N_13302,N_10387,N_10774);
nand U13303 (N_13303,N_10145,N_11749);
nand U13304 (N_13304,N_11150,N_12463);
and U13305 (N_13305,N_10680,N_10372);
nand U13306 (N_13306,N_11733,N_11843);
nand U13307 (N_13307,N_10468,N_12134);
or U13308 (N_13308,N_11807,N_12415);
xnor U13309 (N_13309,N_10195,N_10115);
and U13310 (N_13310,N_10438,N_12270);
nand U13311 (N_13311,N_12158,N_11935);
or U13312 (N_13312,N_11069,N_10513);
nor U13313 (N_13313,N_10728,N_10857);
nor U13314 (N_13314,N_10410,N_12407);
nand U13315 (N_13315,N_12207,N_10470);
nor U13316 (N_13316,N_10952,N_12117);
nor U13317 (N_13317,N_12162,N_12066);
nand U13318 (N_13318,N_11755,N_10568);
or U13319 (N_13319,N_12448,N_10174);
nand U13320 (N_13320,N_11506,N_11713);
nand U13321 (N_13321,N_10949,N_12053);
or U13322 (N_13322,N_11381,N_11972);
xnor U13323 (N_13323,N_12094,N_12210);
nand U13324 (N_13324,N_11071,N_10715);
nor U13325 (N_13325,N_11326,N_10499);
and U13326 (N_13326,N_11946,N_11314);
nor U13327 (N_13327,N_12476,N_11277);
nand U13328 (N_13328,N_10895,N_10874);
or U13329 (N_13329,N_10897,N_10676);
or U13330 (N_13330,N_10189,N_11724);
nor U13331 (N_13331,N_11632,N_12367);
nor U13332 (N_13332,N_10307,N_12257);
or U13333 (N_13333,N_12321,N_11260);
or U13334 (N_13334,N_10950,N_12242);
nor U13335 (N_13335,N_10364,N_10663);
and U13336 (N_13336,N_12274,N_10999);
xor U13337 (N_13337,N_10566,N_10511);
and U13338 (N_13338,N_11393,N_11560);
nor U13339 (N_13339,N_11598,N_11616);
nor U13340 (N_13340,N_12141,N_10155);
xor U13341 (N_13341,N_10252,N_10192);
nor U13342 (N_13342,N_10794,N_10439);
nor U13343 (N_13343,N_11453,N_12225);
nor U13344 (N_13344,N_11011,N_11797);
nand U13345 (N_13345,N_11127,N_10054);
xor U13346 (N_13346,N_11430,N_10579);
or U13347 (N_13347,N_11876,N_11249);
or U13348 (N_13348,N_11884,N_10712);
nor U13349 (N_13349,N_11665,N_11571);
xor U13350 (N_13350,N_10616,N_10678);
and U13351 (N_13351,N_11756,N_12043);
nand U13352 (N_13352,N_11954,N_10132);
or U13353 (N_13353,N_10597,N_10559);
nand U13354 (N_13354,N_10084,N_11092);
nor U13355 (N_13355,N_10097,N_11057);
xor U13356 (N_13356,N_11325,N_11660);
and U13357 (N_13357,N_10637,N_11144);
nor U13358 (N_13358,N_11697,N_10381);
xnor U13359 (N_13359,N_10043,N_10946);
or U13360 (N_13360,N_11298,N_12475);
nand U13361 (N_13361,N_10732,N_11194);
xor U13362 (N_13362,N_10066,N_11780);
or U13363 (N_13363,N_11934,N_10601);
xnor U13364 (N_13364,N_12301,N_11361);
or U13365 (N_13365,N_12462,N_12028);
and U13366 (N_13366,N_10030,N_10380);
nor U13367 (N_13367,N_11773,N_11417);
nor U13368 (N_13368,N_10290,N_12421);
xnor U13369 (N_13369,N_12010,N_10281);
nand U13370 (N_13370,N_11808,N_11380);
xnor U13371 (N_13371,N_10776,N_11709);
or U13372 (N_13372,N_12229,N_10581);
xor U13373 (N_13373,N_10312,N_11933);
nand U13374 (N_13374,N_12149,N_11056);
or U13375 (N_13375,N_10211,N_11702);
nand U13376 (N_13376,N_11845,N_10964);
or U13377 (N_13377,N_11161,N_10303);
nor U13378 (N_13378,N_12004,N_11945);
or U13379 (N_13379,N_12249,N_10332);
nand U13380 (N_13380,N_10963,N_10456);
nand U13381 (N_13381,N_11614,N_10052);
xnor U13382 (N_13382,N_12080,N_10886);
or U13383 (N_13383,N_12491,N_10837);
and U13384 (N_13384,N_12494,N_10069);
nor U13385 (N_13385,N_12063,N_10918);
nand U13386 (N_13386,N_11509,N_11842);
nor U13387 (N_13387,N_10904,N_11651);
xnor U13388 (N_13388,N_10876,N_10553);
nor U13389 (N_13389,N_11059,N_11329);
nor U13390 (N_13390,N_12208,N_10913);
xnor U13391 (N_13391,N_10302,N_11550);
or U13392 (N_13392,N_10201,N_11893);
nor U13393 (N_13393,N_10643,N_11994);
xnor U13394 (N_13394,N_11666,N_10586);
and U13395 (N_13395,N_10242,N_10408);
xor U13396 (N_13396,N_11754,N_12236);
xnor U13397 (N_13397,N_11885,N_10508);
nor U13398 (N_13398,N_10255,N_10576);
and U13399 (N_13399,N_12030,N_11500);
nand U13400 (N_13400,N_11111,N_10543);
and U13401 (N_13401,N_11156,N_11492);
nor U13402 (N_13402,N_10685,N_11498);
and U13403 (N_13403,N_11909,N_11678);
or U13404 (N_13404,N_12011,N_10815);
nand U13405 (N_13405,N_11738,N_10452);
and U13406 (N_13406,N_11347,N_11175);
and U13407 (N_13407,N_11877,N_10026);
nor U13408 (N_13408,N_10367,N_11929);
or U13409 (N_13409,N_12099,N_12055);
nor U13410 (N_13410,N_12255,N_11293);
xor U13411 (N_13411,N_10176,N_10258);
nand U13412 (N_13412,N_10598,N_11918);
and U13413 (N_13413,N_10991,N_10600);
nand U13414 (N_13414,N_11367,N_10366);
xor U13415 (N_13415,N_10485,N_12193);
and U13416 (N_13416,N_10653,N_10257);
and U13417 (N_13417,N_11501,N_11163);
or U13418 (N_13418,N_10335,N_10015);
xor U13419 (N_13419,N_12247,N_11781);
or U13420 (N_13420,N_10249,N_10088);
nand U13421 (N_13421,N_11121,N_10315);
and U13422 (N_13422,N_10165,N_10554);
and U13423 (N_13423,N_11903,N_10003);
xnor U13424 (N_13424,N_11269,N_11154);
xor U13425 (N_13425,N_10237,N_11942);
nor U13426 (N_13426,N_12488,N_10567);
nor U13427 (N_13427,N_11482,N_11911);
nor U13428 (N_13428,N_10206,N_12087);
nand U13429 (N_13429,N_11875,N_10399);
nand U13430 (N_13430,N_11134,N_10489);
nor U13431 (N_13431,N_11589,N_10590);
xor U13432 (N_13432,N_11488,N_11692);
nand U13433 (N_13433,N_12152,N_10495);
nor U13434 (N_13434,N_11316,N_10972);
nor U13435 (N_13435,N_10609,N_12130);
xor U13436 (N_13436,N_11630,N_11402);
nor U13437 (N_13437,N_11533,N_10957);
or U13438 (N_13438,N_11370,N_12081);
xnor U13439 (N_13439,N_11853,N_10750);
xnor U13440 (N_13440,N_10870,N_11544);
xor U13441 (N_13441,N_10391,N_11481);
nand U13442 (N_13442,N_11428,N_10109);
and U13443 (N_13443,N_11187,N_11026);
and U13444 (N_13444,N_10178,N_10865);
nand U13445 (N_13445,N_10926,N_11898);
nor U13446 (N_13446,N_10684,N_11601);
nand U13447 (N_13447,N_10807,N_10769);
nor U13448 (N_13448,N_10208,N_11529);
nor U13449 (N_13449,N_10587,N_10055);
or U13450 (N_13450,N_11228,N_10517);
or U13451 (N_13451,N_11924,N_11649);
nor U13452 (N_13452,N_11081,N_12199);
or U13453 (N_13453,N_10498,N_11006);
or U13454 (N_13454,N_11576,N_10905);
and U13455 (N_13455,N_11076,N_10943);
and U13456 (N_13456,N_10770,N_11818);
nor U13457 (N_13457,N_11307,N_10927);
or U13458 (N_13458,N_11907,N_11941);
and U13459 (N_13459,N_10863,N_11113);
nor U13460 (N_13460,N_10869,N_12318);
and U13461 (N_13461,N_10432,N_10651);
nor U13462 (N_13462,N_11982,N_10140);
xnor U13463 (N_13463,N_11068,N_11388);
and U13464 (N_13464,N_10376,N_11744);
nand U13465 (N_13465,N_10622,N_10747);
xor U13466 (N_13466,N_10293,N_12020);
and U13467 (N_13467,N_10430,N_11303);
nor U13468 (N_13468,N_11688,N_11450);
or U13469 (N_13469,N_11796,N_11330);
xor U13470 (N_13470,N_10640,N_10996);
and U13471 (N_13471,N_11372,N_12156);
nor U13472 (N_13472,N_12161,N_10830);
nand U13473 (N_13473,N_11459,N_11961);
or U13474 (N_13474,N_11420,N_11963);
and U13475 (N_13475,N_10027,N_11554);
nor U13476 (N_13476,N_10823,N_12157);
nor U13477 (N_13477,N_11394,N_12093);
or U13478 (N_13478,N_12350,N_11976);
and U13479 (N_13479,N_11525,N_10212);
xnor U13480 (N_13480,N_11830,N_10777);
or U13481 (N_13481,N_10067,N_10818);
xnor U13482 (N_13482,N_10272,N_12459);
nand U13483 (N_13483,N_10246,N_11839);
or U13484 (N_13484,N_12205,N_11582);
xor U13485 (N_13485,N_11028,N_10867);
or U13486 (N_13486,N_10822,N_10791);
and U13487 (N_13487,N_11168,N_11646);
or U13488 (N_13488,N_10644,N_11446);
xor U13489 (N_13489,N_12203,N_11251);
nor U13490 (N_13490,N_11103,N_10013);
or U13491 (N_13491,N_11118,N_12031);
nor U13492 (N_13492,N_10138,N_11398);
nand U13493 (N_13493,N_11643,N_12062);
nor U13494 (N_13494,N_10574,N_12365);
nand U13495 (N_13495,N_10922,N_11836);
nor U13496 (N_13496,N_11264,N_10979);
or U13497 (N_13497,N_11594,N_10614);
or U13498 (N_13498,N_10571,N_11572);
or U13499 (N_13499,N_11973,N_12439);
xor U13500 (N_13500,N_10259,N_12492);
xor U13501 (N_13501,N_10790,N_12457);
xnor U13502 (N_13502,N_12412,N_10322);
and U13503 (N_13503,N_10758,N_11680);
nor U13504 (N_13504,N_10466,N_11732);
xor U13505 (N_13505,N_11373,N_10661);
nand U13506 (N_13506,N_11360,N_11662);
and U13507 (N_13507,N_10202,N_11826);
or U13508 (N_13508,N_10679,N_10046);
nand U13509 (N_13509,N_11404,N_11823);
xor U13510 (N_13510,N_12315,N_11959);
nor U13511 (N_13511,N_10828,N_10509);
or U13512 (N_13512,N_10748,N_10743);
nand U13513 (N_13513,N_10507,N_11358);
nand U13514 (N_13514,N_10041,N_10570);
and U13515 (N_13515,N_12436,N_11036);
or U13516 (N_13516,N_10146,N_12386);
xnor U13517 (N_13517,N_11117,N_10592);
xnor U13518 (N_13518,N_10838,N_10308);
nand U13519 (N_13519,N_11045,N_11873);
nand U13520 (N_13520,N_11505,N_11489);
xor U13521 (N_13521,N_12276,N_11171);
and U13522 (N_13522,N_12441,N_12282);
nand U13523 (N_13523,N_10040,N_11202);
xnor U13524 (N_13524,N_10510,N_10521);
and U13525 (N_13525,N_11647,N_11166);
or U13526 (N_13526,N_10724,N_10039);
nand U13527 (N_13527,N_11183,N_11165);
and U13528 (N_13528,N_11100,N_12123);
nor U13529 (N_13529,N_10051,N_11179);
nand U13530 (N_13530,N_10966,N_11962);
nor U13531 (N_13531,N_10150,N_10866);
and U13532 (N_13532,N_10453,N_10407);
and U13533 (N_13533,N_10811,N_10906);
or U13534 (N_13534,N_12054,N_12305);
or U13535 (N_13535,N_12022,N_10578);
nor U13536 (N_13536,N_11625,N_10626);
xor U13537 (N_13537,N_11278,N_11454);
xnor U13538 (N_13538,N_10421,N_10698);
and U13539 (N_13539,N_12133,N_12182);
nor U13540 (N_13540,N_12262,N_11199);
xnor U13541 (N_13541,N_11953,N_11193);
nor U13542 (N_13542,N_10226,N_10692);
or U13543 (N_13543,N_12444,N_11112);
and U13544 (N_13544,N_12446,N_10973);
nand U13545 (N_13545,N_10881,N_11944);
and U13546 (N_13546,N_10625,N_11913);
xor U13547 (N_13547,N_11110,N_11177);
nand U13548 (N_13548,N_12021,N_10660);
or U13549 (N_13549,N_10985,N_12045);
xnor U13550 (N_13550,N_10714,N_11499);
nor U13551 (N_13551,N_12374,N_12025);
and U13552 (N_13552,N_10928,N_10434);
and U13553 (N_13553,N_10516,N_11436);
nand U13554 (N_13554,N_11397,N_10021);
nor U13555 (N_13555,N_11335,N_11980);
or U13556 (N_13556,N_11423,N_11413);
or U13557 (N_13557,N_11014,N_11389);
xor U13558 (N_13558,N_11947,N_11810);
nand U13559 (N_13559,N_12285,N_11120);
and U13560 (N_13560,N_12190,N_11541);
nand U13561 (N_13561,N_12175,N_10955);
or U13562 (N_13562,N_11542,N_11205);
and U13563 (N_13563,N_10775,N_10924);
and U13564 (N_13564,N_10292,N_10001);
or U13565 (N_13565,N_11107,N_10726);
or U13566 (N_13566,N_12041,N_11088);
xnor U13567 (N_13567,N_11760,N_11728);
xor U13568 (N_13568,N_12187,N_12191);
and U13569 (N_13569,N_11879,N_12294);
nor U13570 (N_13570,N_11511,N_10058);
nand U13571 (N_13571,N_10095,N_10232);
or U13572 (N_13572,N_10560,N_11145);
nor U13573 (N_13573,N_12173,N_12172);
xnor U13574 (N_13574,N_12345,N_10569);
and U13575 (N_13575,N_11104,N_10506);
or U13576 (N_13576,N_12360,N_10654);
or U13577 (N_13577,N_12154,N_11494);
nor U13578 (N_13578,N_10168,N_10269);
nand U13579 (N_13579,N_11242,N_12387);
nor U13580 (N_13580,N_10236,N_10686);
nor U13581 (N_13581,N_11204,N_11153);
nor U13582 (N_13582,N_11274,N_10024);
nand U13583 (N_13583,N_10827,N_12297);
and U13584 (N_13584,N_11574,N_12404);
nor U13585 (N_13585,N_12216,N_11997);
nand U13586 (N_13586,N_11267,N_10462);
nor U13587 (N_13587,N_12009,N_11331);
and U13588 (N_13588,N_11792,N_11622);
xor U13589 (N_13589,N_10824,N_11868);
nor U13590 (N_13590,N_10958,N_10314);
nor U13591 (N_13591,N_10010,N_12487);
nor U13592 (N_13592,N_10505,N_11722);
nand U13593 (N_13593,N_11475,N_11152);
nor U13594 (N_13594,N_10014,N_11901);
or U13595 (N_13595,N_10706,N_12245);
and U13596 (N_13596,N_11882,N_11765);
and U13597 (N_13597,N_10106,N_10187);
or U13598 (N_13598,N_12267,N_10361);
or U13599 (N_13599,N_11626,N_11474);
xnor U13600 (N_13600,N_10929,N_11979);
nand U13601 (N_13601,N_10851,N_11570);
nand U13602 (N_13602,N_12379,N_12252);
and U13603 (N_13603,N_10004,N_10409);
nor U13604 (N_13604,N_12497,N_10859);
xor U13605 (N_13605,N_11865,N_11222);
nand U13606 (N_13606,N_11138,N_12176);
or U13607 (N_13607,N_11031,N_12024);
nand U13608 (N_13608,N_12393,N_10481);
xor U13609 (N_13609,N_12440,N_12293);
nand U13610 (N_13610,N_10618,N_10848);
xor U13611 (N_13611,N_11266,N_10723);
xor U13612 (N_13612,N_11243,N_11410);
xor U13613 (N_13613,N_11311,N_10780);
or U13614 (N_13614,N_10582,N_10486);
nand U13615 (N_13615,N_12061,N_11369);
or U13616 (N_13616,N_11139,N_10056);
nand U13617 (N_13617,N_12399,N_10225);
xnor U13618 (N_13618,N_12000,N_10887);
xnor U13619 (N_13619,N_10785,N_12112);
nand U13620 (N_13620,N_10328,N_10656);
nand U13621 (N_13621,N_11938,N_12039);
or U13622 (N_13622,N_10181,N_11362);
nand U13623 (N_13623,N_11777,N_12065);
nand U13624 (N_13624,N_12382,N_10083);
nor U13625 (N_13625,N_10369,N_11246);
xnor U13626 (N_13626,N_11751,N_12147);
or U13627 (N_13627,N_11248,N_10483);
or U13628 (N_13628,N_10814,N_12144);
and U13629 (N_13629,N_11520,N_11074);
nand U13630 (N_13630,N_11621,N_11581);
or U13631 (N_13631,N_10423,N_11682);
xnor U13632 (N_13632,N_11521,N_12038);
nor U13633 (N_13633,N_10604,N_10646);
xor U13634 (N_13634,N_10850,N_12008);
nor U13635 (N_13635,N_12477,N_11899);
xor U13636 (N_13636,N_10179,N_10245);
nor U13637 (N_13637,N_11730,N_12101);
xor U13638 (N_13638,N_11714,N_11384);
nor U13639 (N_13639,N_11967,N_11661);
nand U13640 (N_13640,N_11399,N_11999);
nor U13641 (N_13641,N_10691,N_11989);
and U13642 (N_13642,N_11115,N_11783);
nand U13643 (N_13643,N_11191,N_10956);
and U13644 (N_13644,N_11615,N_11442);
nand U13645 (N_13645,N_10713,N_11700);
or U13646 (N_13646,N_11085,N_11534);
xnor U13647 (N_13647,N_10763,N_10683);
nor U13648 (N_13648,N_11435,N_10406);
xnor U13649 (N_13649,N_12265,N_12012);
and U13650 (N_13650,N_12050,N_10227);
nor U13651 (N_13651,N_11155,N_11635);
nand U13652 (N_13652,N_10411,N_12349);
or U13653 (N_13653,N_10797,N_11669);
or U13654 (N_13654,N_11791,N_10710);
nor U13655 (N_13655,N_12427,N_11299);
or U13656 (N_13656,N_11441,N_11764);
or U13657 (N_13657,N_10034,N_12445);
xnor U13658 (N_13658,N_10981,N_10741);
nand U13659 (N_13659,N_12291,N_11971);
xnor U13660 (N_13660,N_10803,N_10762);
and U13661 (N_13661,N_12136,N_12034);
nor U13662 (N_13662,N_10915,N_10060);
xor U13663 (N_13663,N_10351,N_10832);
nand U13664 (N_13664,N_10079,N_10612);
nor U13665 (N_13665,N_11016,N_11346);
and U13666 (N_13666,N_12486,N_11493);
xnor U13667 (N_13667,N_12401,N_10976);
and U13668 (N_13668,N_10695,N_10450);
or U13669 (N_13669,N_11273,N_10538);
nand U13670 (N_13670,N_12196,N_12278);
and U13671 (N_13671,N_10759,N_11690);
or U13672 (N_13672,N_11422,N_11424);
and U13673 (N_13673,N_11671,N_11275);
nand U13674 (N_13674,N_11364,N_11904);
or U13675 (N_13675,N_10503,N_12352);
or U13676 (N_13676,N_12435,N_11216);
nand U13677 (N_13677,N_10593,N_10729);
and U13678 (N_13678,N_11558,N_10720);
nand U13679 (N_13679,N_10273,N_10154);
and U13680 (N_13680,N_12381,N_10898);
nand U13681 (N_13681,N_11672,N_11065);
nand U13682 (N_13682,N_11852,N_12104);
xnor U13683 (N_13683,N_11684,N_10992);
xor U13684 (N_13684,N_10648,N_11342);
nor U13685 (N_13685,N_10256,N_10185);
nand U13686 (N_13686,N_11937,N_11061);
xnor U13687 (N_13687,N_11983,N_12150);
nor U13688 (N_13688,N_11854,N_10251);
nand U13689 (N_13689,N_10118,N_11023);
xnor U13690 (N_13690,N_11125,N_11701);
or U13691 (N_13691,N_11561,N_10533);
xnor U13692 (N_13692,N_11217,N_11445);
and U13693 (N_13693,N_12482,N_11010);
nor U13694 (N_13694,N_12384,N_12019);
nor U13695 (N_13695,N_12092,N_10153);
nand U13696 (N_13696,N_10061,N_11345);
nor U13697 (N_13697,N_11186,N_11096);
nor U13698 (N_13698,N_12334,N_11606);
or U13699 (N_13699,N_10523,N_12040);
nor U13700 (N_13700,N_10833,N_11434);
nor U13701 (N_13701,N_11809,N_10974);
xor U13702 (N_13702,N_12417,N_10300);
or U13703 (N_13703,N_10107,N_10627);
or U13704 (N_13704,N_10659,N_10694);
or U13705 (N_13705,N_12333,N_10029);
nor U13706 (N_13706,N_11712,N_11920);
nor U13707 (N_13707,N_11772,N_11580);
and U13708 (N_13708,N_11291,N_11636);
xnor U13709 (N_13709,N_12396,N_11290);
xor U13710 (N_13710,N_11992,N_11905);
xnor U13711 (N_13711,N_10639,N_10018);
and U13712 (N_13712,N_11072,N_12361);
or U13713 (N_13713,N_10121,N_11086);
nand U13714 (N_13714,N_11197,N_11137);
xnor U13715 (N_13715,N_12111,N_11146);
nor U13716 (N_13716,N_10480,N_11289);
nand U13717 (N_13717,N_10261,N_12108);
or U13718 (N_13718,N_12037,N_10792);
xnor U13719 (N_13719,N_12165,N_10719);
xor U13720 (N_13720,N_12125,N_10667);
and U13721 (N_13721,N_10321,N_12337);
nor U13722 (N_13722,N_12329,N_10497);
nor U13723 (N_13723,N_12429,N_11745);
and U13724 (N_13724,N_10282,N_10998);
and U13725 (N_13725,N_11546,N_11623);
nand U13726 (N_13726,N_11458,N_12437);
xnor U13727 (N_13727,N_12499,N_11043);
xor U13728 (N_13728,N_10441,N_11860);
nand U13729 (N_13729,N_10893,N_12042);
nand U13730 (N_13730,N_12258,N_11109);
and U13731 (N_13731,N_11123,N_11993);
nand U13732 (N_13732,N_10142,N_10883);
xor U13733 (N_13733,N_12102,N_12340);
and U13734 (N_13734,N_10460,N_10173);
or U13735 (N_13735,N_12213,N_10681);
xor U13736 (N_13736,N_10936,N_11244);
nand U13737 (N_13737,N_10944,N_12371);
or U13738 (N_13738,N_11639,N_11310);
and U13739 (N_13739,N_12376,N_10286);
or U13740 (N_13740,N_11174,N_10921);
and U13741 (N_13741,N_10309,N_11094);
and U13742 (N_13742,N_10585,N_11856);
xnor U13743 (N_13743,N_10177,N_11471);
nor U13744 (N_13744,N_10049,N_12269);
nor U13745 (N_13745,N_11637,N_11114);
or U13746 (N_13746,N_10417,N_11776);
xnor U13747 (N_13747,N_10105,N_10858);
or U13748 (N_13748,N_10610,N_11265);
and U13749 (N_13749,N_11261,N_12362);
or U13750 (N_13750,N_11345,N_11019);
or U13751 (N_13751,N_11486,N_12341);
nor U13752 (N_13752,N_10115,N_12005);
or U13753 (N_13753,N_10028,N_11242);
or U13754 (N_13754,N_10724,N_11769);
or U13755 (N_13755,N_10706,N_11783);
xor U13756 (N_13756,N_10193,N_11780);
or U13757 (N_13757,N_12223,N_11536);
or U13758 (N_13758,N_10051,N_12044);
and U13759 (N_13759,N_11057,N_12452);
or U13760 (N_13760,N_12307,N_10220);
or U13761 (N_13761,N_12031,N_10299);
xnor U13762 (N_13762,N_12431,N_11537);
xnor U13763 (N_13763,N_11408,N_12439);
nand U13764 (N_13764,N_10978,N_10301);
nand U13765 (N_13765,N_12330,N_11271);
and U13766 (N_13766,N_12057,N_10105);
or U13767 (N_13767,N_12290,N_11026);
or U13768 (N_13768,N_10479,N_10238);
or U13769 (N_13769,N_10214,N_10760);
xnor U13770 (N_13770,N_12205,N_10808);
xor U13771 (N_13771,N_12249,N_11139);
nand U13772 (N_13772,N_11083,N_11714);
nand U13773 (N_13773,N_10478,N_11601);
nor U13774 (N_13774,N_11317,N_11771);
xor U13775 (N_13775,N_11380,N_11352);
xor U13776 (N_13776,N_10350,N_11489);
nor U13777 (N_13777,N_10591,N_11747);
nor U13778 (N_13778,N_11236,N_12341);
nor U13779 (N_13779,N_11478,N_10627);
or U13780 (N_13780,N_11281,N_11404);
nand U13781 (N_13781,N_10550,N_11209);
or U13782 (N_13782,N_10975,N_12166);
xor U13783 (N_13783,N_11786,N_10335);
nor U13784 (N_13784,N_10523,N_10952);
xnor U13785 (N_13785,N_12074,N_11092);
nand U13786 (N_13786,N_10134,N_10946);
nor U13787 (N_13787,N_11298,N_10517);
nand U13788 (N_13788,N_11047,N_10749);
nor U13789 (N_13789,N_12390,N_11233);
xnor U13790 (N_13790,N_11401,N_10331);
xnor U13791 (N_13791,N_10066,N_11744);
nand U13792 (N_13792,N_11300,N_10191);
nand U13793 (N_13793,N_11953,N_10022);
and U13794 (N_13794,N_11085,N_12066);
xnor U13795 (N_13795,N_10976,N_10662);
nand U13796 (N_13796,N_11257,N_11817);
nor U13797 (N_13797,N_11103,N_11698);
or U13798 (N_13798,N_12360,N_11822);
xnor U13799 (N_13799,N_10929,N_12083);
or U13800 (N_13800,N_10976,N_10854);
and U13801 (N_13801,N_12464,N_10426);
nand U13802 (N_13802,N_11835,N_11372);
nor U13803 (N_13803,N_11264,N_11343);
and U13804 (N_13804,N_11975,N_12415);
nor U13805 (N_13805,N_11213,N_12193);
nor U13806 (N_13806,N_12053,N_11718);
nand U13807 (N_13807,N_10142,N_11691);
and U13808 (N_13808,N_10425,N_12138);
nand U13809 (N_13809,N_10485,N_10444);
or U13810 (N_13810,N_10540,N_11000);
xnor U13811 (N_13811,N_10941,N_10631);
and U13812 (N_13812,N_11601,N_10085);
nor U13813 (N_13813,N_10482,N_10441);
xor U13814 (N_13814,N_12261,N_12287);
xor U13815 (N_13815,N_10116,N_10199);
or U13816 (N_13816,N_11394,N_10941);
nor U13817 (N_13817,N_11844,N_10163);
nand U13818 (N_13818,N_10182,N_11543);
xor U13819 (N_13819,N_10877,N_11840);
and U13820 (N_13820,N_11958,N_12403);
nand U13821 (N_13821,N_10025,N_10764);
nor U13822 (N_13822,N_11425,N_10021);
nand U13823 (N_13823,N_11853,N_11442);
or U13824 (N_13824,N_11179,N_11623);
or U13825 (N_13825,N_11741,N_12365);
and U13826 (N_13826,N_10611,N_12194);
and U13827 (N_13827,N_10733,N_12497);
nand U13828 (N_13828,N_10314,N_12304);
nor U13829 (N_13829,N_11272,N_10937);
or U13830 (N_13830,N_11767,N_10312);
and U13831 (N_13831,N_11904,N_11342);
and U13832 (N_13832,N_10162,N_10197);
and U13833 (N_13833,N_11675,N_10703);
nor U13834 (N_13834,N_11212,N_11754);
and U13835 (N_13835,N_10967,N_10656);
nor U13836 (N_13836,N_12433,N_10737);
nor U13837 (N_13837,N_12413,N_11415);
xnor U13838 (N_13838,N_10470,N_10139);
or U13839 (N_13839,N_12216,N_10966);
xor U13840 (N_13840,N_10117,N_12148);
or U13841 (N_13841,N_11227,N_11584);
nand U13842 (N_13842,N_10277,N_12434);
nor U13843 (N_13843,N_11434,N_11808);
or U13844 (N_13844,N_10006,N_10333);
nor U13845 (N_13845,N_11907,N_11846);
and U13846 (N_13846,N_11307,N_12271);
nor U13847 (N_13847,N_10335,N_12297);
and U13848 (N_13848,N_11280,N_11688);
or U13849 (N_13849,N_11408,N_12451);
and U13850 (N_13850,N_10342,N_12379);
nor U13851 (N_13851,N_10940,N_10758);
and U13852 (N_13852,N_11787,N_11361);
xnor U13853 (N_13853,N_10668,N_11573);
nand U13854 (N_13854,N_12198,N_11743);
nor U13855 (N_13855,N_11092,N_10057);
nor U13856 (N_13856,N_11608,N_11138);
nor U13857 (N_13857,N_11511,N_11058);
or U13858 (N_13858,N_11228,N_10816);
xnor U13859 (N_13859,N_10431,N_12228);
or U13860 (N_13860,N_11863,N_12122);
and U13861 (N_13861,N_12381,N_10689);
nor U13862 (N_13862,N_10779,N_10649);
xor U13863 (N_13863,N_11329,N_11217);
nor U13864 (N_13864,N_12035,N_12136);
or U13865 (N_13865,N_11960,N_11249);
nand U13866 (N_13866,N_10442,N_10703);
nor U13867 (N_13867,N_11374,N_10566);
nor U13868 (N_13868,N_10387,N_11168);
xor U13869 (N_13869,N_10272,N_12101);
nor U13870 (N_13870,N_11824,N_11494);
xnor U13871 (N_13871,N_11625,N_11312);
or U13872 (N_13872,N_11435,N_12307);
and U13873 (N_13873,N_12354,N_10891);
xnor U13874 (N_13874,N_11709,N_11772);
nor U13875 (N_13875,N_11093,N_12090);
nand U13876 (N_13876,N_11109,N_11104);
and U13877 (N_13877,N_11420,N_11238);
nand U13878 (N_13878,N_10565,N_10309);
nor U13879 (N_13879,N_12020,N_11979);
or U13880 (N_13880,N_10264,N_11487);
nor U13881 (N_13881,N_12043,N_10661);
and U13882 (N_13882,N_10405,N_10348);
nand U13883 (N_13883,N_10717,N_11232);
or U13884 (N_13884,N_12490,N_11812);
and U13885 (N_13885,N_10227,N_10925);
or U13886 (N_13886,N_11827,N_11572);
nand U13887 (N_13887,N_11277,N_10978);
xnor U13888 (N_13888,N_11309,N_10333);
and U13889 (N_13889,N_10301,N_11095);
nor U13890 (N_13890,N_10659,N_10118);
and U13891 (N_13891,N_10558,N_11598);
xnor U13892 (N_13892,N_10434,N_10969);
xor U13893 (N_13893,N_10683,N_12073);
or U13894 (N_13894,N_10989,N_11297);
nand U13895 (N_13895,N_11638,N_11125);
nand U13896 (N_13896,N_11009,N_10561);
xnor U13897 (N_13897,N_10496,N_11316);
nand U13898 (N_13898,N_10207,N_11580);
xnor U13899 (N_13899,N_10946,N_11782);
nand U13900 (N_13900,N_10999,N_10112);
nor U13901 (N_13901,N_11156,N_11612);
xnor U13902 (N_13902,N_12183,N_11275);
and U13903 (N_13903,N_12079,N_10315);
nand U13904 (N_13904,N_11449,N_10834);
nor U13905 (N_13905,N_12393,N_10515);
nor U13906 (N_13906,N_10628,N_10119);
and U13907 (N_13907,N_10815,N_11837);
and U13908 (N_13908,N_10222,N_10888);
and U13909 (N_13909,N_11216,N_11352);
nor U13910 (N_13910,N_10120,N_10461);
and U13911 (N_13911,N_11892,N_12375);
and U13912 (N_13912,N_12154,N_10882);
nand U13913 (N_13913,N_11615,N_11978);
or U13914 (N_13914,N_12092,N_12012);
xnor U13915 (N_13915,N_12380,N_11701);
nor U13916 (N_13916,N_11109,N_10022);
or U13917 (N_13917,N_11717,N_11542);
nand U13918 (N_13918,N_11510,N_10434);
nand U13919 (N_13919,N_10075,N_11825);
nand U13920 (N_13920,N_12010,N_12020);
or U13921 (N_13921,N_10921,N_12298);
or U13922 (N_13922,N_12432,N_11029);
nand U13923 (N_13923,N_10240,N_11235);
xor U13924 (N_13924,N_10574,N_11464);
nor U13925 (N_13925,N_10623,N_10770);
and U13926 (N_13926,N_11924,N_11464);
nor U13927 (N_13927,N_10502,N_10814);
and U13928 (N_13928,N_10304,N_12046);
xnor U13929 (N_13929,N_11787,N_10868);
nand U13930 (N_13930,N_11703,N_10400);
and U13931 (N_13931,N_11892,N_10769);
nor U13932 (N_13932,N_12213,N_12146);
and U13933 (N_13933,N_12253,N_11016);
or U13934 (N_13934,N_11234,N_10025);
or U13935 (N_13935,N_10303,N_11854);
nand U13936 (N_13936,N_11013,N_10450);
and U13937 (N_13937,N_12029,N_11351);
and U13938 (N_13938,N_11604,N_10707);
nor U13939 (N_13939,N_11716,N_12384);
xnor U13940 (N_13940,N_11187,N_10172);
or U13941 (N_13941,N_11930,N_11119);
xor U13942 (N_13942,N_11158,N_10775);
nand U13943 (N_13943,N_12090,N_10505);
or U13944 (N_13944,N_11676,N_12282);
or U13945 (N_13945,N_11403,N_10707);
xor U13946 (N_13946,N_11860,N_12208);
and U13947 (N_13947,N_12073,N_11858);
nand U13948 (N_13948,N_10051,N_11636);
or U13949 (N_13949,N_10828,N_11980);
xnor U13950 (N_13950,N_10933,N_11888);
nor U13951 (N_13951,N_11369,N_10556);
nor U13952 (N_13952,N_12254,N_11951);
xor U13953 (N_13953,N_11128,N_10036);
xnor U13954 (N_13954,N_11982,N_10078);
xnor U13955 (N_13955,N_11164,N_10747);
xnor U13956 (N_13956,N_10955,N_10025);
nor U13957 (N_13957,N_10539,N_10350);
or U13958 (N_13958,N_11060,N_12162);
xnor U13959 (N_13959,N_12433,N_10123);
or U13960 (N_13960,N_10316,N_11959);
or U13961 (N_13961,N_11086,N_11213);
nand U13962 (N_13962,N_11060,N_10017);
or U13963 (N_13963,N_11977,N_10118);
xnor U13964 (N_13964,N_12417,N_11519);
nand U13965 (N_13965,N_11648,N_12355);
nand U13966 (N_13966,N_10821,N_10690);
and U13967 (N_13967,N_11857,N_12175);
and U13968 (N_13968,N_11621,N_10156);
and U13969 (N_13969,N_10171,N_11465);
xor U13970 (N_13970,N_10280,N_10313);
or U13971 (N_13971,N_10384,N_12214);
xor U13972 (N_13972,N_11542,N_11435);
and U13973 (N_13973,N_12129,N_10138);
nor U13974 (N_13974,N_10102,N_11823);
nor U13975 (N_13975,N_12492,N_10749);
xor U13976 (N_13976,N_10068,N_11846);
nand U13977 (N_13977,N_12402,N_10458);
nand U13978 (N_13978,N_10681,N_10333);
and U13979 (N_13979,N_10878,N_10957);
or U13980 (N_13980,N_11367,N_10925);
or U13981 (N_13981,N_11184,N_10155);
nand U13982 (N_13982,N_11661,N_12097);
nor U13983 (N_13983,N_11206,N_11284);
xor U13984 (N_13984,N_11903,N_12443);
or U13985 (N_13985,N_11406,N_11634);
xnor U13986 (N_13986,N_10209,N_11969);
nor U13987 (N_13987,N_11971,N_12036);
or U13988 (N_13988,N_10919,N_11597);
and U13989 (N_13989,N_11038,N_11065);
or U13990 (N_13990,N_10225,N_10613);
nand U13991 (N_13991,N_11056,N_11788);
nor U13992 (N_13992,N_11354,N_12167);
xor U13993 (N_13993,N_12253,N_11577);
and U13994 (N_13994,N_11337,N_11798);
or U13995 (N_13995,N_10669,N_10684);
nand U13996 (N_13996,N_10096,N_10732);
nand U13997 (N_13997,N_11458,N_11233);
or U13998 (N_13998,N_10459,N_10805);
nand U13999 (N_13999,N_11817,N_11424);
nor U14000 (N_14000,N_10216,N_10176);
nor U14001 (N_14001,N_10367,N_10209);
xnor U14002 (N_14002,N_11065,N_10070);
or U14003 (N_14003,N_12017,N_11722);
xnor U14004 (N_14004,N_11913,N_11623);
nor U14005 (N_14005,N_11319,N_11200);
nor U14006 (N_14006,N_11148,N_10260);
nand U14007 (N_14007,N_12078,N_11443);
and U14008 (N_14008,N_11152,N_10884);
and U14009 (N_14009,N_10134,N_11844);
nor U14010 (N_14010,N_10910,N_11850);
or U14011 (N_14011,N_10818,N_10642);
or U14012 (N_14012,N_11580,N_11879);
xor U14013 (N_14013,N_10945,N_11554);
and U14014 (N_14014,N_10957,N_11217);
nand U14015 (N_14015,N_10855,N_10890);
nand U14016 (N_14016,N_10958,N_10025);
nand U14017 (N_14017,N_10914,N_11244);
and U14018 (N_14018,N_12493,N_11372);
xnor U14019 (N_14019,N_12202,N_10871);
nor U14020 (N_14020,N_11530,N_11095);
and U14021 (N_14021,N_10571,N_12375);
nand U14022 (N_14022,N_10725,N_10910);
nor U14023 (N_14023,N_11053,N_10597);
nand U14024 (N_14024,N_11004,N_12211);
or U14025 (N_14025,N_11205,N_12345);
nand U14026 (N_14026,N_11932,N_10208);
nand U14027 (N_14027,N_11408,N_10578);
or U14028 (N_14028,N_10849,N_12328);
and U14029 (N_14029,N_11736,N_10048);
xor U14030 (N_14030,N_10221,N_12456);
xnor U14031 (N_14031,N_10081,N_10029);
xor U14032 (N_14032,N_10208,N_12387);
nor U14033 (N_14033,N_10628,N_10228);
or U14034 (N_14034,N_11384,N_11022);
nor U14035 (N_14035,N_12125,N_11612);
xor U14036 (N_14036,N_10593,N_10279);
and U14037 (N_14037,N_11619,N_10775);
xnor U14038 (N_14038,N_10022,N_11294);
nand U14039 (N_14039,N_10385,N_11423);
or U14040 (N_14040,N_12001,N_10325);
or U14041 (N_14041,N_11498,N_10547);
nand U14042 (N_14042,N_10336,N_11770);
nand U14043 (N_14043,N_10155,N_10998);
nor U14044 (N_14044,N_11249,N_11616);
xnor U14045 (N_14045,N_11691,N_11292);
nand U14046 (N_14046,N_11316,N_11475);
nand U14047 (N_14047,N_11942,N_11819);
nor U14048 (N_14048,N_11382,N_11335);
nor U14049 (N_14049,N_10788,N_10019);
nand U14050 (N_14050,N_10715,N_12017);
and U14051 (N_14051,N_10333,N_11608);
xor U14052 (N_14052,N_10963,N_10342);
and U14053 (N_14053,N_12302,N_11286);
or U14054 (N_14054,N_10087,N_11555);
or U14055 (N_14055,N_11787,N_12115);
and U14056 (N_14056,N_11527,N_11363);
nand U14057 (N_14057,N_11854,N_10765);
nor U14058 (N_14058,N_11134,N_10037);
or U14059 (N_14059,N_10504,N_11378);
or U14060 (N_14060,N_10538,N_11314);
nor U14061 (N_14061,N_12215,N_10825);
nand U14062 (N_14062,N_10859,N_11868);
or U14063 (N_14063,N_12049,N_12112);
or U14064 (N_14064,N_10068,N_12323);
and U14065 (N_14065,N_12015,N_11555);
nor U14066 (N_14066,N_10027,N_10927);
nor U14067 (N_14067,N_11431,N_10793);
nand U14068 (N_14068,N_11514,N_11586);
and U14069 (N_14069,N_10882,N_11593);
or U14070 (N_14070,N_10533,N_11663);
or U14071 (N_14071,N_10232,N_12248);
xnor U14072 (N_14072,N_11008,N_12100);
xnor U14073 (N_14073,N_10759,N_10298);
nand U14074 (N_14074,N_12159,N_11965);
nor U14075 (N_14075,N_12311,N_10615);
nor U14076 (N_14076,N_11311,N_11033);
and U14077 (N_14077,N_12224,N_10678);
or U14078 (N_14078,N_10219,N_11514);
and U14079 (N_14079,N_12022,N_10770);
and U14080 (N_14080,N_12228,N_11614);
or U14081 (N_14081,N_10477,N_11021);
xor U14082 (N_14082,N_10720,N_10489);
nand U14083 (N_14083,N_10230,N_10806);
or U14084 (N_14084,N_10935,N_10721);
nor U14085 (N_14085,N_11687,N_10626);
or U14086 (N_14086,N_12456,N_10515);
nand U14087 (N_14087,N_10513,N_11151);
or U14088 (N_14088,N_10936,N_10233);
or U14089 (N_14089,N_10516,N_11119);
nand U14090 (N_14090,N_11644,N_10536);
or U14091 (N_14091,N_11500,N_11723);
and U14092 (N_14092,N_10423,N_11304);
nand U14093 (N_14093,N_12490,N_10229);
and U14094 (N_14094,N_11807,N_11192);
nor U14095 (N_14095,N_10030,N_12011);
or U14096 (N_14096,N_10597,N_10805);
xor U14097 (N_14097,N_10803,N_10240);
or U14098 (N_14098,N_10785,N_11429);
and U14099 (N_14099,N_10380,N_11840);
nor U14100 (N_14100,N_11243,N_11850);
nand U14101 (N_14101,N_10402,N_10997);
xnor U14102 (N_14102,N_10262,N_10851);
xor U14103 (N_14103,N_10747,N_10006);
or U14104 (N_14104,N_11380,N_11874);
or U14105 (N_14105,N_10267,N_12360);
or U14106 (N_14106,N_10928,N_10937);
and U14107 (N_14107,N_10842,N_10494);
and U14108 (N_14108,N_12131,N_11575);
and U14109 (N_14109,N_10430,N_11102);
or U14110 (N_14110,N_10416,N_11885);
nor U14111 (N_14111,N_12209,N_11346);
nor U14112 (N_14112,N_12258,N_12029);
and U14113 (N_14113,N_11731,N_11553);
or U14114 (N_14114,N_11503,N_11539);
nand U14115 (N_14115,N_10491,N_10461);
nand U14116 (N_14116,N_10346,N_10439);
nor U14117 (N_14117,N_11694,N_11054);
nor U14118 (N_14118,N_11156,N_11976);
or U14119 (N_14119,N_12165,N_12290);
or U14120 (N_14120,N_10508,N_11037);
and U14121 (N_14121,N_11320,N_11610);
nor U14122 (N_14122,N_11208,N_10938);
and U14123 (N_14123,N_11626,N_10854);
or U14124 (N_14124,N_10966,N_10086);
nand U14125 (N_14125,N_11500,N_10402);
nand U14126 (N_14126,N_11674,N_10863);
nor U14127 (N_14127,N_11693,N_11620);
and U14128 (N_14128,N_11732,N_11961);
and U14129 (N_14129,N_10488,N_12422);
and U14130 (N_14130,N_10951,N_10923);
xor U14131 (N_14131,N_11855,N_10939);
nand U14132 (N_14132,N_12378,N_11795);
nand U14133 (N_14133,N_10428,N_10691);
nor U14134 (N_14134,N_11878,N_11565);
nor U14135 (N_14135,N_11161,N_11998);
nor U14136 (N_14136,N_11224,N_11196);
nand U14137 (N_14137,N_11566,N_12475);
or U14138 (N_14138,N_10708,N_10644);
xnor U14139 (N_14139,N_11343,N_10911);
or U14140 (N_14140,N_11265,N_12305);
and U14141 (N_14141,N_10886,N_10142);
and U14142 (N_14142,N_10202,N_10149);
nor U14143 (N_14143,N_12190,N_11678);
or U14144 (N_14144,N_12387,N_11994);
nand U14145 (N_14145,N_11041,N_12037);
or U14146 (N_14146,N_10724,N_10567);
nand U14147 (N_14147,N_11305,N_10790);
nor U14148 (N_14148,N_12044,N_10199);
nor U14149 (N_14149,N_11151,N_11401);
nor U14150 (N_14150,N_10318,N_11887);
xnor U14151 (N_14151,N_11173,N_10306);
nor U14152 (N_14152,N_12199,N_11615);
xnor U14153 (N_14153,N_10444,N_10611);
nand U14154 (N_14154,N_11911,N_11728);
or U14155 (N_14155,N_12214,N_11613);
and U14156 (N_14156,N_12224,N_10468);
and U14157 (N_14157,N_11953,N_10315);
xnor U14158 (N_14158,N_10406,N_12040);
nand U14159 (N_14159,N_11490,N_11750);
and U14160 (N_14160,N_10293,N_12035);
or U14161 (N_14161,N_10432,N_11700);
and U14162 (N_14162,N_10293,N_11492);
xor U14163 (N_14163,N_10102,N_10437);
nor U14164 (N_14164,N_10593,N_10734);
xor U14165 (N_14165,N_10619,N_10510);
or U14166 (N_14166,N_10089,N_11006);
and U14167 (N_14167,N_11295,N_10063);
or U14168 (N_14168,N_10092,N_11920);
or U14169 (N_14169,N_11062,N_12247);
xnor U14170 (N_14170,N_10117,N_10865);
xor U14171 (N_14171,N_11459,N_12377);
nand U14172 (N_14172,N_12346,N_10675);
nor U14173 (N_14173,N_11237,N_11996);
nand U14174 (N_14174,N_10557,N_11634);
or U14175 (N_14175,N_10418,N_10517);
xor U14176 (N_14176,N_12471,N_10683);
nand U14177 (N_14177,N_12250,N_11542);
xnor U14178 (N_14178,N_10375,N_10637);
and U14179 (N_14179,N_10092,N_12023);
xor U14180 (N_14180,N_11124,N_11411);
xnor U14181 (N_14181,N_10396,N_10670);
or U14182 (N_14182,N_10115,N_10975);
or U14183 (N_14183,N_10892,N_11837);
nor U14184 (N_14184,N_11481,N_11534);
or U14185 (N_14185,N_12487,N_12140);
xor U14186 (N_14186,N_10778,N_12033);
nand U14187 (N_14187,N_10027,N_10260);
and U14188 (N_14188,N_12493,N_11714);
nand U14189 (N_14189,N_10043,N_11789);
nor U14190 (N_14190,N_10503,N_11311);
and U14191 (N_14191,N_11685,N_12071);
nand U14192 (N_14192,N_11117,N_10812);
nand U14193 (N_14193,N_10127,N_11488);
nand U14194 (N_14194,N_12361,N_10147);
or U14195 (N_14195,N_11540,N_11499);
nor U14196 (N_14196,N_10527,N_10028);
or U14197 (N_14197,N_11407,N_10841);
and U14198 (N_14198,N_11508,N_10804);
or U14199 (N_14199,N_10309,N_11983);
xor U14200 (N_14200,N_10364,N_11085);
xor U14201 (N_14201,N_10211,N_11995);
xor U14202 (N_14202,N_12031,N_12005);
xnor U14203 (N_14203,N_11950,N_11423);
nor U14204 (N_14204,N_11887,N_10560);
or U14205 (N_14205,N_10335,N_11778);
nand U14206 (N_14206,N_11825,N_12188);
and U14207 (N_14207,N_11938,N_12397);
nor U14208 (N_14208,N_12373,N_10662);
nand U14209 (N_14209,N_11372,N_10449);
or U14210 (N_14210,N_11299,N_10630);
xor U14211 (N_14211,N_10715,N_10383);
xnor U14212 (N_14212,N_11013,N_12241);
nand U14213 (N_14213,N_10614,N_10707);
nand U14214 (N_14214,N_10609,N_11893);
nor U14215 (N_14215,N_11219,N_10545);
or U14216 (N_14216,N_11876,N_10230);
or U14217 (N_14217,N_11182,N_10538);
or U14218 (N_14218,N_11579,N_10745);
or U14219 (N_14219,N_11533,N_10092);
and U14220 (N_14220,N_12380,N_11523);
nor U14221 (N_14221,N_10099,N_10682);
xnor U14222 (N_14222,N_11430,N_11795);
or U14223 (N_14223,N_10897,N_10201);
nor U14224 (N_14224,N_10429,N_10420);
nor U14225 (N_14225,N_12233,N_12219);
xnor U14226 (N_14226,N_10146,N_10708);
xor U14227 (N_14227,N_10156,N_11815);
nand U14228 (N_14228,N_11244,N_11874);
and U14229 (N_14229,N_12296,N_10485);
nand U14230 (N_14230,N_10186,N_11086);
nand U14231 (N_14231,N_11247,N_11693);
nor U14232 (N_14232,N_10825,N_11905);
nor U14233 (N_14233,N_11877,N_10484);
and U14234 (N_14234,N_11268,N_11983);
nand U14235 (N_14235,N_12087,N_10858);
and U14236 (N_14236,N_11210,N_11713);
or U14237 (N_14237,N_11750,N_11340);
nor U14238 (N_14238,N_12195,N_10885);
and U14239 (N_14239,N_12188,N_10059);
nand U14240 (N_14240,N_10826,N_11257);
nand U14241 (N_14241,N_10984,N_12060);
or U14242 (N_14242,N_11547,N_10590);
and U14243 (N_14243,N_10570,N_12076);
nor U14244 (N_14244,N_11238,N_10587);
nor U14245 (N_14245,N_10673,N_12371);
nand U14246 (N_14246,N_10764,N_11543);
or U14247 (N_14247,N_10446,N_11866);
or U14248 (N_14248,N_10868,N_11366);
or U14249 (N_14249,N_11497,N_10410);
nor U14250 (N_14250,N_11227,N_11865);
nand U14251 (N_14251,N_10902,N_11286);
or U14252 (N_14252,N_10798,N_12035);
nor U14253 (N_14253,N_11105,N_10917);
nand U14254 (N_14254,N_12308,N_10837);
or U14255 (N_14255,N_10801,N_11852);
xor U14256 (N_14256,N_11399,N_10664);
or U14257 (N_14257,N_11491,N_10993);
nand U14258 (N_14258,N_10774,N_11656);
nor U14259 (N_14259,N_11524,N_10993);
xnor U14260 (N_14260,N_10238,N_11550);
xnor U14261 (N_14261,N_11983,N_11388);
nor U14262 (N_14262,N_11130,N_11686);
nand U14263 (N_14263,N_10468,N_11486);
xor U14264 (N_14264,N_12294,N_10240);
or U14265 (N_14265,N_10423,N_10779);
xor U14266 (N_14266,N_11599,N_10587);
nand U14267 (N_14267,N_12092,N_10794);
nor U14268 (N_14268,N_11429,N_10683);
nor U14269 (N_14269,N_10976,N_11040);
or U14270 (N_14270,N_11506,N_12301);
and U14271 (N_14271,N_12491,N_10181);
or U14272 (N_14272,N_11328,N_10687);
and U14273 (N_14273,N_11027,N_10798);
or U14274 (N_14274,N_12224,N_11947);
xor U14275 (N_14275,N_12240,N_11038);
xnor U14276 (N_14276,N_12292,N_11049);
nor U14277 (N_14277,N_12355,N_12157);
or U14278 (N_14278,N_11669,N_11433);
xor U14279 (N_14279,N_11996,N_12313);
and U14280 (N_14280,N_10050,N_11683);
nor U14281 (N_14281,N_12450,N_10115);
or U14282 (N_14282,N_10248,N_11988);
xor U14283 (N_14283,N_11669,N_10251);
nand U14284 (N_14284,N_12361,N_11341);
nor U14285 (N_14285,N_11287,N_12235);
nand U14286 (N_14286,N_11191,N_12119);
nand U14287 (N_14287,N_10827,N_11310);
and U14288 (N_14288,N_12162,N_12390);
or U14289 (N_14289,N_11066,N_10565);
or U14290 (N_14290,N_10436,N_11623);
nand U14291 (N_14291,N_12345,N_11281);
xor U14292 (N_14292,N_10003,N_11512);
and U14293 (N_14293,N_10215,N_12318);
and U14294 (N_14294,N_10250,N_10418);
or U14295 (N_14295,N_11792,N_11081);
and U14296 (N_14296,N_12252,N_10077);
xor U14297 (N_14297,N_12262,N_12267);
or U14298 (N_14298,N_11049,N_11962);
and U14299 (N_14299,N_11366,N_10685);
xor U14300 (N_14300,N_10407,N_10292);
or U14301 (N_14301,N_11370,N_12109);
or U14302 (N_14302,N_10274,N_12339);
and U14303 (N_14303,N_10787,N_10898);
nor U14304 (N_14304,N_10959,N_11349);
or U14305 (N_14305,N_10636,N_10825);
nor U14306 (N_14306,N_10476,N_12330);
nor U14307 (N_14307,N_12097,N_10150);
or U14308 (N_14308,N_10411,N_12431);
or U14309 (N_14309,N_10079,N_11046);
and U14310 (N_14310,N_10932,N_11373);
xor U14311 (N_14311,N_12277,N_11858);
nand U14312 (N_14312,N_10652,N_11050);
nor U14313 (N_14313,N_11784,N_11160);
nor U14314 (N_14314,N_10414,N_11260);
xor U14315 (N_14315,N_12104,N_10110);
nand U14316 (N_14316,N_11740,N_11107);
and U14317 (N_14317,N_12472,N_10988);
or U14318 (N_14318,N_10886,N_11180);
nand U14319 (N_14319,N_11350,N_10012);
and U14320 (N_14320,N_11166,N_12358);
and U14321 (N_14321,N_10787,N_11099);
or U14322 (N_14322,N_10888,N_10395);
or U14323 (N_14323,N_10733,N_11650);
nand U14324 (N_14324,N_11416,N_12294);
or U14325 (N_14325,N_10781,N_12360);
and U14326 (N_14326,N_11070,N_12445);
or U14327 (N_14327,N_11455,N_10445);
nor U14328 (N_14328,N_11162,N_11671);
nor U14329 (N_14329,N_12440,N_12144);
xor U14330 (N_14330,N_10113,N_10016);
nor U14331 (N_14331,N_10871,N_12094);
and U14332 (N_14332,N_10497,N_11473);
or U14333 (N_14333,N_11423,N_11372);
xor U14334 (N_14334,N_10191,N_12370);
nand U14335 (N_14335,N_12057,N_11847);
nor U14336 (N_14336,N_11035,N_10981);
nand U14337 (N_14337,N_11491,N_12442);
or U14338 (N_14338,N_10200,N_10396);
or U14339 (N_14339,N_10640,N_11457);
xnor U14340 (N_14340,N_11420,N_12171);
nand U14341 (N_14341,N_10324,N_12498);
nand U14342 (N_14342,N_10439,N_10055);
nor U14343 (N_14343,N_11782,N_10242);
or U14344 (N_14344,N_11484,N_11055);
xor U14345 (N_14345,N_10053,N_12327);
xnor U14346 (N_14346,N_10132,N_11835);
and U14347 (N_14347,N_11400,N_10357);
or U14348 (N_14348,N_10682,N_11242);
xor U14349 (N_14349,N_11011,N_11091);
xnor U14350 (N_14350,N_10440,N_10906);
nand U14351 (N_14351,N_12042,N_10835);
nand U14352 (N_14352,N_11743,N_11198);
or U14353 (N_14353,N_11911,N_10468);
or U14354 (N_14354,N_10247,N_10798);
nand U14355 (N_14355,N_10786,N_12256);
and U14356 (N_14356,N_10255,N_12308);
and U14357 (N_14357,N_12010,N_10279);
nand U14358 (N_14358,N_10452,N_12234);
and U14359 (N_14359,N_10170,N_10544);
and U14360 (N_14360,N_10226,N_12137);
nor U14361 (N_14361,N_11545,N_11284);
nor U14362 (N_14362,N_11656,N_10659);
or U14363 (N_14363,N_11723,N_11862);
nand U14364 (N_14364,N_11563,N_12334);
and U14365 (N_14365,N_10454,N_11020);
xnor U14366 (N_14366,N_11208,N_11185);
and U14367 (N_14367,N_11668,N_11715);
and U14368 (N_14368,N_10348,N_10129);
or U14369 (N_14369,N_11134,N_10306);
nor U14370 (N_14370,N_11773,N_10895);
and U14371 (N_14371,N_11522,N_11355);
xor U14372 (N_14372,N_10103,N_11688);
xor U14373 (N_14373,N_10348,N_10122);
and U14374 (N_14374,N_10512,N_10832);
and U14375 (N_14375,N_12017,N_11446);
or U14376 (N_14376,N_11844,N_10922);
or U14377 (N_14377,N_11650,N_11227);
and U14378 (N_14378,N_12213,N_11302);
or U14379 (N_14379,N_11569,N_12259);
or U14380 (N_14380,N_11124,N_12321);
xnor U14381 (N_14381,N_10300,N_12121);
and U14382 (N_14382,N_11024,N_12376);
or U14383 (N_14383,N_10421,N_11176);
and U14384 (N_14384,N_10936,N_10800);
xor U14385 (N_14385,N_11232,N_12003);
xnor U14386 (N_14386,N_10267,N_10625);
and U14387 (N_14387,N_10843,N_10479);
nor U14388 (N_14388,N_10112,N_11871);
nand U14389 (N_14389,N_11741,N_11659);
xnor U14390 (N_14390,N_10821,N_12488);
nand U14391 (N_14391,N_10582,N_11361);
xor U14392 (N_14392,N_12121,N_10263);
or U14393 (N_14393,N_10093,N_10525);
nor U14394 (N_14394,N_11307,N_10906);
or U14395 (N_14395,N_10947,N_10452);
nor U14396 (N_14396,N_10229,N_11650);
or U14397 (N_14397,N_11374,N_11008);
nor U14398 (N_14398,N_12000,N_10040);
or U14399 (N_14399,N_10763,N_10594);
nand U14400 (N_14400,N_11471,N_11413);
xor U14401 (N_14401,N_11428,N_11215);
xnor U14402 (N_14402,N_11891,N_12354);
nor U14403 (N_14403,N_11467,N_10707);
xor U14404 (N_14404,N_12217,N_10752);
or U14405 (N_14405,N_11194,N_10867);
or U14406 (N_14406,N_11816,N_10424);
nand U14407 (N_14407,N_10058,N_11191);
nor U14408 (N_14408,N_12307,N_12499);
or U14409 (N_14409,N_11075,N_11551);
xnor U14410 (N_14410,N_10187,N_11628);
and U14411 (N_14411,N_11133,N_10679);
and U14412 (N_14412,N_11415,N_10054);
nand U14413 (N_14413,N_10019,N_11372);
nor U14414 (N_14414,N_10604,N_12208);
nand U14415 (N_14415,N_11574,N_10502);
nor U14416 (N_14416,N_10092,N_10815);
xnor U14417 (N_14417,N_11406,N_10825);
nor U14418 (N_14418,N_10781,N_10902);
nand U14419 (N_14419,N_12173,N_10747);
nor U14420 (N_14420,N_12370,N_11427);
nor U14421 (N_14421,N_10022,N_10313);
xnor U14422 (N_14422,N_11742,N_11551);
and U14423 (N_14423,N_10438,N_12076);
or U14424 (N_14424,N_10184,N_12284);
xnor U14425 (N_14425,N_10483,N_11205);
or U14426 (N_14426,N_11796,N_11320);
xor U14427 (N_14427,N_10283,N_11551);
nor U14428 (N_14428,N_12032,N_11544);
nand U14429 (N_14429,N_11069,N_11056);
and U14430 (N_14430,N_12410,N_11541);
or U14431 (N_14431,N_10877,N_12087);
and U14432 (N_14432,N_10325,N_11340);
xnor U14433 (N_14433,N_10076,N_10336);
xor U14434 (N_14434,N_10031,N_12366);
xnor U14435 (N_14435,N_11744,N_11827);
and U14436 (N_14436,N_11406,N_11115);
nand U14437 (N_14437,N_10716,N_12101);
or U14438 (N_14438,N_10623,N_11161);
nor U14439 (N_14439,N_12138,N_11277);
or U14440 (N_14440,N_10848,N_12354);
or U14441 (N_14441,N_10503,N_10146);
xor U14442 (N_14442,N_11724,N_11423);
or U14443 (N_14443,N_12408,N_11663);
or U14444 (N_14444,N_10333,N_11741);
and U14445 (N_14445,N_10810,N_10670);
xnor U14446 (N_14446,N_12037,N_12410);
nand U14447 (N_14447,N_10482,N_11539);
nand U14448 (N_14448,N_10697,N_10663);
or U14449 (N_14449,N_12331,N_12251);
nor U14450 (N_14450,N_10150,N_11810);
nor U14451 (N_14451,N_12230,N_10142);
nor U14452 (N_14452,N_12475,N_10164);
nand U14453 (N_14453,N_11307,N_10653);
and U14454 (N_14454,N_12223,N_11544);
nand U14455 (N_14455,N_10265,N_12129);
nor U14456 (N_14456,N_12335,N_10214);
and U14457 (N_14457,N_12261,N_11937);
or U14458 (N_14458,N_10713,N_10539);
and U14459 (N_14459,N_12464,N_11092);
xnor U14460 (N_14460,N_10650,N_12345);
nor U14461 (N_14461,N_12309,N_11971);
and U14462 (N_14462,N_10653,N_10656);
xor U14463 (N_14463,N_11333,N_12083);
and U14464 (N_14464,N_10214,N_11124);
and U14465 (N_14465,N_10781,N_11576);
nand U14466 (N_14466,N_10492,N_10187);
nand U14467 (N_14467,N_10344,N_11842);
nand U14468 (N_14468,N_10222,N_12341);
and U14469 (N_14469,N_11527,N_12069);
and U14470 (N_14470,N_11363,N_12294);
and U14471 (N_14471,N_10626,N_11774);
and U14472 (N_14472,N_10731,N_11299);
xnor U14473 (N_14473,N_11689,N_10107);
nand U14474 (N_14474,N_11476,N_11153);
nor U14475 (N_14475,N_11518,N_12089);
nand U14476 (N_14476,N_12356,N_10952);
or U14477 (N_14477,N_11067,N_12479);
or U14478 (N_14478,N_10555,N_12063);
nor U14479 (N_14479,N_10714,N_10644);
or U14480 (N_14480,N_12368,N_11549);
nor U14481 (N_14481,N_12317,N_10427);
xor U14482 (N_14482,N_11723,N_11635);
nor U14483 (N_14483,N_11812,N_10179);
nor U14484 (N_14484,N_10973,N_11633);
or U14485 (N_14485,N_12231,N_11471);
or U14486 (N_14486,N_11514,N_12336);
or U14487 (N_14487,N_12076,N_12457);
or U14488 (N_14488,N_11278,N_11948);
nand U14489 (N_14489,N_10091,N_11728);
nor U14490 (N_14490,N_11487,N_11049);
xnor U14491 (N_14491,N_11176,N_11537);
nor U14492 (N_14492,N_10303,N_11333);
nand U14493 (N_14493,N_11243,N_10961);
nor U14494 (N_14494,N_11696,N_11555);
and U14495 (N_14495,N_11479,N_11167);
xor U14496 (N_14496,N_12331,N_10654);
nor U14497 (N_14497,N_12244,N_11211);
nor U14498 (N_14498,N_11365,N_10920);
or U14499 (N_14499,N_11993,N_10006);
nor U14500 (N_14500,N_11240,N_11115);
xor U14501 (N_14501,N_11355,N_10063);
xnor U14502 (N_14502,N_10224,N_10778);
or U14503 (N_14503,N_11270,N_10834);
and U14504 (N_14504,N_10089,N_11740);
nor U14505 (N_14505,N_10446,N_12171);
or U14506 (N_14506,N_11278,N_10909);
or U14507 (N_14507,N_10526,N_10867);
xor U14508 (N_14508,N_10302,N_11887);
or U14509 (N_14509,N_10598,N_11663);
xor U14510 (N_14510,N_11658,N_11622);
or U14511 (N_14511,N_10370,N_11924);
nand U14512 (N_14512,N_11265,N_11679);
xor U14513 (N_14513,N_12208,N_12384);
xor U14514 (N_14514,N_10225,N_11001);
nand U14515 (N_14515,N_11487,N_10756);
xnor U14516 (N_14516,N_10644,N_10948);
nand U14517 (N_14517,N_10452,N_10230);
or U14518 (N_14518,N_12077,N_11288);
and U14519 (N_14519,N_11687,N_10984);
xnor U14520 (N_14520,N_10315,N_12021);
xnor U14521 (N_14521,N_10187,N_12174);
and U14522 (N_14522,N_12371,N_10156);
xnor U14523 (N_14523,N_11623,N_11016);
or U14524 (N_14524,N_10212,N_10056);
nand U14525 (N_14525,N_11364,N_11379);
nor U14526 (N_14526,N_12273,N_11988);
xnor U14527 (N_14527,N_10471,N_10623);
nand U14528 (N_14528,N_10798,N_12367);
nand U14529 (N_14529,N_11357,N_11576);
and U14530 (N_14530,N_10493,N_11769);
nand U14531 (N_14531,N_10327,N_11346);
nand U14532 (N_14532,N_10627,N_11767);
and U14533 (N_14533,N_10619,N_10411);
or U14534 (N_14534,N_10839,N_10289);
and U14535 (N_14535,N_11264,N_11814);
xor U14536 (N_14536,N_10728,N_10506);
and U14537 (N_14537,N_11837,N_11758);
nand U14538 (N_14538,N_12028,N_11601);
or U14539 (N_14539,N_10572,N_10149);
nand U14540 (N_14540,N_11959,N_11621);
xnor U14541 (N_14541,N_11671,N_11981);
xor U14542 (N_14542,N_10700,N_11929);
nor U14543 (N_14543,N_11039,N_12047);
xor U14544 (N_14544,N_10357,N_11088);
nor U14545 (N_14545,N_11233,N_11645);
nand U14546 (N_14546,N_12127,N_11604);
and U14547 (N_14547,N_10498,N_10144);
xor U14548 (N_14548,N_11328,N_10540);
nand U14549 (N_14549,N_11135,N_11361);
or U14550 (N_14550,N_10271,N_11135);
or U14551 (N_14551,N_12161,N_10473);
and U14552 (N_14552,N_10425,N_11538);
and U14553 (N_14553,N_11180,N_11979);
nor U14554 (N_14554,N_10005,N_11791);
nand U14555 (N_14555,N_10658,N_10572);
and U14556 (N_14556,N_10200,N_11313);
nor U14557 (N_14557,N_11421,N_10151);
and U14558 (N_14558,N_10808,N_11371);
nor U14559 (N_14559,N_11437,N_12487);
or U14560 (N_14560,N_10664,N_11200);
and U14561 (N_14561,N_11224,N_12293);
xor U14562 (N_14562,N_10746,N_10696);
nor U14563 (N_14563,N_12413,N_11083);
nor U14564 (N_14564,N_11042,N_11523);
and U14565 (N_14565,N_11886,N_10121);
nor U14566 (N_14566,N_12449,N_11652);
and U14567 (N_14567,N_12416,N_11177);
nand U14568 (N_14568,N_10246,N_11072);
nand U14569 (N_14569,N_11532,N_11127);
and U14570 (N_14570,N_12256,N_11916);
xor U14571 (N_14571,N_10134,N_11420);
xnor U14572 (N_14572,N_10930,N_11522);
nand U14573 (N_14573,N_11409,N_11935);
and U14574 (N_14574,N_11958,N_11629);
nor U14575 (N_14575,N_12233,N_11573);
nor U14576 (N_14576,N_10314,N_10354);
and U14577 (N_14577,N_10356,N_12137);
or U14578 (N_14578,N_10943,N_10652);
nor U14579 (N_14579,N_11174,N_11401);
xor U14580 (N_14580,N_10234,N_10859);
and U14581 (N_14581,N_12451,N_12092);
xnor U14582 (N_14582,N_10506,N_12094);
nor U14583 (N_14583,N_12130,N_12157);
nand U14584 (N_14584,N_10121,N_11792);
nor U14585 (N_14585,N_10441,N_10920);
xnor U14586 (N_14586,N_11525,N_10449);
or U14587 (N_14587,N_12143,N_12328);
and U14588 (N_14588,N_11526,N_10066);
and U14589 (N_14589,N_10084,N_12401);
or U14590 (N_14590,N_11273,N_10890);
or U14591 (N_14591,N_11065,N_11596);
xor U14592 (N_14592,N_10478,N_11331);
nor U14593 (N_14593,N_12253,N_10225);
and U14594 (N_14594,N_12036,N_11032);
xnor U14595 (N_14595,N_11038,N_11413);
nor U14596 (N_14596,N_11177,N_11241);
nand U14597 (N_14597,N_10159,N_10588);
nand U14598 (N_14598,N_11705,N_10393);
nand U14599 (N_14599,N_11628,N_11002);
nor U14600 (N_14600,N_11243,N_12246);
and U14601 (N_14601,N_11161,N_11977);
or U14602 (N_14602,N_11312,N_10272);
and U14603 (N_14603,N_11802,N_11204);
or U14604 (N_14604,N_10594,N_10852);
nand U14605 (N_14605,N_10736,N_12165);
nand U14606 (N_14606,N_11369,N_10469);
nand U14607 (N_14607,N_12236,N_11565);
or U14608 (N_14608,N_10327,N_11648);
xnor U14609 (N_14609,N_11742,N_11770);
nor U14610 (N_14610,N_10789,N_12422);
xnor U14611 (N_14611,N_11749,N_10275);
nand U14612 (N_14612,N_11707,N_11425);
and U14613 (N_14613,N_11892,N_11785);
and U14614 (N_14614,N_11463,N_10664);
nand U14615 (N_14615,N_11323,N_10779);
nor U14616 (N_14616,N_10773,N_11237);
xnor U14617 (N_14617,N_11405,N_10842);
nor U14618 (N_14618,N_12178,N_10115);
nor U14619 (N_14619,N_10842,N_11408);
and U14620 (N_14620,N_12224,N_10466);
nor U14621 (N_14621,N_10068,N_10589);
nor U14622 (N_14622,N_10891,N_10384);
xnor U14623 (N_14623,N_10275,N_10110);
or U14624 (N_14624,N_10225,N_11328);
or U14625 (N_14625,N_11027,N_12425);
or U14626 (N_14626,N_11661,N_10359);
and U14627 (N_14627,N_11484,N_10616);
nor U14628 (N_14628,N_11286,N_12062);
or U14629 (N_14629,N_11908,N_11233);
nor U14630 (N_14630,N_12295,N_12333);
nand U14631 (N_14631,N_10541,N_11581);
nand U14632 (N_14632,N_12041,N_10397);
nand U14633 (N_14633,N_11160,N_12490);
nor U14634 (N_14634,N_11871,N_10326);
nand U14635 (N_14635,N_12371,N_12432);
nand U14636 (N_14636,N_10330,N_11069);
nor U14637 (N_14637,N_10484,N_11168);
xnor U14638 (N_14638,N_12240,N_11600);
and U14639 (N_14639,N_11133,N_10014);
nor U14640 (N_14640,N_11231,N_10930);
or U14641 (N_14641,N_10802,N_10542);
or U14642 (N_14642,N_11667,N_11099);
xor U14643 (N_14643,N_11176,N_10642);
nor U14644 (N_14644,N_12107,N_10333);
xor U14645 (N_14645,N_11184,N_12246);
nor U14646 (N_14646,N_10691,N_11265);
xnor U14647 (N_14647,N_12424,N_11489);
and U14648 (N_14648,N_11467,N_11672);
nor U14649 (N_14649,N_10682,N_10958);
or U14650 (N_14650,N_12146,N_12095);
nand U14651 (N_14651,N_11123,N_11221);
or U14652 (N_14652,N_10455,N_11496);
or U14653 (N_14653,N_10664,N_10997);
nor U14654 (N_14654,N_11282,N_11418);
or U14655 (N_14655,N_10786,N_11187);
or U14656 (N_14656,N_11361,N_10103);
xor U14657 (N_14657,N_11965,N_11550);
and U14658 (N_14658,N_11286,N_12350);
and U14659 (N_14659,N_10305,N_10592);
xnor U14660 (N_14660,N_12164,N_11457);
and U14661 (N_14661,N_10707,N_10738);
xor U14662 (N_14662,N_11420,N_11312);
xnor U14663 (N_14663,N_10673,N_12476);
and U14664 (N_14664,N_11452,N_10478);
and U14665 (N_14665,N_11179,N_10002);
nor U14666 (N_14666,N_11006,N_11699);
or U14667 (N_14667,N_12251,N_10852);
xnor U14668 (N_14668,N_10405,N_10102);
or U14669 (N_14669,N_10872,N_12015);
and U14670 (N_14670,N_11737,N_12012);
and U14671 (N_14671,N_12406,N_10653);
xnor U14672 (N_14672,N_11152,N_12015);
xor U14673 (N_14673,N_12247,N_10437);
nor U14674 (N_14674,N_12290,N_11267);
and U14675 (N_14675,N_11593,N_11018);
or U14676 (N_14676,N_10363,N_12410);
or U14677 (N_14677,N_11200,N_12314);
xnor U14678 (N_14678,N_10323,N_11399);
nand U14679 (N_14679,N_10535,N_10439);
xor U14680 (N_14680,N_11926,N_10403);
xor U14681 (N_14681,N_12043,N_11124);
nor U14682 (N_14682,N_12116,N_12287);
xor U14683 (N_14683,N_10050,N_11828);
and U14684 (N_14684,N_10628,N_10421);
and U14685 (N_14685,N_12393,N_12403);
nand U14686 (N_14686,N_10906,N_10662);
nor U14687 (N_14687,N_10852,N_10453);
and U14688 (N_14688,N_12300,N_10824);
and U14689 (N_14689,N_10443,N_12056);
nor U14690 (N_14690,N_10685,N_12137);
or U14691 (N_14691,N_12093,N_12049);
and U14692 (N_14692,N_10766,N_11291);
and U14693 (N_14693,N_12139,N_12464);
xnor U14694 (N_14694,N_11066,N_11664);
and U14695 (N_14695,N_11701,N_11579);
nand U14696 (N_14696,N_12406,N_12012);
and U14697 (N_14697,N_11499,N_11927);
and U14698 (N_14698,N_10612,N_10616);
xor U14699 (N_14699,N_12022,N_12069);
xor U14700 (N_14700,N_12019,N_11196);
and U14701 (N_14701,N_11518,N_11939);
nor U14702 (N_14702,N_10245,N_11069);
or U14703 (N_14703,N_10879,N_12029);
nor U14704 (N_14704,N_12319,N_11410);
nand U14705 (N_14705,N_11593,N_11515);
and U14706 (N_14706,N_11395,N_11473);
nor U14707 (N_14707,N_10553,N_12126);
and U14708 (N_14708,N_11698,N_11133);
or U14709 (N_14709,N_10449,N_10143);
xnor U14710 (N_14710,N_11851,N_10538);
and U14711 (N_14711,N_10373,N_11281);
nor U14712 (N_14712,N_12366,N_12160);
or U14713 (N_14713,N_12033,N_12177);
xnor U14714 (N_14714,N_11043,N_12366);
or U14715 (N_14715,N_10631,N_12196);
or U14716 (N_14716,N_11226,N_10366);
xnor U14717 (N_14717,N_11355,N_11364);
nand U14718 (N_14718,N_10449,N_12395);
nand U14719 (N_14719,N_10538,N_11889);
nand U14720 (N_14720,N_10945,N_10488);
and U14721 (N_14721,N_10024,N_10515);
or U14722 (N_14722,N_10539,N_11872);
nand U14723 (N_14723,N_10011,N_11622);
and U14724 (N_14724,N_11729,N_10830);
or U14725 (N_14725,N_10258,N_11725);
nor U14726 (N_14726,N_12087,N_12439);
nor U14727 (N_14727,N_10844,N_11956);
nor U14728 (N_14728,N_11670,N_11839);
nor U14729 (N_14729,N_11269,N_11400);
or U14730 (N_14730,N_11520,N_10753);
nor U14731 (N_14731,N_11440,N_12030);
or U14732 (N_14732,N_10506,N_11398);
xnor U14733 (N_14733,N_10929,N_12322);
and U14734 (N_14734,N_10582,N_10251);
xor U14735 (N_14735,N_10929,N_11175);
or U14736 (N_14736,N_10975,N_10092);
nand U14737 (N_14737,N_10606,N_10905);
or U14738 (N_14738,N_10626,N_10370);
and U14739 (N_14739,N_11736,N_10022);
nor U14740 (N_14740,N_12065,N_10257);
or U14741 (N_14741,N_10339,N_10209);
or U14742 (N_14742,N_11102,N_10821);
xor U14743 (N_14743,N_11140,N_10280);
xor U14744 (N_14744,N_11968,N_10970);
xnor U14745 (N_14745,N_10092,N_11152);
nor U14746 (N_14746,N_11813,N_11561);
xor U14747 (N_14747,N_10222,N_11473);
nor U14748 (N_14748,N_11820,N_12198);
or U14749 (N_14749,N_11400,N_12002);
xor U14750 (N_14750,N_11312,N_11848);
xnor U14751 (N_14751,N_11725,N_11831);
or U14752 (N_14752,N_10337,N_11498);
nand U14753 (N_14753,N_12389,N_10785);
nor U14754 (N_14754,N_12442,N_11173);
xor U14755 (N_14755,N_12134,N_12027);
or U14756 (N_14756,N_10878,N_10016);
and U14757 (N_14757,N_10831,N_12336);
nor U14758 (N_14758,N_10281,N_11820);
and U14759 (N_14759,N_11991,N_11356);
or U14760 (N_14760,N_11547,N_12445);
nand U14761 (N_14761,N_10028,N_11514);
or U14762 (N_14762,N_11775,N_10234);
nand U14763 (N_14763,N_10988,N_12011);
and U14764 (N_14764,N_11493,N_10703);
and U14765 (N_14765,N_10039,N_10438);
nor U14766 (N_14766,N_10603,N_10850);
nand U14767 (N_14767,N_11694,N_11329);
nand U14768 (N_14768,N_11737,N_10110);
nor U14769 (N_14769,N_12363,N_10862);
or U14770 (N_14770,N_12259,N_10904);
xnor U14771 (N_14771,N_10392,N_11826);
xnor U14772 (N_14772,N_11523,N_10103);
or U14773 (N_14773,N_11253,N_10349);
and U14774 (N_14774,N_11468,N_11282);
nor U14775 (N_14775,N_12174,N_10273);
nand U14776 (N_14776,N_10085,N_12141);
nand U14777 (N_14777,N_11239,N_10939);
and U14778 (N_14778,N_11476,N_11009);
nor U14779 (N_14779,N_11268,N_12494);
or U14780 (N_14780,N_11533,N_10158);
nor U14781 (N_14781,N_12013,N_11618);
nand U14782 (N_14782,N_11082,N_11548);
and U14783 (N_14783,N_11534,N_11711);
and U14784 (N_14784,N_10934,N_10630);
nand U14785 (N_14785,N_11141,N_10811);
xor U14786 (N_14786,N_11536,N_11198);
xnor U14787 (N_14787,N_11469,N_12302);
nor U14788 (N_14788,N_10086,N_11378);
nor U14789 (N_14789,N_11234,N_11786);
or U14790 (N_14790,N_12162,N_12271);
nand U14791 (N_14791,N_10495,N_11294);
xnor U14792 (N_14792,N_11543,N_10217);
nor U14793 (N_14793,N_11688,N_12131);
nor U14794 (N_14794,N_11284,N_10198);
nand U14795 (N_14795,N_10997,N_11005);
nor U14796 (N_14796,N_11864,N_11301);
or U14797 (N_14797,N_12365,N_10907);
xor U14798 (N_14798,N_11919,N_10391);
and U14799 (N_14799,N_11206,N_11900);
and U14800 (N_14800,N_11493,N_12304);
nor U14801 (N_14801,N_10131,N_11844);
and U14802 (N_14802,N_12390,N_10953);
nand U14803 (N_14803,N_10130,N_12237);
xnor U14804 (N_14804,N_11714,N_11450);
nor U14805 (N_14805,N_11351,N_10076);
nor U14806 (N_14806,N_10572,N_10301);
or U14807 (N_14807,N_11933,N_12251);
xnor U14808 (N_14808,N_11756,N_10919);
and U14809 (N_14809,N_11304,N_12439);
and U14810 (N_14810,N_12470,N_10639);
nor U14811 (N_14811,N_12455,N_11630);
or U14812 (N_14812,N_10001,N_10040);
xnor U14813 (N_14813,N_11158,N_11938);
nor U14814 (N_14814,N_11116,N_11640);
or U14815 (N_14815,N_12085,N_10032);
nand U14816 (N_14816,N_10257,N_10180);
or U14817 (N_14817,N_10570,N_10734);
nor U14818 (N_14818,N_11703,N_12061);
xor U14819 (N_14819,N_10309,N_11722);
nand U14820 (N_14820,N_12193,N_11356);
nor U14821 (N_14821,N_10054,N_10531);
nand U14822 (N_14822,N_11698,N_10576);
nand U14823 (N_14823,N_12435,N_11109);
and U14824 (N_14824,N_10417,N_10812);
and U14825 (N_14825,N_11500,N_11445);
xor U14826 (N_14826,N_10937,N_10226);
nand U14827 (N_14827,N_11662,N_10300);
or U14828 (N_14828,N_10769,N_11998);
nor U14829 (N_14829,N_10929,N_11302);
or U14830 (N_14830,N_12463,N_10538);
nor U14831 (N_14831,N_10240,N_10294);
nor U14832 (N_14832,N_11795,N_10565);
or U14833 (N_14833,N_11544,N_12061);
and U14834 (N_14834,N_10920,N_10176);
or U14835 (N_14835,N_11386,N_10329);
and U14836 (N_14836,N_10576,N_10428);
and U14837 (N_14837,N_11430,N_11632);
and U14838 (N_14838,N_11991,N_10986);
nand U14839 (N_14839,N_11845,N_10771);
xor U14840 (N_14840,N_11209,N_10870);
nor U14841 (N_14841,N_10658,N_11001);
and U14842 (N_14842,N_12302,N_12119);
or U14843 (N_14843,N_10117,N_11341);
xnor U14844 (N_14844,N_12491,N_10549);
and U14845 (N_14845,N_10812,N_11670);
nand U14846 (N_14846,N_12339,N_10914);
nand U14847 (N_14847,N_11736,N_10903);
and U14848 (N_14848,N_12319,N_10992);
nand U14849 (N_14849,N_12392,N_11979);
nand U14850 (N_14850,N_10075,N_12229);
and U14851 (N_14851,N_10937,N_10759);
or U14852 (N_14852,N_11321,N_10800);
nand U14853 (N_14853,N_12320,N_11226);
and U14854 (N_14854,N_10033,N_11960);
nor U14855 (N_14855,N_10852,N_11561);
nor U14856 (N_14856,N_10766,N_11505);
and U14857 (N_14857,N_10105,N_11863);
xor U14858 (N_14858,N_10368,N_11393);
or U14859 (N_14859,N_11947,N_12247);
or U14860 (N_14860,N_10514,N_11045);
nand U14861 (N_14861,N_10823,N_11370);
xnor U14862 (N_14862,N_11843,N_12237);
or U14863 (N_14863,N_10924,N_11346);
nor U14864 (N_14864,N_12485,N_10253);
and U14865 (N_14865,N_11987,N_11679);
nor U14866 (N_14866,N_11749,N_10865);
or U14867 (N_14867,N_10835,N_11319);
or U14868 (N_14868,N_11687,N_12308);
and U14869 (N_14869,N_10366,N_12334);
or U14870 (N_14870,N_10603,N_11917);
and U14871 (N_14871,N_11011,N_12187);
xnor U14872 (N_14872,N_10565,N_10308);
and U14873 (N_14873,N_11067,N_12218);
or U14874 (N_14874,N_10770,N_10062);
xor U14875 (N_14875,N_11140,N_11533);
nand U14876 (N_14876,N_12026,N_10693);
or U14877 (N_14877,N_10169,N_11449);
or U14878 (N_14878,N_11498,N_10727);
and U14879 (N_14879,N_11040,N_10879);
xnor U14880 (N_14880,N_11397,N_11941);
xor U14881 (N_14881,N_11476,N_10734);
and U14882 (N_14882,N_10700,N_10503);
nand U14883 (N_14883,N_12058,N_12119);
xor U14884 (N_14884,N_11710,N_10355);
nand U14885 (N_14885,N_10677,N_12189);
or U14886 (N_14886,N_10176,N_10934);
or U14887 (N_14887,N_10924,N_11187);
xnor U14888 (N_14888,N_11230,N_10819);
xnor U14889 (N_14889,N_10529,N_10414);
and U14890 (N_14890,N_11478,N_10015);
nor U14891 (N_14891,N_11960,N_12369);
nor U14892 (N_14892,N_11027,N_12499);
or U14893 (N_14893,N_12232,N_10649);
or U14894 (N_14894,N_11602,N_11927);
nor U14895 (N_14895,N_10332,N_12419);
nand U14896 (N_14896,N_10499,N_11354);
nor U14897 (N_14897,N_10549,N_11744);
xnor U14898 (N_14898,N_11182,N_11253);
or U14899 (N_14899,N_12066,N_11430);
and U14900 (N_14900,N_12382,N_11993);
and U14901 (N_14901,N_12049,N_11495);
and U14902 (N_14902,N_12083,N_10490);
nand U14903 (N_14903,N_12247,N_10503);
nand U14904 (N_14904,N_10270,N_11916);
nand U14905 (N_14905,N_12498,N_10968);
or U14906 (N_14906,N_11971,N_11782);
or U14907 (N_14907,N_10190,N_11352);
nand U14908 (N_14908,N_11988,N_10987);
or U14909 (N_14909,N_11293,N_12281);
nor U14910 (N_14910,N_12286,N_11006);
and U14911 (N_14911,N_11642,N_11253);
and U14912 (N_14912,N_12360,N_11824);
or U14913 (N_14913,N_10416,N_11970);
and U14914 (N_14914,N_11164,N_12148);
and U14915 (N_14915,N_10216,N_11295);
and U14916 (N_14916,N_11353,N_12179);
xnor U14917 (N_14917,N_12274,N_10421);
or U14918 (N_14918,N_10371,N_11233);
or U14919 (N_14919,N_12122,N_12150);
nor U14920 (N_14920,N_11247,N_10237);
nand U14921 (N_14921,N_11712,N_10837);
nor U14922 (N_14922,N_11964,N_10975);
or U14923 (N_14923,N_11296,N_11120);
and U14924 (N_14924,N_10477,N_10580);
nor U14925 (N_14925,N_12163,N_10658);
xnor U14926 (N_14926,N_12229,N_12175);
xnor U14927 (N_14927,N_10418,N_11014);
nor U14928 (N_14928,N_10639,N_10320);
xnor U14929 (N_14929,N_10554,N_10321);
nor U14930 (N_14930,N_11959,N_11770);
xnor U14931 (N_14931,N_10475,N_11781);
nor U14932 (N_14932,N_11284,N_11290);
nand U14933 (N_14933,N_11910,N_11842);
nand U14934 (N_14934,N_12188,N_12009);
nand U14935 (N_14935,N_10347,N_11358);
nand U14936 (N_14936,N_10438,N_12457);
and U14937 (N_14937,N_10475,N_10180);
and U14938 (N_14938,N_11462,N_12339);
xnor U14939 (N_14939,N_12211,N_11811);
nand U14940 (N_14940,N_11752,N_10184);
and U14941 (N_14941,N_11031,N_12114);
nor U14942 (N_14942,N_10139,N_12477);
xnor U14943 (N_14943,N_10421,N_11249);
xor U14944 (N_14944,N_10184,N_11615);
nand U14945 (N_14945,N_11258,N_10903);
xor U14946 (N_14946,N_10164,N_11320);
nor U14947 (N_14947,N_11490,N_10210);
nand U14948 (N_14948,N_11622,N_10422);
and U14949 (N_14949,N_11091,N_10454);
nand U14950 (N_14950,N_10174,N_10340);
xnor U14951 (N_14951,N_12187,N_10291);
xnor U14952 (N_14952,N_10763,N_11855);
xnor U14953 (N_14953,N_12493,N_11572);
xor U14954 (N_14954,N_10394,N_11195);
nand U14955 (N_14955,N_10010,N_10678);
xnor U14956 (N_14956,N_10885,N_12218);
nand U14957 (N_14957,N_11632,N_11839);
xnor U14958 (N_14958,N_11832,N_11731);
xor U14959 (N_14959,N_10569,N_11402);
xor U14960 (N_14960,N_12402,N_11444);
and U14961 (N_14961,N_11801,N_10211);
or U14962 (N_14962,N_12074,N_10930);
and U14963 (N_14963,N_10160,N_10808);
nand U14964 (N_14964,N_10984,N_11422);
and U14965 (N_14965,N_12057,N_10267);
nand U14966 (N_14966,N_11130,N_12370);
and U14967 (N_14967,N_11226,N_10578);
nand U14968 (N_14968,N_11701,N_12176);
nor U14969 (N_14969,N_10625,N_11038);
nor U14970 (N_14970,N_11287,N_10411);
nor U14971 (N_14971,N_10328,N_10844);
or U14972 (N_14972,N_11273,N_11036);
or U14973 (N_14973,N_10276,N_11070);
nand U14974 (N_14974,N_10222,N_10252);
xnor U14975 (N_14975,N_10497,N_10154);
and U14976 (N_14976,N_10428,N_11574);
or U14977 (N_14977,N_11306,N_11571);
or U14978 (N_14978,N_12095,N_10379);
nor U14979 (N_14979,N_12436,N_10366);
nor U14980 (N_14980,N_11649,N_10555);
or U14981 (N_14981,N_11050,N_11691);
xnor U14982 (N_14982,N_12122,N_10584);
nor U14983 (N_14983,N_11269,N_12019);
nor U14984 (N_14984,N_11507,N_12189);
and U14985 (N_14985,N_11179,N_10381);
xor U14986 (N_14986,N_10173,N_10839);
nand U14987 (N_14987,N_10669,N_10692);
and U14988 (N_14988,N_10272,N_10141);
xor U14989 (N_14989,N_10763,N_11657);
xor U14990 (N_14990,N_11982,N_11119);
xnor U14991 (N_14991,N_12480,N_12201);
and U14992 (N_14992,N_10203,N_11996);
and U14993 (N_14993,N_10262,N_10728);
nand U14994 (N_14994,N_12357,N_11290);
nand U14995 (N_14995,N_11676,N_11988);
or U14996 (N_14996,N_10989,N_10496);
and U14997 (N_14997,N_10981,N_10010);
or U14998 (N_14998,N_12046,N_10510);
and U14999 (N_14999,N_12323,N_11384);
or U15000 (N_15000,N_13229,N_12896);
nor U15001 (N_15001,N_14225,N_14911);
nor U15002 (N_15002,N_13387,N_13970);
nor U15003 (N_15003,N_14916,N_14704);
or U15004 (N_15004,N_14637,N_12568);
xnor U15005 (N_15005,N_13655,N_13090);
nand U15006 (N_15006,N_12541,N_13384);
or U15007 (N_15007,N_14381,N_13945);
or U15008 (N_15008,N_12737,N_13890);
xor U15009 (N_15009,N_13081,N_12687);
nand U15010 (N_15010,N_13550,N_14746);
nand U15011 (N_15011,N_14332,N_13809);
and U15012 (N_15012,N_13286,N_13064);
nor U15013 (N_15013,N_13589,N_13623);
nor U15014 (N_15014,N_14183,N_14780);
nor U15015 (N_15015,N_13715,N_14005);
xor U15016 (N_15016,N_14794,N_12834);
nor U15017 (N_15017,N_14923,N_13603);
nor U15018 (N_15018,N_13089,N_12999);
xnor U15019 (N_15019,N_13086,N_13857);
nor U15020 (N_15020,N_12923,N_14173);
and U15021 (N_15021,N_14051,N_13175);
nor U15022 (N_15022,N_14272,N_14833);
or U15023 (N_15023,N_12703,N_14206);
and U15024 (N_15024,N_14847,N_14751);
nor U15025 (N_15025,N_14857,N_12680);
or U15026 (N_15026,N_12612,N_14126);
nor U15027 (N_15027,N_13453,N_13687);
or U15028 (N_15028,N_12567,N_13088);
and U15029 (N_15029,N_13368,N_12935);
nor U15030 (N_15030,N_14514,N_14256);
xnor U15031 (N_15031,N_13129,N_14761);
nor U15032 (N_15032,N_13183,N_12509);
or U15033 (N_15033,N_13518,N_14934);
xor U15034 (N_15034,N_12547,N_14830);
nor U15035 (N_15035,N_13997,N_13803);
nand U15036 (N_15036,N_13959,N_12694);
and U15037 (N_15037,N_12786,N_14157);
or U15038 (N_15038,N_13869,N_12854);
nor U15039 (N_15039,N_12513,N_12552);
and U15040 (N_15040,N_13745,N_14900);
nand U15041 (N_15041,N_14499,N_12977);
nand U15042 (N_15042,N_14523,N_13922);
and U15043 (N_15043,N_14233,N_14975);
or U15044 (N_15044,N_13202,N_12936);
or U15045 (N_15045,N_12549,N_12996);
or U15046 (N_15046,N_14615,N_13549);
nand U15047 (N_15047,N_14583,N_13590);
xor U15048 (N_15048,N_13782,N_12589);
xnor U15049 (N_15049,N_14550,N_13796);
or U15050 (N_15050,N_13271,N_14047);
or U15051 (N_15051,N_14141,N_12898);
xor U15052 (N_15052,N_14049,N_14677);
nor U15053 (N_15053,N_12879,N_14396);
nor U15054 (N_15054,N_13405,N_13801);
and U15055 (N_15055,N_13167,N_13134);
and U15056 (N_15056,N_14928,N_12783);
nor U15057 (N_15057,N_14376,N_14714);
xor U15058 (N_15058,N_12527,N_13901);
or U15059 (N_15059,N_13486,N_13475);
and U15060 (N_15060,N_12553,N_14188);
nor U15061 (N_15061,N_14216,N_14698);
nor U15062 (N_15062,N_14625,N_13921);
xor U15063 (N_15063,N_14007,N_12722);
nand U15064 (N_15064,N_14924,N_14255);
xor U15065 (N_15065,N_12662,N_13818);
nor U15066 (N_15066,N_14706,N_14019);
xor U15067 (N_15067,N_14419,N_14565);
nand U15068 (N_15068,N_12658,N_13893);
nor U15069 (N_15069,N_13908,N_12610);
nand U15070 (N_15070,N_14449,N_14184);
and U15071 (N_15071,N_14506,N_12685);
nand U15072 (N_15072,N_14388,N_13057);
and U15073 (N_15073,N_12798,N_14441);
xnor U15074 (N_15074,N_12821,N_14367);
nor U15075 (N_15075,N_14720,N_13231);
and U15076 (N_15076,N_14628,N_13885);
and U15077 (N_15077,N_12664,N_13833);
nand U15078 (N_15078,N_12802,N_13325);
xnor U15079 (N_15079,N_13932,N_14631);
nor U15080 (N_15080,N_14581,N_13267);
nand U15081 (N_15081,N_13630,N_13858);
xnor U15082 (N_15082,N_14021,N_13353);
or U15083 (N_15083,N_13190,N_12624);
or U15084 (N_15084,N_14164,N_13262);
or U15085 (N_15085,N_14525,N_12913);
xor U15086 (N_15086,N_13751,N_13826);
nand U15087 (N_15087,N_12950,N_14180);
xnor U15088 (N_15088,N_13334,N_14545);
xnor U15089 (N_15089,N_13663,N_12503);
nand U15090 (N_15090,N_13709,N_13701);
or U15091 (N_15091,N_13144,N_13240);
nand U15092 (N_15092,N_13128,N_14518);
or U15093 (N_15093,N_13697,N_14319);
nand U15094 (N_15094,N_13160,N_12533);
and U15095 (N_15095,N_14241,N_12741);
xnor U15096 (N_15096,N_14354,N_14868);
or U15097 (N_15097,N_13537,N_12570);
or U15098 (N_15098,N_14703,N_14351);
and U15099 (N_15099,N_14674,N_13112);
xnor U15100 (N_15100,N_14635,N_14828);
or U15101 (N_15101,N_13258,N_14234);
nand U15102 (N_15102,N_12960,N_14682);
xor U15103 (N_15103,N_14827,N_13422);
nand U15104 (N_15104,N_12794,N_13768);
nand U15105 (N_15105,N_14410,N_14080);
nand U15106 (N_15106,N_12609,N_13142);
nand U15107 (N_15107,N_14754,N_13668);
or U15108 (N_15108,N_12519,N_14789);
and U15109 (N_15109,N_13395,N_14564);
xnor U15110 (N_15110,N_14008,N_13054);
xor U15111 (N_15111,N_14786,N_13487);
nand U15112 (N_15112,N_12908,N_13068);
nor U15113 (N_15113,N_14147,N_14885);
nand U15114 (N_15114,N_13702,N_14987);
nand U15115 (N_15115,N_12683,N_13503);
xnor U15116 (N_15116,N_13980,N_13835);
nand U15117 (N_15117,N_13181,N_13130);
nor U15118 (N_15118,N_13681,N_14105);
or U15119 (N_15119,N_13667,N_12766);
xnor U15120 (N_15120,N_13032,N_14066);
or U15121 (N_15121,N_12708,N_12837);
nor U15122 (N_15122,N_12791,N_13410);
or U15123 (N_15123,N_12998,N_14323);
nand U15124 (N_15124,N_14731,N_14087);
nor U15125 (N_15125,N_14774,N_14311);
nor U15126 (N_15126,N_13497,N_13771);
or U15127 (N_15127,N_13637,N_13673);
nor U15128 (N_15128,N_12600,N_13974);
xnor U15129 (N_15129,N_13149,N_12730);
xor U15130 (N_15130,N_13252,N_13888);
xor U15131 (N_15131,N_13052,N_12666);
nand U15132 (N_15132,N_13562,N_12593);
or U15133 (N_15133,N_14578,N_13926);
or U15134 (N_15134,N_13005,N_13241);
nand U15135 (N_15135,N_13509,N_13610);
xnor U15136 (N_15136,N_14237,N_13923);
nand U15137 (N_15137,N_14996,N_13641);
nand U15138 (N_15138,N_13688,N_13958);
nand U15139 (N_15139,N_12508,N_14922);
nand U15140 (N_15140,N_14958,N_13101);
and U15141 (N_15141,N_14520,N_13306);
nor U15142 (N_15142,N_14544,N_13010);
nor U15143 (N_15143,N_14197,N_14334);
xor U15144 (N_15144,N_12877,N_13331);
xnor U15145 (N_15145,N_14891,N_12842);
xnor U15146 (N_15146,N_13582,N_14722);
and U15147 (N_15147,N_13498,N_13444);
nand U15148 (N_15148,N_13783,N_14957);
and U15149 (N_15149,N_12551,N_14296);
or U15150 (N_15150,N_13233,N_12506);
nor U15151 (N_15151,N_13140,N_13627);
nand U15152 (N_15152,N_14070,N_14215);
xor U15153 (N_15153,N_14328,N_14344);
and U15154 (N_15154,N_14551,N_13883);
nand U15155 (N_15155,N_13686,N_14403);
nand U15156 (N_15156,N_14816,N_13520);
nor U15157 (N_15157,N_14025,N_14022);
xnor U15158 (N_15158,N_14063,N_14364);
nor U15159 (N_15159,N_14824,N_13659);
or U15160 (N_15160,N_14909,N_12653);
xnor U15161 (N_15161,N_13047,N_14547);
and U15162 (N_15162,N_14515,N_14616);
and U15163 (N_15163,N_12966,N_13021);
nand U15164 (N_15164,N_13062,N_13332);
and U15165 (N_15165,N_14430,N_14997);
nand U15166 (N_15166,N_13247,N_12546);
nand U15167 (N_15167,N_14863,N_13515);
xor U15168 (N_15168,N_13541,N_14309);
xnor U15169 (N_15169,N_12673,N_13018);
or U15170 (N_15170,N_14114,N_14370);
nand U15171 (N_15171,N_14340,N_13730);
or U15172 (N_15172,N_14196,N_13127);
nor U15173 (N_15173,N_13947,N_14042);
xnor U15174 (N_15174,N_14522,N_13457);
nand U15175 (N_15175,N_14003,N_14929);
nand U15176 (N_15176,N_12857,N_14490);
nor U15177 (N_15177,N_12542,N_14552);
nor U15178 (N_15178,N_13208,N_14756);
nor U15179 (N_15179,N_14718,N_14651);
nand U15180 (N_15180,N_14737,N_12693);
nor U15181 (N_15181,N_14765,N_12720);
or U15182 (N_15182,N_13098,N_12771);
xor U15183 (N_15183,N_13555,N_13053);
or U15184 (N_15184,N_13171,N_13735);
or U15185 (N_15185,N_14355,N_12828);
nor U15186 (N_15186,N_14799,N_14093);
or U15187 (N_15187,N_14684,N_13371);
and U15188 (N_15188,N_14163,N_13810);
nand U15189 (N_15189,N_14336,N_14809);
and U15190 (N_15190,N_12539,N_13107);
or U15191 (N_15191,N_13085,N_13600);
nor U15192 (N_15192,N_13824,N_14558);
or U15193 (N_15193,N_13626,N_13693);
nand U15194 (N_15194,N_13558,N_13392);
xor U15195 (N_15195,N_13911,N_14588);
and U15196 (N_15196,N_12918,N_12814);
xor U15197 (N_15197,N_14038,N_14012);
nor U15198 (N_15198,N_13312,N_12599);
xnor U15199 (N_15199,N_13689,N_13408);
nor U15200 (N_15200,N_13789,N_12986);
and U15201 (N_15201,N_13205,N_13987);
nand U15202 (N_15202,N_13133,N_13812);
xor U15203 (N_15203,N_14989,N_13711);
nor U15204 (N_15204,N_12819,N_13639);
nand U15205 (N_15205,N_14853,N_14011);
xor U15206 (N_15206,N_14166,N_13419);
or U15207 (N_15207,N_13277,N_13532);
and U15208 (N_15208,N_13114,N_12691);
xor U15209 (N_15209,N_12543,N_12699);
xnor U15210 (N_15210,N_13184,N_13882);
and U15211 (N_15211,N_12630,N_14527);
and U15212 (N_15212,N_13454,N_13349);
xnor U15213 (N_15213,N_14366,N_12822);
xnor U15214 (N_15214,N_14643,N_14293);
nand U15215 (N_15215,N_12782,N_12907);
or U15216 (N_15216,N_14448,N_14901);
xnor U15217 (N_15217,N_13712,N_12606);
nand U15218 (N_15218,N_12592,N_14779);
nand U15219 (N_15219,N_14471,N_13827);
nor U15220 (N_15220,N_14102,N_13988);
nor U15221 (N_15221,N_13850,N_14017);
or U15222 (N_15222,N_12564,N_14401);
and U15223 (N_15223,N_14738,N_14873);
or U15224 (N_15224,N_14646,N_13083);
nor U15225 (N_15225,N_14866,N_14856);
nor U15226 (N_15226,N_14519,N_13095);
nand U15227 (N_15227,N_14962,N_14251);
or U15228 (N_15228,N_14266,N_14264);
or U15229 (N_15229,N_13842,N_14443);
nor U15230 (N_15230,N_14100,N_13607);
or U15231 (N_15231,N_14084,N_14505);
or U15232 (N_15232,N_13415,N_14421);
nor U15233 (N_15233,N_13399,N_13654);
and U15234 (N_15234,N_12604,N_13716);
or U15235 (N_15235,N_13120,N_13717);
xnor U15236 (N_15236,N_12897,N_12677);
and U15237 (N_15237,N_14742,N_14150);
and U15238 (N_15238,N_12629,N_14397);
and U15239 (N_15239,N_14465,N_13588);
xor U15240 (N_15240,N_13939,N_13268);
or U15241 (N_15241,N_13206,N_12975);
and U15242 (N_15242,N_12944,N_14154);
xnor U15243 (N_15243,N_13478,N_12949);
or U15244 (N_15244,N_13676,N_13618);
and U15245 (N_15245,N_14723,N_14733);
nor U15246 (N_15246,N_12895,N_14329);
xor U15247 (N_15247,N_12514,N_13030);
or U15248 (N_15248,N_12726,N_12672);
nor U15249 (N_15249,N_12816,N_12811);
nor U15250 (N_15250,N_13055,N_12670);
or U15251 (N_15251,N_13377,N_13892);
nor U15252 (N_15252,N_13283,N_13015);
or U15253 (N_15253,N_12698,N_14678);
nor U15254 (N_15254,N_12682,N_14463);
nand U15255 (N_15255,N_14835,N_13212);
xor U15256 (N_15256,N_13157,N_12689);
xnor U15257 (N_15257,N_14318,N_14645);
xnor U15258 (N_15258,N_14877,N_14158);
nor U15259 (N_15259,N_12957,N_14852);
nor U15260 (N_15260,N_14555,N_13458);
xor U15261 (N_15261,N_14026,N_13971);
nand U15262 (N_15262,N_14249,N_14963);
nand U15263 (N_15263,N_13597,N_13841);
and U15264 (N_15264,N_14613,N_13916);
nand U15265 (N_15265,N_13027,N_13910);
nand U15266 (N_15266,N_13502,N_12572);
and U15267 (N_15267,N_13544,N_13075);
nor U15268 (N_15268,N_14207,N_13311);
nand U15269 (N_15269,N_13466,N_12587);
nand U15270 (N_15270,N_12563,N_12550);
nor U15271 (N_15271,N_13522,N_14808);
nand U15272 (N_15272,N_13770,N_13289);
and U15273 (N_15273,N_14956,N_14055);
nor U15274 (N_15274,N_14338,N_12660);
nand U15275 (N_15275,N_13321,N_14906);
and U15276 (N_15276,N_13216,N_13757);
nor U15277 (N_15277,N_12953,N_13372);
and U15278 (N_15278,N_13418,N_12707);
or U15279 (N_15279,N_12853,N_12845);
or U15280 (N_15280,N_13747,N_13942);
nand U15281 (N_15281,N_13675,N_14825);
or U15282 (N_15282,N_13536,N_14161);
xnor U15283 (N_15283,N_14748,N_13265);
and U15284 (N_15284,N_14998,N_13438);
and U15285 (N_15285,N_12871,N_13861);
xor U15286 (N_15286,N_12988,N_13867);
xnor U15287 (N_15287,N_14730,N_13437);
xor U15288 (N_15288,N_13944,N_13665);
xnor U15289 (N_15289,N_13937,N_14287);
nand U15290 (N_15290,N_13889,N_12626);
xor U15291 (N_15291,N_14569,N_13200);
and U15292 (N_15292,N_14585,N_13426);
xnor U15293 (N_15293,N_14298,N_12595);
xnor U15294 (N_15294,N_13664,N_14400);
xnor U15295 (N_15295,N_14858,N_12806);
xor U15296 (N_15296,N_14680,N_13256);
and U15297 (N_15297,N_13042,N_14258);
nand U15298 (N_15298,N_14894,N_13708);
xnor U15299 (N_15299,N_13228,N_13699);
nor U15300 (N_15300,N_14438,N_13766);
or U15301 (N_15301,N_14424,N_13952);
xor U15302 (N_15302,N_14407,N_14124);
nor U15303 (N_15303,N_14069,N_14123);
nor U15304 (N_15304,N_14362,N_14728);
nand U15305 (N_15305,N_14314,N_13093);
or U15306 (N_15306,N_13749,N_12915);
nor U15307 (N_15307,N_14317,N_14701);
nor U15308 (N_15308,N_14895,N_13351);
xnor U15309 (N_15309,N_13461,N_13906);
nor U15310 (N_15310,N_13656,N_13388);
xnor U15311 (N_15311,N_14693,N_14120);
or U15312 (N_15312,N_12756,N_14152);
or U15313 (N_15313,N_13403,N_13797);
xor U15314 (N_15314,N_14115,N_13574);
or U15315 (N_15315,N_14553,N_13188);
or U15316 (N_15316,N_13998,N_14959);
and U15317 (N_15317,N_12777,N_14666);
nand U15318 (N_15318,N_13674,N_12789);
nand U15319 (N_15319,N_14044,N_14371);
xor U15320 (N_15320,N_13225,N_13559);
and U15321 (N_15321,N_13614,N_14601);
nand U15322 (N_15322,N_13723,N_12878);
nor U15323 (N_15323,N_13741,N_13425);
nor U15324 (N_15324,N_14431,N_13602);
and U15325 (N_15325,N_14846,N_12761);
or U15326 (N_15326,N_13039,N_14342);
nand U15327 (N_15327,N_12537,N_14411);
or U15328 (N_15328,N_13421,N_13315);
or U15329 (N_15329,N_14171,N_13084);
nand U15330 (N_15330,N_13397,N_13428);
and U15331 (N_15331,N_14935,N_14634);
and U15332 (N_15332,N_12676,N_14095);
nand U15333 (N_15333,N_13568,N_12731);
xor U15334 (N_15334,N_14148,N_13007);
nor U15335 (N_15335,N_13904,N_14591);
xor U15336 (N_15336,N_14942,N_14944);
nor U15337 (N_15337,N_14876,N_12968);
or U15338 (N_15338,N_14524,N_14488);
nand U15339 (N_15339,N_14450,N_13337);
or U15340 (N_15340,N_13807,N_14002);
xnor U15341 (N_15341,N_13727,N_14949);
or U15342 (N_15342,N_13777,N_13424);
and U15343 (N_15343,N_14927,N_14322);
and U15344 (N_15344,N_13155,N_14712);
xnor U15345 (N_15345,N_14380,N_14791);
nand U15346 (N_15346,N_14758,N_12721);
and U15347 (N_15347,N_13103,N_12757);
nor U15348 (N_15348,N_14033,N_13163);
xor U15349 (N_15349,N_14969,N_13746);
nor U15350 (N_15350,N_12535,N_12750);
and U15351 (N_15351,N_12869,N_13754);
nand U15352 (N_15352,N_13976,N_14999);
nor U15353 (N_15353,N_12881,N_14139);
xnor U15354 (N_15354,N_14755,N_13837);
nand U15355 (N_15355,N_14104,N_13058);
nand U15356 (N_15356,N_12554,N_13196);
and U15357 (N_15357,N_14579,N_14494);
xor U15358 (N_15358,N_13452,N_14775);
or U15359 (N_15359,N_14849,N_13379);
nand U15360 (N_15360,N_14881,N_12964);
and U15361 (N_15361,N_13963,N_14820);
nand U15362 (N_15362,N_13401,N_14392);
and U15363 (N_15363,N_14162,N_13924);
xor U15364 (N_15364,N_14676,N_12544);
xnor U15365 (N_15365,N_14213,N_13378);
and U15366 (N_15366,N_12608,N_13391);
nor U15367 (N_15367,N_14052,N_13625);
nor U15368 (N_15368,N_13002,N_13104);
nand U15369 (N_15369,N_13448,N_13553);
or U15370 (N_15370,N_13385,N_13613);
and U15371 (N_15371,N_14548,N_13806);
or U15372 (N_15372,N_12651,N_14566);
nor U15373 (N_15373,N_14377,N_13992);
xnor U15374 (N_15374,N_14202,N_14890);
or U15375 (N_15375,N_14357,N_13648);
xnor U15376 (N_15376,N_14530,N_12706);
and U15377 (N_15377,N_13570,N_13412);
or U15378 (N_15378,N_13977,N_12585);
and U15379 (N_15379,N_14467,N_14222);
or U15380 (N_15380,N_14284,N_14811);
nor U15381 (N_15381,N_13760,N_13534);
or U15382 (N_15382,N_12690,N_13006);
or U15383 (N_15383,N_14930,N_14302);
and U15384 (N_15384,N_13305,N_14994);
and U15385 (N_15385,N_14694,N_14594);
or U15386 (N_15386,N_13117,N_14734);
nor U15387 (N_15387,N_12919,N_12765);
nand U15388 (N_15388,N_13631,N_14598);
nor U15389 (N_15389,N_14554,N_14750);
or U15390 (N_15390,N_14608,N_13594);
nor U15391 (N_15391,N_13523,N_13748);
xnor U15392 (N_15392,N_14982,N_13821);
or U15393 (N_15393,N_14667,N_13158);
xnor U15394 (N_15394,N_12669,N_13302);
or U15395 (N_15395,N_14130,N_12874);
and U15396 (N_15396,N_14321,N_13473);
nor U15397 (N_15397,N_13413,N_14889);
nor U15398 (N_15398,N_14784,N_14574);
nand U15399 (N_15399,N_14778,N_12695);
nor U15400 (N_15400,N_12729,N_12529);
or U15401 (N_15401,N_14313,N_12588);
xnor U15402 (N_15402,N_14976,N_13650);
or U15403 (N_15403,N_13740,N_14903);
nand U15404 (N_15404,N_13925,N_12674);
xor U15405 (N_15405,N_13038,N_13822);
and U15406 (N_15406,N_13929,N_12911);
and U15407 (N_15407,N_13174,N_12917);
or U15408 (N_15408,N_12793,N_13634);
xor U15409 (N_15409,N_14316,N_14539);
nand U15410 (N_15410,N_13617,N_12663);
nor U15411 (N_15411,N_13825,N_12701);
and U15412 (N_15412,N_14621,N_13336);
xor U15413 (N_15413,N_13226,N_13622);
nor U15414 (N_15414,N_13245,N_14481);
and U15415 (N_15415,N_13930,N_12574);
nand U15416 (N_15416,N_14771,N_13940);
or U15417 (N_15417,N_14729,N_14509);
nand U15418 (N_15418,N_14306,N_12538);
or U15419 (N_15419,N_13074,N_13710);
nor U15420 (N_15420,N_14368,N_13877);
nor U15421 (N_15421,N_14270,N_14943);
and U15422 (N_15422,N_12888,N_14268);
nand U15423 (N_15423,N_12616,N_14373);
or U15424 (N_15424,N_13215,N_13313);
xnor U15425 (N_15425,N_14263,N_12643);
nor U15426 (N_15426,N_13843,N_12640);
or U15427 (N_15427,N_14285,N_13100);
and U15428 (N_15428,N_13489,N_13565);
or U15429 (N_15429,N_14968,N_12951);
nor U15430 (N_15430,N_14947,N_13270);
or U15431 (N_15431,N_13170,N_13137);
xor U15432 (N_15432,N_13433,N_14727);
or U15433 (N_15433,N_14918,N_14023);
and U15434 (N_15434,N_13019,N_14653);
xor U15435 (N_15435,N_14172,N_14468);
nor U15436 (N_15436,N_13577,N_14821);
or U15437 (N_15437,N_14016,N_14422);
nor U15438 (N_15438,N_13671,N_12607);
and U15439 (N_15439,N_12619,N_14456);
nand U15440 (N_15440,N_14262,N_14446);
and U15441 (N_15441,N_13649,N_14337);
and U15442 (N_15442,N_13141,N_13572);
and U15443 (N_15443,N_13722,N_12884);
or U15444 (N_15444,N_14869,N_12686);
xor U15445 (N_15445,N_12856,N_13986);
nand U15446 (N_15446,N_13927,N_12779);
nand U15447 (N_15447,N_14785,N_12784);
and U15448 (N_15448,N_13762,N_14977);
xnor U15449 (N_15449,N_13776,N_13177);
or U15450 (N_15450,N_12921,N_13920);
and U15451 (N_15451,N_13968,N_14193);
and U15452 (N_15452,N_13257,N_14609);
or U15453 (N_15453,N_12916,N_14090);
nor U15454 (N_15454,N_14304,N_14269);
xnor U15455 (N_15455,N_14437,N_12767);
nand U15456 (N_15456,N_12679,N_14109);
xor U15457 (N_15457,N_14851,N_14587);
or U15458 (N_15458,N_13773,N_13737);
nand U15459 (N_15459,N_13836,N_12652);
xnor U15460 (N_15460,N_12956,N_13364);
nand U15461 (N_15461,N_14528,N_13640);
xnor U15462 (N_15462,N_14133,N_14879);
xnor U15463 (N_15463,N_12773,N_14662);
nor U15464 (N_15464,N_14806,N_14767);
nor U15465 (N_15465,N_12545,N_13300);
nand U15466 (N_15466,N_13266,N_13679);
xor U15467 (N_15467,N_12763,N_14412);
nand U15468 (N_15468,N_13838,N_14436);
nand U15469 (N_15469,N_12696,N_13099);
or U15470 (N_15470,N_14295,N_14705);
and U15471 (N_15471,N_12644,N_14349);
nand U15472 (N_15472,N_13774,N_12532);
or U15473 (N_15473,N_13862,N_14681);
and U15474 (N_15474,N_14516,N_13529);
nor U15475 (N_15475,N_14155,N_14228);
xnor U15476 (N_15476,N_12905,N_13147);
or U15477 (N_15477,N_14217,N_12808);
and U15478 (N_15478,N_14178,N_13347);
xor U15479 (N_15479,N_13314,N_14174);
or U15480 (N_15480,N_12559,N_14736);
and U15481 (N_15481,N_13434,N_13344);
xnor U15482 (N_15482,N_12555,N_13767);
nand U15483 (N_15483,N_12634,N_13872);
or U15484 (N_15484,N_12823,N_13380);
and U15485 (N_15485,N_12515,N_14657);
and U15486 (N_15486,N_14119,N_14904);
and U15487 (N_15487,N_13703,N_13899);
and U15488 (N_15488,N_14966,N_12650);
nor U15489 (N_15489,N_13192,N_14000);
or U15490 (N_15490,N_14980,N_13035);
or U15491 (N_15491,N_13109,N_13635);
nor U15492 (N_15492,N_13474,N_12873);
xor U15493 (N_15493,N_12523,N_14198);
nand U15494 (N_15494,N_12831,N_13269);
xnor U15495 (N_15495,N_12702,N_12678);
xnor U15496 (N_15496,N_12863,N_13012);
xor U15497 (N_15497,N_14083,N_13587);
xnor U15498 (N_15498,N_13513,N_14605);
xor U15499 (N_15499,N_13180,N_12681);
or U15500 (N_15500,N_13666,N_14076);
xnor U15501 (N_15501,N_13615,N_13514);
and U15502 (N_15502,N_14589,N_14290);
and U15503 (N_15503,N_14797,N_14632);
or U15504 (N_15504,N_13660,N_12776);
xnor U15505 (N_15505,N_13382,N_14138);
xor U15506 (N_15506,N_14053,N_14972);
nand U15507 (N_15507,N_14834,N_12985);
nand U15508 (N_15508,N_13828,N_14654);
and U15509 (N_15509,N_13645,N_12939);
or U15510 (N_15510,N_14711,N_14614);
xor U15511 (N_15511,N_13191,N_13599);
and U15512 (N_15512,N_13193,N_14724);
xnor U15513 (N_15513,N_13991,N_14819);
nor U15514 (N_15514,N_13209,N_13725);
nand U15515 (N_15515,N_13878,N_14195);
nand U15516 (N_15516,N_14971,N_14001);
and U15517 (N_15517,N_14507,N_14747);
and U15518 (N_15518,N_14470,N_14485);
nand U15519 (N_15519,N_13545,N_13456);
nor U15520 (N_15520,N_13243,N_13333);
nand U15521 (N_15521,N_13606,N_12892);
or U15522 (N_15522,N_13898,N_13902);
and U15523 (N_15523,N_13094,N_13624);
nand U15524 (N_15524,N_14359,N_13324);
nor U15525 (N_15525,N_14802,N_12938);
nand U15526 (N_15526,N_13595,N_13786);
or U15527 (N_15527,N_13285,N_13865);
nor U15528 (N_15528,N_14117,N_13790);
nor U15529 (N_15529,N_13001,N_12995);
nor U15530 (N_15530,N_13483,N_14946);
nor U15531 (N_15531,N_13586,N_13046);
nor U15532 (N_15532,N_13159,N_14391);
nor U15533 (N_15533,N_14492,N_13148);
nor U15534 (N_15534,N_14493,N_14305);
nand U15535 (N_15535,N_13683,N_14086);
or U15536 (N_15536,N_12890,N_14253);
and U15537 (N_15537,N_14699,N_13355);
and U15538 (N_15538,N_13652,N_14642);
and U15539 (N_15539,N_13763,N_12739);
or U15540 (N_15540,N_12684,N_14428);
nor U15541 (N_15541,N_13446,N_12976);
nand U15542 (N_15542,N_14630,N_12705);
nor U15543 (N_15543,N_12826,N_12927);
and U15544 (N_15544,N_13082,N_12627);
and U15545 (N_15545,N_13919,N_12768);
xnor U15546 (N_15546,N_14014,N_14379);
and U15547 (N_15547,N_13420,N_13966);
and U15548 (N_15548,N_12796,N_14458);
or U15549 (N_15549,N_12972,N_14577);
xnor U15550 (N_15550,N_14983,N_13863);
nor U15551 (N_15551,N_13780,N_13967);
and U15552 (N_15552,N_14369,N_12924);
nand U15553 (N_15553,N_14027,N_12586);
or U15554 (N_15554,N_14659,N_14116);
or U15555 (N_15555,N_14844,N_13435);
nor U15556 (N_15556,N_12772,N_12575);
nand U15557 (N_15557,N_13034,N_12832);
and U15558 (N_15558,N_14415,N_13447);
nand U15559 (N_15559,N_14619,N_13077);
and U15560 (N_15560,N_13414,N_13009);
and U15561 (N_15561,N_12521,N_13736);
xor U15562 (N_15562,N_14259,N_12920);
nand U15563 (N_15563,N_13417,N_13296);
xor U15564 (N_15564,N_12954,N_13221);
nand U15565 (N_15565,N_12979,N_13831);
or U15566 (N_15566,N_14658,N_12645);
nor U15567 (N_15567,N_13815,N_13759);
or U15568 (N_15568,N_14236,N_14170);
nor U15569 (N_15569,N_14500,N_13696);
nand U15570 (N_15570,N_14513,N_13501);
nor U15571 (N_15571,N_12556,N_14078);
or U15572 (N_15572,N_14590,N_14035);
xor U15573 (N_15573,N_12751,N_14872);
and U15574 (N_15574,N_12569,N_14773);
xor U15575 (N_15575,N_13122,N_12862);
or U15576 (N_15576,N_13427,N_12583);
and U15577 (N_15577,N_12914,N_14964);
xor U15578 (N_15578,N_14144,N_14965);
xnor U15579 (N_15579,N_14107,N_14843);
xor U15580 (N_15580,N_14503,N_13376);
nand U15581 (N_15581,N_14006,N_14131);
nand U15582 (N_15582,N_14793,N_14804);
and U15583 (N_15583,N_13016,N_13956);
xnor U15584 (N_15584,N_12661,N_13264);
or U15585 (N_15585,N_12571,N_14433);
and U15586 (N_15586,N_14898,N_14768);
nand U15587 (N_15587,N_12597,N_12566);
and U15588 (N_15588,N_13189,N_14214);
nor U15589 (N_15589,N_14762,N_14464);
nand U15590 (N_15590,N_13928,N_13278);
nand U15591 (N_15591,N_13049,N_13896);
nor U15592 (N_15592,N_13304,N_14960);
and U15593 (N_15593,N_13450,N_13407);
nor U15594 (N_15594,N_13143,N_12578);
or U15595 (N_15595,N_13800,N_14219);
nor U15596 (N_15596,N_13028,N_13996);
nand U15597 (N_15597,N_12928,N_13350);
xor U15598 (N_15598,N_13358,N_14740);
nor U15599 (N_15599,N_13611,N_12785);
nand U15600 (N_15600,N_13207,N_14345);
or U15601 (N_15601,N_13662,N_12809);
xnor U15602 (N_15602,N_14136,N_14884);
and U15603 (N_15603,N_14826,N_13535);
or U15604 (N_15604,N_14886,N_13579);
or U15605 (N_15605,N_13309,N_14413);
and U15606 (N_15606,N_12781,N_13330);
or U15607 (N_15607,N_14427,N_12734);
and U15608 (N_15608,N_12959,N_12889);
nor U15609 (N_15609,N_14647,N_13829);
and U15610 (N_15610,N_13477,N_13479);
or U15611 (N_15611,N_14510,N_13633);
or U15612 (N_15612,N_14878,N_13950);
xnor U15613 (N_15613,N_13432,N_14897);
nor U15614 (N_15614,N_14991,N_14713);
or U15615 (N_15615,N_14837,N_13472);
nor U15616 (N_15616,N_14240,N_13844);
xnor U15617 (N_15617,N_14288,N_12620);
or U15618 (N_15618,N_13097,N_14838);
xor U15619 (N_15619,N_14089,N_12611);
or U15620 (N_15620,N_12632,N_13538);
and U15621 (N_15621,N_14082,N_14361);
nor U15622 (N_15622,N_14636,N_13451);
nand U15623 (N_15623,N_14627,N_14867);
xnor U15624 (N_15624,N_14810,N_14719);
xor U15625 (N_15625,N_12971,N_13162);
and U15626 (N_15626,N_12692,N_13521);
and U15627 (N_15627,N_13752,N_14453);
nor U15628 (N_15628,N_13070,N_14444);
nand U15629 (N_15629,N_13979,N_14273);
nand U15630 (N_15630,N_13348,N_13164);
or U15631 (N_15631,N_13287,N_13319);
or U15632 (N_15632,N_14297,N_14840);
and U15633 (N_15633,N_13576,N_14672);
xor U15634 (N_15634,N_13000,N_13775);
xor U15635 (N_15635,N_12598,N_13557);
and U15636 (N_15636,N_12868,N_14466);
nor U15637 (N_15637,N_13416,N_13698);
and U15638 (N_15638,N_13530,N_12628);
nor U15639 (N_15639,N_13169,N_14325);
nor U15640 (N_15640,N_13840,N_14717);
or U15641 (N_15641,N_13374,N_14146);
and U15642 (N_15642,N_12885,N_14860);
nand U15643 (N_15643,N_14875,N_13185);
or U15644 (N_15644,N_13684,N_13692);
xnor U15645 (N_15645,N_13322,N_13238);
or U15646 (N_15646,N_12711,N_12754);
and U15647 (N_15647,N_12840,N_12736);
or U15648 (N_15648,N_14232,N_13485);
nor U15649 (N_15649,N_12992,N_12820);
or U15650 (N_15650,N_13554,N_13551);
and U15651 (N_15651,N_13999,N_13166);
nand U15652 (N_15652,N_14326,N_13860);
and U15653 (N_15653,N_12967,N_13700);
nor U15654 (N_15654,N_14064,N_13578);
nor U15655 (N_15655,N_13061,N_12830);
xor U15656 (N_15656,N_14504,N_12803);
nor U15657 (N_15657,N_14482,N_13248);
nor U15658 (N_15658,N_12524,N_14024);
nor U15659 (N_15659,N_12675,N_14386);
and U15660 (N_15660,N_14417,N_13299);
nand U15661 (N_15661,N_14378,N_13915);
and U15662 (N_15662,N_14156,N_14883);
xnor U15663 (N_15663,N_14781,N_14915);
or U15664 (N_15664,N_12531,N_14685);
nand U15665 (N_15665,N_14831,N_13632);
xor U15666 (N_15666,N_14593,N_12940);
nand U15667 (N_15667,N_14660,N_13508);
or U15668 (N_15668,N_14708,N_14990);
or U15669 (N_15669,N_14281,N_14250);
or U15670 (N_15670,N_12500,N_14426);
or U15671 (N_15671,N_13873,N_14936);
xor U15672 (N_15672,N_14384,N_13744);
or U15673 (N_15673,N_14291,N_14445);
xor U15674 (N_15674,N_13394,N_12648);
and U15675 (N_15675,N_13151,N_12667);
xor U15676 (N_15676,N_12901,N_14099);
nor U15677 (N_15677,N_12507,N_14938);
nor U15678 (N_15678,N_13500,N_13685);
nand U15679 (N_15679,N_13292,N_14352);
and U15680 (N_15680,N_14871,N_14057);
nand U15681 (N_15681,N_12655,N_13008);
nand U15682 (N_15682,N_13646,N_14611);
nand U15683 (N_15683,N_13031,N_13476);
nand U15684 (N_15684,N_14920,N_14562);
and U15685 (N_15685,N_13533,N_13195);
or U15686 (N_15686,N_14185,N_14167);
xor U15687 (N_15687,N_14181,N_14988);
nand U15688 (N_15688,N_13168,N_13756);
nor U15689 (N_15689,N_14735,N_12591);
xnor U15690 (N_15690,N_12899,N_13552);
and U15691 (N_15691,N_13628,N_14310);
nand U15692 (N_15692,N_12654,N_14054);
nor U15693 (N_15693,N_14501,N_13469);
xor U15694 (N_15694,N_14655,N_14489);
and U15695 (N_15695,N_14480,N_14557);
nand U15696 (N_15696,N_13323,N_12839);
and U15697 (N_15697,N_13217,N_14294);
nor U15698 (N_15698,N_14549,N_13680);
or U15699 (N_15699,N_13505,N_14612);
or U15700 (N_15700,N_13575,N_12635);
xor U15701 (N_15701,N_14125,N_13063);
or U15702 (N_15702,N_13609,N_13251);
or U15703 (N_15703,N_13604,N_13480);
and U15704 (N_15704,N_14425,N_14650);
nand U15705 (N_15705,N_13020,N_14801);
and U15706 (N_15706,N_13290,N_14476);
and U15707 (N_15707,N_13275,N_13516);
and U15708 (N_15708,N_13118,N_13024);
nand U15709 (N_15709,N_13496,N_14508);
or U15710 (N_15710,N_12562,N_14818);
or U15711 (N_15711,N_13912,N_14874);
and U15712 (N_15712,N_14058,N_12900);
and U15713 (N_15713,N_14537,N_13363);
or U15714 (N_15714,N_14399,N_13584);
nand U15715 (N_15715,N_14230,N_13962);
nor U15716 (N_15716,N_14521,N_13381);
nand U15717 (N_15717,N_14995,N_13040);
xnor U15718 (N_15718,N_12557,N_13440);
or U15719 (N_15719,N_12812,N_12636);
nand U15720 (N_15720,N_14169,N_12980);
nor U15721 (N_15721,N_12740,N_12774);
nor U15722 (N_15722,N_13581,N_13830);
xor U15723 (N_15723,N_12605,N_14335);
and U15724 (N_15724,N_14910,N_14040);
nor U15725 (N_15725,N_14981,N_13138);
or U15726 (N_15726,N_13484,N_12713);
or U15727 (N_15727,N_14633,N_14452);
and U15728 (N_15728,N_14113,N_13638);
and U15729 (N_15729,N_13092,N_13179);
nand U15730 (N_15730,N_13907,N_14226);
xnor U15731 (N_15731,N_13983,N_13161);
and U15732 (N_15732,N_14725,N_14211);
nor U15733 (N_15733,N_12891,N_14970);
xnor U15734 (N_15734,N_14191,N_12937);
nand U15735 (N_15735,N_14015,N_12994);
xnor U15736 (N_15736,N_13848,N_14045);
and U15737 (N_15737,N_14143,N_14056);
nor U15738 (N_15738,N_13273,N_14542);
nor U15739 (N_15739,N_13172,N_13732);
nor U15740 (N_15740,N_13605,N_14247);
or U15741 (N_15741,N_14248,N_14429);
and U15742 (N_15742,N_12790,N_12780);
xnor U15743 (N_15743,N_12815,N_14541);
xnor U15744 (N_15744,N_13261,N_14275);
xor U15745 (N_15745,N_12866,N_14763);
and U15746 (N_15746,N_12973,N_12710);
nor U15747 (N_15747,N_13900,N_12880);
nand U15748 (N_15748,N_13023,N_14688);
and U15749 (N_15749,N_12723,N_14252);
nor U15750 (N_15750,N_14279,N_12955);
xor U15751 (N_15751,N_13994,N_12850);
nor U15752 (N_15752,N_12659,N_14393);
nand U15753 (N_15753,N_13430,N_13339);
and U15754 (N_15754,N_14091,N_14300);
nand U15755 (N_15755,N_13792,N_13393);
nor U15756 (N_15756,N_13326,N_14788);
nand U15757 (N_15757,N_13852,N_14744);
nand U15758 (N_15758,N_13022,N_13993);
xnor U15759 (N_15759,N_14394,N_13295);
nor U15760 (N_15760,N_13670,N_12510);
nand U15761 (N_15761,N_13072,N_14940);
and U15762 (N_15762,N_13218,N_13423);
nand U15763 (N_15763,N_14743,N_13682);
or U15764 (N_15764,N_13139,N_13653);
nor U15765 (N_15765,N_14348,N_14029);
nor U15766 (N_15766,N_14599,N_13591);
xnor U15767 (N_15767,N_13547,N_14813);
nor U15768 (N_15768,N_14661,N_12565);
nand U15769 (N_15769,N_13526,N_13990);
nand U15770 (N_15770,N_14122,N_13936);
or U15771 (N_15771,N_13441,N_14993);
and U15772 (N_15772,N_13059,N_12727);
xor U15773 (N_15773,N_13855,N_14622);
nand U15774 (N_15774,N_14223,N_13369);
nor U15775 (N_15775,N_12930,N_14870);
and U15776 (N_15776,N_13619,N_14640);
nor U15777 (N_15777,N_13755,N_13881);
nand U15778 (N_15778,N_14716,N_12755);
nor U15779 (N_15779,N_12870,N_12805);
and U15780 (N_15780,N_13135,N_13854);
and U15781 (N_15781,N_12844,N_13025);
xnor U15782 (N_15782,N_13328,N_13259);
nand U15783 (N_15783,N_13957,N_13203);
or U15784 (N_15784,N_14239,N_14586);
nor U15785 (N_15785,N_13705,N_12700);
xor U15786 (N_15786,N_14560,N_14331);
nand U15787 (N_15787,N_14358,N_13909);
and U15788 (N_15788,N_13227,N_12728);
and U15789 (N_15789,N_14795,N_14696);
or U15790 (N_15790,N_12540,N_14908);
nor U15791 (N_15791,N_12633,N_13404);
or U15792 (N_15792,N_13846,N_13620);
xnor U15793 (N_15793,N_13037,N_13329);
nand U15794 (N_15794,N_13778,N_13495);
or U15795 (N_15795,N_12801,N_12797);
or U15796 (N_15796,N_14495,N_14312);
xnor U15797 (N_15797,N_14032,N_13781);
and U15798 (N_15798,N_14350,N_13345);
or U15799 (N_15799,N_13647,N_14546);
nand U15800 (N_15800,N_12893,N_14420);
nand U15801 (N_15801,N_12560,N_13282);
or U15802 (N_15802,N_13156,N_13583);
nand U15803 (N_15803,N_14805,N_13386);
nor U15804 (N_15804,N_14405,N_13677);
nand U15805 (N_15805,N_14108,N_12746);
nor U15806 (N_15806,N_14836,N_13078);
xor U15807 (N_15807,N_14985,N_12982);
xor U15808 (N_15808,N_14899,N_12576);
and U15809 (N_15809,N_14347,N_13621);
and U15810 (N_15810,N_12526,N_14543);
nor U15811 (N_15811,N_13352,N_14303);
xnor U15812 (N_15812,N_12558,N_14986);
nand U15813 (N_15813,N_13431,N_14447);
or U15814 (N_15814,N_13733,N_12518);
nor U15815 (N_15815,N_13561,N_14855);
or U15816 (N_15816,N_12852,N_12825);
or U15817 (N_15817,N_14383,N_13069);
xor U15818 (N_15818,N_14277,N_14210);
and U15819 (N_15819,N_13894,N_14638);
nor U15820 (N_15820,N_12887,N_13237);
nor U15821 (N_15821,N_13820,N_12594);
and U15822 (N_15822,N_14356,N_14073);
xor U15823 (N_15823,N_14907,N_13954);
and U15824 (N_15824,N_12733,N_13298);
xor U15825 (N_15825,N_13356,N_14941);
or U15826 (N_15826,N_13969,N_14992);
and U15827 (N_15827,N_14048,N_14404);
xor U15828 (N_15828,N_14030,N_14602);
nand U15829 (N_15829,N_14343,N_14953);
or U15830 (N_15830,N_13995,N_14639);
xnor U15831 (N_15831,N_12997,N_13931);
nand U15832 (N_15832,N_13704,N_12525);
xor U15833 (N_15833,N_14194,N_13464);
and U15834 (N_15834,N_13965,N_14931);
nor U15835 (N_15835,N_14571,N_14176);
or U15836 (N_15836,N_13294,N_13729);
nor U15837 (N_15837,N_13481,N_14671);
nor U15838 (N_15838,N_13320,N_14790);
xnor U15839 (N_15839,N_12621,N_13488);
or U15840 (N_15840,N_13360,N_14861);
nor U15841 (N_15841,N_13884,N_14865);
nand U15842 (N_15842,N_13897,N_12516);
xor U15843 (N_15843,N_12787,N_12875);
and U15844 (N_15844,N_14265,N_12981);
and U15845 (N_15845,N_13669,N_13948);
nand U15846 (N_15846,N_12958,N_13110);
and U15847 (N_15847,N_13455,N_12993);
nor U15848 (N_15848,N_13303,N_13492);
xor U15849 (N_15849,N_12617,N_14346);
nor U15850 (N_15850,N_13201,N_14709);
nand U15851 (N_15851,N_14668,N_14267);
and U15852 (N_15852,N_14135,N_13220);
nand U15853 (N_15853,N_13519,N_13224);
nand U15854 (N_15854,N_12987,N_14149);
or U15855 (N_15855,N_13043,N_13004);
and U15856 (N_15856,N_13935,N_12709);
xor U15857 (N_15857,N_13887,N_14597);
nor U15858 (N_15858,N_12858,N_13366);
and U15859 (N_15859,N_13003,N_12580);
and U15860 (N_15860,N_12748,N_12818);
or U15861 (N_15861,N_14974,N_13013);
nor U15862 (N_15862,N_13108,N_14896);
xnor U15863 (N_15863,N_12775,N_13080);
nor U15864 (N_15864,N_13864,N_14526);
xnor U15865 (N_15865,N_12827,N_13787);
or U15866 (N_15866,N_14606,N_14556);
xor U15867 (N_15867,N_13764,N_12804);
nand U15868 (N_15868,N_12932,N_13814);
nor U15869 (N_15869,N_13367,N_13548);
or U15870 (N_15870,N_12738,N_14592);
or U15871 (N_15871,N_13341,N_14031);
or U15872 (N_15872,N_13504,N_13462);
xnor U15873 (N_15873,N_13242,N_14967);
xnor U15874 (N_15874,N_14280,N_13802);
nand U15875 (N_15875,N_12596,N_12894);
and U15876 (N_15876,N_13512,N_14770);
xor U15877 (N_15877,N_13131,N_13145);
or U15878 (N_15878,N_14402,N_13197);
and U15879 (N_15879,N_14697,N_14039);
and U15880 (N_15880,N_13678,N_13491);
nand U15881 (N_15881,N_12665,N_14829);
nor U15882 (N_15882,N_12745,N_14111);
xnor U15883 (N_15883,N_14656,N_14914);
nor U15884 (N_15884,N_13886,N_14776);
and U15885 (N_15885,N_14081,N_14620);
xnor U15886 (N_15886,N_13571,N_14205);
nor U15887 (N_15887,N_14473,N_14330);
and U15888 (N_15888,N_14626,N_13851);
xor U15889 (N_15889,N_14561,N_14618);
and U15890 (N_15890,N_12942,N_14046);
xnor U15891 (N_15891,N_14732,N_14165);
nand U15892 (N_15892,N_13734,N_14460);
nor U15893 (N_15893,N_12714,N_14902);
nand U15894 (N_15894,N_12851,N_12799);
nor U15895 (N_15895,N_14559,N_14200);
and U15896 (N_15896,N_14098,N_13517);
and U15897 (N_15897,N_12502,N_14531);
xnor U15898 (N_15898,N_14192,N_13186);
or U15899 (N_15899,N_14979,N_13527);
xnor U15900 (N_15900,N_13494,N_12613);
xnor U15901 (N_15901,N_12925,N_13279);
or U15902 (N_15902,N_12501,N_13091);
xnor U15903 (N_15903,N_14018,N_13236);
nor U15904 (N_15904,N_13657,N_14221);
nand U15905 (N_15905,N_14919,N_13359);
xnor U15906 (N_15906,N_14892,N_13753);
or U15907 (N_15907,N_12838,N_14439);
xor U15908 (N_15908,N_13531,N_13354);
nand U15909 (N_15909,N_13178,N_13914);
and U15910 (N_15910,N_13876,N_13409);
nand U15911 (N_15911,N_13194,N_12912);
nand U15912 (N_15912,N_14695,N_13244);
nand U15913 (N_15913,N_13816,N_14472);
or U15914 (N_15914,N_13695,N_14061);
and U15915 (N_15915,N_14652,N_13439);
or U15916 (N_15916,N_14862,N_14491);
nand U15917 (N_15917,N_14333,N_12984);
and U15918 (N_15918,N_14796,N_13011);
xor U15919 (N_15919,N_13540,N_14692);
or U15920 (N_15920,N_12704,N_14766);
xnor U15921 (N_15921,N_12716,N_13779);
and U15922 (N_15922,N_13580,N_13389);
nor U15923 (N_15923,N_13116,N_14600);
nor U15924 (N_15924,N_14289,N_13985);
nor U15925 (N_15925,N_12579,N_13281);
xnor U15926 (N_15926,N_13274,N_13280);
or U15927 (N_15927,N_13868,N_13411);
or U15928 (N_15928,N_13400,N_12788);
and U15929 (N_15929,N_13340,N_14092);
xor U15930 (N_15930,N_12697,N_12732);
nand U15931 (N_15931,N_14406,N_14137);
nand U15932 (N_15932,N_14009,N_12836);
or U15933 (N_15933,N_13346,N_13941);
and U15934 (N_15934,N_12872,N_14845);
and U15935 (N_15935,N_12848,N_12841);
nor U15936 (N_15936,N_13567,N_14529);
and U15937 (N_15937,N_14435,N_13546);
nand U15938 (N_15938,N_14097,N_14454);
nor U15939 (N_15939,N_13460,N_13585);
or U15940 (N_15940,N_12947,N_13234);
and U15941 (N_15941,N_12603,N_13933);
xor U15942 (N_15942,N_14839,N_13106);
nand U15943 (N_15943,N_12778,N_14110);
and U15944 (N_15944,N_12522,N_12910);
or U15945 (N_15945,N_13875,N_13795);
xnor U15946 (N_15946,N_14913,N_14199);
nand U15947 (N_15947,N_12631,N_13317);
nand U15948 (N_15948,N_13493,N_13563);
or U15949 (N_15949,N_12867,N_13060);
nand U15950 (N_15950,N_14118,N_12948);
nand U15951 (N_15951,N_14315,N_13199);
or U15952 (N_15952,N_14575,N_14954);
xor U15953 (N_15953,N_14572,N_14408);
and U15954 (N_15954,N_12860,N_12941);
xnor U15955 (N_15955,N_13784,N_14595);
nand U15956 (N_15956,N_14301,N_13173);
nand U15957 (N_15957,N_13813,N_14085);
nor U15958 (N_15958,N_14151,N_14246);
or U15959 (N_15959,N_14912,N_13598);
or U15960 (N_15960,N_13525,N_14663);
or U15961 (N_15961,N_12614,N_14010);
and U15962 (N_15962,N_14563,N_14822);
xor U15963 (N_15963,N_14283,N_14961);
or U15964 (N_15964,N_13573,N_13297);
xnor U15965 (N_15965,N_14307,N_13342);
nor U15966 (N_15966,N_12963,N_13566);
xnor U15967 (N_15967,N_12945,N_14101);
nand U15968 (N_15968,N_12641,N_14372);
nand U15969 (N_15969,N_13973,N_13539);
or U15970 (N_15970,N_12859,N_14208);
nor U15971 (N_15971,N_12715,N_13934);
and U15972 (N_15972,N_14782,N_13528);
xor U15973 (N_15973,N_14570,N_13714);
nor U15974 (N_15974,N_14823,N_12876);
nor U15975 (N_15975,N_14121,N_12792);
xnor U15976 (N_15976,N_14683,N_14568);
xor U15977 (N_15977,N_13463,N_13239);
nand U15978 (N_15978,N_13791,N_12943);
nand U15979 (N_15979,N_14715,N_13799);
nor U15980 (N_15980,N_14434,N_14757);
or U15981 (N_15981,N_13429,N_14375);
or U15982 (N_15982,N_12962,N_12512);
and U15983 (N_15983,N_12970,N_14179);
nand U15984 (N_15984,N_13724,N_13406);
and U15985 (N_15985,N_14932,N_13960);
nand U15986 (N_15986,N_14414,N_14418);
and U15987 (N_15987,N_12536,N_14669);
xor U15988 (N_15988,N_14382,N_12807);
and U15989 (N_15989,N_13249,N_14075);
and U15990 (N_15990,N_14036,N_13045);
xnor U15991 (N_15991,N_14363,N_14043);
and U15992 (N_15992,N_14741,N_14739);
nor U15993 (N_15993,N_12800,N_14041);
or U15994 (N_15994,N_13246,N_13235);
xor U15995 (N_15995,N_12904,N_12835);
and U15996 (N_15996,N_14534,N_14687);
or U15997 (N_15997,N_13198,N_14299);
nor U15998 (N_15998,N_14059,N_13307);
or U15999 (N_15999,N_13154,N_12577);
or U16000 (N_16000,N_12528,N_14538);
nand U16001 (N_16001,N_13096,N_12886);
nor U16002 (N_16002,N_13230,N_13905);
xnor U16003 (N_16003,N_12759,N_14390);
and U16004 (N_16004,N_14573,N_12622);
and U16005 (N_16005,N_14074,N_14353);
nor U16006 (N_16006,N_14817,N_12753);
and U16007 (N_16007,N_14478,N_12933);
or U16008 (N_16008,N_12601,N_13866);
nand U16009 (N_16009,N_12883,N_13132);
or U16010 (N_16010,N_14065,N_14229);
or U16011 (N_16011,N_13593,N_12829);
nor U16012 (N_16012,N_12647,N_13612);
or U16013 (N_16013,N_14067,N_14227);
and U16014 (N_16014,N_13543,N_13014);
xor U16015 (N_16015,N_14511,N_14159);
nand U16016 (N_16016,N_13026,N_13785);
and U16017 (N_16017,N_13975,N_12770);
nor U16018 (N_16018,N_14798,N_13981);
xor U16019 (N_16019,N_12561,N_14186);
or U16020 (N_16020,N_13316,N_14457);
nand U16021 (N_16021,N_14973,N_13511);
nor U16022 (N_16022,N_14224,N_14841);
nor U16023 (N_16023,N_14800,N_13373);
or U16024 (N_16024,N_13255,N_13955);
nor U16025 (N_16025,N_14432,N_13470);
xnor U16026 (N_16026,N_14596,N_14679);
nor U16027 (N_16027,N_14567,N_13608);
or U16028 (N_16028,N_14764,N_12646);
and U16029 (N_16029,N_12764,N_13071);
or U16030 (N_16030,N_13338,N_14341);
and U16031 (N_16031,N_13951,N_13643);
nand U16032 (N_16032,N_12965,N_14760);
nor U16033 (N_16033,N_14160,N_14013);
or U16034 (N_16034,N_14459,N_13616);
or U16035 (N_16035,N_14020,N_13165);
nor U16036 (N_16036,N_13938,N_12926);
xor U16037 (N_16037,N_14629,N_13482);
nor U16038 (N_16038,N_12989,N_13065);
or U16039 (N_16039,N_13718,N_13375);
nor U16040 (N_16040,N_14689,N_14477);
nand U16041 (N_16041,N_12505,N_14201);
and U16042 (N_16042,N_13569,N_14604);
nor U16043 (N_16043,N_13232,N_12929);
and U16044 (N_16044,N_14260,N_14673);
nand U16045 (N_16045,N_12649,N_14242);
nor U16046 (N_16046,N_14068,N_14320);
xnor U16047 (N_16047,N_14175,N_13467);
and U16048 (N_16048,N_14254,N_14339);
nand U16049 (N_16049,N_13819,N_14772);
nand U16050 (N_16050,N_13223,N_14937);
and U16051 (N_16051,N_13370,N_14243);
and U16052 (N_16052,N_13402,N_12991);
nand U16053 (N_16053,N_13284,N_13125);
nor U16054 (N_16054,N_13706,N_14182);
and U16055 (N_16055,N_13293,N_13308);
and U16056 (N_16056,N_13765,N_13123);
or U16057 (N_16057,N_14177,N_14238);
or U16058 (N_16058,N_14807,N_14753);
and U16059 (N_16059,N_14385,N_14759);
and U16060 (N_16060,N_13288,N_14536);
nor U16061 (N_16061,N_14416,N_13879);
and U16062 (N_16062,N_13465,N_14231);
nor U16063 (N_16063,N_14455,N_13742);
and U16064 (N_16064,N_13119,N_13343);
nand U16065 (N_16065,N_12712,N_13596);
or U16066 (N_16066,N_13601,N_14533);
and U16067 (N_16067,N_12758,N_13041);
nor U16068 (N_16068,N_13989,N_14203);
or U16069 (N_16069,N_13642,N_14327);
nor U16070 (N_16070,N_13335,N_12902);
nand U16071 (N_16071,N_13592,N_13832);
nor U16072 (N_16072,N_14540,N_13721);
nor U16073 (N_16073,N_13442,N_14783);
xor U16074 (N_16074,N_14153,N_13153);
nor U16075 (N_16075,N_13272,N_12590);
nor U16076 (N_16076,N_13691,N_12623);
xor U16077 (N_16077,N_13121,N_14497);
nor U16078 (N_16078,N_12952,N_13719);
xor U16079 (N_16079,N_13211,N_13443);
or U16080 (N_16080,N_14442,N_14721);
nor U16081 (N_16081,N_14502,N_14644);
xor U16082 (N_16082,N_13964,N_14088);
nor U16083 (N_16083,N_12520,N_13276);
or U16084 (N_16084,N_12824,N_13794);
xnor U16085 (N_16085,N_14387,N_12903);
xor U16086 (N_16086,N_13029,N_12762);
or U16087 (N_16087,N_13253,N_13847);
nand U16088 (N_16088,N_13943,N_14952);
nand U16089 (N_16089,N_14933,N_13644);
nor U16090 (N_16090,N_12946,N_14278);
xnor U16091 (N_16091,N_14864,N_14951);
and U16092 (N_16092,N_13672,N_14603);
nor U16093 (N_16093,N_12864,N_14486);
or U16094 (N_16094,N_13357,N_14893);
xnor U16095 (N_16095,N_13720,N_14244);
nand U16096 (N_16096,N_14094,N_14532);
and U16097 (N_16097,N_13219,N_12581);
and U16098 (N_16098,N_13661,N_14848);
nor U16099 (N_16099,N_13301,N_14710);
and U16100 (N_16100,N_13365,N_12849);
nand U16101 (N_16101,N_14880,N_14815);
nor U16102 (N_16102,N_13213,N_14365);
nor U16103 (N_16103,N_13728,N_14324);
and U16104 (N_16104,N_12744,N_13769);
xor U16105 (N_16105,N_13449,N_14245);
and U16106 (N_16106,N_13972,N_13817);
nand U16107 (N_16107,N_14440,N_14882);
xor U16108 (N_16108,N_14512,N_14461);
nor U16109 (N_16109,N_12668,N_13506);
nand U16110 (N_16110,N_13126,N_13761);
and U16111 (N_16111,N_14854,N_14905);
nor U16112 (N_16112,N_13560,N_14925);
or U16113 (N_16113,N_12743,N_13459);
xnor U16114 (N_16114,N_13073,N_13903);
nand U16115 (N_16115,N_12504,N_13291);
xor U16116 (N_16116,N_13758,N_13361);
nor U16117 (N_16117,N_14469,N_14584);
and U16118 (N_16118,N_14803,N_12846);
and U16119 (N_16119,N_14670,N_13859);
and U16120 (N_16120,N_12724,N_14034);
nor U16121 (N_16121,N_14792,N_12747);
and U16122 (N_16122,N_12922,N_12833);
xor U16123 (N_16123,N_14580,N_12961);
nor U16124 (N_16124,N_13845,N_12718);
nor U16125 (N_16125,N_14218,N_12752);
nand U16126 (N_16126,N_12548,N_14409);
or U16127 (N_16127,N_14451,N_13849);
and U16128 (N_16128,N_13044,N_14939);
xor U16129 (N_16129,N_13629,N_14132);
xor U16130 (N_16130,N_12618,N_13250);
or U16131 (N_16131,N_12688,N_14462);
nand U16132 (N_16132,N_12637,N_13362);
nor U16133 (N_16133,N_13871,N_13111);
and U16134 (N_16134,N_12843,N_13204);
nor U16135 (N_16135,N_13214,N_14624);
xnor U16136 (N_16136,N_14129,N_12573);
nand U16137 (N_16137,N_13913,N_13136);
xor U16138 (N_16138,N_13870,N_13383);
nand U16139 (N_16139,N_12735,N_12906);
or U16140 (N_16140,N_12656,N_12974);
nand U16141 (N_16141,N_14071,N_13651);
nor U16142 (N_16142,N_12602,N_13146);
or U16143 (N_16143,N_14276,N_13874);
nor U16144 (N_16144,N_14978,N_14261);
nand U16145 (N_16145,N_13048,N_12638);
or U16146 (N_16146,N_14700,N_13731);
nand U16147 (N_16147,N_14103,N_14145);
nor U16148 (N_16148,N_14398,N_13811);
nand U16149 (N_16149,N_13067,N_13254);
nand U16150 (N_16150,N_14582,N_14360);
nand U16151 (N_16151,N_13187,N_13853);
nor U16152 (N_16152,N_13056,N_13694);
nand U16153 (N_16153,N_13102,N_13263);
or U16154 (N_16154,N_14945,N_13507);
and U16155 (N_16155,N_12931,N_13499);
nor U16156 (N_16156,N_14077,N_14950);
nor U16157 (N_16157,N_14777,N_14484);
nor U16158 (N_16158,N_14128,N_14308);
and U16159 (N_16159,N_14112,N_12584);
xor U16160 (N_16160,N_14850,N_14106);
nor U16161 (N_16161,N_13808,N_14664);
nor U16162 (N_16162,N_13918,N_13804);
nand U16163 (N_16163,N_14271,N_13471);
or U16164 (N_16164,N_13793,N_13390);
nor U16165 (N_16165,N_14374,N_13895);
nor U16166 (N_16166,N_14483,N_14060);
xnor U16167 (N_16167,N_14955,N_14475);
nand U16168 (N_16168,N_13150,N_14423);
nand U16169 (N_16169,N_13105,N_14189);
nand U16170 (N_16170,N_13880,N_12769);
nor U16171 (N_16171,N_12717,N_13490);
or U16172 (N_16172,N_14292,N_13182);
xnor U16173 (N_16173,N_13542,N_12760);
xnor U16174 (N_16174,N_14142,N_13839);
nand U16175 (N_16175,N_12969,N_14607);
or U16176 (N_16176,N_14888,N_13436);
xnor U16177 (N_16177,N_14209,N_13949);
nand U16178 (N_16178,N_13739,N_13396);
nand U16179 (N_16179,N_14395,N_13564);
xnor U16180 (N_16180,N_13524,N_12934);
or U16181 (N_16181,N_13445,N_12847);
xor U16182 (N_16182,N_13318,N_12671);
xnor U16183 (N_16183,N_14517,N_14140);
or U16184 (N_16184,N_13124,N_14690);
or U16185 (N_16185,N_13788,N_13176);
and U16186 (N_16186,N_14745,N_14623);
and U16187 (N_16187,N_14072,N_14096);
xor U16188 (N_16188,N_14062,N_13152);
xnor U16189 (N_16189,N_14220,N_14274);
nand U16190 (N_16190,N_14842,N_13260);
nor U16191 (N_16191,N_14127,N_12534);
and U16192 (N_16192,N_13556,N_14389);
xnor U16193 (N_16193,N_12978,N_13017);
xor U16194 (N_16194,N_14787,N_12882);
nand U16195 (N_16195,N_14887,N_14726);
nand U16196 (N_16196,N_14190,N_13222);
and U16197 (N_16197,N_13033,N_14859);
nand U16198 (N_16198,N_13891,N_14617);
or U16199 (N_16199,N_14921,N_14648);
and U16200 (N_16200,N_13087,N_13978);
nor U16201 (N_16201,N_14079,N_13750);
or U16202 (N_16202,N_13946,N_12813);
and U16203 (N_16203,N_12909,N_13310);
xnor U16204 (N_16204,N_13658,N_14675);
xor U16205 (N_16205,N_14286,N_12865);
nand U16206 (N_16206,N_13468,N_12795);
or U16207 (N_16207,N_12719,N_12983);
or U16208 (N_16208,N_13856,N_13834);
or U16209 (N_16209,N_13953,N_14498);
nor U16210 (N_16210,N_13707,N_12517);
nor U16211 (N_16211,N_14235,N_14917);
xor U16212 (N_16212,N_12615,N_12625);
nor U16213 (N_16213,N_13398,N_14641);
nor U16214 (N_16214,N_14050,N_12657);
xnor U16215 (N_16215,N_14487,N_12639);
nor U16216 (N_16216,N_13051,N_13036);
xor U16217 (N_16217,N_12725,N_12810);
xor U16218 (N_16218,N_13113,N_12749);
xor U16219 (N_16219,N_14749,N_13079);
nand U16220 (N_16220,N_14134,N_13961);
nor U16221 (N_16221,N_14665,N_13115);
nor U16222 (N_16222,N_14832,N_13076);
xor U16223 (N_16223,N_13984,N_13066);
xor U16224 (N_16224,N_12855,N_14535);
or U16225 (N_16225,N_13327,N_14926);
and U16226 (N_16226,N_14702,N_14168);
nor U16227 (N_16227,N_12582,N_12990);
and U16228 (N_16228,N_13805,N_14752);
xnor U16229 (N_16229,N_14212,N_14004);
nand U16230 (N_16230,N_13636,N_14707);
xor U16231 (N_16231,N_14204,N_14769);
or U16232 (N_16232,N_14812,N_14187);
nor U16233 (N_16233,N_14984,N_14257);
xnor U16234 (N_16234,N_14282,N_14474);
xor U16235 (N_16235,N_14496,N_13738);
or U16236 (N_16236,N_13798,N_13726);
and U16237 (N_16237,N_12742,N_13743);
nand U16238 (N_16238,N_13823,N_14948);
nand U16239 (N_16239,N_14686,N_13713);
and U16240 (N_16240,N_12817,N_14691);
and U16241 (N_16241,N_14649,N_14610);
or U16242 (N_16242,N_13690,N_13982);
xor U16243 (N_16243,N_12861,N_14479);
xor U16244 (N_16244,N_13210,N_14576);
xnor U16245 (N_16245,N_14814,N_13510);
and U16246 (N_16246,N_12642,N_14037);
nor U16247 (N_16247,N_14028,N_13772);
xor U16248 (N_16248,N_13917,N_13050);
or U16249 (N_16249,N_12530,N_12511);
nor U16250 (N_16250,N_13712,N_12698);
and U16251 (N_16251,N_14418,N_14460);
nand U16252 (N_16252,N_14619,N_14220);
or U16253 (N_16253,N_12827,N_14340);
nand U16254 (N_16254,N_13883,N_13479);
and U16255 (N_16255,N_14410,N_14898);
and U16256 (N_16256,N_13139,N_14401);
nand U16257 (N_16257,N_13777,N_13784);
nor U16258 (N_16258,N_14374,N_12537);
xor U16259 (N_16259,N_14377,N_12645);
xor U16260 (N_16260,N_13520,N_12679);
nand U16261 (N_16261,N_13801,N_14501);
nor U16262 (N_16262,N_13474,N_12595);
or U16263 (N_16263,N_12826,N_13035);
xor U16264 (N_16264,N_13880,N_13591);
nand U16265 (N_16265,N_14721,N_14513);
or U16266 (N_16266,N_14424,N_12899);
or U16267 (N_16267,N_14946,N_13611);
or U16268 (N_16268,N_13588,N_13681);
nor U16269 (N_16269,N_14059,N_12618);
nand U16270 (N_16270,N_13185,N_13511);
xor U16271 (N_16271,N_13559,N_14364);
and U16272 (N_16272,N_14934,N_12505);
and U16273 (N_16273,N_12945,N_14700);
and U16274 (N_16274,N_12569,N_13023);
and U16275 (N_16275,N_12751,N_13496);
nor U16276 (N_16276,N_13196,N_14290);
nor U16277 (N_16277,N_13237,N_12667);
or U16278 (N_16278,N_14418,N_12515);
nand U16279 (N_16279,N_14285,N_14305);
nor U16280 (N_16280,N_12850,N_12525);
nand U16281 (N_16281,N_14883,N_13977);
and U16282 (N_16282,N_14956,N_12565);
nor U16283 (N_16283,N_13841,N_13567);
and U16284 (N_16284,N_12948,N_13788);
or U16285 (N_16285,N_13616,N_14299);
and U16286 (N_16286,N_14161,N_13711);
nand U16287 (N_16287,N_13212,N_13879);
nand U16288 (N_16288,N_13393,N_14870);
nor U16289 (N_16289,N_13932,N_12745);
xnor U16290 (N_16290,N_13285,N_14385);
nand U16291 (N_16291,N_13621,N_14849);
nand U16292 (N_16292,N_13526,N_14729);
nor U16293 (N_16293,N_14565,N_12947);
or U16294 (N_16294,N_14543,N_12828);
or U16295 (N_16295,N_13002,N_14644);
xnor U16296 (N_16296,N_14512,N_14193);
nand U16297 (N_16297,N_13767,N_14486);
or U16298 (N_16298,N_12670,N_13302);
and U16299 (N_16299,N_13619,N_13676);
nand U16300 (N_16300,N_14155,N_13225);
or U16301 (N_16301,N_13987,N_14939);
or U16302 (N_16302,N_13520,N_13662);
xor U16303 (N_16303,N_13777,N_14369);
nor U16304 (N_16304,N_14565,N_14264);
nor U16305 (N_16305,N_14046,N_14195);
and U16306 (N_16306,N_12663,N_13720);
and U16307 (N_16307,N_12925,N_12666);
and U16308 (N_16308,N_14157,N_14049);
nor U16309 (N_16309,N_14568,N_13164);
and U16310 (N_16310,N_13288,N_14291);
and U16311 (N_16311,N_14232,N_14087);
nor U16312 (N_16312,N_14795,N_13494);
or U16313 (N_16313,N_14453,N_12571);
nor U16314 (N_16314,N_14470,N_14793);
xor U16315 (N_16315,N_13048,N_12646);
or U16316 (N_16316,N_14501,N_14946);
nor U16317 (N_16317,N_13277,N_14288);
nor U16318 (N_16318,N_14951,N_14771);
xor U16319 (N_16319,N_14204,N_14326);
nand U16320 (N_16320,N_13682,N_13760);
nor U16321 (N_16321,N_13602,N_13169);
and U16322 (N_16322,N_13440,N_14524);
and U16323 (N_16323,N_13444,N_13118);
or U16324 (N_16324,N_13835,N_14467);
xnor U16325 (N_16325,N_12951,N_13612);
and U16326 (N_16326,N_13051,N_14535);
nor U16327 (N_16327,N_12910,N_14637);
xor U16328 (N_16328,N_14501,N_12526);
or U16329 (N_16329,N_13930,N_13502);
nand U16330 (N_16330,N_14724,N_13585);
nand U16331 (N_16331,N_12944,N_13944);
nand U16332 (N_16332,N_14937,N_12754);
xor U16333 (N_16333,N_14136,N_14454);
nand U16334 (N_16334,N_13612,N_14130);
or U16335 (N_16335,N_12587,N_13972);
nand U16336 (N_16336,N_13683,N_14003);
or U16337 (N_16337,N_14811,N_13486);
nand U16338 (N_16338,N_13098,N_14477);
and U16339 (N_16339,N_13503,N_13115);
xnor U16340 (N_16340,N_12895,N_13135);
nand U16341 (N_16341,N_14552,N_14765);
xnor U16342 (N_16342,N_14535,N_13794);
xor U16343 (N_16343,N_13312,N_13562);
xnor U16344 (N_16344,N_14534,N_12848);
or U16345 (N_16345,N_14226,N_13085);
and U16346 (N_16346,N_13299,N_13520);
or U16347 (N_16347,N_14463,N_13900);
nand U16348 (N_16348,N_14671,N_13243);
or U16349 (N_16349,N_12658,N_13861);
or U16350 (N_16350,N_13050,N_12840);
or U16351 (N_16351,N_14841,N_13766);
nor U16352 (N_16352,N_13180,N_12820);
nor U16353 (N_16353,N_14865,N_14622);
or U16354 (N_16354,N_14770,N_13410);
or U16355 (N_16355,N_14848,N_12734);
xnor U16356 (N_16356,N_12551,N_14364);
and U16357 (N_16357,N_13300,N_13462);
or U16358 (N_16358,N_14239,N_13426);
or U16359 (N_16359,N_14950,N_13106);
and U16360 (N_16360,N_14350,N_12770);
or U16361 (N_16361,N_14832,N_12556);
xnor U16362 (N_16362,N_13427,N_12594);
or U16363 (N_16363,N_12555,N_13985);
nand U16364 (N_16364,N_14865,N_13945);
nor U16365 (N_16365,N_12600,N_14392);
and U16366 (N_16366,N_13166,N_12984);
nand U16367 (N_16367,N_12920,N_12661);
and U16368 (N_16368,N_13982,N_13326);
nand U16369 (N_16369,N_13260,N_14848);
or U16370 (N_16370,N_14087,N_14909);
and U16371 (N_16371,N_14980,N_12843);
xnor U16372 (N_16372,N_12758,N_13039);
nand U16373 (N_16373,N_14636,N_12670);
nand U16374 (N_16374,N_12748,N_14680);
xor U16375 (N_16375,N_13166,N_14246);
xnor U16376 (N_16376,N_14501,N_12586);
nand U16377 (N_16377,N_14689,N_13264);
xor U16378 (N_16378,N_14932,N_14879);
nand U16379 (N_16379,N_14463,N_14752);
nand U16380 (N_16380,N_13207,N_13768);
nor U16381 (N_16381,N_14038,N_14450);
nor U16382 (N_16382,N_12554,N_14883);
xor U16383 (N_16383,N_14218,N_12537);
and U16384 (N_16384,N_13393,N_13296);
xor U16385 (N_16385,N_13793,N_14451);
xor U16386 (N_16386,N_12816,N_13664);
nand U16387 (N_16387,N_13000,N_12659);
xor U16388 (N_16388,N_14221,N_13387);
xor U16389 (N_16389,N_14120,N_13763);
nand U16390 (N_16390,N_13293,N_13809);
and U16391 (N_16391,N_14255,N_14977);
nand U16392 (N_16392,N_13037,N_13603);
and U16393 (N_16393,N_12887,N_12971);
xor U16394 (N_16394,N_13912,N_12795);
or U16395 (N_16395,N_14903,N_12947);
nand U16396 (N_16396,N_12854,N_14144);
nor U16397 (N_16397,N_14683,N_14859);
and U16398 (N_16398,N_14114,N_12714);
nor U16399 (N_16399,N_12644,N_14028);
and U16400 (N_16400,N_14104,N_14246);
nand U16401 (N_16401,N_13071,N_14262);
or U16402 (N_16402,N_12632,N_13113);
xor U16403 (N_16403,N_13750,N_14013);
nor U16404 (N_16404,N_13027,N_13196);
xnor U16405 (N_16405,N_14901,N_12724);
nand U16406 (N_16406,N_14293,N_13617);
or U16407 (N_16407,N_13231,N_13131);
xnor U16408 (N_16408,N_13814,N_13695);
xor U16409 (N_16409,N_13121,N_12681);
xnor U16410 (N_16410,N_14213,N_14719);
and U16411 (N_16411,N_14751,N_13733);
or U16412 (N_16412,N_13476,N_12614);
and U16413 (N_16413,N_12650,N_14770);
nor U16414 (N_16414,N_14025,N_12506);
nor U16415 (N_16415,N_12786,N_14820);
or U16416 (N_16416,N_13652,N_13373);
nor U16417 (N_16417,N_13661,N_12845);
nor U16418 (N_16418,N_14416,N_13842);
xor U16419 (N_16419,N_14566,N_12652);
nand U16420 (N_16420,N_12899,N_12592);
and U16421 (N_16421,N_13766,N_14654);
nor U16422 (N_16422,N_13479,N_13862);
nand U16423 (N_16423,N_13807,N_14934);
nand U16424 (N_16424,N_13824,N_14824);
xor U16425 (N_16425,N_13374,N_14602);
and U16426 (N_16426,N_14607,N_14219);
nand U16427 (N_16427,N_13867,N_13873);
nor U16428 (N_16428,N_13856,N_13683);
and U16429 (N_16429,N_13518,N_14622);
xor U16430 (N_16430,N_12644,N_13204);
nand U16431 (N_16431,N_13383,N_14771);
xor U16432 (N_16432,N_12637,N_13052);
and U16433 (N_16433,N_12932,N_13753);
xnor U16434 (N_16434,N_13818,N_14984);
xnor U16435 (N_16435,N_13839,N_14876);
xor U16436 (N_16436,N_14262,N_13302);
xnor U16437 (N_16437,N_13379,N_14809);
nand U16438 (N_16438,N_14438,N_13078);
or U16439 (N_16439,N_14221,N_14301);
and U16440 (N_16440,N_13906,N_14336);
nand U16441 (N_16441,N_14289,N_14373);
nor U16442 (N_16442,N_14716,N_12804);
nand U16443 (N_16443,N_14110,N_12658);
xor U16444 (N_16444,N_13299,N_13060);
and U16445 (N_16445,N_14712,N_14684);
or U16446 (N_16446,N_14166,N_13460);
nand U16447 (N_16447,N_14777,N_14252);
nand U16448 (N_16448,N_12979,N_13235);
xor U16449 (N_16449,N_12717,N_14932);
xor U16450 (N_16450,N_12846,N_14170);
nor U16451 (N_16451,N_13859,N_13027);
or U16452 (N_16452,N_14891,N_13719);
nor U16453 (N_16453,N_14095,N_14358);
or U16454 (N_16454,N_14134,N_13924);
nand U16455 (N_16455,N_13329,N_13446);
and U16456 (N_16456,N_13515,N_14077);
nand U16457 (N_16457,N_12600,N_13376);
xnor U16458 (N_16458,N_13118,N_14692);
or U16459 (N_16459,N_14397,N_14200);
xor U16460 (N_16460,N_12788,N_13510);
xor U16461 (N_16461,N_13077,N_12763);
xnor U16462 (N_16462,N_14743,N_14291);
xnor U16463 (N_16463,N_12637,N_14081);
nand U16464 (N_16464,N_12835,N_13040);
xor U16465 (N_16465,N_14685,N_12746);
nand U16466 (N_16466,N_13312,N_14047);
nand U16467 (N_16467,N_14286,N_13240);
nand U16468 (N_16468,N_14209,N_12798);
xor U16469 (N_16469,N_13265,N_14891);
nand U16470 (N_16470,N_14154,N_14034);
xnor U16471 (N_16471,N_13250,N_14981);
nor U16472 (N_16472,N_12785,N_13286);
xnor U16473 (N_16473,N_12516,N_13239);
nor U16474 (N_16474,N_13334,N_13074);
xor U16475 (N_16475,N_14985,N_13518);
nand U16476 (N_16476,N_13065,N_13952);
or U16477 (N_16477,N_14753,N_14313);
nand U16478 (N_16478,N_12954,N_13320);
or U16479 (N_16479,N_14989,N_13901);
nor U16480 (N_16480,N_13405,N_14798);
nor U16481 (N_16481,N_13129,N_14131);
nand U16482 (N_16482,N_14102,N_13372);
xor U16483 (N_16483,N_14608,N_14421);
or U16484 (N_16484,N_14309,N_13223);
nor U16485 (N_16485,N_13374,N_14823);
xor U16486 (N_16486,N_14580,N_14847);
and U16487 (N_16487,N_12933,N_14654);
nand U16488 (N_16488,N_14425,N_14718);
or U16489 (N_16489,N_12558,N_14505);
or U16490 (N_16490,N_14376,N_14147);
and U16491 (N_16491,N_12983,N_14718);
nor U16492 (N_16492,N_14213,N_13977);
nand U16493 (N_16493,N_14952,N_14970);
or U16494 (N_16494,N_14372,N_13004);
or U16495 (N_16495,N_13154,N_12814);
nor U16496 (N_16496,N_14437,N_12899);
or U16497 (N_16497,N_12615,N_13994);
nand U16498 (N_16498,N_12858,N_14566);
nand U16499 (N_16499,N_13360,N_13549);
or U16500 (N_16500,N_13122,N_12516);
and U16501 (N_16501,N_14207,N_13402);
xor U16502 (N_16502,N_13919,N_13943);
nand U16503 (N_16503,N_13879,N_14539);
or U16504 (N_16504,N_14582,N_14755);
nor U16505 (N_16505,N_13337,N_14936);
nor U16506 (N_16506,N_14234,N_13785);
nand U16507 (N_16507,N_12758,N_14530);
xnor U16508 (N_16508,N_12989,N_13368);
nor U16509 (N_16509,N_14607,N_14776);
xnor U16510 (N_16510,N_13027,N_14305);
or U16511 (N_16511,N_14827,N_14078);
and U16512 (N_16512,N_12524,N_12698);
and U16513 (N_16513,N_12887,N_12525);
nor U16514 (N_16514,N_13389,N_14191);
nand U16515 (N_16515,N_14880,N_13679);
xor U16516 (N_16516,N_14379,N_14545);
nor U16517 (N_16517,N_14804,N_12976);
xnor U16518 (N_16518,N_14228,N_13332);
nand U16519 (N_16519,N_12744,N_12788);
nor U16520 (N_16520,N_13058,N_13266);
nor U16521 (N_16521,N_13438,N_13088);
nor U16522 (N_16522,N_13131,N_12890);
or U16523 (N_16523,N_13991,N_12550);
or U16524 (N_16524,N_14607,N_14397);
xor U16525 (N_16525,N_12790,N_14774);
xor U16526 (N_16526,N_14817,N_13910);
xor U16527 (N_16527,N_14007,N_13655);
or U16528 (N_16528,N_14286,N_14188);
nand U16529 (N_16529,N_14222,N_14164);
or U16530 (N_16530,N_13048,N_14090);
or U16531 (N_16531,N_13307,N_12520);
and U16532 (N_16532,N_13858,N_13663);
nand U16533 (N_16533,N_13054,N_14167);
nor U16534 (N_16534,N_12512,N_14525);
or U16535 (N_16535,N_13028,N_13645);
xnor U16536 (N_16536,N_14776,N_14018);
or U16537 (N_16537,N_13597,N_12878);
xnor U16538 (N_16538,N_14723,N_13481);
or U16539 (N_16539,N_14564,N_13665);
nor U16540 (N_16540,N_12585,N_13779);
nand U16541 (N_16541,N_14126,N_14699);
xor U16542 (N_16542,N_14979,N_13851);
and U16543 (N_16543,N_13410,N_13310);
xnor U16544 (N_16544,N_13297,N_12559);
and U16545 (N_16545,N_14665,N_13036);
and U16546 (N_16546,N_12705,N_12577);
nor U16547 (N_16547,N_13046,N_14171);
nand U16548 (N_16548,N_12889,N_12756);
and U16549 (N_16549,N_13359,N_14444);
nor U16550 (N_16550,N_13006,N_12800);
or U16551 (N_16551,N_13336,N_12823);
nand U16552 (N_16552,N_13905,N_13671);
or U16553 (N_16553,N_14561,N_12709);
nor U16554 (N_16554,N_13014,N_13549);
nor U16555 (N_16555,N_14317,N_14146);
or U16556 (N_16556,N_14123,N_14109);
and U16557 (N_16557,N_14567,N_14547);
and U16558 (N_16558,N_14026,N_13825);
xnor U16559 (N_16559,N_14807,N_12827);
xnor U16560 (N_16560,N_14474,N_13730);
nand U16561 (N_16561,N_13326,N_13679);
and U16562 (N_16562,N_12590,N_13842);
or U16563 (N_16563,N_13144,N_14620);
xnor U16564 (N_16564,N_14022,N_14452);
or U16565 (N_16565,N_13765,N_13674);
nor U16566 (N_16566,N_12519,N_14169);
nand U16567 (N_16567,N_14626,N_14049);
or U16568 (N_16568,N_13394,N_14930);
nor U16569 (N_16569,N_14617,N_13464);
nor U16570 (N_16570,N_13569,N_14042);
and U16571 (N_16571,N_13152,N_12921);
xor U16572 (N_16572,N_13451,N_13498);
nand U16573 (N_16573,N_14048,N_14686);
and U16574 (N_16574,N_13507,N_12764);
or U16575 (N_16575,N_14082,N_14288);
nor U16576 (N_16576,N_13822,N_12904);
nand U16577 (N_16577,N_13156,N_12572);
nor U16578 (N_16578,N_13229,N_14323);
nand U16579 (N_16579,N_13821,N_12914);
and U16580 (N_16580,N_13423,N_14949);
or U16581 (N_16581,N_14861,N_14367);
and U16582 (N_16582,N_14683,N_13803);
or U16583 (N_16583,N_14073,N_14308);
or U16584 (N_16584,N_13553,N_13131);
and U16585 (N_16585,N_12863,N_13628);
xnor U16586 (N_16586,N_14745,N_14097);
nor U16587 (N_16587,N_14039,N_13145);
nand U16588 (N_16588,N_14203,N_14858);
nand U16589 (N_16589,N_13349,N_14457);
nor U16590 (N_16590,N_13387,N_13454);
nor U16591 (N_16591,N_14212,N_13131);
nand U16592 (N_16592,N_14835,N_13584);
xnor U16593 (N_16593,N_13987,N_14978);
nand U16594 (N_16594,N_12757,N_12741);
nor U16595 (N_16595,N_13566,N_12829);
xor U16596 (N_16596,N_12991,N_14700);
or U16597 (N_16597,N_14728,N_13832);
and U16598 (N_16598,N_14993,N_14127);
or U16599 (N_16599,N_14576,N_14917);
and U16600 (N_16600,N_14788,N_12861);
or U16601 (N_16601,N_14615,N_14433);
or U16602 (N_16602,N_13464,N_14318);
nor U16603 (N_16603,N_14300,N_14834);
xnor U16604 (N_16604,N_12876,N_14041);
and U16605 (N_16605,N_13089,N_14802);
and U16606 (N_16606,N_13065,N_13764);
xor U16607 (N_16607,N_13601,N_13390);
nor U16608 (N_16608,N_14369,N_14045);
or U16609 (N_16609,N_13366,N_12899);
and U16610 (N_16610,N_14897,N_13431);
xor U16611 (N_16611,N_13061,N_12800);
nor U16612 (N_16612,N_13321,N_14763);
xor U16613 (N_16613,N_13354,N_14078);
or U16614 (N_16614,N_14057,N_12946);
nor U16615 (N_16615,N_13066,N_13957);
nand U16616 (N_16616,N_12822,N_12880);
nand U16617 (N_16617,N_12903,N_13888);
nor U16618 (N_16618,N_13456,N_12555);
or U16619 (N_16619,N_13401,N_13767);
xnor U16620 (N_16620,N_13788,N_13130);
or U16621 (N_16621,N_13400,N_14655);
nor U16622 (N_16622,N_13487,N_13875);
or U16623 (N_16623,N_13209,N_14877);
nor U16624 (N_16624,N_13819,N_14683);
and U16625 (N_16625,N_12547,N_13141);
nand U16626 (N_16626,N_14213,N_14437);
and U16627 (N_16627,N_14705,N_14288);
and U16628 (N_16628,N_14417,N_14975);
and U16629 (N_16629,N_13110,N_13890);
or U16630 (N_16630,N_12700,N_14465);
xnor U16631 (N_16631,N_14563,N_12998);
nor U16632 (N_16632,N_13425,N_13626);
nand U16633 (N_16633,N_14111,N_14456);
nor U16634 (N_16634,N_14276,N_14699);
and U16635 (N_16635,N_14061,N_14032);
nor U16636 (N_16636,N_14401,N_13452);
nor U16637 (N_16637,N_14710,N_14285);
nand U16638 (N_16638,N_14749,N_13021);
xor U16639 (N_16639,N_13316,N_14955);
xnor U16640 (N_16640,N_14397,N_12601);
nand U16641 (N_16641,N_14582,N_13262);
and U16642 (N_16642,N_14728,N_14834);
nand U16643 (N_16643,N_13916,N_12574);
xnor U16644 (N_16644,N_13813,N_14449);
and U16645 (N_16645,N_12892,N_14895);
nor U16646 (N_16646,N_14436,N_12920);
nand U16647 (N_16647,N_13397,N_14414);
or U16648 (N_16648,N_13518,N_13230);
or U16649 (N_16649,N_13373,N_12746);
nor U16650 (N_16650,N_14956,N_12829);
nand U16651 (N_16651,N_12534,N_14533);
and U16652 (N_16652,N_13915,N_14697);
xnor U16653 (N_16653,N_13134,N_13513);
nand U16654 (N_16654,N_13107,N_12543);
and U16655 (N_16655,N_13545,N_13276);
or U16656 (N_16656,N_12723,N_13774);
nand U16657 (N_16657,N_14069,N_14037);
xnor U16658 (N_16658,N_12861,N_12978);
nand U16659 (N_16659,N_14160,N_14168);
nor U16660 (N_16660,N_13176,N_14091);
nand U16661 (N_16661,N_14949,N_12883);
xnor U16662 (N_16662,N_12508,N_13577);
or U16663 (N_16663,N_14825,N_12922);
or U16664 (N_16664,N_13391,N_14472);
xor U16665 (N_16665,N_12627,N_13453);
or U16666 (N_16666,N_13936,N_12882);
xor U16667 (N_16667,N_14265,N_13307);
or U16668 (N_16668,N_14836,N_12738);
nand U16669 (N_16669,N_14753,N_13772);
nand U16670 (N_16670,N_14291,N_13552);
xor U16671 (N_16671,N_12776,N_13894);
nand U16672 (N_16672,N_14007,N_14561);
nand U16673 (N_16673,N_13083,N_13514);
or U16674 (N_16674,N_13410,N_12851);
xnor U16675 (N_16675,N_13135,N_13116);
xor U16676 (N_16676,N_12937,N_13228);
nor U16677 (N_16677,N_13053,N_13373);
nand U16678 (N_16678,N_12564,N_13743);
xor U16679 (N_16679,N_12606,N_13154);
nor U16680 (N_16680,N_14749,N_13546);
xor U16681 (N_16681,N_14647,N_13474);
nand U16682 (N_16682,N_14642,N_13298);
or U16683 (N_16683,N_12646,N_14796);
nand U16684 (N_16684,N_13190,N_12670);
or U16685 (N_16685,N_12959,N_12955);
xor U16686 (N_16686,N_13937,N_14543);
nor U16687 (N_16687,N_13081,N_12833);
or U16688 (N_16688,N_12970,N_13243);
nand U16689 (N_16689,N_12813,N_13252);
nor U16690 (N_16690,N_14919,N_12757);
xnor U16691 (N_16691,N_13502,N_13397);
nor U16692 (N_16692,N_14460,N_14350);
or U16693 (N_16693,N_13110,N_12511);
nand U16694 (N_16694,N_14692,N_13566);
xor U16695 (N_16695,N_13136,N_13954);
and U16696 (N_16696,N_13709,N_12701);
xor U16697 (N_16697,N_14911,N_12667);
and U16698 (N_16698,N_14078,N_13876);
or U16699 (N_16699,N_13985,N_12832);
xor U16700 (N_16700,N_13089,N_13348);
or U16701 (N_16701,N_12531,N_13933);
nand U16702 (N_16702,N_13497,N_14602);
nor U16703 (N_16703,N_12524,N_13421);
nor U16704 (N_16704,N_13412,N_14429);
xnor U16705 (N_16705,N_13352,N_13056);
xnor U16706 (N_16706,N_13158,N_13648);
or U16707 (N_16707,N_13512,N_12571);
or U16708 (N_16708,N_14570,N_13597);
nand U16709 (N_16709,N_14697,N_13179);
nand U16710 (N_16710,N_13425,N_13647);
or U16711 (N_16711,N_14074,N_14327);
xor U16712 (N_16712,N_14025,N_12805);
nor U16713 (N_16713,N_13750,N_13667);
nor U16714 (N_16714,N_14430,N_14192);
xor U16715 (N_16715,N_14141,N_14770);
or U16716 (N_16716,N_14687,N_13756);
and U16717 (N_16717,N_14613,N_14701);
xor U16718 (N_16718,N_13906,N_14636);
or U16719 (N_16719,N_14869,N_13585);
nand U16720 (N_16720,N_12787,N_14652);
nor U16721 (N_16721,N_12963,N_13934);
nand U16722 (N_16722,N_13245,N_13576);
nor U16723 (N_16723,N_14695,N_13050);
xnor U16724 (N_16724,N_13647,N_13173);
nor U16725 (N_16725,N_14300,N_12829);
xnor U16726 (N_16726,N_12819,N_14927);
nand U16727 (N_16727,N_12910,N_13159);
nand U16728 (N_16728,N_14459,N_14490);
and U16729 (N_16729,N_13804,N_14616);
nand U16730 (N_16730,N_14712,N_14928);
xor U16731 (N_16731,N_12570,N_12984);
and U16732 (N_16732,N_14913,N_14225);
nor U16733 (N_16733,N_14013,N_14392);
and U16734 (N_16734,N_12950,N_14529);
xor U16735 (N_16735,N_14090,N_13082);
nand U16736 (N_16736,N_12938,N_13031);
and U16737 (N_16737,N_14740,N_14427);
and U16738 (N_16738,N_13320,N_14561);
nor U16739 (N_16739,N_14387,N_14017);
xor U16740 (N_16740,N_13444,N_13090);
or U16741 (N_16741,N_13248,N_13913);
nor U16742 (N_16742,N_13064,N_12914);
nand U16743 (N_16743,N_13124,N_13363);
and U16744 (N_16744,N_14233,N_14144);
xor U16745 (N_16745,N_13314,N_13903);
nor U16746 (N_16746,N_12824,N_14385);
nand U16747 (N_16747,N_12784,N_13106);
or U16748 (N_16748,N_13048,N_14284);
nor U16749 (N_16749,N_13212,N_13806);
xnor U16750 (N_16750,N_12662,N_13727);
xor U16751 (N_16751,N_13175,N_13531);
and U16752 (N_16752,N_14980,N_12585);
and U16753 (N_16753,N_13948,N_13082);
xnor U16754 (N_16754,N_13068,N_12823);
and U16755 (N_16755,N_14641,N_12753);
or U16756 (N_16756,N_14913,N_14943);
nor U16757 (N_16757,N_12556,N_13283);
and U16758 (N_16758,N_14259,N_13758);
and U16759 (N_16759,N_13205,N_13269);
nand U16760 (N_16760,N_14982,N_14026);
and U16761 (N_16761,N_14668,N_13907);
nand U16762 (N_16762,N_13946,N_14803);
or U16763 (N_16763,N_12828,N_14965);
nand U16764 (N_16764,N_13345,N_12535);
or U16765 (N_16765,N_13413,N_13302);
nor U16766 (N_16766,N_14232,N_13302);
nor U16767 (N_16767,N_14510,N_12610);
or U16768 (N_16768,N_13876,N_13349);
nand U16769 (N_16769,N_13716,N_14802);
xnor U16770 (N_16770,N_12737,N_14905);
nand U16771 (N_16771,N_13995,N_12624);
or U16772 (N_16772,N_12547,N_14032);
nand U16773 (N_16773,N_14538,N_12833);
and U16774 (N_16774,N_12569,N_12604);
and U16775 (N_16775,N_13578,N_13227);
xnor U16776 (N_16776,N_14899,N_13323);
nor U16777 (N_16777,N_13595,N_14165);
nand U16778 (N_16778,N_13601,N_14528);
xor U16779 (N_16779,N_14536,N_12756);
nand U16780 (N_16780,N_14112,N_12707);
xnor U16781 (N_16781,N_12995,N_12785);
or U16782 (N_16782,N_12767,N_13603);
nor U16783 (N_16783,N_14355,N_14784);
and U16784 (N_16784,N_14816,N_14143);
and U16785 (N_16785,N_14717,N_12710);
xor U16786 (N_16786,N_13738,N_14324);
or U16787 (N_16787,N_13511,N_12638);
or U16788 (N_16788,N_13336,N_13684);
nand U16789 (N_16789,N_12656,N_14751);
xor U16790 (N_16790,N_12648,N_14768);
nor U16791 (N_16791,N_14584,N_14101);
nor U16792 (N_16792,N_14894,N_13207);
nand U16793 (N_16793,N_12846,N_14829);
and U16794 (N_16794,N_14887,N_14928);
and U16795 (N_16795,N_12876,N_12594);
nand U16796 (N_16796,N_13034,N_13700);
nand U16797 (N_16797,N_14481,N_13208);
or U16798 (N_16798,N_12656,N_13213);
or U16799 (N_16799,N_12597,N_12542);
and U16800 (N_16800,N_13614,N_13592);
nand U16801 (N_16801,N_14442,N_14658);
or U16802 (N_16802,N_14265,N_14099);
nor U16803 (N_16803,N_14847,N_13606);
nand U16804 (N_16804,N_14338,N_13085);
and U16805 (N_16805,N_14447,N_14979);
or U16806 (N_16806,N_14850,N_13424);
and U16807 (N_16807,N_13682,N_13324);
and U16808 (N_16808,N_14560,N_12976);
nand U16809 (N_16809,N_14642,N_14761);
or U16810 (N_16810,N_14784,N_13743);
nor U16811 (N_16811,N_13815,N_14630);
nand U16812 (N_16812,N_14950,N_14356);
xnor U16813 (N_16813,N_14426,N_13738);
nand U16814 (N_16814,N_12786,N_14456);
nor U16815 (N_16815,N_14066,N_14471);
nor U16816 (N_16816,N_14888,N_13609);
xor U16817 (N_16817,N_14500,N_14544);
nand U16818 (N_16818,N_14018,N_13561);
nor U16819 (N_16819,N_12781,N_14400);
xnor U16820 (N_16820,N_14632,N_13430);
and U16821 (N_16821,N_14764,N_13466);
nand U16822 (N_16822,N_12649,N_14802);
nand U16823 (N_16823,N_13297,N_13326);
or U16824 (N_16824,N_12581,N_13170);
or U16825 (N_16825,N_12518,N_14456);
or U16826 (N_16826,N_12689,N_14638);
xnor U16827 (N_16827,N_13748,N_14300);
xor U16828 (N_16828,N_13980,N_14282);
xor U16829 (N_16829,N_13891,N_13089);
nor U16830 (N_16830,N_13428,N_14788);
xnor U16831 (N_16831,N_14113,N_12689);
xnor U16832 (N_16832,N_14606,N_13597);
nand U16833 (N_16833,N_13342,N_13196);
xnor U16834 (N_16834,N_14232,N_13205);
nand U16835 (N_16835,N_12873,N_13858);
or U16836 (N_16836,N_13826,N_13246);
nor U16837 (N_16837,N_13662,N_14512);
or U16838 (N_16838,N_14094,N_13630);
xor U16839 (N_16839,N_13068,N_14795);
nand U16840 (N_16840,N_13287,N_13709);
or U16841 (N_16841,N_14401,N_14241);
or U16842 (N_16842,N_14916,N_12794);
or U16843 (N_16843,N_14254,N_14943);
nor U16844 (N_16844,N_14517,N_13524);
nand U16845 (N_16845,N_14512,N_12898);
nand U16846 (N_16846,N_14006,N_13701);
nor U16847 (N_16847,N_14778,N_14002);
and U16848 (N_16848,N_12812,N_13756);
nand U16849 (N_16849,N_14593,N_12600);
xor U16850 (N_16850,N_13675,N_12548);
nand U16851 (N_16851,N_12522,N_14021);
or U16852 (N_16852,N_14464,N_12698);
nand U16853 (N_16853,N_14974,N_14336);
or U16854 (N_16854,N_13407,N_14130);
and U16855 (N_16855,N_13347,N_13949);
nand U16856 (N_16856,N_13038,N_12525);
or U16857 (N_16857,N_14199,N_13857);
nor U16858 (N_16858,N_14836,N_14689);
and U16859 (N_16859,N_12978,N_14623);
or U16860 (N_16860,N_14734,N_13262);
xnor U16861 (N_16861,N_12914,N_12908);
nor U16862 (N_16862,N_13408,N_13842);
nor U16863 (N_16863,N_14432,N_14259);
xnor U16864 (N_16864,N_13623,N_13307);
nand U16865 (N_16865,N_12504,N_12809);
nor U16866 (N_16866,N_13128,N_14780);
nor U16867 (N_16867,N_12561,N_14635);
or U16868 (N_16868,N_14779,N_13817);
nand U16869 (N_16869,N_13110,N_13276);
xor U16870 (N_16870,N_14689,N_12687);
nor U16871 (N_16871,N_13005,N_13338);
xor U16872 (N_16872,N_13434,N_13107);
and U16873 (N_16873,N_13457,N_14769);
nand U16874 (N_16874,N_13635,N_14626);
and U16875 (N_16875,N_12720,N_13430);
nor U16876 (N_16876,N_13726,N_14870);
or U16877 (N_16877,N_13992,N_13352);
and U16878 (N_16878,N_14027,N_12708);
and U16879 (N_16879,N_13780,N_14990);
nor U16880 (N_16880,N_13162,N_13135);
nor U16881 (N_16881,N_13570,N_12699);
nand U16882 (N_16882,N_12610,N_13482);
and U16883 (N_16883,N_13942,N_13202);
and U16884 (N_16884,N_12549,N_13065);
and U16885 (N_16885,N_14416,N_13045);
and U16886 (N_16886,N_13063,N_14917);
and U16887 (N_16887,N_13444,N_13237);
and U16888 (N_16888,N_14640,N_14583);
nor U16889 (N_16889,N_14888,N_14273);
or U16890 (N_16890,N_14850,N_13043);
nor U16891 (N_16891,N_13725,N_14530);
xnor U16892 (N_16892,N_14518,N_13728);
nor U16893 (N_16893,N_14361,N_13914);
or U16894 (N_16894,N_12936,N_13372);
and U16895 (N_16895,N_13037,N_14895);
and U16896 (N_16896,N_12846,N_12907);
or U16897 (N_16897,N_14428,N_13323);
and U16898 (N_16898,N_14162,N_14876);
xor U16899 (N_16899,N_14637,N_14351);
xor U16900 (N_16900,N_14032,N_13522);
nor U16901 (N_16901,N_13985,N_13215);
and U16902 (N_16902,N_14802,N_13380);
nand U16903 (N_16903,N_12996,N_13977);
nor U16904 (N_16904,N_12543,N_14921);
and U16905 (N_16905,N_14142,N_14565);
nor U16906 (N_16906,N_13110,N_14762);
and U16907 (N_16907,N_13474,N_12560);
and U16908 (N_16908,N_13834,N_12525);
or U16909 (N_16909,N_14279,N_12744);
xnor U16910 (N_16910,N_14663,N_14908);
nor U16911 (N_16911,N_14800,N_13215);
nor U16912 (N_16912,N_14865,N_14326);
and U16913 (N_16913,N_14079,N_13176);
xnor U16914 (N_16914,N_13239,N_14496);
xnor U16915 (N_16915,N_13719,N_13225);
and U16916 (N_16916,N_13096,N_13803);
nor U16917 (N_16917,N_14483,N_14387);
or U16918 (N_16918,N_13063,N_14065);
and U16919 (N_16919,N_12555,N_14590);
nand U16920 (N_16920,N_12549,N_13433);
xor U16921 (N_16921,N_13156,N_14881);
or U16922 (N_16922,N_13399,N_13335);
and U16923 (N_16923,N_14345,N_14890);
xor U16924 (N_16924,N_13315,N_12514);
and U16925 (N_16925,N_14471,N_14708);
and U16926 (N_16926,N_13293,N_12871);
and U16927 (N_16927,N_14858,N_13738);
and U16928 (N_16928,N_14810,N_14679);
nand U16929 (N_16929,N_14377,N_13579);
and U16930 (N_16930,N_13471,N_14259);
nand U16931 (N_16931,N_13801,N_13841);
nand U16932 (N_16932,N_13801,N_12805);
or U16933 (N_16933,N_14911,N_13529);
and U16934 (N_16934,N_14388,N_14807);
and U16935 (N_16935,N_14717,N_13408);
or U16936 (N_16936,N_14223,N_13819);
and U16937 (N_16937,N_14670,N_14379);
nand U16938 (N_16938,N_12990,N_14575);
nor U16939 (N_16939,N_13203,N_13311);
nand U16940 (N_16940,N_14999,N_13867);
xor U16941 (N_16941,N_13087,N_14575);
nand U16942 (N_16942,N_14110,N_14180);
nor U16943 (N_16943,N_13598,N_13784);
nor U16944 (N_16944,N_14612,N_13034);
and U16945 (N_16945,N_13571,N_13166);
xnor U16946 (N_16946,N_14174,N_14883);
nor U16947 (N_16947,N_13992,N_14842);
nand U16948 (N_16948,N_13156,N_13440);
nor U16949 (N_16949,N_12595,N_14939);
nor U16950 (N_16950,N_12757,N_14326);
and U16951 (N_16951,N_13828,N_13985);
xnor U16952 (N_16952,N_14771,N_13846);
and U16953 (N_16953,N_13282,N_13936);
or U16954 (N_16954,N_13223,N_13464);
nor U16955 (N_16955,N_13377,N_14009);
nor U16956 (N_16956,N_12856,N_14373);
xor U16957 (N_16957,N_12914,N_12529);
or U16958 (N_16958,N_14903,N_12826);
nor U16959 (N_16959,N_12916,N_14796);
nand U16960 (N_16960,N_13679,N_13415);
nand U16961 (N_16961,N_14058,N_13636);
nor U16962 (N_16962,N_13072,N_14454);
xor U16963 (N_16963,N_12803,N_13751);
or U16964 (N_16964,N_14066,N_13789);
xor U16965 (N_16965,N_12968,N_13026);
nor U16966 (N_16966,N_13152,N_14734);
or U16967 (N_16967,N_14839,N_13122);
nor U16968 (N_16968,N_12717,N_14418);
nor U16969 (N_16969,N_14436,N_12600);
or U16970 (N_16970,N_14266,N_14416);
or U16971 (N_16971,N_13132,N_12566);
and U16972 (N_16972,N_14366,N_14571);
nor U16973 (N_16973,N_13061,N_13793);
or U16974 (N_16974,N_14554,N_13662);
or U16975 (N_16975,N_13056,N_12685);
nand U16976 (N_16976,N_12892,N_14019);
nor U16977 (N_16977,N_14473,N_13425);
or U16978 (N_16978,N_14295,N_12726);
nor U16979 (N_16979,N_13967,N_13905);
nor U16980 (N_16980,N_14705,N_12746);
nor U16981 (N_16981,N_14528,N_14187);
xor U16982 (N_16982,N_13328,N_14279);
and U16983 (N_16983,N_14672,N_13913);
nand U16984 (N_16984,N_14330,N_13759);
nand U16985 (N_16985,N_13422,N_14802);
nor U16986 (N_16986,N_14796,N_13353);
nand U16987 (N_16987,N_13576,N_14325);
and U16988 (N_16988,N_13618,N_14877);
and U16989 (N_16989,N_12918,N_12730);
nand U16990 (N_16990,N_14156,N_14040);
or U16991 (N_16991,N_13104,N_13042);
xor U16992 (N_16992,N_14695,N_12677);
nor U16993 (N_16993,N_13939,N_14930);
nor U16994 (N_16994,N_14525,N_13700);
nand U16995 (N_16995,N_13570,N_14563);
nand U16996 (N_16996,N_13166,N_13606);
or U16997 (N_16997,N_12783,N_13161);
and U16998 (N_16998,N_14874,N_14418);
and U16999 (N_16999,N_13555,N_13317);
or U17000 (N_17000,N_13518,N_14864);
or U17001 (N_17001,N_13673,N_14999);
and U17002 (N_17002,N_14557,N_12654);
nor U17003 (N_17003,N_13911,N_13611);
xor U17004 (N_17004,N_14553,N_13048);
or U17005 (N_17005,N_13047,N_13625);
or U17006 (N_17006,N_13784,N_14275);
nor U17007 (N_17007,N_14714,N_14899);
xor U17008 (N_17008,N_14385,N_13434);
xnor U17009 (N_17009,N_14471,N_13804);
nor U17010 (N_17010,N_13050,N_14330);
nor U17011 (N_17011,N_13196,N_14889);
and U17012 (N_17012,N_14047,N_12875);
or U17013 (N_17013,N_14246,N_12801);
xnor U17014 (N_17014,N_13623,N_14171);
xnor U17015 (N_17015,N_13312,N_13468);
or U17016 (N_17016,N_13877,N_14952);
and U17017 (N_17017,N_14968,N_13274);
nor U17018 (N_17018,N_14970,N_14819);
xnor U17019 (N_17019,N_14338,N_14804);
and U17020 (N_17020,N_12659,N_14640);
and U17021 (N_17021,N_12889,N_12781);
xnor U17022 (N_17022,N_13426,N_14892);
nor U17023 (N_17023,N_14098,N_13815);
xnor U17024 (N_17024,N_14449,N_14027);
or U17025 (N_17025,N_13868,N_13374);
xnor U17026 (N_17026,N_13163,N_13666);
nor U17027 (N_17027,N_14083,N_12960);
nand U17028 (N_17028,N_13071,N_14206);
nor U17029 (N_17029,N_12619,N_14421);
or U17030 (N_17030,N_14886,N_12709);
xnor U17031 (N_17031,N_13663,N_13741);
or U17032 (N_17032,N_13452,N_13852);
or U17033 (N_17033,N_14644,N_14847);
or U17034 (N_17034,N_12922,N_13770);
or U17035 (N_17035,N_12820,N_14170);
nand U17036 (N_17036,N_14396,N_13635);
xnor U17037 (N_17037,N_12850,N_14657);
nor U17038 (N_17038,N_14944,N_14112);
and U17039 (N_17039,N_13688,N_14260);
nor U17040 (N_17040,N_13928,N_13975);
nor U17041 (N_17041,N_13770,N_14166);
and U17042 (N_17042,N_13766,N_14312);
or U17043 (N_17043,N_13748,N_12879);
nor U17044 (N_17044,N_14142,N_13665);
or U17045 (N_17045,N_13885,N_14900);
xnor U17046 (N_17046,N_13344,N_13128);
and U17047 (N_17047,N_14060,N_14451);
nand U17048 (N_17048,N_13248,N_12570);
nor U17049 (N_17049,N_12896,N_13762);
nand U17050 (N_17050,N_14950,N_13743);
xor U17051 (N_17051,N_13228,N_13031);
or U17052 (N_17052,N_13245,N_13546);
and U17053 (N_17053,N_14506,N_13031);
xor U17054 (N_17054,N_12743,N_13577);
nand U17055 (N_17055,N_14837,N_12559);
and U17056 (N_17056,N_12768,N_12961);
or U17057 (N_17057,N_13844,N_14760);
and U17058 (N_17058,N_14074,N_12714);
nand U17059 (N_17059,N_14799,N_14150);
or U17060 (N_17060,N_14138,N_13118);
and U17061 (N_17061,N_13964,N_13179);
nand U17062 (N_17062,N_14764,N_14893);
and U17063 (N_17063,N_14665,N_13896);
nor U17064 (N_17064,N_14609,N_14025);
and U17065 (N_17065,N_14825,N_13303);
or U17066 (N_17066,N_13708,N_13399);
nor U17067 (N_17067,N_12526,N_14170);
or U17068 (N_17068,N_14952,N_13539);
xor U17069 (N_17069,N_14349,N_13315);
or U17070 (N_17070,N_13701,N_14088);
and U17071 (N_17071,N_14315,N_13912);
nand U17072 (N_17072,N_12640,N_13077);
nor U17073 (N_17073,N_13554,N_12518);
or U17074 (N_17074,N_13468,N_13115);
xor U17075 (N_17075,N_13330,N_13928);
xor U17076 (N_17076,N_14183,N_14617);
nor U17077 (N_17077,N_13319,N_14907);
or U17078 (N_17078,N_14547,N_14838);
and U17079 (N_17079,N_14939,N_13014);
and U17080 (N_17080,N_12650,N_14871);
nand U17081 (N_17081,N_13254,N_12516);
or U17082 (N_17082,N_13997,N_13277);
nand U17083 (N_17083,N_13067,N_12563);
or U17084 (N_17084,N_13528,N_14275);
and U17085 (N_17085,N_14665,N_14354);
nand U17086 (N_17086,N_12986,N_13060);
and U17087 (N_17087,N_14229,N_13948);
xor U17088 (N_17088,N_13680,N_13816);
or U17089 (N_17089,N_13945,N_13654);
nor U17090 (N_17090,N_12802,N_13717);
nor U17091 (N_17091,N_12950,N_14064);
and U17092 (N_17092,N_14152,N_12805);
nor U17093 (N_17093,N_14704,N_13257);
nor U17094 (N_17094,N_14688,N_13402);
xnor U17095 (N_17095,N_13195,N_14472);
and U17096 (N_17096,N_14988,N_12671);
nand U17097 (N_17097,N_14874,N_13217);
xnor U17098 (N_17098,N_13369,N_12895);
nor U17099 (N_17099,N_13386,N_14036);
nor U17100 (N_17100,N_14113,N_14632);
xor U17101 (N_17101,N_14562,N_13455);
or U17102 (N_17102,N_14278,N_13213);
nor U17103 (N_17103,N_12684,N_14403);
or U17104 (N_17104,N_12533,N_14460);
or U17105 (N_17105,N_14017,N_14404);
nand U17106 (N_17106,N_12575,N_13104);
or U17107 (N_17107,N_13571,N_13044);
nor U17108 (N_17108,N_13801,N_13036);
nand U17109 (N_17109,N_14447,N_14850);
nand U17110 (N_17110,N_12619,N_13294);
and U17111 (N_17111,N_14165,N_14189);
nand U17112 (N_17112,N_14677,N_13047);
and U17113 (N_17113,N_13252,N_14466);
and U17114 (N_17114,N_13310,N_12893);
or U17115 (N_17115,N_13722,N_13870);
xor U17116 (N_17116,N_13220,N_13589);
nand U17117 (N_17117,N_14682,N_13751);
or U17118 (N_17118,N_12549,N_12943);
nand U17119 (N_17119,N_12734,N_14938);
xnor U17120 (N_17120,N_13825,N_12718);
nand U17121 (N_17121,N_14234,N_14997);
xnor U17122 (N_17122,N_14673,N_13545);
xor U17123 (N_17123,N_12751,N_14891);
and U17124 (N_17124,N_13012,N_13259);
or U17125 (N_17125,N_13337,N_13495);
xnor U17126 (N_17126,N_13419,N_13195);
nor U17127 (N_17127,N_14758,N_14651);
and U17128 (N_17128,N_12715,N_13546);
or U17129 (N_17129,N_14539,N_13398);
nand U17130 (N_17130,N_13005,N_13463);
and U17131 (N_17131,N_14409,N_14819);
xor U17132 (N_17132,N_13103,N_13690);
nand U17133 (N_17133,N_13565,N_12983);
nor U17134 (N_17134,N_14512,N_14097);
or U17135 (N_17135,N_12906,N_13566);
nor U17136 (N_17136,N_14255,N_13474);
and U17137 (N_17137,N_14817,N_14209);
or U17138 (N_17138,N_14711,N_13535);
nor U17139 (N_17139,N_12717,N_14902);
or U17140 (N_17140,N_12878,N_14495);
xnor U17141 (N_17141,N_13081,N_14111);
nand U17142 (N_17142,N_14769,N_13546);
xnor U17143 (N_17143,N_13298,N_12850);
xnor U17144 (N_17144,N_14515,N_13311);
nand U17145 (N_17145,N_14369,N_13389);
nand U17146 (N_17146,N_14203,N_14560);
nand U17147 (N_17147,N_14285,N_14673);
and U17148 (N_17148,N_13498,N_12729);
or U17149 (N_17149,N_13902,N_12711);
xor U17150 (N_17150,N_14737,N_13679);
or U17151 (N_17151,N_12715,N_12872);
and U17152 (N_17152,N_12772,N_13442);
or U17153 (N_17153,N_14788,N_12617);
nor U17154 (N_17154,N_12502,N_12855);
or U17155 (N_17155,N_14744,N_14683);
nand U17156 (N_17156,N_12532,N_14186);
and U17157 (N_17157,N_13494,N_13067);
and U17158 (N_17158,N_13640,N_12779);
or U17159 (N_17159,N_13997,N_14603);
nor U17160 (N_17160,N_14931,N_13625);
or U17161 (N_17161,N_13472,N_13580);
and U17162 (N_17162,N_12861,N_14328);
and U17163 (N_17163,N_12672,N_13327);
nand U17164 (N_17164,N_12772,N_14069);
nor U17165 (N_17165,N_13190,N_13873);
nor U17166 (N_17166,N_14893,N_14087);
or U17167 (N_17167,N_13742,N_13792);
nand U17168 (N_17168,N_14574,N_13639);
nand U17169 (N_17169,N_13071,N_13929);
nand U17170 (N_17170,N_14123,N_14534);
nor U17171 (N_17171,N_13657,N_14261);
nor U17172 (N_17172,N_12646,N_14627);
or U17173 (N_17173,N_12872,N_12595);
nand U17174 (N_17174,N_13833,N_14725);
nand U17175 (N_17175,N_13448,N_14407);
nor U17176 (N_17176,N_14838,N_14016);
nor U17177 (N_17177,N_13413,N_13317);
nor U17178 (N_17178,N_13103,N_12547);
nor U17179 (N_17179,N_14955,N_14933);
nor U17180 (N_17180,N_13769,N_13347);
xnor U17181 (N_17181,N_13481,N_13119);
and U17182 (N_17182,N_14271,N_14800);
nand U17183 (N_17183,N_13419,N_12861);
xor U17184 (N_17184,N_13973,N_14620);
xnor U17185 (N_17185,N_12853,N_14497);
xnor U17186 (N_17186,N_14157,N_13170);
nand U17187 (N_17187,N_12645,N_13460);
nand U17188 (N_17188,N_13432,N_14255);
nor U17189 (N_17189,N_13072,N_14036);
or U17190 (N_17190,N_14093,N_12760);
nand U17191 (N_17191,N_14379,N_12638);
xnor U17192 (N_17192,N_14915,N_14173);
and U17193 (N_17193,N_13139,N_13865);
or U17194 (N_17194,N_13542,N_13902);
or U17195 (N_17195,N_13207,N_13834);
nand U17196 (N_17196,N_14042,N_13823);
nor U17197 (N_17197,N_13505,N_14099);
xnor U17198 (N_17198,N_13883,N_14431);
nand U17199 (N_17199,N_13634,N_14123);
xnor U17200 (N_17200,N_14990,N_14189);
or U17201 (N_17201,N_13877,N_14435);
or U17202 (N_17202,N_13221,N_13266);
nand U17203 (N_17203,N_14548,N_14081);
or U17204 (N_17204,N_14774,N_14139);
and U17205 (N_17205,N_14161,N_13199);
xnor U17206 (N_17206,N_13085,N_12513);
or U17207 (N_17207,N_13439,N_13447);
xor U17208 (N_17208,N_13424,N_14267);
xor U17209 (N_17209,N_12546,N_14596);
xor U17210 (N_17210,N_13672,N_12762);
nor U17211 (N_17211,N_14006,N_14476);
and U17212 (N_17212,N_13543,N_12698);
nor U17213 (N_17213,N_13566,N_13101);
nand U17214 (N_17214,N_14960,N_14838);
nor U17215 (N_17215,N_13427,N_14981);
and U17216 (N_17216,N_13518,N_13091);
nand U17217 (N_17217,N_12557,N_14612);
nand U17218 (N_17218,N_14274,N_14700);
nor U17219 (N_17219,N_14188,N_14458);
or U17220 (N_17220,N_13495,N_14551);
or U17221 (N_17221,N_14069,N_13118);
xor U17222 (N_17222,N_14443,N_14944);
xor U17223 (N_17223,N_14239,N_14404);
nor U17224 (N_17224,N_12787,N_13322);
xor U17225 (N_17225,N_12710,N_12522);
nor U17226 (N_17226,N_13333,N_12587);
nand U17227 (N_17227,N_14587,N_14037);
nand U17228 (N_17228,N_13060,N_13821);
nor U17229 (N_17229,N_13576,N_13254);
xnor U17230 (N_17230,N_13672,N_13921);
nand U17231 (N_17231,N_14414,N_12680);
or U17232 (N_17232,N_13799,N_14176);
and U17233 (N_17233,N_14012,N_13353);
or U17234 (N_17234,N_12735,N_13006);
nor U17235 (N_17235,N_12560,N_13700);
nand U17236 (N_17236,N_14170,N_12834);
nand U17237 (N_17237,N_14664,N_12749);
and U17238 (N_17238,N_12962,N_14757);
nor U17239 (N_17239,N_13995,N_13880);
xnor U17240 (N_17240,N_12796,N_14106);
nand U17241 (N_17241,N_14490,N_14691);
and U17242 (N_17242,N_12534,N_12689);
nor U17243 (N_17243,N_14788,N_12521);
nor U17244 (N_17244,N_12604,N_13661);
and U17245 (N_17245,N_13839,N_14738);
or U17246 (N_17246,N_14757,N_13613);
and U17247 (N_17247,N_14865,N_13046);
or U17248 (N_17248,N_13191,N_14241);
nand U17249 (N_17249,N_13092,N_13818);
xnor U17250 (N_17250,N_12935,N_13228);
or U17251 (N_17251,N_14943,N_12616);
and U17252 (N_17252,N_14771,N_12673);
nor U17253 (N_17253,N_14674,N_14123);
xor U17254 (N_17254,N_14151,N_14898);
xor U17255 (N_17255,N_14441,N_14920);
or U17256 (N_17256,N_12745,N_14692);
nand U17257 (N_17257,N_13072,N_13111);
nand U17258 (N_17258,N_14022,N_14151);
nand U17259 (N_17259,N_12752,N_14069);
nand U17260 (N_17260,N_14274,N_13368);
or U17261 (N_17261,N_13043,N_13974);
nand U17262 (N_17262,N_12957,N_13782);
and U17263 (N_17263,N_14731,N_14459);
xnor U17264 (N_17264,N_14075,N_14480);
and U17265 (N_17265,N_13419,N_14169);
nand U17266 (N_17266,N_12723,N_13396);
nand U17267 (N_17267,N_14939,N_13451);
nor U17268 (N_17268,N_14949,N_14127);
nand U17269 (N_17269,N_14211,N_13958);
nor U17270 (N_17270,N_13629,N_14379);
nor U17271 (N_17271,N_14830,N_14438);
nand U17272 (N_17272,N_14498,N_13863);
or U17273 (N_17273,N_12937,N_12855);
nor U17274 (N_17274,N_12507,N_14035);
or U17275 (N_17275,N_14607,N_14775);
or U17276 (N_17276,N_13606,N_14802);
xnor U17277 (N_17277,N_12641,N_13181);
or U17278 (N_17278,N_14259,N_12941);
nand U17279 (N_17279,N_12610,N_14884);
or U17280 (N_17280,N_13410,N_13383);
xor U17281 (N_17281,N_13041,N_14786);
and U17282 (N_17282,N_12558,N_14868);
xnor U17283 (N_17283,N_12738,N_14142);
nor U17284 (N_17284,N_14284,N_14381);
nand U17285 (N_17285,N_13081,N_13987);
xor U17286 (N_17286,N_12925,N_13952);
nor U17287 (N_17287,N_13211,N_13120);
and U17288 (N_17288,N_13917,N_13456);
xnor U17289 (N_17289,N_12849,N_13733);
nor U17290 (N_17290,N_14935,N_14036);
nand U17291 (N_17291,N_12726,N_12887);
and U17292 (N_17292,N_12794,N_12574);
nand U17293 (N_17293,N_13764,N_13031);
nand U17294 (N_17294,N_13881,N_14256);
and U17295 (N_17295,N_14474,N_14999);
nand U17296 (N_17296,N_12922,N_13261);
xor U17297 (N_17297,N_13183,N_12827);
nand U17298 (N_17298,N_12683,N_14317);
xnor U17299 (N_17299,N_14356,N_14896);
nor U17300 (N_17300,N_14098,N_13787);
nor U17301 (N_17301,N_14611,N_12583);
or U17302 (N_17302,N_14734,N_14082);
nor U17303 (N_17303,N_12963,N_14022);
and U17304 (N_17304,N_13047,N_13416);
or U17305 (N_17305,N_13202,N_12907);
nor U17306 (N_17306,N_14456,N_14469);
nor U17307 (N_17307,N_13005,N_13458);
nor U17308 (N_17308,N_14349,N_13625);
nor U17309 (N_17309,N_14128,N_14571);
or U17310 (N_17310,N_14339,N_12576);
and U17311 (N_17311,N_14688,N_12749);
nand U17312 (N_17312,N_13194,N_14424);
nor U17313 (N_17313,N_14158,N_13904);
nor U17314 (N_17314,N_13422,N_14322);
nand U17315 (N_17315,N_13285,N_14867);
and U17316 (N_17316,N_13508,N_12522);
nor U17317 (N_17317,N_13310,N_14298);
nand U17318 (N_17318,N_14801,N_14713);
nand U17319 (N_17319,N_14758,N_12857);
and U17320 (N_17320,N_14366,N_13216);
and U17321 (N_17321,N_13464,N_13645);
xnor U17322 (N_17322,N_14246,N_13043);
nand U17323 (N_17323,N_14433,N_14052);
and U17324 (N_17324,N_13073,N_14098);
or U17325 (N_17325,N_14941,N_12547);
nand U17326 (N_17326,N_12676,N_14833);
and U17327 (N_17327,N_13675,N_12575);
or U17328 (N_17328,N_13110,N_13280);
nand U17329 (N_17329,N_13009,N_12748);
nor U17330 (N_17330,N_12963,N_12879);
and U17331 (N_17331,N_12749,N_14820);
xnor U17332 (N_17332,N_13003,N_13588);
xnor U17333 (N_17333,N_13229,N_13022);
nand U17334 (N_17334,N_14739,N_12883);
nand U17335 (N_17335,N_14426,N_13342);
nand U17336 (N_17336,N_12913,N_12565);
and U17337 (N_17337,N_13291,N_14984);
xor U17338 (N_17338,N_13853,N_14156);
xnor U17339 (N_17339,N_13790,N_12510);
and U17340 (N_17340,N_12877,N_14447);
nand U17341 (N_17341,N_12514,N_12696);
and U17342 (N_17342,N_14702,N_14801);
or U17343 (N_17343,N_14251,N_12905);
nand U17344 (N_17344,N_12884,N_13201);
or U17345 (N_17345,N_12899,N_13084);
xor U17346 (N_17346,N_14091,N_12882);
nand U17347 (N_17347,N_14291,N_14894);
or U17348 (N_17348,N_14019,N_12641);
or U17349 (N_17349,N_14420,N_14126);
xnor U17350 (N_17350,N_14895,N_13749);
or U17351 (N_17351,N_14998,N_13146);
nor U17352 (N_17352,N_14361,N_12971);
xor U17353 (N_17353,N_13202,N_13511);
or U17354 (N_17354,N_14997,N_13064);
nand U17355 (N_17355,N_12532,N_12902);
xor U17356 (N_17356,N_12578,N_14051);
and U17357 (N_17357,N_14458,N_14154);
nor U17358 (N_17358,N_14805,N_13171);
nand U17359 (N_17359,N_14150,N_14777);
and U17360 (N_17360,N_13256,N_12842);
xor U17361 (N_17361,N_13633,N_13047);
xnor U17362 (N_17362,N_14277,N_12747);
and U17363 (N_17363,N_12761,N_14548);
nor U17364 (N_17364,N_13312,N_12689);
nand U17365 (N_17365,N_14231,N_13922);
xnor U17366 (N_17366,N_14337,N_12660);
nor U17367 (N_17367,N_14616,N_13346);
xnor U17368 (N_17368,N_13385,N_13839);
or U17369 (N_17369,N_12991,N_14034);
and U17370 (N_17370,N_14262,N_14952);
or U17371 (N_17371,N_14143,N_13647);
and U17372 (N_17372,N_12894,N_14079);
xor U17373 (N_17373,N_13513,N_14930);
nor U17374 (N_17374,N_14062,N_14699);
nor U17375 (N_17375,N_14440,N_14998);
and U17376 (N_17376,N_14171,N_14798);
nor U17377 (N_17377,N_12630,N_12721);
nand U17378 (N_17378,N_12846,N_13962);
nand U17379 (N_17379,N_13632,N_13995);
and U17380 (N_17380,N_13179,N_14128);
or U17381 (N_17381,N_14449,N_14659);
nor U17382 (N_17382,N_14614,N_12664);
xor U17383 (N_17383,N_12765,N_12953);
xor U17384 (N_17384,N_13810,N_14515);
nor U17385 (N_17385,N_14169,N_13563);
nand U17386 (N_17386,N_12589,N_14979);
and U17387 (N_17387,N_13136,N_13752);
or U17388 (N_17388,N_13482,N_13020);
xnor U17389 (N_17389,N_13901,N_14769);
or U17390 (N_17390,N_13641,N_12603);
and U17391 (N_17391,N_12559,N_14903);
nand U17392 (N_17392,N_12802,N_13372);
nor U17393 (N_17393,N_14724,N_13551);
and U17394 (N_17394,N_14629,N_13401);
xnor U17395 (N_17395,N_14689,N_14389);
or U17396 (N_17396,N_13435,N_13340);
or U17397 (N_17397,N_13943,N_13821);
nor U17398 (N_17398,N_13335,N_14816);
nand U17399 (N_17399,N_14677,N_13051);
or U17400 (N_17400,N_14103,N_14693);
or U17401 (N_17401,N_12732,N_13854);
and U17402 (N_17402,N_12906,N_13261);
nor U17403 (N_17403,N_14901,N_14273);
and U17404 (N_17404,N_14355,N_14667);
and U17405 (N_17405,N_14547,N_13510);
nor U17406 (N_17406,N_13958,N_13080);
xnor U17407 (N_17407,N_14845,N_14001);
nor U17408 (N_17408,N_14127,N_13259);
nor U17409 (N_17409,N_13990,N_13596);
xnor U17410 (N_17410,N_13997,N_14541);
nand U17411 (N_17411,N_13776,N_13903);
xnor U17412 (N_17412,N_13887,N_14375);
and U17413 (N_17413,N_14482,N_13244);
and U17414 (N_17414,N_14421,N_12627);
nor U17415 (N_17415,N_14274,N_14513);
and U17416 (N_17416,N_12935,N_14682);
and U17417 (N_17417,N_13218,N_13621);
or U17418 (N_17418,N_14858,N_13051);
xor U17419 (N_17419,N_14451,N_13296);
or U17420 (N_17420,N_13842,N_14050);
nand U17421 (N_17421,N_13645,N_14523);
nand U17422 (N_17422,N_14446,N_13173);
or U17423 (N_17423,N_14645,N_13594);
nor U17424 (N_17424,N_14267,N_14346);
xnor U17425 (N_17425,N_14319,N_13237);
and U17426 (N_17426,N_14806,N_13577);
and U17427 (N_17427,N_13243,N_14831);
nor U17428 (N_17428,N_13480,N_13818);
or U17429 (N_17429,N_14251,N_14333);
or U17430 (N_17430,N_14414,N_13758);
nand U17431 (N_17431,N_14833,N_14606);
xnor U17432 (N_17432,N_14506,N_13514);
nor U17433 (N_17433,N_14484,N_13184);
xor U17434 (N_17434,N_13712,N_14172);
xor U17435 (N_17435,N_14422,N_14910);
nand U17436 (N_17436,N_14226,N_14485);
and U17437 (N_17437,N_14574,N_12826);
or U17438 (N_17438,N_13857,N_14275);
nor U17439 (N_17439,N_14264,N_13586);
nand U17440 (N_17440,N_12735,N_13929);
nand U17441 (N_17441,N_12580,N_13150);
or U17442 (N_17442,N_14373,N_13419);
nand U17443 (N_17443,N_14669,N_14251);
and U17444 (N_17444,N_14876,N_14120);
and U17445 (N_17445,N_13968,N_14366);
nor U17446 (N_17446,N_14182,N_12834);
nand U17447 (N_17447,N_14157,N_13176);
nand U17448 (N_17448,N_12784,N_13776);
nand U17449 (N_17449,N_12898,N_12580);
nor U17450 (N_17450,N_12932,N_13967);
nor U17451 (N_17451,N_13804,N_12790);
nor U17452 (N_17452,N_14731,N_12695);
xor U17453 (N_17453,N_13727,N_13744);
nor U17454 (N_17454,N_13212,N_14642);
nand U17455 (N_17455,N_14735,N_13028);
nand U17456 (N_17456,N_14787,N_14750);
and U17457 (N_17457,N_12567,N_13077);
nand U17458 (N_17458,N_13963,N_14061);
xor U17459 (N_17459,N_14474,N_14536);
nand U17460 (N_17460,N_13240,N_14432);
or U17461 (N_17461,N_12974,N_12964);
and U17462 (N_17462,N_13504,N_14267);
or U17463 (N_17463,N_14770,N_13735);
nor U17464 (N_17464,N_13124,N_13740);
xor U17465 (N_17465,N_13721,N_14646);
nor U17466 (N_17466,N_13942,N_12859);
xnor U17467 (N_17467,N_13626,N_14845);
xor U17468 (N_17468,N_14259,N_14605);
xnor U17469 (N_17469,N_13035,N_13845);
or U17470 (N_17470,N_14217,N_12749);
or U17471 (N_17471,N_13952,N_13457);
nand U17472 (N_17472,N_14159,N_13768);
and U17473 (N_17473,N_13791,N_13648);
or U17474 (N_17474,N_13480,N_13120);
nand U17475 (N_17475,N_14206,N_12873);
nand U17476 (N_17476,N_13973,N_13016);
xnor U17477 (N_17477,N_12932,N_13619);
nor U17478 (N_17478,N_14809,N_13812);
or U17479 (N_17479,N_13815,N_13991);
nor U17480 (N_17480,N_13270,N_13236);
and U17481 (N_17481,N_13982,N_13150);
nand U17482 (N_17482,N_14345,N_13570);
xor U17483 (N_17483,N_14556,N_13915);
and U17484 (N_17484,N_14232,N_14755);
nand U17485 (N_17485,N_13657,N_14411);
nor U17486 (N_17486,N_13440,N_14839);
xnor U17487 (N_17487,N_12531,N_14795);
nand U17488 (N_17488,N_14257,N_13632);
xor U17489 (N_17489,N_13928,N_13571);
xor U17490 (N_17490,N_12968,N_13372);
nor U17491 (N_17491,N_14822,N_13174);
nand U17492 (N_17492,N_13665,N_13626);
nor U17493 (N_17493,N_12675,N_13857);
nor U17494 (N_17494,N_14682,N_14127);
xor U17495 (N_17495,N_13571,N_12505);
or U17496 (N_17496,N_13066,N_13380);
nand U17497 (N_17497,N_14463,N_14945);
xnor U17498 (N_17498,N_13387,N_13486);
and U17499 (N_17499,N_13760,N_13427);
and U17500 (N_17500,N_15893,N_15691);
and U17501 (N_17501,N_15423,N_16523);
or U17502 (N_17502,N_15080,N_16245);
or U17503 (N_17503,N_15505,N_15849);
or U17504 (N_17504,N_16151,N_16954);
xnor U17505 (N_17505,N_15156,N_17214);
or U17506 (N_17506,N_15330,N_16915);
xnor U17507 (N_17507,N_16207,N_15494);
or U17508 (N_17508,N_15420,N_15935);
nor U17509 (N_17509,N_15746,N_15334);
and U17510 (N_17510,N_15899,N_16462);
nand U17511 (N_17511,N_16440,N_17114);
nor U17512 (N_17512,N_17475,N_15525);
or U17513 (N_17513,N_15234,N_17010);
and U17514 (N_17514,N_16555,N_16347);
or U17515 (N_17515,N_15223,N_16810);
and U17516 (N_17516,N_15078,N_15013);
nor U17517 (N_17517,N_15023,N_16020);
and U17518 (N_17518,N_17182,N_17153);
and U17519 (N_17519,N_16794,N_17276);
xor U17520 (N_17520,N_16087,N_16456);
nand U17521 (N_17521,N_17086,N_16983);
and U17522 (N_17522,N_15747,N_16909);
or U17523 (N_17523,N_15296,N_15391);
or U17524 (N_17524,N_16789,N_16150);
xnor U17525 (N_17525,N_16904,N_16211);
nor U17526 (N_17526,N_16468,N_16529);
nand U17527 (N_17527,N_16684,N_15952);
nor U17528 (N_17528,N_16861,N_16977);
xor U17529 (N_17529,N_15966,N_17316);
nor U17530 (N_17530,N_15780,N_15671);
nand U17531 (N_17531,N_15121,N_17148);
and U17532 (N_17532,N_16885,N_16390);
nor U17533 (N_17533,N_16569,N_16683);
and U17534 (N_17534,N_15909,N_16773);
nand U17535 (N_17535,N_16765,N_16549);
nand U17536 (N_17536,N_15698,N_15866);
nand U17537 (N_17537,N_15610,N_15016);
nand U17538 (N_17538,N_16689,N_16632);
xor U17539 (N_17539,N_16221,N_17160);
nand U17540 (N_17540,N_17179,N_17071);
xor U17541 (N_17541,N_16469,N_16856);
and U17542 (N_17542,N_15255,N_15421);
and U17543 (N_17543,N_16295,N_15553);
nand U17544 (N_17544,N_15073,N_17038);
or U17545 (N_17545,N_15493,N_16346);
xor U17546 (N_17546,N_17423,N_15516);
or U17547 (N_17547,N_17391,N_15695);
nand U17548 (N_17548,N_15247,N_17430);
or U17549 (N_17549,N_15193,N_15020);
or U17550 (N_17550,N_17385,N_15620);
and U17551 (N_17551,N_17116,N_15167);
or U17552 (N_17552,N_15171,N_15678);
or U17553 (N_17553,N_15715,N_16050);
nor U17554 (N_17554,N_15536,N_15635);
xnor U17555 (N_17555,N_16329,N_16966);
xnor U17556 (N_17556,N_15004,N_16835);
or U17557 (N_17557,N_15157,N_17396);
nand U17558 (N_17558,N_15809,N_16545);
nor U17559 (N_17559,N_17446,N_17079);
or U17560 (N_17560,N_15065,N_15586);
nand U17561 (N_17561,N_16598,N_15875);
and U17562 (N_17562,N_15528,N_15649);
xor U17563 (N_17563,N_16970,N_15408);
nand U17564 (N_17564,N_17091,N_16460);
nand U17565 (N_17565,N_15645,N_17226);
xor U17566 (N_17566,N_15384,N_16158);
nor U17567 (N_17567,N_15266,N_16760);
or U17568 (N_17568,N_15922,N_15377);
and U17569 (N_17569,N_17386,N_17296);
and U17570 (N_17570,N_17237,N_17189);
and U17571 (N_17571,N_17485,N_16265);
or U17572 (N_17572,N_15018,N_17095);
nor U17573 (N_17573,N_16627,N_17335);
nand U17574 (N_17574,N_16613,N_15769);
xnor U17575 (N_17575,N_15965,N_16302);
and U17576 (N_17576,N_16908,N_15794);
xnor U17577 (N_17577,N_17378,N_15317);
or U17578 (N_17578,N_16105,N_15870);
xnor U17579 (N_17579,N_16359,N_16444);
nor U17580 (N_17580,N_16369,N_16233);
and U17581 (N_17581,N_16512,N_16715);
and U17582 (N_17582,N_16036,N_16212);
nor U17583 (N_17583,N_17104,N_16363);
xnor U17584 (N_17584,N_15179,N_17497);
xor U17585 (N_17585,N_16941,N_15636);
or U17586 (N_17586,N_16644,N_16338);
nand U17587 (N_17587,N_16406,N_15279);
or U17588 (N_17588,N_17108,N_15478);
nor U17589 (N_17589,N_17286,N_15168);
and U17590 (N_17590,N_16923,N_16143);
xnor U17591 (N_17591,N_15109,N_17305);
xor U17592 (N_17592,N_15934,N_16799);
or U17593 (N_17593,N_16645,N_15075);
nand U17594 (N_17594,N_16649,N_17201);
xor U17595 (N_17595,N_16039,N_17422);
nor U17596 (N_17596,N_16771,N_15342);
nor U17597 (N_17597,N_16099,N_17344);
or U17598 (N_17598,N_16337,N_17339);
or U17599 (N_17599,N_15214,N_17245);
or U17600 (N_17600,N_16592,N_16677);
nand U17601 (N_17601,N_16565,N_15693);
nand U17602 (N_17602,N_15859,N_16030);
nor U17603 (N_17603,N_16046,N_16232);
nor U17604 (N_17604,N_17431,N_16074);
xnor U17605 (N_17605,N_17209,N_15000);
or U17606 (N_17606,N_16426,N_15361);
nor U17607 (N_17607,N_15322,N_17013);
nand U17608 (N_17608,N_15598,N_16957);
nand U17609 (N_17609,N_16052,N_16690);
and U17610 (N_17610,N_16774,N_16292);
nand U17611 (N_17611,N_17025,N_16993);
nand U17612 (N_17612,N_15521,N_15430);
nand U17613 (N_17613,N_16628,N_15680);
or U17614 (N_17614,N_17399,N_16678);
and U17615 (N_17615,N_15010,N_17440);
nor U17616 (N_17616,N_15422,N_15900);
xnor U17617 (N_17617,N_15164,N_16193);
nor U17618 (N_17618,N_17051,N_15951);
and U17619 (N_17619,N_17046,N_16669);
and U17620 (N_17620,N_17055,N_15136);
xnor U17621 (N_17621,N_17483,N_15450);
xnor U17622 (N_17622,N_16668,N_16717);
nand U17623 (N_17623,N_17195,N_15512);
nand U17624 (N_17624,N_15545,N_15520);
nand U17625 (N_17625,N_15947,N_16559);
and U17626 (N_17626,N_16167,N_15704);
or U17627 (N_17627,N_15412,N_17068);
or U17628 (N_17628,N_17176,N_15486);
xnor U17629 (N_17629,N_15881,N_17081);
and U17630 (N_17630,N_17297,N_16186);
and U17631 (N_17631,N_16484,N_15537);
and U17632 (N_17632,N_16521,N_15352);
and U17633 (N_17633,N_15338,N_16542);
and U17634 (N_17634,N_15379,N_17194);
nand U17635 (N_17635,N_15030,N_16612);
and U17636 (N_17636,N_15385,N_15655);
nand U17637 (N_17637,N_16222,N_15631);
or U17638 (N_17638,N_17458,N_16951);
or U17639 (N_17639,N_17227,N_17023);
nand U17640 (N_17640,N_15263,N_15467);
nand U17641 (N_17641,N_15582,N_17368);
nand U17642 (N_17642,N_15823,N_15395);
xor U17643 (N_17643,N_15217,N_15551);
nor U17644 (N_17644,N_17034,N_15064);
and U17645 (N_17645,N_16253,N_16134);
or U17646 (N_17646,N_15916,N_15974);
xor U17647 (N_17647,N_17005,N_15788);
nor U17648 (N_17648,N_15927,N_15465);
or U17649 (N_17649,N_15890,N_16790);
and U17650 (N_17650,N_17419,N_16382);
and U17651 (N_17651,N_17269,N_16162);
and U17652 (N_17652,N_16621,N_17230);
or U17653 (N_17653,N_17318,N_15891);
and U17654 (N_17654,N_15574,N_17451);
and U17655 (N_17655,N_15968,N_17383);
and U17656 (N_17656,N_15772,N_17124);
xor U17657 (N_17657,N_15448,N_15535);
or U17658 (N_17658,N_16558,N_15288);
nor U17659 (N_17659,N_16439,N_15058);
nor U17660 (N_17660,N_16452,N_15803);
and U17661 (N_17661,N_17438,N_16284);
nor U17662 (N_17662,N_15487,N_16088);
nand U17663 (N_17663,N_17345,N_17494);
and U17664 (N_17664,N_15211,N_16383);
and U17665 (N_17665,N_16311,N_17122);
and U17666 (N_17666,N_15414,N_16935);
nand U17667 (N_17667,N_16213,N_17033);
nor U17668 (N_17668,N_16631,N_15653);
nand U17669 (N_17669,N_16059,N_16492);
nand U17670 (N_17670,N_15290,N_15656);
and U17671 (N_17671,N_17340,N_16504);
xor U17672 (N_17672,N_17328,N_17224);
and U17673 (N_17673,N_16886,N_16584);
xor U17674 (N_17674,N_15964,N_15542);
and U17675 (N_17675,N_15221,N_16758);
or U17676 (N_17676,N_15611,N_15957);
nand U17677 (N_17677,N_16356,N_16179);
nor U17678 (N_17678,N_15576,N_16917);
or U17679 (N_17679,N_15049,N_16409);
xnor U17680 (N_17680,N_15730,N_17084);
nand U17681 (N_17681,N_16032,N_16630);
and U17682 (N_17682,N_17078,N_15640);
and U17683 (N_17683,N_15009,N_15481);
and U17684 (N_17684,N_16783,N_16463);
xor U17685 (N_17685,N_16495,N_17463);
nand U17686 (N_17686,N_16890,N_16092);
xnor U17687 (N_17687,N_16842,N_16287);
and U17688 (N_17688,N_16833,N_16428);
and U17689 (N_17689,N_16424,N_15496);
nor U17690 (N_17690,N_17354,N_15345);
xnor U17691 (N_17691,N_15667,N_15741);
xnor U17692 (N_17692,N_15212,N_16125);
nand U17693 (N_17693,N_16729,N_15273);
nor U17694 (N_17694,N_15274,N_15751);
and U17695 (N_17695,N_16129,N_15034);
and U17696 (N_17696,N_15912,N_17246);
nand U17697 (N_17697,N_15941,N_15407);
or U17698 (N_17698,N_16664,N_16705);
xor U17699 (N_17699,N_17466,N_16898);
and U17700 (N_17700,N_16417,N_15309);
xor U17701 (N_17701,N_17498,N_16096);
or U17702 (N_17702,N_15284,N_17044);
nand U17703 (N_17703,N_17253,N_16914);
xnor U17704 (N_17704,N_15988,N_15222);
and U17705 (N_17705,N_16724,N_15261);
nor U17706 (N_17706,N_15089,N_15775);
nand U17707 (N_17707,N_17304,N_15235);
or U17708 (N_17708,N_16175,N_15679);
and U17709 (N_17709,N_15626,N_15059);
or U17710 (N_17710,N_15682,N_15443);
or U17711 (N_17711,N_15606,N_16570);
xnor U17712 (N_17712,N_16508,N_15464);
xor U17713 (N_17713,N_15427,N_15014);
or U17714 (N_17714,N_17303,N_15372);
or U17715 (N_17715,N_16198,N_17107);
nor U17716 (N_17716,N_15419,N_17394);
nor U17717 (N_17717,N_16474,N_17076);
nand U17718 (N_17718,N_16879,N_16285);
nor U17719 (N_17719,N_16522,N_16980);
and U17720 (N_17720,N_15527,N_16601);
nand U17721 (N_17721,N_15150,N_15683);
nor U17722 (N_17722,N_15474,N_16071);
nand U17723 (N_17723,N_16061,N_15958);
nor U17724 (N_17724,N_16307,N_15661);
nand U17725 (N_17725,N_17447,N_15477);
and U17726 (N_17726,N_16070,N_16499);
or U17727 (N_17727,N_16636,N_16293);
xnor U17728 (N_17728,N_16275,N_15027);
or U17729 (N_17729,N_17175,N_15623);
or U17730 (N_17730,N_16078,N_15699);
nor U17731 (N_17731,N_17395,N_16988);
nand U17732 (N_17732,N_16192,N_15457);
or U17733 (N_17733,N_15758,N_17263);
nor U17734 (N_17734,N_15128,N_17319);
xor U17735 (N_17735,N_16454,N_16183);
nand U17736 (N_17736,N_16738,N_15650);
xnor U17737 (N_17737,N_15652,N_16012);
nand U17738 (N_17738,N_17093,N_16647);
or U17739 (N_17739,N_15728,N_16118);
or U17740 (N_17740,N_16323,N_17143);
nand U17741 (N_17741,N_16726,N_15170);
nor U17742 (N_17742,N_17472,N_16297);
and U17743 (N_17743,N_15711,N_16402);
xnor U17744 (N_17744,N_15216,N_15019);
and U17745 (N_17745,N_15142,N_16163);
nand U17746 (N_17746,N_16610,N_16906);
nor U17747 (N_17747,N_16986,N_15953);
nand U17748 (N_17748,N_15461,N_15604);
nand U17749 (N_17749,N_17418,N_17457);
nand U17750 (N_17750,N_15973,N_16916);
or U17751 (N_17751,N_17356,N_17390);
nor U17752 (N_17752,N_16116,N_17198);
or U17753 (N_17753,N_15458,N_16401);
nand U17754 (N_17754,N_16985,N_16698);
and U17755 (N_17755,N_16814,N_17434);
nor U17756 (N_17756,N_16816,N_15830);
nor U17757 (N_17757,N_17113,N_15602);
nand U17758 (N_17758,N_15603,N_15524);
and U17759 (N_17759,N_16498,N_15618);
xor U17760 (N_17760,N_17247,N_15921);
nand U17761 (N_17761,N_16240,N_17141);
and U17762 (N_17762,N_15822,N_15697);
or U17763 (N_17763,N_17105,N_15703);
nand U17764 (N_17764,N_16004,N_17006);
or U17765 (N_17765,N_15425,N_17311);
xnor U17766 (N_17766,N_15318,N_15463);
nor U17767 (N_17767,N_16742,N_16018);
xor U17768 (N_17768,N_16526,N_16485);
nand U17769 (N_17769,N_15798,N_16617);
nand U17770 (N_17770,N_15720,N_17031);
and U17771 (N_17771,N_17257,N_17417);
nand U17772 (N_17772,N_15845,N_17347);
nor U17773 (N_17773,N_17210,N_15111);
nand U17774 (N_17774,N_17101,N_15329);
nand U17775 (N_17775,N_17073,N_16748);
nor U17776 (N_17776,N_16140,N_15702);
and U17777 (N_17777,N_15569,N_15184);
nor U17778 (N_17778,N_15785,N_15841);
and U17779 (N_17779,N_17052,N_16478);
and U17780 (N_17780,N_16778,N_15585);
nand U17781 (N_17781,N_15116,N_15763);
xor U17782 (N_17782,N_16837,N_15144);
and U17783 (N_17783,N_16527,N_16869);
and U17784 (N_17784,N_15575,N_17471);
xnor U17785 (N_17785,N_16712,N_16351);
or U17786 (N_17786,N_16900,N_16546);
or U17787 (N_17787,N_16502,N_16852);
nor U17788 (N_17788,N_15155,N_16342);
xnor U17789 (N_17789,N_16614,N_17089);
nor U17790 (N_17790,N_15475,N_17097);
nor U17791 (N_17791,N_15654,N_15275);
or U17792 (N_17792,N_15031,N_16234);
or U17793 (N_17793,N_16016,N_15094);
xor U17794 (N_17794,N_16793,N_15162);
and U17795 (N_17795,N_15066,N_17490);
nor U17796 (N_17796,N_15928,N_16656);
and U17797 (N_17797,N_17461,N_15307);
or U17798 (N_17798,N_15539,N_15861);
xor U17799 (N_17799,N_16365,N_16676);
nor U17800 (N_17800,N_15021,N_15087);
xor U17801 (N_17801,N_15596,N_17222);
xor U17802 (N_17802,N_15908,N_15681);
or U17803 (N_17803,N_15584,N_16196);
or U17804 (N_17804,N_16568,N_15624);
xor U17805 (N_17805,N_16655,N_16739);
nand U17806 (N_17806,N_17039,N_16892);
xnor U17807 (N_17807,N_16769,N_16539);
nand U17808 (N_17808,N_15931,N_15901);
nor U17809 (N_17809,N_15637,N_17350);
nor U17810 (N_17810,N_15858,N_15605);
or U17811 (N_17811,N_17302,N_17402);
or U17812 (N_17812,N_15490,N_16024);
or U17813 (N_17813,N_17439,N_15955);
nor U17814 (N_17814,N_15036,N_17443);
nor U17815 (N_17815,N_16608,N_15375);
or U17816 (N_17816,N_15300,N_17301);
and U17817 (N_17817,N_16579,N_15709);
or U17818 (N_17818,N_17281,N_15615);
or U17819 (N_17819,N_15340,N_15839);
xnor U17820 (N_17820,N_16375,N_16379);
or U17821 (N_17821,N_17118,N_16421);
or U17822 (N_17822,N_15335,N_16550);
xnor U17823 (N_17823,N_16146,N_17489);
and U17824 (N_17824,N_15436,N_16557);
xnor U17825 (N_17825,N_15978,N_16663);
nand U17826 (N_17826,N_16832,N_15236);
nor U17827 (N_17827,N_16261,N_16776);
nor U17828 (N_17828,N_16397,N_15660);
nor U17829 (N_17829,N_16770,N_15426);
xor U17830 (N_17830,N_16761,N_17070);
xor U17831 (N_17831,N_16376,N_17215);
or U17832 (N_17832,N_15657,N_16662);
or U17833 (N_17833,N_15595,N_17487);
and U17834 (N_17834,N_16552,N_17331);
and U17835 (N_17835,N_15095,N_16947);
xnor U17836 (N_17836,N_17037,N_15373);
and U17837 (N_17837,N_15359,N_15100);
and U17838 (N_17838,N_15821,N_15440);
nor U17839 (N_17839,N_16034,N_16465);
or U17840 (N_17840,N_16380,N_16824);
nand U17841 (N_17841,N_16675,N_15028);
and U17842 (N_17842,N_15942,N_17479);
xnor U17843 (N_17843,N_17282,N_17330);
or U17844 (N_17844,N_15903,N_15745);
or U17845 (N_17845,N_16476,N_15882);
and U17846 (N_17846,N_16405,N_15756);
nor U17847 (N_17847,N_16755,N_15444);
and U17848 (N_17848,N_16272,N_15376);
nor U17849 (N_17849,N_15970,N_17341);
xor U17850 (N_17850,N_16144,N_17000);
or U17851 (N_17851,N_16325,N_17480);
or U17852 (N_17852,N_15755,N_16423);
nor U17853 (N_17853,N_15812,N_16108);
xor U17854 (N_17854,N_16160,N_16511);
nor U17855 (N_17855,N_16625,N_15497);
or U17856 (N_17856,N_17449,N_15990);
and U17857 (N_17857,N_16560,N_16149);
xor U17858 (N_17858,N_15489,N_15400);
nand U17859 (N_17859,N_17059,N_16797);
nor U17860 (N_17860,N_15024,N_16894);
nand U17861 (N_17861,N_17169,N_16795);
and U17862 (N_17862,N_16944,N_17348);
nand U17863 (N_17863,N_17491,N_17199);
nand U17864 (N_17864,N_17380,N_15616);
or U17865 (N_17865,N_15191,N_15685);
nor U17866 (N_17866,N_16387,N_16849);
and U17867 (N_17867,N_17022,N_15540);
nor U17868 (N_17868,N_17426,N_16102);
nor U17869 (N_17869,N_16355,N_15999);
nand U17870 (N_17870,N_15339,N_15555);
nand U17871 (N_17871,N_16236,N_15945);
xnor U17872 (N_17872,N_16870,N_16360);
or U17873 (N_17873,N_15905,N_15301);
and U17874 (N_17874,N_17370,N_15271);
nor U17875 (N_17875,N_15668,N_15165);
and U17876 (N_17876,N_16590,N_16964);
xor U17877 (N_17877,N_16072,N_15259);
and U17878 (N_17878,N_16800,N_15081);
nor U17879 (N_17879,N_16249,N_17203);
and U17880 (N_17880,N_16562,N_16115);
nor U17881 (N_17881,N_16348,N_15280);
nor U17882 (N_17882,N_16930,N_15374);
nor U17883 (N_17883,N_16194,N_16638);
xnor U17884 (N_17884,N_16195,N_15765);
nor U17885 (N_17885,N_17142,N_16073);
xnor U17886 (N_17886,N_16425,N_16180);
nand U17887 (N_17887,N_16844,N_15848);
nor U17888 (N_17888,N_15435,N_15153);
and U17889 (N_17889,N_16173,N_16496);
or U17890 (N_17890,N_17250,N_15151);
xnor U17891 (N_17891,N_17362,N_15178);
nand U17892 (N_17892,N_15272,N_17047);
nor U17893 (N_17893,N_16114,N_16594);
or U17894 (N_17894,N_15079,N_17064);
and U17895 (N_17895,N_15690,N_15328);
and U17896 (N_17896,N_15718,N_15726);
xor U17897 (N_17897,N_16691,N_15517);
and U17898 (N_17898,N_17040,N_16001);
and U17899 (N_17899,N_16999,N_15675);
and U17900 (N_17900,N_16704,N_17236);
or U17901 (N_17901,N_17292,N_15091);
xor U17902 (N_17902,N_15612,N_16026);
nand U17903 (N_17903,N_15197,N_16839);
xor U17904 (N_17904,N_15559,N_15907);
nand U17905 (N_17905,N_16315,N_16939);
and U17906 (N_17906,N_16708,N_15969);
nand U17907 (N_17907,N_15158,N_16533);
nor U17908 (N_17908,N_15133,N_15950);
nand U17909 (N_17909,N_17112,N_16056);
nor U17910 (N_17910,N_16730,N_16576);
nand U17911 (N_17911,N_17163,N_16699);
nor U17912 (N_17912,N_17015,N_15006);
nand U17913 (N_17913,N_15177,N_15914);
xor U17914 (N_17914,N_17058,N_16124);
nor U17915 (N_17915,N_17453,N_15348);
and U17916 (N_17916,N_15954,N_16670);
or U17917 (N_17917,N_16399,N_17481);
nor U17918 (N_17918,N_16728,N_16553);
nor U17919 (N_17919,N_16956,N_16161);
or U17920 (N_17920,N_15642,N_17420);
nand U17921 (N_17921,N_17054,N_16962);
nand U17922 (N_17922,N_17244,N_16182);
or U17923 (N_17923,N_15411,N_15045);
nand U17924 (N_17924,N_16419,N_17377);
or U17925 (N_17925,N_16803,N_16455);
xor U17926 (N_17926,N_15415,N_16696);
or U17927 (N_17927,N_16170,N_15082);
nand U17928 (N_17928,N_16224,N_17149);
nand U17929 (N_17929,N_15090,N_17026);
xor U17930 (N_17930,N_16357,N_16880);
nand U17931 (N_17931,N_17220,N_15738);
or U17932 (N_17932,N_16414,N_15131);
or U17933 (N_17933,N_17008,N_17499);
xnor U17934 (N_17934,N_15114,N_15783);
nor U17935 (N_17935,N_15306,N_16178);
and U17936 (N_17936,N_16220,N_15192);
and U17937 (N_17937,N_16754,N_15913);
nand U17938 (N_17938,N_15560,N_17233);
or U17939 (N_17939,N_15919,N_17320);
or U17940 (N_17940,N_17315,N_17181);
nand U17941 (N_17941,N_16318,N_17492);
and U17942 (N_17942,N_16543,N_16332);
nand U17943 (N_17943,N_15710,N_15231);
xor U17944 (N_17944,N_17048,N_15813);
xnor U17945 (N_17945,N_16829,N_16327);
nand U17946 (N_17946,N_15557,N_16585);
and U17947 (N_17947,N_16745,N_15061);
nor U17948 (N_17948,N_15451,N_16106);
nand U17949 (N_17949,N_15337,N_17359);
nand U17950 (N_17950,N_16741,N_15552);
nor U17951 (N_17951,N_15257,N_16480);
or U17952 (N_17952,N_17248,N_15062);
and U17953 (N_17953,N_15252,N_16659);
nand U17954 (N_17954,N_16219,N_15868);
nand U17955 (N_17955,N_16159,N_17096);
xnor U17956 (N_17956,N_16047,N_15506);
or U17957 (N_17957,N_16117,N_15993);
nor U17958 (N_17958,N_16933,N_16660);
nand U17959 (N_17959,N_16710,N_16267);
xnor U17960 (N_17960,N_16244,N_17464);
nand U17961 (N_17961,N_15714,N_15840);
xnor U17962 (N_17962,N_17208,N_16801);
and U17963 (N_17963,N_16350,N_17404);
nand U17964 (N_17964,N_16391,N_15991);
xor U17965 (N_17965,N_16961,N_16051);
xor U17966 (N_17966,N_15692,N_16720);
nor U17967 (N_17967,N_16174,N_17355);
or U17968 (N_17968,N_15773,N_15103);
nand U17969 (N_17969,N_16386,N_15251);
nor U17970 (N_17970,N_15563,N_16817);
xor U17971 (N_17971,N_15688,N_15514);
and U17972 (N_17972,N_16226,N_16006);
nand U17973 (N_17973,N_15500,N_17225);
xor U17974 (N_17974,N_17366,N_15015);
xor U17975 (N_17975,N_15378,N_15701);
or U17976 (N_17976,N_17465,N_16203);
and U17977 (N_17977,N_17478,N_16063);
and U17978 (N_17978,N_16633,N_15824);
nand U17979 (N_17979,N_17062,N_15005);
and U17980 (N_17980,N_16927,N_15470);
nor U17981 (N_17981,N_17140,N_15209);
nand U17982 (N_17982,N_17152,N_17277);
nor U17983 (N_17983,N_16208,N_15282);
nor U17984 (N_17984,N_16561,N_17150);
nor U17985 (N_17985,N_15292,N_16023);
nand U17986 (N_17986,N_15092,N_16103);
and U17987 (N_17987,N_16945,N_17098);
or U17988 (N_17988,N_16687,N_17083);
xor U17989 (N_17989,N_15872,N_17389);
xor U17990 (N_17990,N_17428,N_15573);
nor U17991 (N_17991,N_15737,N_16412);
nor U17992 (N_17992,N_15892,N_16946);
nand U17993 (N_17993,N_15298,N_15396);
nand U17994 (N_17994,N_15353,N_16813);
and U17995 (N_17995,N_17205,N_15739);
nor U17996 (N_17996,N_16075,N_15172);
xnor U17997 (N_17997,N_16085,N_17258);
or U17998 (N_17998,N_16788,N_16320);
xnor U17999 (N_17999,N_15621,N_15482);
nor U18000 (N_18000,N_15105,N_15382);
and U18001 (N_18001,N_16674,N_15268);
and U18002 (N_18002,N_16091,N_16657);
nor U18003 (N_18003,N_16459,N_17147);
or U18004 (N_18004,N_15124,N_15827);
or U18005 (N_18005,N_16525,N_16850);
nor U18006 (N_18006,N_15351,N_17184);
or U18007 (N_18007,N_17484,N_15233);
or U18008 (N_18008,N_15294,N_15689);
xor U18009 (N_18009,N_15409,N_16230);
nand U18010 (N_18010,N_16291,N_16926);
and U18011 (N_18011,N_17030,N_15220);
and U18012 (N_18012,N_16768,N_15101);
nor U18013 (N_18013,N_15399,N_17011);
or U18014 (N_18014,N_16273,N_17482);
nor U18015 (N_18015,N_17336,N_16666);
and U18016 (N_18016,N_16959,N_16786);
or U18017 (N_18017,N_15123,N_17060);
nand U18018 (N_18018,N_15753,N_15072);
or U18019 (N_18019,N_16022,N_15227);
xnor U18020 (N_18020,N_16268,N_16807);
nor U18021 (N_18021,N_15161,N_16693);
and U18022 (N_18022,N_15441,N_15519);
xnor U18023 (N_18023,N_17075,N_15046);
or U18024 (N_18024,N_16882,N_16466);
nor U18025 (N_18025,N_16005,N_16781);
and U18026 (N_18026,N_16334,N_15293);
and U18027 (N_18027,N_16599,N_16700);
nand U18028 (N_18028,N_17298,N_16671);
nand U18029 (N_18029,N_15911,N_16040);
or U18030 (N_18030,N_16873,N_15588);
xor U18031 (N_18031,N_16766,N_16054);
xor U18032 (N_18032,N_16353,N_15855);
xnor U18033 (N_18033,N_16002,N_15589);
nand U18034 (N_18034,N_16665,N_15202);
xor U18035 (N_18035,N_15975,N_15902);
and U18036 (N_18036,N_17177,N_16467);
nor U18037 (N_18037,N_15587,N_17159);
nor U18038 (N_18038,N_16418,N_16041);
nor U18039 (N_18039,N_16011,N_16931);
xnor U18040 (N_18040,N_17343,N_15801);
and U18041 (N_18041,N_16464,N_16593);
nor U18042 (N_18042,N_16218,N_15666);
or U18043 (N_18043,N_15592,N_16912);
and U18044 (N_18044,N_15933,N_15835);
or U18045 (N_18045,N_15764,N_17429);
or U18046 (N_18046,N_15404,N_17229);
xor U18047 (N_18047,N_17240,N_16097);
or U18048 (N_18048,N_16845,N_15771);
xor U18049 (N_18049,N_15476,N_15850);
or U18050 (N_18050,N_15245,N_15146);
nand U18051 (N_18051,N_15532,N_16806);
nand U18052 (N_18052,N_16600,N_17036);
xor U18053 (N_18053,N_17357,N_15976);
nand U18054 (N_18054,N_15321,N_15776);
nor U18055 (N_18055,N_17351,N_15283);
or U18056 (N_18056,N_16377,N_17312);
or U18057 (N_18057,N_16126,N_16731);
and U18058 (N_18058,N_17400,N_16176);
nand U18059 (N_18059,N_15989,N_15898);
nand U18060 (N_18060,N_15185,N_16457);
or U18061 (N_18061,N_15159,N_16887);
and U18062 (N_18062,N_15196,N_15388);
or U18063 (N_18063,N_16872,N_16235);
xnor U18064 (N_18064,N_16202,N_15805);
nand U18065 (N_18065,N_15724,N_15043);
nor U18066 (N_18066,N_16330,N_15897);
nor U18067 (N_18067,N_15357,N_16566);
xnor U18068 (N_18068,N_15547,N_16303);
or U18069 (N_18069,N_17032,N_16537);
nand U18070 (N_18070,N_16257,N_16152);
xnor U18071 (N_18071,N_16473,N_15176);
nor U18072 (N_18072,N_16922,N_16378);
nor U18073 (N_18073,N_16436,N_15413);
nor U18074 (N_18074,N_16308,N_15132);
nand U18075 (N_18075,N_15117,N_15088);
nand U18076 (N_18076,N_15740,N_16540);
nand U18077 (N_18077,N_15838,N_16619);
xor U18078 (N_18078,N_16981,N_16156);
nor U18079 (N_18079,N_15609,N_16934);
or U18080 (N_18080,N_16831,N_16119);
xor U18081 (N_18081,N_16107,N_16828);
xor U18082 (N_18082,N_16242,N_16811);
xor U18083 (N_18083,N_15232,N_15308);
xor U18084 (N_18084,N_16408,N_15860);
xnor U18085 (N_18085,N_15672,N_15096);
nor U18086 (N_18086,N_15705,N_15686);
xnor U18087 (N_18087,N_16121,N_15056);
or U18088 (N_18088,N_16122,N_15979);
nor U18089 (N_18089,N_16101,N_16431);
nand U18090 (N_18090,N_15639,N_16732);
nand U18091 (N_18091,N_15053,N_15925);
and U18092 (N_18092,N_16111,N_15508);
nand U18093 (N_18093,N_15906,N_15175);
nand U18094 (N_18094,N_15940,N_16990);
nor U18095 (N_18095,N_16701,N_16500);
nand U18096 (N_18096,N_15387,N_16069);
nand U18097 (N_18097,N_15314,N_16722);
nand U18098 (N_18098,N_15276,N_15052);
nand U18099 (N_18099,N_16201,N_15208);
xnor U18100 (N_18100,N_17460,N_17146);
or U18101 (N_18101,N_17126,N_17409);
nor U18102 (N_18102,N_16148,N_16475);
xor U18103 (N_18103,N_16635,N_15828);
and U18104 (N_18104,N_16210,N_17077);
nand U18105 (N_18105,N_17206,N_15743);
xnor U18106 (N_18106,N_16197,N_16709);
nor U18107 (N_18107,N_16756,N_16711);
xnor U18108 (N_18108,N_15389,N_17130);
xnor U18109 (N_18109,N_17136,N_15791);
nor U18110 (N_18110,N_16451,N_17121);
nand U18111 (N_18111,N_15786,N_16893);
nor U18112 (N_18112,N_16834,N_16538);
nor U18113 (N_18113,N_16974,N_15808);
and U18114 (N_18114,N_16975,N_15438);
nor U18115 (N_18115,N_17427,N_15883);
xnor U18116 (N_18116,N_16634,N_16458);
nand U18117 (N_18117,N_15397,N_15434);
nor U18118 (N_18118,N_16996,N_15924);
or U18119 (N_18119,N_16015,N_16973);
and U18120 (N_18120,N_15270,N_17115);
nor U18121 (N_18121,N_15981,N_17332);
and U18122 (N_18122,N_17200,N_17267);
xor U18123 (N_18123,N_16306,N_16798);
xnor U18124 (N_18124,N_15278,N_15843);
nor U18125 (N_18125,N_15041,N_16181);
and U18126 (N_18126,N_16932,N_15139);
xor U18127 (N_18127,N_17406,N_15894);
and U18128 (N_18128,N_16972,N_16857);
nand U18129 (N_18129,N_17452,N_17352);
and U18130 (N_18130,N_15719,N_15944);
nor U18131 (N_18131,N_17290,N_16086);
or U18132 (N_18132,N_17322,N_15145);
nor U18133 (N_18133,N_15207,N_16784);
or U18134 (N_18134,N_15749,N_17382);
nand U18135 (N_18135,N_16191,N_16309);
and U18136 (N_18136,N_17174,N_17080);
xor U18137 (N_18137,N_17109,N_16736);
xor U18138 (N_18138,N_15960,N_15304);
or U18139 (N_18139,N_15187,N_15663);
or U18140 (N_18140,N_15323,N_15138);
or U18141 (N_18141,N_15936,N_17135);
nand U18142 (N_18142,N_16147,N_16217);
nor U18143 (N_18143,N_16535,N_16936);
xor U18144 (N_18144,N_17242,N_15429);
or U18145 (N_18145,N_15242,N_17238);
nor U18146 (N_18146,N_15670,N_17413);
or U18147 (N_18147,N_15394,N_16867);
or U18148 (N_18148,N_17398,N_15237);
xor U18149 (N_18149,N_17256,N_16727);
and U18150 (N_18150,N_16846,N_17448);
and U18151 (N_18151,N_15070,N_17067);
xnor U18152 (N_18152,N_16187,N_15001);
or U18153 (N_18153,N_15929,N_15354);
xnor U18154 (N_18154,N_17334,N_15885);
nor U18155 (N_18155,N_15507,N_15198);
nand U18156 (N_18156,N_16725,N_16752);
or U18157 (N_18157,N_15483,N_16301);
and U18158 (N_18158,N_15137,N_16853);
or U18159 (N_18159,N_16580,N_16646);
xnor U18160 (N_18160,N_16910,N_17120);
xor U18161 (N_18161,N_16746,N_17001);
and U18162 (N_18162,N_15086,N_15331);
xnor U18163 (N_18163,N_16411,N_16780);
and U18164 (N_18164,N_17454,N_15572);
nand U18165 (N_18165,N_16978,N_16658);
or U18166 (N_18166,N_15533,N_16013);
xor U18167 (N_18167,N_15938,N_17323);
or U18168 (N_18168,N_16639,N_16289);
nor U18169 (N_18169,N_16616,N_17165);
xor U18170 (N_18170,N_16836,N_16281);
nand U18171 (N_18171,N_16694,N_15188);
nand U18172 (N_18172,N_15511,N_17333);
or U18173 (N_18173,N_15853,N_15961);
and U18174 (N_18174,N_15854,N_15879);
or U18175 (N_18175,N_16838,N_16400);
and U18176 (N_18176,N_16274,N_15987);
or U18177 (N_18177,N_15915,N_17279);
xnor U18178 (N_18178,N_16595,N_16155);
and U18179 (N_18179,N_16427,N_16924);
nor U18180 (N_18180,N_16358,N_15807);
xor U18181 (N_18181,N_16503,N_17228);
nor U18182 (N_18182,N_17265,N_16481);
xor U18183 (N_18183,N_15135,N_16506);
nand U18184 (N_18184,N_15877,N_16603);
nand U18185 (N_18185,N_15846,N_15468);
xor U18186 (N_18186,N_15313,N_15967);
xnor U18187 (N_18187,N_17094,N_17041);
or U18188 (N_18188,N_16131,N_15878);
and U18189 (N_18189,N_16682,N_15398);
and U18190 (N_18190,N_17158,N_16567);
and U18191 (N_18191,N_16920,N_16895);
or U18192 (N_18192,N_15503,N_15638);
nand U18193 (N_18193,N_16573,N_16637);
xor U18194 (N_18194,N_16516,N_16667);
xor U18195 (N_18195,N_17441,N_17468);
and U18196 (N_18196,N_15986,N_16381);
and U18197 (N_18197,N_15713,N_16703);
nor U18198 (N_18198,N_16928,N_15152);
or U18199 (N_18199,N_16536,N_17278);
or U18200 (N_18200,N_15760,N_15126);
nand U18201 (N_18201,N_15792,N_17295);
nor U18202 (N_18202,N_15319,N_15416);
and U18203 (N_18203,N_16821,N_16520);
and U18204 (N_18204,N_16991,N_17361);
xor U18205 (N_18205,N_15147,N_16053);
nand U18206 (N_18206,N_15356,N_15926);
xor U18207 (N_18207,N_16588,N_15108);
or U18208 (N_18208,N_15039,N_16483);
nor U18209 (N_18209,N_15995,N_16902);
nand U18210 (N_18210,N_16204,N_16650);
xnor U18211 (N_18211,N_16749,N_17474);
and U18212 (N_18212,N_16989,N_15037);
or U18213 (N_18213,N_15658,N_17065);
nor U18214 (N_18214,N_15515,N_15369);
xor U18215 (N_18215,N_16413,N_16582);
nand U18216 (N_18216,N_15327,N_16875);
nand U18217 (N_18217,N_16000,N_15549);
and U18218 (N_18218,N_16128,N_16461);
xnor U18219 (N_18219,N_16058,N_15593);
and U18220 (N_18220,N_15732,N_15962);
nor U18221 (N_18221,N_15541,N_15643);
xnor U18222 (N_18222,N_16290,N_15556);
nor U18223 (N_18223,N_17369,N_15346);
nand U18224 (N_18224,N_16429,N_17092);
nand U18225 (N_18225,N_16333,N_17125);
xor U18226 (N_18226,N_15051,N_16394);
nor U18227 (N_18227,N_15365,N_15723);
nand U18228 (N_18228,N_17053,N_15768);
nand U18229 (N_18229,N_16950,N_15205);
nor U18230 (N_18230,N_16841,N_15215);
nor U18231 (N_18231,N_15782,N_15534);
nand U18232 (N_18232,N_15889,N_16326);
nor U18233 (N_18233,N_17218,N_15632);
xnor U18234 (N_18234,N_15097,N_16597);
and U18235 (N_18235,N_15099,N_15665);
or U18236 (N_18236,N_16921,N_17016);
xnor U18237 (N_18237,N_16266,N_16057);
xor U18238 (N_18238,N_15200,N_16955);
nand U18239 (N_18239,N_15816,N_16317);
and U18240 (N_18240,N_15386,N_17243);
or U18241 (N_18241,N_15644,N_16596);
and U18242 (N_18242,N_15580,N_17241);
xor U18243 (N_18243,N_15554,N_17410);
nor U18244 (N_18244,N_17180,N_16300);
and U18245 (N_18245,N_15863,N_15431);
and U18246 (N_18246,N_16688,N_15518);
nor U18247 (N_18247,N_15820,N_16368);
nor U18248 (N_18248,N_17259,N_16393);
nand U18249 (N_18249,N_15561,N_16734);
and U18250 (N_18250,N_17212,N_15366);
nor U18251 (N_18251,N_15057,N_15032);
xnor U18252 (N_18252,N_17183,N_17255);
nand U18253 (N_18253,N_15862,N_17131);
xor U18254 (N_18254,N_17239,N_15368);
xor U18255 (N_18255,N_15083,N_17360);
nor U18256 (N_18256,N_15044,N_17346);
or U18257 (N_18257,N_17166,N_16185);
nand U18258 (N_18258,N_15946,N_16142);
or U18259 (N_18259,N_15316,N_15543);
or U18260 (N_18260,N_16624,N_16138);
and U18261 (N_18261,N_15757,N_15834);
and U18262 (N_18262,N_15129,N_17190);
and U18263 (N_18263,N_16336,N_15700);
nand U18264 (N_18264,N_15622,N_15244);
and U18265 (N_18265,N_15836,N_15648);
and U18266 (N_18266,N_15996,N_16531);
nand U18267 (N_18267,N_15277,N_15106);
and U18268 (N_18268,N_16037,N_17433);
or U18269 (N_18269,N_16681,N_15498);
and U18270 (N_18270,N_16157,N_16958);
and U18271 (N_18271,N_15538,N_16952);
or U18272 (N_18272,N_16241,N_16294);
or U18273 (N_18273,N_17191,N_15035);
or U18274 (N_18274,N_16029,N_15362);
nand U18275 (N_18275,N_16282,N_15864);
nor U18276 (N_18276,N_16606,N_15026);
or U18277 (N_18277,N_15852,N_16165);
xnor U18278 (N_18278,N_16008,N_16296);
nor U18279 (N_18279,N_17128,N_16490);
and U18280 (N_18280,N_15169,N_15662);
or U18281 (N_18281,N_17435,N_17127);
or U18282 (N_18282,N_17424,N_16497);
nand U18283 (N_18283,N_17476,N_16033);
and U18284 (N_18284,N_15285,N_16344);
nor U18285 (N_18285,N_15871,N_16035);
nor U18286 (N_18286,N_17309,N_16943);
and U18287 (N_18287,N_15502,N_15047);
and U18288 (N_18288,N_16792,N_16010);
and U18289 (N_18289,N_15579,N_17217);
and U18290 (N_18290,N_15281,N_16283);
nor U18291 (N_18291,N_16721,N_15148);
or U18292 (N_18292,N_16918,N_15302);
or U18293 (N_18293,N_15829,N_16479);
nand U18294 (N_18294,N_16995,N_15183);
nor U18295 (N_18295,N_16448,N_16827);
xor U18296 (N_18296,N_16199,N_17139);
nand U18297 (N_18297,N_16661,N_15530);
nand U18298 (N_18298,N_15286,N_15910);
nor U18299 (N_18299,N_16823,N_15819);
xnor U18300 (N_18300,N_16276,N_17477);
nor U18301 (N_18301,N_17285,N_16470);
or U18302 (N_18302,N_16472,N_16740);
nand U18303 (N_18303,N_17273,N_15779);
nor U18304 (N_18304,N_16055,N_17467);
xor U18305 (N_18305,N_16432,N_15949);
xnor U18306 (N_18306,N_16982,N_16605);
and U18307 (N_18307,N_15315,N_15774);
or U18308 (N_18308,N_15055,N_16530);
nor U18309 (N_18309,N_15888,N_16877);
and U18310 (N_18310,N_16277,N_15815);
xnor U18311 (N_18311,N_16697,N_17310);
and U18312 (N_18312,N_17132,N_16361);
nand U18313 (N_18313,N_16438,N_15744);
nand U18314 (N_18314,N_17459,N_16747);
nor U18315 (N_18315,N_15851,N_16809);
xnor U18316 (N_18316,N_15256,N_15529);
and U18317 (N_18317,N_16911,N_16025);
nand U18318 (N_18318,N_16680,N_16651);
nor U18319 (N_18319,N_17495,N_16779);
nand U18320 (N_18320,N_17063,N_16855);
or U18321 (N_18321,N_16169,N_15250);
or U18322 (N_18322,N_15341,N_16782);
xnor U18323 (N_18323,N_17003,N_16713);
xnor U18324 (N_18324,N_15433,N_15664);
xnor U18325 (N_18325,N_15752,N_17027);
xnor U18326 (N_18326,N_16913,N_15669);
nand U18327 (N_18327,N_15761,N_17444);
and U18328 (N_18328,N_16404,N_16802);
nor U18329 (N_18329,N_16494,N_17469);
nor U18330 (N_18330,N_16642,N_15558);
and U18331 (N_18331,N_15759,N_15608);
nor U18332 (N_18332,N_16979,N_15325);
xnor U18333 (N_18333,N_16312,N_15814);
xor U18334 (N_18334,N_17012,N_15360);
or U18335 (N_18335,N_16441,N_16563);
xnor U18336 (N_18336,N_16532,N_15630);
nor U18337 (N_18337,N_17168,N_15115);
nor U18338 (N_18338,N_16864,N_17202);
or U18339 (N_18339,N_15349,N_16443);
xor U18340 (N_18340,N_15501,N_16534);
or U18341 (N_18341,N_16139,N_15880);
and U18342 (N_18342,N_17145,N_15708);
xnor U18343 (N_18343,N_17045,N_16009);
nor U18344 (N_18344,N_16586,N_15797);
and U18345 (N_18345,N_15817,N_17407);
and U18346 (N_18346,N_16239,N_16043);
and U18347 (N_18347,N_16737,N_16611);
nor U18348 (N_18348,N_15923,N_17293);
nor U18349 (N_18349,N_17188,N_15591);
nand U18350 (N_18350,N_16751,N_16066);
nand U18351 (N_18351,N_15364,N_15789);
and U18352 (N_18352,N_16279,N_17110);
nand U18353 (N_18353,N_17488,N_15886);
nand U18354 (N_18354,N_17170,N_16544);
nor U18355 (N_18355,N_16305,N_16820);
or U18356 (N_18356,N_15847,N_15796);
and U18357 (N_18357,N_15446,N_16733);
nand U18358 (N_18358,N_15007,N_17119);
nand U18359 (N_18359,N_15696,N_15856);
or U18360 (N_18360,N_16410,N_15320);
and U18361 (N_18361,N_15590,N_15122);
nor U18362 (N_18362,N_15844,N_15778);
nand U18363 (N_18363,N_15484,N_16987);
xor U18364 (N_18364,N_15613,N_16370);
xor U18365 (N_18365,N_16620,N_15358);
nand U18366 (N_18366,N_15410,N_17035);
xnor U18367 (N_18367,N_15895,N_16591);
and U18368 (N_18368,N_16104,N_17028);
or U18369 (N_18369,N_15994,N_16453);
and U18370 (N_18370,N_16618,N_17384);
or U18371 (N_18371,N_17138,N_16450);
xor U18372 (N_18372,N_15344,N_17057);
xnor U18373 (N_18373,N_16019,N_17392);
or U18374 (N_18374,N_15712,N_17358);
nand U18375 (N_18375,N_15731,N_16044);
and U18376 (N_18376,N_15295,N_15210);
nor U18377 (N_18377,N_15067,N_16089);
or U18378 (N_18378,N_15127,N_16714);
nor U18379 (N_18379,N_16446,N_17372);
nor U18380 (N_18380,N_16269,N_15017);
and U18381 (N_18381,N_17326,N_15303);
nand U18382 (N_18382,N_15226,N_16518);
nand U18383 (N_18383,N_15800,N_15206);
nor U18384 (N_18384,N_17099,N_15832);
xor U18385 (N_18385,N_17117,N_16515);
and U18386 (N_18386,N_17196,N_17111);
and U18387 (N_18387,N_17155,N_17019);
or U18388 (N_18388,N_16963,N_17042);
xor U18389 (N_18389,N_15204,N_16818);
xnor U18390 (N_18390,N_17473,N_15918);
nor U18391 (N_18391,N_15119,N_15904);
nand U18392 (N_18392,N_15201,N_17462);
nand U18393 (N_18393,N_16716,N_15401);
xor U18394 (N_18394,N_16848,N_16876);
or U18395 (N_18395,N_16863,N_16062);
nor U18396 (N_18396,N_16607,N_15312);
or U18397 (N_18397,N_15381,N_16971);
xnor U18398 (N_18398,N_15186,N_15600);
and U18399 (N_18399,N_16866,N_16435);
or U18400 (N_18400,N_15617,N_17002);
nand U18401 (N_18401,N_16299,N_17069);
xnor U18402 (N_18402,N_15424,N_15867);
nand U18403 (N_18403,N_16654,N_17161);
or U18404 (N_18404,N_15833,N_15544);
or U18405 (N_18405,N_16859,N_16064);
or U18406 (N_18406,N_15040,N_17020);
nand U18407 (N_18407,N_15071,N_15956);
nand U18408 (N_18408,N_16082,N_15479);
xor U18409 (N_18409,N_16808,N_17103);
and U18410 (N_18410,N_17284,N_17193);
nand U18411 (N_18411,N_16723,N_15254);
xor U18412 (N_18412,N_17411,N_15766);
nand U18413 (N_18413,N_16127,N_16889);
nand U18414 (N_18414,N_15546,N_16190);
nor U18415 (N_18415,N_16209,N_16477);
nand U18416 (N_18416,N_15673,N_16992);
xor U18417 (N_18417,N_16577,N_15876);
xor U18418 (N_18418,N_15195,N_16328);
nand U18419 (N_18419,N_17221,N_17186);
nor U18420 (N_18420,N_15799,N_16398);
nor U18421 (N_18421,N_15790,N_15068);
xor U18422 (N_18422,N_16090,N_17397);
xor U18423 (N_18423,N_15432,N_17129);
or U18424 (N_18424,N_15011,N_16153);
xor U18425 (N_18425,N_15332,N_15143);
or U18426 (N_18426,N_17436,N_17100);
and U18427 (N_18427,N_15228,N_15513);
nand U18428 (N_18428,N_17167,N_16247);
xor U18429 (N_18429,N_17017,N_16238);
xor U18430 (N_18430,N_16112,N_15628);
or U18431 (N_18431,N_15550,N_15577);
xnor U18432 (N_18432,N_15371,N_15707);
and U18433 (N_18433,N_17349,N_15983);
or U18434 (N_18434,N_16079,N_16145);
xnor U18435 (N_18435,N_15459,N_15455);
xnor U18436 (N_18436,N_16785,N_17123);
nand U18437 (N_18437,N_15219,N_16164);
nor U18438 (N_18438,N_15837,N_15594);
xor U18439 (N_18439,N_15326,N_15449);
xor U18440 (N_18440,N_17074,N_16743);
nor U18441 (N_18441,N_16007,N_16270);
or U18442 (N_18442,N_15674,N_16519);
nand U18443 (N_18443,N_15291,N_16629);
and U18444 (N_18444,N_17421,N_17299);
and U18445 (N_18445,N_15526,N_15029);
xnor U18446 (N_18446,N_17365,N_16604);
or U18447 (N_18447,N_15163,N_15225);
or U18448 (N_18448,N_17353,N_16488);
or U18449 (N_18449,N_16324,N_16255);
and U18450 (N_18450,N_16416,N_16367);
or U18451 (N_18451,N_16897,N_16706);
nand U18452 (N_18452,N_15454,N_17283);
xnor U18453 (N_18453,N_15980,N_16819);
xnor U18454 (N_18454,N_15181,N_15417);
and U18455 (N_18455,N_16100,N_16260);
or U18456 (N_18456,N_15734,N_16083);
nor U18457 (N_18457,N_16960,N_16486);
nand U18458 (N_18458,N_17450,N_16396);
or U18459 (N_18459,N_17403,N_15240);
nor U18460 (N_18460,N_15042,N_16392);
or U18461 (N_18461,N_16648,N_16822);
and U18462 (N_18462,N_15390,N_15717);
nand U18463 (N_18463,N_16501,N_16038);
nand U18464 (N_18464,N_17280,N_16707);
nand U18465 (N_18465,N_16938,N_17308);
xnor U18466 (N_18466,N_17412,N_15182);
nor U18467 (N_18467,N_15920,N_15118);
and U18468 (N_18468,N_16551,N_15149);
nand U18469 (N_18469,N_16750,N_15218);
xnor U18470 (N_18470,N_17393,N_17379);
xnor U18471 (N_18471,N_15022,N_16385);
xnor U18472 (N_18472,N_17401,N_15033);
xnor U18473 (N_18473,N_15581,N_15460);
xor U18474 (N_18474,N_17072,N_16548);
xnor U18475 (N_18475,N_16719,N_15239);
or U18476 (N_18476,N_16076,N_15048);
xor U18477 (N_18477,N_17324,N_15997);
xnor U18478 (N_18478,N_15229,N_15625);
and U18479 (N_18479,N_16757,N_15818);
and U18480 (N_18480,N_16858,N_15442);
or U18481 (N_18481,N_15437,N_15098);
nand U18482 (N_18482,N_15076,N_16762);
or U18483 (N_18483,N_16442,N_16258);
nand U18484 (N_18484,N_17266,N_15722);
xnor U18485 (N_18485,N_15629,N_16965);
xor U18486 (N_18486,N_16847,N_16349);
or U18487 (N_18487,N_17102,N_16223);
or U18488 (N_18488,N_17364,N_16903);
nand U18489 (N_18489,N_16331,N_15190);
or U18490 (N_18490,N_15112,N_16137);
xnor U18491 (N_18491,N_16449,N_16447);
nand U18492 (N_18492,N_15393,N_17162);
xnor U18493 (N_18493,N_16571,N_16017);
xnor U18494 (N_18494,N_15447,N_15472);
nor U18495 (N_18495,N_16804,N_17133);
and U18496 (N_18496,N_15647,N_15523);
nor U18497 (N_18497,N_16278,N_15742);
and U18498 (N_18498,N_16685,N_15619);
or U18499 (N_18499,N_15736,N_15984);
xor U18500 (N_18500,N_17251,N_15963);
nand U18501 (N_18501,N_15473,N_15246);
nor U18502 (N_18502,N_15258,N_15120);
or U18503 (N_18503,N_15264,N_16251);
nor U18504 (N_18504,N_17232,N_15627);
xor U18505 (N_18505,N_16587,N_16339);
xor U18506 (N_18506,N_16901,N_16335);
nor U18507 (N_18507,N_16014,N_15865);
nand U18508 (N_18508,N_17088,N_16113);
nand U18509 (N_18509,N_17274,N_17307);
or U18510 (N_18510,N_16354,N_17291);
xor U18511 (N_18511,N_15733,N_17050);
nand U18512 (N_18512,N_15959,N_15355);
nor U18513 (N_18513,N_17219,N_15917);
nor U18514 (N_18514,N_16940,N_17197);
nor U18515 (N_18515,N_16206,N_15887);
nor U18516 (N_18516,N_16489,N_16554);
or U18517 (N_18517,N_16581,N_15977);
nor U18518 (N_18518,N_15939,N_16969);
or U18519 (N_18519,N_17275,N_16214);
and U18520 (N_18520,N_17171,N_17388);
or U18521 (N_18521,N_15992,N_17405);
and U18522 (N_18522,N_17231,N_17021);
or U18523 (N_18523,N_15485,N_15060);
xor U18524 (N_18524,N_16437,N_15160);
nor U18525 (N_18525,N_16547,N_16815);
xor U18526 (N_18526,N_15085,N_15583);
and U18527 (N_18527,N_15311,N_15402);
xnor U18528 (N_18528,N_15930,N_15370);
and U18529 (N_18529,N_16825,N_16578);
and U18530 (N_18530,N_15721,N_16564);
nor U18531 (N_18531,N_16049,N_15050);
or U18532 (N_18532,N_17049,N_16288);
or U18533 (N_18533,N_16888,N_15659);
nand U18534 (N_18534,N_16865,N_16130);
or U18535 (N_18535,N_15488,N_15937);
nor U18536 (N_18536,N_17432,N_15305);
and U18537 (N_18537,N_17018,N_17260);
nor U18538 (N_18538,N_16166,N_17164);
xor U18539 (N_18539,N_17288,N_17387);
and U18540 (N_18540,N_16120,N_17272);
nor U18541 (N_18541,N_16919,N_15874);
nor U18542 (N_18542,N_15597,N_17329);
xnor U18543 (N_18543,N_15224,N_15012);
nand U18544 (N_18544,N_17327,N_17178);
and U18545 (N_18545,N_16171,N_15857);
and U18546 (N_18546,N_15777,N_15363);
nor U18547 (N_18547,N_15998,N_16840);
nand U18548 (N_18548,N_15077,N_16851);
xor U18549 (N_18549,N_16254,N_16364);
or U18550 (N_18550,N_16136,N_17374);
and U18551 (N_18551,N_16110,N_15793);
or U18552 (N_18552,N_16775,N_15727);
xnor U18553 (N_18553,N_16200,N_16487);
or U18554 (N_18554,N_16574,N_17144);
nor U18555 (N_18555,N_15336,N_15787);
xnor U18556 (N_18556,N_15367,N_15767);
xnor U18557 (N_18557,N_15491,N_16878);
nor U18558 (N_18558,N_17216,N_16759);
and U18559 (N_18559,N_17056,N_16514);
xor U18560 (N_18560,N_16572,N_15826);
xor U18561 (N_18561,N_16248,N_15564);
xnor U18562 (N_18562,N_16172,N_16976);
xor U18563 (N_18563,N_15194,N_16322);
and U18564 (N_18564,N_16271,N_17300);
and U18565 (N_18565,N_15565,N_15462);
nor U18566 (N_18566,N_17381,N_15694);
nand U18567 (N_18567,N_16686,N_16237);
nand U18568 (N_18568,N_15350,N_15578);
and U18569 (N_18569,N_15748,N_16081);
or U18570 (N_18570,N_16925,N_15495);
nor U18571 (N_18571,N_16679,N_15262);
nor U18572 (N_18572,N_16899,N_17325);
xnor U18573 (N_18573,N_16905,N_16896);
nand U18574 (N_18574,N_15522,N_16123);
and U18575 (N_18575,N_16994,N_15562);
xnor U18576 (N_18576,N_16310,N_16482);
xor U18577 (N_18577,N_15510,N_15260);
or U18578 (N_18578,N_16652,N_15297);
and U18579 (N_18579,N_16264,N_17087);
xnor U18580 (N_18580,N_15825,N_15729);
and U18581 (N_18581,N_17371,N_15418);
nand U18582 (N_18582,N_17437,N_15614);
nor U18583 (N_18583,N_16626,N_16188);
xor U18584 (N_18584,N_15253,N_17151);
and U18585 (N_18585,N_17235,N_16854);
nor U18586 (N_18586,N_15199,N_15676);
nand U18587 (N_18587,N_16718,N_15735);
nand U18588 (N_18588,N_17192,N_16942);
nor U18589 (N_18589,N_16109,N_16874);
or U18590 (N_18590,N_17261,N_15428);
nand U18591 (N_18591,N_17185,N_15310);
and U18592 (N_18592,N_15677,N_17321);
nor U18593 (N_18593,N_15238,N_17043);
nand U18594 (N_18594,N_16060,N_17342);
and U18595 (N_18595,N_16984,N_15750);
or U18596 (N_18596,N_17363,N_16027);
or U18597 (N_18597,N_16430,N_15248);
nand U18598 (N_18598,N_16313,N_15125);
nand U18599 (N_18599,N_15243,N_17425);
xnor U18600 (N_18600,N_16524,N_16953);
or U18601 (N_18601,N_16826,N_15471);
and U18602 (N_18602,N_16389,N_17271);
and U18603 (N_18603,N_17337,N_15174);
xor U18604 (N_18604,N_15504,N_15831);
nand U18605 (N_18605,N_17173,N_16407);
nand U18606 (N_18606,N_16640,N_16352);
nand U18607 (N_18607,N_15982,N_16225);
or U18608 (N_18608,N_15811,N_16045);
and U18609 (N_18609,N_15972,N_16843);
and U18610 (N_18610,N_16507,N_15599);
or U18611 (N_18611,N_16243,N_17455);
and U18612 (N_18612,N_16509,N_15943);
xor U18613 (N_18613,N_16095,N_16493);
nand U18614 (N_18614,N_17306,N_16623);
nor U18615 (N_18615,N_17289,N_15107);
or U18616 (N_18616,N_16228,N_16777);
nand U18617 (N_18617,N_16345,N_15230);
or U18618 (N_18618,N_16341,N_15985);
nor U18619 (N_18619,N_16068,N_16316);
nor U18620 (N_18620,N_16763,N_16884);
and U18621 (N_18621,N_17007,N_17496);
nor U18622 (N_18622,N_16702,N_15166);
nor U18623 (N_18623,N_16362,N_16787);
nor U18624 (N_18624,N_15896,N_15392);
nand U18625 (N_18625,N_16491,N_17338);
nor U18626 (N_18626,N_16575,N_15063);
xnor U18627 (N_18627,N_15025,N_17134);
nand U18628 (N_18628,N_15804,N_15002);
nand U18629 (N_18629,N_16373,N_16067);
xor U18630 (N_18630,N_16862,N_15453);
and U18631 (N_18631,N_15568,N_15452);
xnor U18632 (N_18632,N_15971,N_16395);
nand U18633 (N_18633,N_15469,N_15347);
nand U18634 (N_18634,N_15762,N_16948);
nor U18635 (N_18635,N_15781,N_15180);
nand U18636 (N_18636,N_16132,N_17029);
nand U18637 (N_18637,N_16135,N_17154);
xor U18638 (N_18638,N_17223,N_16077);
nand U18639 (N_18639,N_15267,N_15104);
and U18640 (N_18640,N_15684,N_17262);
xor U18641 (N_18641,N_17270,N_15113);
nand U18642 (N_18642,N_15633,N_15601);
xor U18643 (N_18643,N_16615,N_15130);
or U18644 (N_18644,N_15716,N_15403);
xnor U18645 (N_18645,N_15333,N_17367);
nand U18646 (N_18646,N_15289,N_15008);
nor U18647 (N_18647,N_16881,N_17106);
or U18648 (N_18648,N_16510,N_15383);
nor U18649 (N_18649,N_16177,N_15287);
xor U18650 (N_18650,N_17249,N_16929);
nand U18651 (N_18651,N_16216,N_16998);
nand U18652 (N_18652,N_16764,N_16319);
nor U18653 (N_18653,N_16505,N_15439);
nand U18654 (N_18654,N_16042,N_17024);
xnor U18655 (N_18655,N_16215,N_17375);
and U18656 (N_18656,N_15499,N_15509);
or U18657 (N_18657,N_15932,N_16304);
or U18658 (N_18658,N_16517,N_17470);
nor U18659 (N_18659,N_17204,N_17252);
and U18660 (N_18660,N_15842,N_16868);
xnor U18661 (N_18661,N_17486,N_16280);
or U18662 (N_18662,N_17082,N_16968);
or U18663 (N_18663,N_15406,N_15795);
nor U18664 (N_18664,N_16028,N_16871);
or U18665 (N_18665,N_15869,N_17415);
xnor U18666 (N_18666,N_15456,N_15038);
and U18667 (N_18667,N_17254,N_16434);
nor U18668 (N_18668,N_16168,N_15173);
nand U18669 (N_18669,N_15249,N_15566);
and U18670 (N_18670,N_16321,N_16263);
nor U18671 (N_18671,N_17317,N_15269);
and U18672 (N_18672,N_16250,N_16184);
nor U18673 (N_18673,N_16366,N_16812);
nor U18674 (N_18674,N_16791,N_17408);
xnor U18675 (N_18675,N_17090,N_17294);
and U18676 (N_18676,N_17442,N_16583);
nand U18677 (N_18677,N_16883,N_17004);
nor U18678 (N_18678,N_16528,N_15084);
xnor U18679 (N_18679,N_15299,N_16003);
nor U18680 (N_18680,N_16259,N_16262);
and U18681 (N_18681,N_16415,N_16949);
or U18682 (N_18682,N_15324,N_16695);
nor U18683 (N_18683,N_16080,N_16692);
xor U18684 (N_18684,N_15141,N_15948);
or U18685 (N_18685,N_15203,N_16673);
or U18686 (N_18686,N_15571,N_15480);
nor U18687 (N_18687,N_16048,N_15110);
nand U18688 (N_18688,N_15806,N_16189);
or U18689 (N_18689,N_16513,N_16622);
nand U18690 (N_18690,N_15003,N_15492);
nand U18691 (N_18691,N_17414,N_16094);
nand U18692 (N_18692,N_15754,N_15343);
nand U18693 (N_18693,N_16830,N_15548);
xnor U18694 (N_18694,N_16602,N_15140);
and U18695 (N_18695,N_15651,N_16433);
nor U18696 (N_18696,N_15873,N_17187);
nor U18697 (N_18697,N_17157,N_17416);
xnor U18698 (N_18698,N_15567,N_15646);
nand U18699 (N_18699,N_16937,N_17234);
and U18700 (N_18700,N_15102,N_17493);
nand U18701 (N_18701,N_16796,N_17456);
nand U18702 (N_18702,N_15884,N_16031);
nor U18703 (N_18703,N_17314,N_15810);
nor U18704 (N_18704,N_17373,N_16556);
or U18705 (N_18705,N_16374,N_16246);
nand U18706 (N_18706,N_17156,N_15570);
nor U18707 (N_18707,N_16084,N_16231);
nor U18708 (N_18708,N_15069,N_15213);
and U18709 (N_18709,N_15093,N_15054);
nor U18710 (N_18710,N_16422,N_16609);
and U18711 (N_18711,N_16805,N_16653);
xnor U18712 (N_18712,N_17213,N_16298);
nor U18713 (N_18713,N_15154,N_17376);
and U18714 (N_18714,N_16445,N_16907);
xnor U18715 (N_18715,N_16471,N_15641);
nor U18716 (N_18716,N_16641,N_15687);
and U18717 (N_18717,N_16133,N_16227);
xor U18718 (N_18718,N_16967,N_16314);
nor U18719 (N_18719,N_17207,N_15725);
nand U18720 (N_18720,N_16154,N_16256);
and U18721 (N_18721,N_17287,N_16541);
nand U18722 (N_18722,N_16860,N_15445);
and U18723 (N_18723,N_16735,N_16205);
nor U18724 (N_18724,N_15134,N_16372);
nor U18725 (N_18725,N_17264,N_15770);
xnor U18726 (N_18726,N_16065,N_15241);
nor U18727 (N_18727,N_17061,N_16141);
and U18728 (N_18728,N_16286,N_15802);
xor U18729 (N_18729,N_17172,N_15784);
nor U18730 (N_18730,N_17268,N_15466);
and U18731 (N_18731,N_16891,N_16252);
or U18732 (N_18732,N_16021,N_16229);
xor U18733 (N_18733,N_16371,N_15189);
and U18734 (N_18734,N_15074,N_16093);
nor U18735 (N_18735,N_16589,N_16420);
xor U18736 (N_18736,N_15607,N_16672);
nand U18737 (N_18737,N_17009,N_15706);
or U18738 (N_18738,N_16340,N_15531);
and U18739 (N_18739,N_15380,N_15265);
or U18740 (N_18740,N_16403,N_16343);
or U18741 (N_18741,N_16388,N_16384);
nor U18742 (N_18742,N_17137,N_17313);
or U18743 (N_18743,N_15634,N_16744);
or U18744 (N_18744,N_17085,N_16767);
xor U18745 (N_18745,N_16997,N_16098);
and U18746 (N_18746,N_15405,N_17445);
and U18747 (N_18747,N_17014,N_16643);
nand U18748 (N_18748,N_16772,N_16753);
xnor U18749 (N_18749,N_17211,N_17066);
or U18750 (N_18750,N_15086,N_16499);
xnor U18751 (N_18751,N_16536,N_15629);
or U18752 (N_18752,N_16549,N_17249);
xor U18753 (N_18753,N_17419,N_15259);
and U18754 (N_18754,N_17085,N_17103);
xnor U18755 (N_18755,N_16348,N_16636);
xor U18756 (N_18756,N_15552,N_15940);
nand U18757 (N_18757,N_16575,N_15382);
xnor U18758 (N_18758,N_15214,N_16149);
or U18759 (N_18759,N_15546,N_15635);
nand U18760 (N_18760,N_15680,N_17100);
nand U18761 (N_18761,N_17442,N_15368);
nand U18762 (N_18762,N_15702,N_16491);
xnor U18763 (N_18763,N_16810,N_16408);
xor U18764 (N_18764,N_17445,N_16376);
xnor U18765 (N_18765,N_16815,N_16182);
nor U18766 (N_18766,N_15944,N_17051);
and U18767 (N_18767,N_15586,N_16540);
xnor U18768 (N_18768,N_17246,N_15609);
nand U18769 (N_18769,N_15333,N_17120);
and U18770 (N_18770,N_16375,N_17186);
xnor U18771 (N_18771,N_15950,N_15462);
xnor U18772 (N_18772,N_15949,N_15672);
nor U18773 (N_18773,N_15132,N_17462);
and U18774 (N_18774,N_15147,N_15596);
nor U18775 (N_18775,N_15213,N_15992);
nand U18776 (N_18776,N_16325,N_17363);
xor U18777 (N_18777,N_16292,N_17425);
or U18778 (N_18778,N_16204,N_15237);
or U18779 (N_18779,N_16480,N_16690);
xor U18780 (N_18780,N_17392,N_17395);
nor U18781 (N_18781,N_15116,N_16843);
or U18782 (N_18782,N_15956,N_16147);
xnor U18783 (N_18783,N_17127,N_15526);
nor U18784 (N_18784,N_16035,N_15046);
and U18785 (N_18785,N_15021,N_15718);
xor U18786 (N_18786,N_17155,N_15649);
xor U18787 (N_18787,N_17367,N_16479);
nand U18788 (N_18788,N_17464,N_17335);
nor U18789 (N_18789,N_15165,N_16883);
and U18790 (N_18790,N_15853,N_16685);
xnor U18791 (N_18791,N_17082,N_16158);
or U18792 (N_18792,N_15844,N_16115);
and U18793 (N_18793,N_17307,N_15608);
nor U18794 (N_18794,N_17002,N_15076);
nand U18795 (N_18795,N_17062,N_16307);
and U18796 (N_18796,N_17164,N_15098);
and U18797 (N_18797,N_15552,N_15257);
xor U18798 (N_18798,N_16677,N_15172);
nor U18799 (N_18799,N_15267,N_17136);
and U18800 (N_18800,N_15588,N_16447);
or U18801 (N_18801,N_16053,N_15328);
nor U18802 (N_18802,N_15654,N_15269);
or U18803 (N_18803,N_15561,N_15201);
nor U18804 (N_18804,N_15930,N_16344);
or U18805 (N_18805,N_16768,N_16343);
xnor U18806 (N_18806,N_15694,N_15159);
or U18807 (N_18807,N_16403,N_15287);
nand U18808 (N_18808,N_16358,N_15871);
xor U18809 (N_18809,N_15098,N_15598);
xor U18810 (N_18810,N_16231,N_15985);
or U18811 (N_18811,N_16420,N_16951);
xor U18812 (N_18812,N_15416,N_16915);
or U18813 (N_18813,N_15661,N_16709);
nor U18814 (N_18814,N_17023,N_17318);
and U18815 (N_18815,N_17216,N_16197);
nor U18816 (N_18816,N_16869,N_17235);
xor U18817 (N_18817,N_16723,N_16044);
or U18818 (N_18818,N_16988,N_16931);
or U18819 (N_18819,N_15597,N_17142);
nor U18820 (N_18820,N_17308,N_15642);
xor U18821 (N_18821,N_15475,N_15312);
xor U18822 (N_18822,N_15316,N_15280);
or U18823 (N_18823,N_16930,N_15191);
nor U18824 (N_18824,N_16702,N_16684);
and U18825 (N_18825,N_17357,N_16609);
and U18826 (N_18826,N_15152,N_16864);
xor U18827 (N_18827,N_15111,N_17442);
and U18828 (N_18828,N_15100,N_16103);
nor U18829 (N_18829,N_15428,N_16535);
nor U18830 (N_18830,N_15622,N_15725);
or U18831 (N_18831,N_16868,N_17009);
nor U18832 (N_18832,N_15311,N_16190);
xor U18833 (N_18833,N_15812,N_15742);
or U18834 (N_18834,N_16282,N_17321);
nor U18835 (N_18835,N_15619,N_15728);
nor U18836 (N_18836,N_16667,N_15862);
nor U18837 (N_18837,N_16342,N_17435);
xor U18838 (N_18838,N_16305,N_17488);
or U18839 (N_18839,N_16892,N_15239);
and U18840 (N_18840,N_15267,N_16935);
xor U18841 (N_18841,N_15516,N_16861);
nor U18842 (N_18842,N_17282,N_16193);
nand U18843 (N_18843,N_16125,N_16602);
and U18844 (N_18844,N_16526,N_15073);
nor U18845 (N_18845,N_16564,N_15322);
and U18846 (N_18846,N_15673,N_16433);
nand U18847 (N_18847,N_17493,N_17245);
and U18848 (N_18848,N_15508,N_16567);
xnor U18849 (N_18849,N_16704,N_16580);
and U18850 (N_18850,N_17172,N_15687);
or U18851 (N_18851,N_17106,N_15658);
or U18852 (N_18852,N_15573,N_16568);
xnor U18853 (N_18853,N_15505,N_16505);
or U18854 (N_18854,N_17018,N_16750);
nor U18855 (N_18855,N_15608,N_16426);
nand U18856 (N_18856,N_16992,N_15469);
and U18857 (N_18857,N_16486,N_16164);
xor U18858 (N_18858,N_15097,N_15254);
nand U18859 (N_18859,N_16483,N_17027);
nand U18860 (N_18860,N_16185,N_16031);
or U18861 (N_18861,N_16075,N_15068);
xnor U18862 (N_18862,N_16729,N_16724);
nand U18863 (N_18863,N_16259,N_15121);
xnor U18864 (N_18864,N_16943,N_15604);
or U18865 (N_18865,N_15787,N_15716);
nor U18866 (N_18866,N_16547,N_15932);
and U18867 (N_18867,N_15631,N_15562);
or U18868 (N_18868,N_16164,N_17341);
nand U18869 (N_18869,N_15486,N_16094);
and U18870 (N_18870,N_16753,N_16101);
xor U18871 (N_18871,N_15369,N_16893);
nor U18872 (N_18872,N_17218,N_15736);
xor U18873 (N_18873,N_15891,N_15350);
xnor U18874 (N_18874,N_17228,N_16543);
xor U18875 (N_18875,N_17409,N_16326);
or U18876 (N_18876,N_16048,N_15092);
xor U18877 (N_18877,N_16974,N_15168);
xnor U18878 (N_18878,N_15436,N_15163);
nor U18879 (N_18879,N_17034,N_16090);
or U18880 (N_18880,N_17132,N_15678);
or U18881 (N_18881,N_17464,N_16236);
xor U18882 (N_18882,N_17188,N_15768);
nor U18883 (N_18883,N_15198,N_15124);
or U18884 (N_18884,N_15583,N_15339);
nor U18885 (N_18885,N_15976,N_16653);
and U18886 (N_18886,N_15051,N_17479);
or U18887 (N_18887,N_16941,N_16324);
xnor U18888 (N_18888,N_17171,N_15282);
nor U18889 (N_18889,N_15001,N_16578);
nand U18890 (N_18890,N_15181,N_16217);
or U18891 (N_18891,N_17235,N_15887);
nor U18892 (N_18892,N_15294,N_15506);
xor U18893 (N_18893,N_15292,N_16099);
and U18894 (N_18894,N_16983,N_15628);
nand U18895 (N_18895,N_15424,N_16059);
xnor U18896 (N_18896,N_15400,N_16161);
and U18897 (N_18897,N_15223,N_16337);
nor U18898 (N_18898,N_15625,N_16654);
nand U18899 (N_18899,N_16058,N_15003);
and U18900 (N_18900,N_16353,N_15171);
and U18901 (N_18901,N_15741,N_16088);
or U18902 (N_18902,N_15887,N_15440);
nand U18903 (N_18903,N_16157,N_16694);
nor U18904 (N_18904,N_16753,N_16378);
xor U18905 (N_18905,N_16090,N_15535);
and U18906 (N_18906,N_15834,N_15395);
nand U18907 (N_18907,N_16724,N_17342);
nor U18908 (N_18908,N_15438,N_15919);
and U18909 (N_18909,N_16821,N_16877);
and U18910 (N_18910,N_16964,N_15686);
and U18911 (N_18911,N_15995,N_15913);
xnor U18912 (N_18912,N_16773,N_16136);
xor U18913 (N_18913,N_15068,N_16974);
and U18914 (N_18914,N_17273,N_17242);
nand U18915 (N_18915,N_15344,N_17129);
xor U18916 (N_18916,N_15191,N_15370);
nand U18917 (N_18917,N_15344,N_17437);
nor U18918 (N_18918,N_17051,N_16022);
or U18919 (N_18919,N_16627,N_15899);
or U18920 (N_18920,N_17269,N_15859);
nor U18921 (N_18921,N_16562,N_15214);
nor U18922 (N_18922,N_15903,N_15703);
nor U18923 (N_18923,N_15654,N_15632);
nand U18924 (N_18924,N_16968,N_16563);
nor U18925 (N_18925,N_15452,N_16300);
nor U18926 (N_18926,N_15556,N_15070);
and U18927 (N_18927,N_16949,N_16377);
xnor U18928 (N_18928,N_16987,N_17333);
nor U18929 (N_18929,N_16874,N_17256);
or U18930 (N_18930,N_15646,N_15537);
or U18931 (N_18931,N_17382,N_15170);
xnor U18932 (N_18932,N_15792,N_15483);
nand U18933 (N_18933,N_16594,N_16099);
xor U18934 (N_18934,N_17344,N_15684);
nor U18935 (N_18935,N_16807,N_15808);
xor U18936 (N_18936,N_16260,N_16418);
nand U18937 (N_18937,N_17136,N_16095);
or U18938 (N_18938,N_17473,N_16264);
nor U18939 (N_18939,N_17296,N_15634);
or U18940 (N_18940,N_17155,N_15485);
nor U18941 (N_18941,N_15039,N_17302);
nor U18942 (N_18942,N_16718,N_16407);
xor U18943 (N_18943,N_15020,N_15622);
nor U18944 (N_18944,N_16594,N_17369);
or U18945 (N_18945,N_15322,N_15100);
nand U18946 (N_18946,N_16095,N_15419);
nor U18947 (N_18947,N_16777,N_15190);
nand U18948 (N_18948,N_17032,N_15427);
nor U18949 (N_18949,N_16077,N_16387);
xor U18950 (N_18950,N_15627,N_16676);
nor U18951 (N_18951,N_15083,N_16816);
and U18952 (N_18952,N_15221,N_17091);
xnor U18953 (N_18953,N_15444,N_15447);
or U18954 (N_18954,N_15114,N_17007);
and U18955 (N_18955,N_15993,N_17085);
and U18956 (N_18956,N_16113,N_16718);
and U18957 (N_18957,N_15876,N_15976);
or U18958 (N_18958,N_16389,N_16957);
or U18959 (N_18959,N_17298,N_15837);
and U18960 (N_18960,N_16324,N_16220);
and U18961 (N_18961,N_16792,N_15646);
xor U18962 (N_18962,N_16974,N_15411);
and U18963 (N_18963,N_15080,N_15620);
or U18964 (N_18964,N_15630,N_15619);
xor U18965 (N_18965,N_16532,N_16676);
and U18966 (N_18966,N_15892,N_17245);
nand U18967 (N_18967,N_17413,N_16633);
nor U18968 (N_18968,N_17118,N_17433);
nor U18969 (N_18969,N_15587,N_15605);
xor U18970 (N_18970,N_15709,N_15475);
nand U18971 (N_18971,N_16414,N_17377);
or U18972 (N_18972,N_17178,N_17341);
or U18973 (N_18973,N_15535,N_17285);
nand U18974 (N_18974,N_16035,N_17331);
or U18975 (N_18975,N_15530,N_15553);
nor U18976 (N_18976,N_16335,N_17007);
xor U18977 (N_18977,N_15627,N_16237);
nand U18978 (N_18978,N_16705,N_15425);
nand U18979 (N_18979,N_16527,N_16125);
xor U18980 (N_18980,N_17455,N_15993);
and U18981 (N_18981,N_16891,N_16472);
nor U18982 (N_18982,N_15040,N_17365);
xnor U18983 (N_18983,N_15462,N_17159);
or U18984 (N_18984,N_17312,N_16244);
nand U18985 (N_18985,N_16231,N_17011);
nand U18986 (N_18986,N_16361,N_16815);
or U18987 (N_18987,N_16988,N_15753);
or U18988 (N_18988,N_17465,N_17332);
or U18989 (N_18989,N_15540,N_15904);
or U18990 (N_18990,N_15935,N_15564);
xnor U18991 (N_18991,N_15250,N_16344);
nand U18992 (N_18992,N_16693,N_17231);
nor U18993 (N_18993,N_17446,N_17118);
nor U18994 (N_18994,N_17419,N_16019);
and U18995 (N_18995,N_17163,N_17476);
nor U18996 (N_18996,N_16923,N_16522);
xnor U18997 (N_18997,N_17365,N_16008);
or U18998 (N_18998,N_16642,N_17218);
nor U18999 (N_18999,N_17152,N_17243);
and U19000 (N_19000,N_17394,N_16423);
nor U19001 (N_19001,N_15288,N_15602);
xnor U19002 (N_19002,N_16176,N_15538);
nor U19003 (N_19003,N_16462,N_15645);
xor U19004 (N_19004,N_16981,N_15085);
nor U19005 (N_19005,N_16843,N_17267);
nor U19006 (N_19006,N_17105,N_15440);
xnor U19007 (N_19007,N_17351,N_17459);
xor U19008 (N_19008,N_16119,N_17213);
nor U19009 (N_19009,N_15086,N_15828);
nand U19010 (N_19010,N_16204,N_15014);
or U19011 (N_19011,N_17031,N_15757);
and U19012 (N_19012,N_16000,N_15505);
nor U19013 (N_19013,N_17267,N_15290);
nor U19014 (N_19014,N_16548,N_15907);
or U19015 (N_19015,N_16209,N_15061);
xnor U19016 (N_19016,N_15592,N_16546);
nor U19017 (N_19017,N_16114,N_15637);
and U19018 (N_19018,N_16844,N_16367);
or U19019 (N_19019,N_17064,N_15046);
nand U19020 (N_19020,N_15331,N_15305);
or U19021 (N_19021,N_15841,N_16265);
nor U19022 (N_19022,N_15303,N_16617);
nand U19023 (N_19023,N_16451,N_16253);
xor U19024 (N_19024,N_17405,N_16015);
and U19025 (N_19025,N_16754,N_16900);
nor U19026 (N_19026,N_17280,N_15349);
or U19027 (N_19027,N_15784,N_15993);
xor U19028 (N_19028,N_15078,N_17186);
nand U19029 (N_19029,N_16404,N_15111);
or U19030 (N_19030,N_17319,N_15667);
nand U19031 (N_19031,N_16281,N_17129);
nor U19032 (N_19032,N_16365,N_15036);
or U19033 (N_19033,N_15136,N_15720);
nor U19034 (N_19034,N_15386,N_15055);
and U19035 (N_19035,N_16163,N_16337);
xor U19036 (N_19036,N_15385,N_16737);
or U19037 (N_19037,N_16046,N_15121);
or U19038 (N_19038,N_16469,N_15228);
nor U19039 (N_19039,N_15087,N_17093);
and U19040 (N_19040,N_15366,N_15596);
and U19041 (N_19041,N_15650,N_17264);
xor U19042 (N_19042,N_17040,N_15070);
and U19043 (N_19043,N_16248,N_16845);
xnor U19044 (N_19044,N_15171,N_17072);
or U19045 (N_19045,N_15933,N_15404);
or U19046 (N_19046,N_15257,N_15869);
nand U19047 (N_19047,N_15243,N_17103);
and U19048 (N_19048,N_15637,N_16718);
xnor U19049 (N_19049,N_15483,N_15793);
nor U19050 (N_19050,N_16171,N_15405);
nand U19051 (N_19051,N_17064,N_15214);
and U19052 (N_19052,N_15094,N_15439);
or U19053 (N_19053,N_15729,N_15581);
nand U19054 (N_19054,N_16634,N_16174);
nand U19055 (N_19055,N_15359,N_15210);
nor U19056 (N_19056,N_16324,N_16640);
xor U19057 (N_19057,N_17387,N_15304);
or U19058 (N_19058,N_15348,N_17049);
nor U19059 (N_19059,N_17438,N_16805);
nand U19060 (N_19060,N_15802,N_16789);
and U19061 (N_19061,N_15965,N_17459);
xor U19062 (N_19062,N_15053,N_15499);
xnor U19063 (N_19063,N_15440,N_17322);
nand U19064 (N_19064,N_15179,N_15072);
nand U19065 (N_19065,N_16945,N_15425);
or U19066 (N_19066,N_16526,N_15400);
xor U19067 (N_19067,N_15641,N_16788);
xor U19068 (N_19068,N_16420,N_15742);
nor U19069 (N_19069,N_17113,N_16824);
xnor U19070 (N_19070,N_15779,N_16556);
nor U19071 (N_19071,N_15769,N_16461);
or U19072 (N_19072,N_15403,N_15224);
xnor U19073 (N_19073,N_16327,N_15711);
and U19074 (N_19074,N_15184,N_15952);
or U19075 (N_19075,N_16883,N_16439);
nand U19076 (N_19076,N_15473,N_16415);
xor U19077 (N_19077,N_15145,N_16644);
nand U19078 (N_19078,N_16584,N_16741);
or U19079 (N_19079,N_16141,N_17079);
xnor U19080 (N_19080,N_16217,N_16621);
xor U19081 (N_19081,N_17156,N_17390);
and U19082 (N_19082,N_16486,N_16974);
xor U19083 (N_19083,N_15118,N_16087);
or U19084 (N_19084,N_15085,N_15477);
nand U19085 (N_19085,N_17127,N_15585);
or U19086 (N_19086,N_16028,N_16652);
xor U19087 (N_19087,N_17267,N_15978);
and U19088 (N_19088,N_15932,N_16266);
xor U19089 (N_19089,N_16072,N_15130);
nor U19090 (N_19090,N_16360,N_16807);
or U19091 (N_19091,N_16008,N_16821);
or U19092 (N_19092,N_16713,N_16710);
nor U19093 (N_19093,N_15222,N_16382);
xor U19094 (N_19094,N_15961,N_16958);
or U19095 (N_19095,N_15135,N_16916);
xor U19096 (N_19096,N_17465,N_15404);
nand U19097 (N_19097,N_16928,N_15709);
or U19098 (N_19098,N_17184,N_16050);
or U19099 (N_19099,N_16735,N_17356);
nor U19100 (N_19100,N_15701,N_16597);
nor U19101 (N_19101,N_15784,N_16174);
or U19102 (N_19102,N_16375,N_15194);
xor U19103 (N_19103,N_15503,N_16138);
and U19104 (N_19104,N_16536,N_15626);
nor U19105 (N_19105,N_16941,N_15558);
or U19106 (N_19106,N_15317,N_17149);
nor U19107 (N_19107,N_15965,N_15368);
and U19108 (N_19108,N_15247,N_15085);
xor U19109 (N_19109,N_16218,N_17223);
xnor U19110 (N_19110,N_16045,N_16406);
or U19111 (N_19111,N_15904,N_16861);
nor U19112 (N_19112,N_15841,N_17095);
nor U19113 (N_19113,N_16191,N_15624);
nor U19114 (N_19114,N_16835,N_16226);
and U19115 (N_19115,N_15793,N_16897);
nand U19116 (N_19116,N_16682,N_16032);
and U19117 (N_19117,N_15401,N_15028);
nor U19118 (N_19118,N_15539,N_16024);
or U19119 (N_19119,N_15221,N_15144);
and U19120 (N_19120,N_17115,N_15515);
or U19121 (N_19121,N_15177,N_15153);
nor U19122 (N_19122,N_15390,N_16542);
and U19123 (N_19123,N_17048,N_15098);
or U19124 (N_19124,N_17025,N_16846);
nand U19125 (N_19125,N_16108,N_16115);
nand U19126 (N_19126,N_17182,N_16312);
or U19127 (N_19127,N_16948,N_15673);
or U19128 (N_19128,N_16218,N_15292);
nand U19129 (N_19129,N_16110,N_16918);
or U19130 (N_19130,N_15545,N_17114);
nand U19131 (N_19131,N_15561,N_17181);
nor U19132 (N_19132,N_16799,N_16898);
and U19133 (N_19133,N_17118,N_17131);
or U19134 (N_19134,N_16658,N_16370);
nor U19135 (N_19135,N_15161,N_16754);
nand U19136 (N_19136,N_16634,N_17236);
xor U19137 (N_19137,N_15721,N_17381);
and U19138 (N_19138,N_15741,N_15767);
xor U19139 (N_19139,N_16466,N_16819);
and U19140 (N_19140,N_15352,N_15422);
or U19141 (N_19141,N_15496,N_15823);
nor U19142 (N_19142,N_16688,N_15454);
nand U19143 (N_19143,N_15215,N_16798);
and U19144 (N_19144,N_16219,N_16648);
nand U19145 (N_19145,N_16595,N_15711);
xor U19146 (N_19146,N_15249,N_15935);
nand U19147 (N_19147,N_16722,N_16741);
nand U19148 (N_19148,N_15697,N_16480);
nor U19149 (N_19149,N_16151,N_15911);
xnor U19150 (N_19150,N_15845,N_15347);
xor U19151 (N_19151,N_15619,N_16834);
nor U19152 (N_19152,N_15828,N_16435);
xnor U19153 (N_19153,N_16766,N_16713);
xor U19154 (N_19154,N_17059,N_15348);
or U19155 (N_19155,N_15610,N_17043);
nand U19156 (N_19156,N_17202,N_15074);
nor U19157 (N_19157,N_15921,N_15287);
and U19158 (N_19158,N_17015,N_17252);
or U19159 (N_19159,N_15885,N_17160);
and U19160 (N_19160,N_15838,N_15755);
nor U19161 (N_19161,N_16051,N_16513);
nand U19162 (N_19162,N_16876,N_15584);
nor U19163 (N_19163,N_15304,N_17057);
and U19164 (N_19164,N_17447,N_17385);
nand U19165 (N_19165,N_15502,N_17097);
xor U19166 (N_19166,N_16691,N_15908);
nor U19167 (N_19167,N_17452,N_15552);
xnor U19168 (N_19168,N_17049,N_15291);
and U19169 (N_19169,N_15852,N_17255);
nor U19170 (N_19170,N_17082,N_17194);
nor U19171 (N_19171,N_17404,N_16361);
and U19172 (N_19172,N_16989,N_17172);
and U19173 (N_19173,N_17104,N_17154);
xor U19174 (N_19174,N_17344,N_16883);
xor U19175 (N_19175,N_15038,N_16320);
and U19176 (N_19176,N_16196,N_16694);
or U19177 (N_19177,N_17282,N_15101);
or U19178 (N_19178,N_16779,N_16063);
xor U19179 (N_19179,N_15079,N_15130);
and U19180 (N_19180,N_15968,N_16756);
nor U19181 (N_19181,N_15147,N_16901);
xor U19182 (N_19182,N_17149,N_17090);
and U19183 (N_19183,N_16642,N_16657);
nor U19184 (N_19184,N_17328,N_15754);
nor U19185 (N_19185,N_16826,N_16685);
xnor U19186 (N_19186,N_15704,N_17044);
xnor U19187 (N_19187,N_17412,N_15359);
or U19188 (N_19188,N_16207,N_15450);
and U19189 (N_19189,N_16092,N_15741);
nand U19190 (N_19190,N_16505,N_16837);
and U19191 (N_19191,N_16921,N_15369);
and U19192 (N_19192,N_15421,N_16807);
nand U19193 (N_19193,N_16866,N_15152);
or U19194 (N_19194,N_16443,N_16709);
and U19195 (N_19195,N_16330,N_16115);
nand U19196 (N_19196,N_16886,N_15632);
and U19197 (N_19197,N_17036,N_17206);
xnor U19198 (N_19198,N_17024,N_17418);
nor U19199 (N_19199,N_15678,N_17199);
and U19200 (N_19200,N_17049,N_16846);
nor U19201 (N_19201,N_17048,N_16525);
and U19202 (N_19202,N_17412,N_15981);
xnor U19203 (N_19203,N_16347,N_16769);
xnor U19204 (N_19204,N_15617,N_15641);
nand U19205 (N_19205,N_16860,N_16274);
xor U19206 (N_19206,N_16905,N_16020);
xor U19207 (N_19207,N_15554,N_15548);
or U19208 (N_19208,N_17371,N_15338);
or U19209 (N_19209,N_16318,N_17481);
nor U19210 (N_19210,N_15206,N_16535);
or U19211 (N_19211,N_17329,N_16269);
nor U19212 (N_19212,N_17289,N_17385);
nor U19213 (N_19213,N_17345,N_15627);
nor U19214 (N_19214,N_17125,N_16060);
xnor U19215 (N_19215,N_17422,N_16680);
and U19216 (N_19216,N_16399,N_15273);
or U19217 (N_19217,N_15431,N_16942);
or U19218 (N_19218,N_15803,N_15057);
or U19219 (N_19219,N_17215,N_16176);
nand U19220 (N_19220,N_16913,N_15564);
xor U19221 (N_19221,N_15415,N_17491);
and U19222 (N_19222,N_16040,N_15144);
and U19223 (N_19223,N_16576,N_15420);
nand U19224 (N_19224,N_16568,N_15461);
or U19225 (N_19225,N_16866,N_17327);
xnor U19226 (N_19226,N_15428,N_16615);
and U19227 (N_19227,N_16585,N_15219);
xor U19228 (N_19228,N_17205,N_15694);
nand U19229 (N_19229,N_15128,N_17163);
and U19230 (N_19230,N_15846,N_16410);
and U19231 (N_19231,N_15298,N_15398);
xor U19232 (N_19232,N_17013,N_17460);
nor U19233 (N_19233,N_17126,N_16756);
nand U19234 (N_19234,N_16175,N_16180);
or U19235 (N_19235,N_17148,N_15918);
nor U19236 (N_19236,N_15636,N_16868);
nand U19237 (N_19237,N_17282,N_15324);
xor U19238 (N_19238,N_17177,N_15766);
nand U19239 (N_19239,N_15181,N_15239);
and U19240 (N_19240,N_17296,N_17000);
nand U19241 (N_19241,N_15238,N_15026);
xnor U19242 (N_19242,N_16769,N_16524);
or U19243 (N_19243,N_17119,N_16852);
nor U19244 (N_19244,N_16951,N_17278);
xor U19245 (N_19245,N_17288,N_16073);
or U19246 (N_19246,N_17220,N_16932);
xnor U19247 (N_19247,N_15540,N_15360);
xor U19248 (N_19248,N_17402,N_16144);
nor U19249 (N_19249,N_16929,N_16239);
and U19250 (N_19250,N_15134,N_15769);
and U19251 (N_19251,N_16586,N_17023);
nand U19252 (N_19252,N_15520,N_17218);
nand U19253 (N_19253,N_15769,N_16016);
xor U19254 (N_19254,N_15298,N_16492);
and U19255 (N_19255,N_16087,N_15580);
xor U19256 (N_19256,N_16184,N_17480);
or U19257 (N_19257,N_16418,N_16035);
and U19258 (N_19258,N_16024,N_15891);
or U19259 (N_19259,N_16071,N_15639);
or U19260 (N_19260,N_17079,N_16276);
nand U19261 (N_19261,N_15958,N_15953);
nand U19262 (N_19262,N_15086,N_16975);
and U19263 (N_19263,N_15631,N_16420);
or U19264 (N_19264,N_15652,N_16592);
or U19265 (N_19265,N_15432,N_15721);
xnor U19266 (N_19266,N_17126,N_16449);
nand U19267 (N_19267,N_15194,N_16251);
nor U19268 (N_19268,N_16434,N_16183);
xor U19269 (N_19269,N_16802,N_17004);
xor U19270 (N_19270,N_16124,N_16300);
or U19271 (N_19271,N_17338,N_15680);
nand U19272 (N_19272,N_15942,N_16997);
and U19273 (N_19273,N_16185,N_15341);
nand U19274 (N_19274,N_16243,N_15072);
xnor U19275 (N_19275,N_15493,N_16579);
or U19276 (N_19276,N_15551,N_16089);
xnor U19277 (N_19277,N_15014,N_16247);
xnor U19278 (N_19278,N_17246,N_16421);
or U19279 (N_19279,N_17034,N_15689);
and U19280 (N_19280,N_17265,N_15897);
xnor U19281 (N_19281,N_16858,N_17272);
nand U19282 (N_19282,N_17140,N_15054);
nor U19283 (N_19283,N_16503,N_15989);
nand U19284 (N_19284,N_17179,N_17379);
xor U19285 (N_19285,N_16885,N_15892);
and U19286 (N_19286,N_15810,N_16358);
nand U19287 (N_19287,N_16545,N_16420);
or U19288 (N_19288,N_17072,N_16387);
and U19289 (N_19289,N_16441,N_16837);
and U19290 (N_19290,N_17235,N_17443);
or U19291 (N_19291,N_16973,N_16716);
and U19292 (N_19292,N_17375,N_17218);
or U19293 (N_19293,N_16197,N_16140);
nor U19294 (N_19294,N_16265,N_16713);
nor U19295 (N_19295,N_17041,N_15113);
or U19296 (N_19296,N_16137,N_17342);
or U19297 (N_19297,N_15069,N_17325);
or U19298 (N_19298,N_16742,N_17036);
nand U19299 (N_19299,N_17498,N_17413);
nor U19300 (N_19300,N_16990,N_15881);
xor U19301 (N_19301,N_15061,N_15098);
and U19302 (N_19302,N_17405,N_15644);
nor U19303 (N_19303,N_16833,N_15198);
or U19304 (N_19304,N_17357,N_15734);
nor U19305 (N_19305,N_16536,N_17205);
or U19306 (N_19306,N_15638,N_15327);
or U19307 (N_19307,N_17065,N_17332);
and U19308 (N_19308,N_17139,N_16163);
xnor U19309 (N_19309,N_15540,N_16333);
nand U19310 (N_19310,N_15266,N_17179);
xnor U19311 (N_19311,N_15487,N_17471);
and U19312 (N_19312,N_17412,N_15086);
nand U19313 (N_19313,N_16269,N_15847);
nor U19314 (N_19314,N_15752,N_15766);
nor U19315 (N_19315,N_15845,N_16581);
nor U19316 (N_19316,N_16830,N_15659);
nor U19317 (N_19317,N_16522,N_17108);
nor U19318 (N_19318,N_15551,N_17138);
nor U19319 (N_19319,N_17327,N_16177);
xor U19320 (N_19320,N_15775,N_17106);
xnor U19321 (N_19321,N_16971,N_16315);
or U19322 (N_19322,N_16330,N_15498);
xnor U19323 (N_19323,N_15548,N_17311);
and U19324 (N_19324,N_16543,N_17116);
and U19325 (N_19325,N_17140,N_15083);
xnor U19326 (N_19326,N_15002,N_16677);
nand U19327 (N_19327,N_15140,N_16265);
nand U19328 (N_19328,N_17289,N_17252);
or U19329 (N_19329,N_17397,N_15680);
xnor U19330 (N_19330,N_17346,N_15642);
and U19331 (N_19331,N_16612,N_16052);
xor U19332 (N_19332,N_15001,N_15434);
nand U19333 (N_19333,N_15819,N_17478);
nor U19334 (N_19334,N_17319,N_17088);
xnor U19335 (N_19335,N_16206,N_15978);
or U19336 (N_19336,N_15653,N_15981);
and U19337 (N_19337,N_15080,N_17307);
nand U19338 (N_19338,N_17309,N_15492);
and U19339 (N_19339,N_16673,N_16004);
or U19340 (N_19340,N_16339,N_16983);
xor U19341 (N_19341,N_17372,N_15149);
nor U19342 (N_19342,N_16359,N_16350);
xnor U19343 (N_19343,N_15771,N_17043);
nand U19344 (N_19344,N_16763,N_15877);
or U19345 (N_19345,N_16979,N_17343);
nand U19346 (N_19346,N_16149,N_16048);
or U19347 (N_19347,N_16188,N_15824);
nor U19348 (N_19348,N_17307,N_17372);
and U19349 (N_19349,N_15755,N_16269);
nor U19350 (N_19350,N_15578,N_16536);
nand U19351 (N_19351,N_16797,N_17167);
nor U19352 (N_19352,N_15644,N_15587);
nand U19353 (N_19353,N_16691,N_15494);
nor U19354 (N_19354,N_16077,N_16501);
or U19355 (N_19355,N_15479,N_15833);
xor U19356 (N_19356,N_15210,N_16444);
nor U19357 (N_19357,N_16282,N_15622);
xor U19358 (N_19358,N_15233,N_15677);
and U19359 (N_19359,N_15312,N_17414);
xnor U19360 (N_19360,N_16425,N_16653);
nor U19361 (N_19361,N_17242,N_17057);
and U19362 (N_19362,N_16430,N_17051);
xor U19363 (N_19363,N_15161,N_17177);
nor U19364 (N_19364,N_15070,N_17097);
and U19365 (N_19365,N_15681,N_16186);
nor U19366 (N_19366,N_17285,N_16807);
nor U19367 (N_19367,N_17444,N_17187);
nor U19368 (N_19368,N_16839,N_15173);
nand U19369 (N_19369,N_15821,N_15934);
nor U19370 (N_19370,N_16650,N_16964);
xnor U19371 (N_19371,N_15567,N_16282);
and U19372 (N_19372,N_15793,N_17081);
or U19373 (N_19373,N_17178,N_16196);
xnor U19374 (N_19374,N_16178,N_17206);
or U19375 (N_19375,N_15523,N_15568);
or U19376 (N_19376,N_16901,N_16875);
or U19377 (N_19377,N_16157,N_15457);
nand U19378 (N_19378,N_16716,N_17340);
and U19379 (N_19379,N_16284,N_15732);
xor U19380 (N_19380,N_16400,N_16194);
nor U19381 (N_19381,N_15938,N_16445);
xor U19382 (N_19382,N_15611,N_15117);
and U19383 (N_19383,N_16701,N_16429);
or U19384 (N_19384,N_15721,N_16718);
or U19385 (N_19385,N_17313,N_17486);
nand U19386 (N_19386,N_15886,N_15709);
and U19387 (N_19387,N_15987,N_16086);
nand U19388 (N_19388,N_17166,N_15973);
or U19389 (N_19389,N_15312,N_15837);
nand U19390 (N_19390,N_15684,N_16313);
nand U19391 (N_19391,N_16072,N_15048);
xnor U19392 (N_19392,N_16075,N_15655);
and U19393 (N_19393,N_15944,N_15027);
nor U19394 (N_19394,N_15258,N_16651);
nand U19395 (N_19395,N_15669,N_17170);
and U19396 (N_19396,N_15621,N_15052);
nand U19397 (N_19397,N_16777,N_17136);
nand U19398 (N_19398,N_15621,N_15253);
or U19399 (N_19399,N_15541,N_16349);
nand U19400 (N_19400,N_15951,N_15417);
nor U19401 (N_19401,N_15156,N_15297);
and U19402 (N_19402,N_16059,N_16149);
xor U19403 (N_19403,N_16594,N_15418);
and U19404 (N_19404,N_16977,N_16813);
or U19405 (N_19405,N_15371,N_17462);
nor U19406 (N_19406,N_15565,N_15169);
and U19407 (N_19407,N_15640,N_16569);
nor U19408 (N_19408,N_17235,N_16958);
or U19409 (N_19409,N_15383,N_15507);
nand U19410 (N_19410,N_17217,N_15591);
nor U19411 (N_19411,N_16561,N_16281);
nor U19412 (N_19412,N_17417,N_17305);
or U19413 (N_19413,N_15565,N_16978);
and U19414 (N_19414,N_16940,N_16995);
nand U19415 (N_19415,N_15648,N_16338);
nand U19416 (N_19416,N_15233,N_15054);
xnor U19417 (N_19417,N_16810,N_16194);
nand U19418 (N_19418,N_16723,N_17298);
xnor U19419 (N_19419,N_17411,N_16468);
and U19420 (N_19420,N_16938,N_17015);
nand U19421 (N_19421,N_16461,N_15567);
and U19422 (N_19422,N_15186,N_15230);
nand U19423 (N_19423,N_15615,N_15619);
nand U19424 (N_19424,N_15204,N_16169);
or U19425 (N_19425,N_16140,N_15410);
and U19426 (N_19426,N_16836,N_15070);
nor U19427 (N_19427,N_16755,N_17232);
xor U19428 (N_19428,N_17171,N_17274);
and U19429 (N_19429,N_16734,N_15778);
xor U19430 (N_19430,N_15278,N_16336);
xnor U19431 (N_19431,N_17180,N_15141);
xnor U19432 (N_19432,N_16197,N_15819);
xor U19433 (N_19433,N_15078,N_15755);
and U19434 (N_19434,N_15776,N_15628);
and U19435 (N_19435,N_17036,N_16898);
and U19436 (N_19436,N_16836,N_16949);
and U19437 (N_19437,N_15263,N_16003);
nor U19438 (N_19438,N_15039,N_17419);
xnor U19439 (N_19439,N_17301,N_16287);
nor U19440 (N_19440,N_16472,N_15683);
xor U19441 (N_19441,N_16234,N_17167);
nor U19442 (N_19442,N_15964,N_15185);
and U19443 (N_19443,N_15378,N_16378);
or U19444 (N_19444,N_17440,N_17225);
nand U19445 (N_19445,N_16171,N_15509);
nor U19446 (N_19446,N_16977,N_16552);
and U19447 (N_19447,N_15757,N_17183);
and U19448 (N_19448,N_16864,N_16919);
nor U19449 (N_19449,N_15819,N_16773);
xor U19450 (N_19450,N_17146,N_17227);
or U19451 (N_19451,N_15005,N_16265);
xor U19452 (N_19452,N_15792,N_16263);
nor U19453 (N_19453,N_16499,N_16406);
nand U19454 (N_19454,N_15231,N_17489);
nand U19455 (N_19455,N_16893,N_16024);
and U19456 (N_19456,N_15868,N_15748);
and U19457 (N_19457,N_17336,N_15352);
or U19458 (N_19458,N_17435,N_15104);
or U19459 (N_19459,N_15958,N_17370);
and U19460 (N_19460,N_16071,N_15392);
nor U19461 (N_19461,N_16808,N_17051);
nand U19462 (N_19462,N_17153,N_15633);
xor U19463 (N_19463,N_15747,N_16469);
nor U19464 (N_19464,N_16990,N_15266);
nand U19465 (N_19465,N_15127,N_15803);
nor U19466 (N_19466,N_17126,N_15310);
nand U19467 (N_19467,N_15889,N_15494);
nor U19468 (N_19468,N_15304,N_16316);
nor U19469 (N_19469,N_17387,N_15014);
or U19470 (N_19470,N_17037,N_16555);
xnor U19471 (N_19471,N_16322,N_16469);
or U19472 (N_19472,N_15683,N_17167);
or U19473 (N_19473,N_15476,N_16845);
xor U19474 (N_19474,N_16559,N_16353);
and U19475 (N_19475,N_15185,N_16249);
xnor U19476 (N_19476,N_15530,N_15207);
nand U19477 (N_19477,N_16894,N_16033);
and U19478 (N_19478,N_15611,N_16484);
and U19479 (N_19479,N_15287,N_15657);
xnor U19480 (N_19480,N_16842,N_15889);
nor U19481 (N_19481,N_15006,N_17422);
or U19482 (N_19482,N_16482,N_17205);
nand U19483 (N_19483,N_15967,N_16110);
nor U19484 (N_19484,N_16145,N_15633);
or U19485 (N_19485,N_17021,N_16491);
and U19486 (N_19486,N_15377,N_16559);
nor U19487 (N_19487,N_15182,N_16448);
nand U19488 (N_19488,N_16620,N_15526);
nor U19489 (N_19489,N_15795,N_15445);
and U19490 (N_19490,N_15598,N_15118);
xnor U19491 (N_19491,N_16096,N_16918);
nand U19492 (N_19492,N_15182,N_16292);
nor U19493 (N_19493,N_15967,N_15106);
xnor U19494 (N_19494,N_15913,N_16436);
nor U19495 (N_19495,N_16906,N_16585);
and U19496 (N_19496,N_16691,N_16091);
nand U19497 (N_19497,N_15483,N_16300);
xor U19498 (N_19498,N_16933,N_16410);
nand U19499 (N_19499,N_16907,N_16646);
and U19500 (N_19500,N_15547,N_16647);
nor U19501 (N_19501,N_17349,N_17298);
nor U19502 (N_19502,N_16755,N_16426);
nor U19503 (N_19503,N_15114,N_16172);
xor U19504 (N_19504,N_15739,N_15029);
or U19505 (N_19505,N_16562,N_17353);
nand U19506 (N_19506,N_17124,N_16249);
or U19507 (N_19507,N_16150,N_16262);
xor U19508 (N_19508,N_15142,N_16687);
nor U19509 (N_19509,N_15817,N_17107);
or U19510 (N_19510,N_15033,N_17360);
xnor U19511 (N_19511,N_15543,N_17341);
xnor U19512 (N_19512,N_15666,N_15585);
nor U19513 (N_19513,N_16614,N_16831);
and U19514 (N_19514,N_15406,N_15941);
nor U19515 (N_19515,N_17216,N_16685);
xnor U19516 (N_19516,N_16268,N_16967);
xor U19517 (N_19517,N_16411,N_15678);
nand U19518 (N_19518,N_17094,N_15406);
or U19519 (N_19519,N_16364,N_16402);
xor U19520 (N_19520,N_15426,N_17374);
xnor U19521 (N_19521,N_16807,N_15233);
nor U19522 (N_19522,N_16375,N_16446);
xnor U19523 (N_19523,N_16296,N_16278);
nand U19524 (N_19524,N_15026,N_15162);
nor U19525 (N_19525,N_15755,N_17012);
or U19526 (N_19526,N_16693,N_16014);
and U19527 (N_19527,N_15621,N_15870);
nand U19528 (N_19528,N_16690,N_15550);
or U19529 (N_19529,N_15707,N_16519);
or U19530 (N_19530,N_15803,N_16021);
xor U19531 (N_19531,N_15870,N_15290);
and U19532 (N_19532,N_16848,N_15656);
and U19533 (N_19533,N_16288,N_16439);
or U19534 (N_19534,N_16605,N_16475);
and U19535 (N_19535,N_15786,N_16954);
nor U19536 (N_19536,N_16677,N_16338);
nor U19537 (N_19537,N_17211,N_16560);
or U19538 (N_19538,N_16807,N_15746);
xnor U19539 (N_19539,N_15878,N_16935);
nor U19540 (N_19540,N_15084,N_16512);
or U19541 (N_19541,N_15527,N_15354);
or U19542 (N_19542,N_15379,N_15796);
xnor U19543 (N_19543,N_16344,N_16515);
and U19544 (N_19544,N_15098,N_16919);
xor U19545 (N_19545,N_17068,N_16590);
or U19546 (N_19546,N_17397,N_16751);
nor U19547 (N_19547,N_15974,N_16170);
and U19548 (N_19548,N_16536,N_16658);
nand U19549 (N_19549,N_16823,N_15970);
or U19550 (N_19550,N_16522,N_16093);
nor U19551 (N_19551,N_15780,N_16922);
and U19552 (N_19552,N_17003,N_15196);
or U19553 (N_19553,N_15050,N_15250);
xnor U19554 (N_19554,N_16782,N_16837);
xor U19555 (N_19555,N_16422,N_16401);
xor U19556 (N_19556,N_17312,N_15809);
or U19557 (N_19557,N_15184,N_17230);
nor U19558 (N_19558,N_17468,N_15620);
or U19559 (N_19559,N_15765,N_17063);
or U19560 (N_19560,N_15909,N_16201);
xnor U19561 (N_19561,N_17145,N_15644);
nand U19562 (N_19562,N_16079,N_16064);
nand U19563 (N_19563,N_16326,N_15964);
nor U19564 (N_19564,N_17477,N_15514);
or U19565 (N_19565,N_15972,N_16382);
nor U19566 (N_19566,N_15221,N_15301);
xnor U19567 (N_19567,N_16937,N_16212);
nand U19568 (N_19568,N_17408,N_15579);
nor U19569 (N_19569,N_15509,N_15405);
or U19570 (N_19570,N_17079,N_17236);
or U19571 (N_19571,N_16751,N_16898);
and U19572 (N_19572,N_16970,N_15256);
nor U19573 (N_19573,N_17028,N_15264);
nor U19574 (N_19574,N_15554,N_15494);
or U19575 (N_19575,N_15973,N_15791);
or U19576 (N_19576,N_15664,N_15838);
and U19577 (N_19577,N_16608,N_15188);
and U19578 (N_19578,N_15591,N_16661);
and U19579 (N_19579,N_15856,N_15615);
nor U19580 (N_19580,N_16450,N_16128);
xnor U19581 (N_19581,N_15870,N_15841);
and U19582 (N_19582,N_16121,N_15211);
or U19583 (N_19583,N_17001,N_16321);
and U19584 (N_19584,N_15233,N_17088);
nand U19585 (N_19585,N_15262,N_17486);
nand U19586 (N_19586,N_16878,N_16119);
nor U19587 (N_19587,N_15653,N_16879);
nand U19588 (N_19588,N_15365,N_16639);
or U19589 (N_19589,N_17026,N_16581);
and U19590 (N_19590,N_16662,N_15700);
or U19591 (N_19591,N_17210,N_15457);
and U19592 (N_19592,N_15982,N_15050);
xor U19593 (N_19593,N_15703,N_16795);
xnor U19594 (N_19594,N_16852,N_15539);
nor U19595 (N_19595,N_16695,N_16541);
and U19596 (N_19596,N_15137,N_15983);
xnor U19597 (N_19597,N_16504,N_16828);
or U19598 (N_19598,N_16902,N_15255);
nand U19599 (N_19599,N_17233,N_16394);
nand U19600 (N_19600,N_16779,N_16079);
or U19601 (N_19601,N_15508,N_16559);
xor U19602 (N_19602,N_15970,N_17383);
nand U19603 (N_19603,N_15869,N_15785);
or U19604 (N_19604,N_17289,N_16700);
or U19605 (N_19605,N_15911,N_17069);
and U19606 (N_19606,N_17336,N_17257);
nor U19607 (N_19607,N_15920,N_16070);
nor U19608 (N_19608,N_17019,N_15698);
nor U19609 (N_19609,N_15116,N_15660);
or U19610 (N_19610,N_15300,N_15699);
nor U19611 (N_19611,N_15699,N_16252);
and U19612 (N_19612,N_16780,N_16644);
xor U19613 (N_19613,N_16954,N_17317);
xor U19614 (N_19614,N_16385,N_17214);
nand U19615 (N_19615,N_16301,N_16531);
and U19616 (N_19616,N_17131,N_16139);
xor U19617 (N_19617,N_15673,N_16716);
and U19618 (N_19618,N_15580,N_15526);
nor U19619 (N_19619,N_16906,N_15323);
nor U19620 (N_19620,N_15647,N_17005);
nand U19621 (N_19621,N_15222,N_16263);
and U19622 (N_19622,N_16132,N_15707);
and U19623 (N_19623,N_16449,N_17066);
nand U19624 (N_19624,N_16930,N_17331);
or U19625 (N_19625,N_16447,N_15851);
nor U19626 (N_19626,N_16192,N_15909);
nand U19627 (N_19627,N_15958,N_15076);
nand U19628 (N_19628,N_15140,N_15940);
and U19629 (N_19629,N_16020,N_16042);
xnor U19630 (N_19630,N_15333,N_16942);
xnor U19631 (N_19631,N_16170,N_16765);
or U19632 (N_19632,N_16932,N_16899);
nor U19633 (N_19633,N_17196,N_16981);
and U19634 (N_19634,N_15087,N_15357);
nor U19635 (N_19635,N_15516,N_17127);
xnor U19636 (N_19636,N_16776,N_15907);
xnor U19637 (N_19637,N_16523,N_17204);
or U19638 (N_19638,N_17263,N_16613);
xor U19639 (N_19639,N_16692,N_16068);
xor U19640 (N_19640,N_15498,N_16662);
nand U19641 (N_19641,N_15861,N_16480);
or U19642 (N_19642,N_16747,N_15819);
nor U19643 (N_19643,N_17487,N_16436);
nand U19644 (N_19644,N_15405,N_16405);
or U19645 (N_19645,N_16536,N_17036);
nand U19646 (N_19646,N_15038,N_17412);
xnor U19647 (N_19647,N_15943,N_15503);
nand U19648 (N_19648,N_15738,N_15617);
and U19649 (N_19649,N_16805,N_15736);
or U19650 (N_19650,N_15605,N_16783);
nor U19651 (N_19651,N_17179,N_16797);
or U19652 (N_19652,N_16116,N_16266);
nor U19653 (N_19653,N_15048,N_16156);
or U19654 (N_19654,N_15053,N_17278);
xor U19655 (N_19655,N_15559,N_15442);
or U19656 (N_19656,N_17011,N_17087);
and U19657 (N_19657,N_17088,N_16315);
nor U19658 (N_19658,N_15464,N_15229);
nor U19659 (N_19659,N_15881,N_16618);
or U19660 (N_19660,N_15204,N_15369);
xor U19661 (N_19661,N_16263,N_16220);
and U19662 (N_19662,N_15252,N_16456);
or U19663 (N_19663,N_17395,N_15601);
nand U19664 (N_19664,N_16363,N_16022);
nor U19665 (N_19665,N_16496,N_16414);
and U19666 (N_19666,N_17365,N_16899);
nand U19667 (N_19667,N_17380,N_15460);
nor U19668 (N_19668,N_15529,N_17303);
nor U19669 (N_19669,N_17313,N_15784);
xnor U19670 (N_19670,N_17031,N_15355);
nor U19671 (N_19671,N_16057,N_15773);
or U19672 (N_19672,N_15838,N_16403);
and U19673 (N_19673,N_15148,N_15651);
nand U19674 (N_19674,N_15157,N_15744);
xnor U19675 (N_19675,N_16731,N_16137);
xor U19676 (N_19676,N_16090,N_15989);
nand U19677 (N_19677,N_16277,N_17058);
nor U19678 (N_19678,N_16728,N_17444);
xnor U19679 (N_19679,N_15784,N_16031);
xnor U19680 (N_19680,N_16854,N_15522);
and U19681 (N_19681,N_15033,N_17115);
or U19682 (N_19682,N_15184,N_17161);
or U19683 (N_19683,N_17165,N_15506);
or U19684 (N_19684,N_15535,N_17088);
nand U19685 (N_19685,N_16491,N_16100);
nand U19686 (N_19686,N_16685,N_17337);
nor U19687 (N_19687,N_17398,N_16512);
nand U19688 (N_19688,N_15945,N_15772);
nand U19689 (N_19689,N_16006,N_15783);
nand U19690 (N_19690,N_15172,N_16911);
and U19691 (N_19691,N_16405,N_16812);
xor U19692 (N_19692,N_16836,N_16776);
or U19693 (N_19693,N_15486,N_15954);
or U19694 (N_19694,N_15416,N_16366);
nand U19695 (N_19695,N_17146,N_15542);
xor U19696 (N_19696,N_16230,N_15249);
nand U19697 (N_19697,N_16969,N_15309);
and U19698 (N_19698,N_17340,N_15974);
nand U19699 (N_19699,N_16717,N_15537);
nor U19700 (N_19700,N_15479,N_16234);
nand U19701 (N_19701,N_16132,N_15521);
nand U19702 (N_19702,N_16124,N_15778);
and U19703 (N_19703,N_16581,N_15452);
or U19704 (N_19704,N_15654,N_17318);
nand U19705 (N_19705,N_15306,N_16564);
nand U19706 (N_19706,N_17444,N_16024);
nand U19707 (N_19707,N_16470,N_15756);
or U19708 (N_19708,N_15213,N_16096);
xor U19709 (N_19709,N_15908,N_15967);
and U19710 (N_19710,N_16973,N_15920);
xnor U19711 (N_19711,N_17135,N_17009);
and U19712 (N_19712,N_17062,N_16385);
or U19713 (N_19713,N_17006,N_16708);
and U19714 (N_19714,N_15928,N_16544);
nor U19715 (N_19715,N_15374,N_16436);
nand U19716 (N_19716,N_16009,N_15906);
xor U19717 (N_19717,N_17093,N_15173);
xor U19718 (N_19718,N_15576,N_15551);
and U19719 (N_19719,N_16237,N_16503);
and U19720 (N_19720,N_16956,N_16460);
nand U19721 (N_19721,N_15081,N_16858);
xor U19722 (N_19722,N_16402,N_15555);
nand U19723 (N_19723,N_15207,N_17167);
or U19724 (N_19724,N_15543,N_15809);
and U19725 (N_19725,N_15804,N_15150);
nor U19726 (N_19726,N_16099,N_15661);
xor U19727 (N_19727,N_15096,N_16942);
nand U19728 (N_19728,N_16317,N_16829);
and U19729 (N_19729,N_15320,N_17128);
and U19730 (N_19730,N_16152,N_15746);
and U19731 (N_19731,N_16495,N_15722);
or U19732 (N_19732,N_15175,N_16030);
and U19733 (N_19733,N_15628,N_16716);
or U19734 (N_19734,N_16297,N_17312);
nand U19735 (N_19735,N_15372,N_16297);
nor U19736 (N_19736,N_16443,N_16618);
or U19737 (N_19737,N_15010,N_17179);
or U19738 (N_19738,N_16643,N_17074);
xor U19739 (N_19739,N_17302,N_16406);
xor U19740 (N_19740,N_15864,N_15818);
or U19741 (N_19741,N_15621,N_16536);
and U19742 (N_19742,N_17265,N_17314);
xnor U19743 (N_19743,N_15816,N_15694);
and U19744 (N_19744,N_16104,N_15226);
or U19745 (N_19745,N_15845,N_15373);
nor U19746 (N_19746,N_15291,N_16525);
nor U19747 (N_19747,N_17392,N_16310);
or U19748 (N_19748,N_15542,N_16121);
and U19749 (N_19749,N_15315,N_17225);
xnor U19750 (N_19750,N_15492,N_16123);
nand U19751 (N_19751,N_17411,N_16039);
nor U19752 (N_19752,N_15939,N_15012);
nand U19753 (N_19753,N_17007,N_16889);
xnor U19754 (N_19754,N_16645,N_16869);
nor U19755 (N_19755,N_16180,N_16027);
nor U19756 (N_19756,N_16559,N_15304);
nand U19757 (N_19757,N_15978,N_16091);
and U19758 (N_19758,N_17304,N_16459);
nor U19759 (N_19759,N_16216,N_16934);
nor U19760 (N_19760,N_17388,N_17262);
or U19761 (N_19761,N_16617,N_15138);
nand U19762 (N_19762,N_16268,N_15098);
and U19763 (N_19763,N_16586,N_15154);
nor U19764 (N_19764,N_17309,N_15598);
nor U19765 (N_19765,N_16214,N_16578);
xor U19766 (N_19766,N_16963,N_17297);
xnor U19767 (N_19767,N_17253,N_17277);
nand U19768 (N_19768,N_15603,N_16114);
or U19769 (N_19769,N_16041,N_17193);
and U19770 (N_19770,N_16042,N_16586);
and U19771 (N_19771,N_17090,N_15058);
nor U19772 (N_19772,N_15209,N_17403);
nor U19773 (N_19773,N_16302,N_16086);
nand U19774 (N_19774,N_16213,N_15296);
nor U19775 (N_19775,N_17030,N_17254);
and U19776 (N_19776,N_15024,N_16132);
xnor U19777 (N_19777,N_17278,N_15103);
or U19778 (N_19778,N_17068,N_17383);
nor U19779 (N_19779,N_16806,N_17082);
xnor U19780 (N_19780,N_17247,N_17170);
xor U19781 (N_19781,N_15106,N_17184);
nor U19782 (N_19782,N_15665,N_15459);
nor U19783 (N_19783,N_16053,N_16489);
and U19784 (N_19784,N_15281,N_17055);
and U19785 (N_19785,N_15875,N_15817);
nor U19786 (N_19786,N_16305,N_16884);
nor U19787 (N_19787,N_15669,N_17169);
nand U19788 (N_19788,N_16863,N_16321);
xnor U19789 (N_19789,N_16316,N_17200);
xnor U19790 (N_19790,N_16334,N_17462);
or U19791 (N_19791,N_16811,N_15667);
or U19792 (N_19792,N_15891,N_16282);
or U19793 (N_19793,N_16497,N_17343);
and U19794 (N_19794,N_16883,N_16480);
and U19795 (N_19795,N_17390,N_16658);
or U19796 (N_19796,N_17097,N_17395);
and U19797 (N_19797,N_15062,N_15564);
nor U19798 (N_19798,N_15841,N_15328);
and U19799 (N_19799,N_15093,N_16630);
xor U19800 (N_19800,N_15716,N_15588);
or U19801 (N_19801,N_16928,N_15497);
nand U19802 (N_19802,N_16669,N_15902);
and U19803 (N_19803,N_16939,N_16958);
or U19804 (N_19804,N_16130,N_15281);
nand U19805 (N_19805,N_15798,N_15825);
and U19806 (N_19806,N_15150,N_17394);
nand U19807 (N_19807,N_15756,N_16437);
or U19808 (N_19808,N_17135,N_15698);
and U19809 (N_19809,N_15860,N_15918);
nor U19810 (N_19810,N_15305,N_15531);
nor U19811 (N_19811,N_15141,N_15823);
nor U19812 (N_19812,N_15918,N_16953);
nor U19813 (N_19813,N_17124,N_15920);
xnor U19814 (N_19814,N_15426,N_16607);
nand U19815 (N_19815,N_16012,N_16693);
or U19816 (N_19816,N_15153,N_16963);
nand U19817 (N_19817,N_15954,N_16780);
and U19818 (N_19818,N_17148,N_15829);
and U19819 (N_19819,N_15054,N_16324);
nor U19820 (N_19820,N_15027,N_15491);
and U19821 (N_19821,N_16560,N_17065);
xor U19822 (N_19822,N_15758,N_17184);
nor U19823 (N_19823,N_15217,N_17179);
nand U19824 (N_19824,N_16888,N_16923);
and U19825 (N_19825,N_17443,N_16604);
xor U19826 (N_19826,N_17232,N_16354);
xor U19827 (N_19827,N_17002,N_15424);
nand U19828 (N_19828,N_16228,N_17150);
nand U19829 (N_19829,N_15322,N_15056);
or U19830 (N_19830,N_15539,N_15564);
xor U19831 (N_19831,N_16099,N_17047);
nand U19832 (N_19832,N_15095,N_17318);
and U19833 (N_19833,N_17122,N_16658);
or U19834 (N_19834,N_15321,N_16661);
nand U19835 (N_19835,N_16302,N_15113);
xor U19836 (N_19836,N_15445,N_16775);
nor U19837 (N_19837,N_16146,N_15039);
and U19838 (N_19838,N_17398,N_16291);
or U19839 (N_19839,N_17284,N_17472);
nor U19840 (N_19840,N_16385,N_15898);
xnor U19841 (N_19841,N_16876,N_16050);
or U19842 (N_19842,N_15612,N_16396);
and U19843 (N_19843,N_16507,N_16805);
xor U19844 (N_19844,N_15311,N_15108);
nor U19845 (N_19845,N_16810,N_16149);
or U19846 (N_19846,N_15103,N_16668);
xor U19847 (N_19847,N_16027,N_15310);
nor U19848 (N_19848,N_15865,N_15034);
nand U19849 (N_19849,N_16418,N_15726);
xor U19850 (N_19850,N_16289,N_16202);
xnor U19851 (N_19851,N_17490,N_16741);
or U19852 (N_19852,N_15525,N_15573);
or U19853 (N_19853,N_17119,N_16606);
nand U19854 (N_19854,N_15980,N_16467);
nor U19855 (N_19855,N_15288,N_16597);
and U19856 (N_19856,N_17176,N_16473);
and U19857 (N_19857,N_16605,N_16192);
nor U19858 (N_19858,N_16128,N_16635);
or U19859 (N_19859,N_17147,N_15146);
nor U19860 (N_19860,N_17231,N_16867);
xor U19861 (N_19861,N_16649,N_15920);
nand U19862 (N_19862,N_17028,N_16042);
and U19863 (N_19863,N_17462,N_17128);
and U19864 (N_19864,N_16672,N_16093);
or U19865 (N_19865,N_16685,N_15700);
xnor U19866 (N_19866,N_15834,N_15434);
or U19867 (N_19867,N_15349,N_16842);
nor U19868 (N_19868,N_16682,N_16401);
nor U19869 (N_19869,N_15602,N_15848);
nand U19870 (N_19870,N_16355,N_16678);
nand U19871 (N_19871,N_16228,N_17304);
xor U19872 (N_19872,N_16463,N_17040);
and U19873 (N_19873,N_15690,N_16483);
or U19874 (N_19874,N_16233,N_17038);
xor U19875 (N_19875,N_17405,N_15134);
and U19876 (N_19876,N_16108,N_16859);
xnor U19877 (N_19877,N_15114,N_16851);
xnor U19878 (N_19878,N_15216,N_16662);
or U19879 (N_19879,N_16235,N_16853);
nand U19880 (N_19880,N_17214,N_15111);
or U19881 (N_19881,N_15373,N_15484);
nor U19882 (N_19882,N_16038,N_15744);
and U19883 (N_19883,N_17046,N_16918);
or U19884 (N_19884,N_15145,N_15925);
and U19885 (N_19885,N_16882,N_17199);
nor U19886 (N_19886,N_16895,N_17316);
nand U19887 (N_19887,N_16870,N_16169);
nand U19888 (N_19888,N_17376,N_15628);
nand U19889 (N_19889,N_15908,N_17199);
nor U19890 (N_19890,N_16938,N_16373);
nor U19891 (N_19891,N_15871,N_16796);
or U19892 (N_19892,N_16615,N_17117);
and U19893 (N_19893,N_15408,N_15753);
xor U19894 (N_19894,N_15741,N_15877);
and U19895 (N_19895,N_16465,N_16484);
nand U19896 (N_19896,N_16167,N_15501);
xnor U19897 (N_19897,N_15004,N_16335);
xor U19898 (N_19898,N_16520,N_17077);
nand U19899 (N_19899,N_17441,N_17190);
nor U19900 (N_19900,N_16328,N_16816);
nand U19901 (N_19901,N_15253,N_16236);
or U19902 (N_19902,N_15865,N_15636);
nor U19903 (N_19903,N_17121,N_16977);
xnor U19904 (N_19904,N_17485,N_17314);
and U19905 (N_19905,N_15666,N_17021);
nand U19906 (N_19906,N_15604,N_15198);
nand U19907 (N_19907,N_16162,N_16910);
or U19908 (N_19908,N_16552,N_16771);
and U19909 (N_19909,N_16666,N_15723);
and U19910 (N_19910,N_16530,N_16273);
and U19911 (N_19911,N_17263,N_15051);
nand U19912 (N_19912,N_15534,N_15207);
or U19913 (N_19913,N_16276,N_15060);
or U19914 (N_19914,N_15721,N_17435);
nand U19915 (N_19915,N_15011,N_15035);
and U19916 (N_19916,N_16914,N_15064);
xor U19917 (N_19917,N_17052,N_15878);
xor U19918 (N_19918,N_15838,N_15236);
or U19919 (N_19919,N_17200,N_16718);
or U19920 (N_19920,N_17490,N_15775);
xnor U19921 (N_19921,N_17154,N_15352);
xor U19922 (N_19922,N_15993,N_15498);
nor U19923 (N_19923,N_15786,N_15872);
xor U19924 (N_19924,N_15965,N_15615);
nor U19925 (N_19925,N_15095,N_17422);
nor U19926 (N_19926,N_16593,N_15260);
nand U19927 (N_19927,N_16409,N_16983);
xnor U19928 (N_19928,N_16896,N_16904);
or U19929 (N_19929,N_16450,N_16060);
xnor U19930 (N_19930,N_16309,N_15109);
nand U19931 (N_19931,N_15247,N_15037);
xnor U19932 (N_19932,N_17083,N_15459);
nor U19933 (N_19933,N_16673,N_15612);
or U19934 (N_19934,N_17081,N_17041);
and U19935 (N_19935,N_17183,N_15543);
nand U19936 (N_19936,N_16779,N_15515);
nand U19937 (N_19937,N_17345,N_15231);
or U19938 (N_19938,N_15553,N_15567);
or U19939 (N_19939,N_17470,N_16205);
or U19940 (N_19940,N_15768,N_15279);
or U19941 (N_19941,N_16528,N_15024);
or U19942 (N_19942,N_16179,N_16564);
and U19943 (N_19943,N_17280,N_16753);
nand U19944 (N_19944,N_16209,N_17079);
nor U19945 (N_19945,N_16841,N_15978);
nor U19946 (N_19946,N_16403,N_15334);
xor U19947 (N_19947,N_17137,N_15037);
or U19948 (N_19948,N_17158,N_17054);
xor U19949 (N_19949,N_15984,N_15758);
and U19950 (N_19950,N_16321,N_16832);
xnor U19951 (N_19951,N_16181,N_16828);
nand U19952 (N_19952,N_17385,N_16913);
nand U19953 (N_19953,N_17145,N_15135);
and U19954 (N_19954,N_16578,N_15686);
and U19955 (N_19955,N_15378,N_15200);
nor U19956 (N_19956,N_16632,N_16715);
xnor U19957 (N_19957,N_17384,N_15844);
xnor U19958 (N_19958,N_15417,N_17062);
xnor U19959 (N_19959,N_17442,N_15750);
or U19960 (N_19960,N_16711,N_16584);
nor U19961 (N_19961,N_17302,N_16549);
nor U19962 (N_19962,N_17164,N_15398);
and U19963 (N_19963,N_15861,N_15659);
xnor U19964 (N_19964,N_16170,N_15600);
xor U19965 (N_19965,N_16318,N_16749);
or U19966 (N_19966,N_15305,N_15742);
nor U19967 (N_19967,N_15302,N_16416);
and U19968 (N_19968,N_15073,N_17438);
or U19969 (N_19969,N_16366,N_16346);
or U19970 (N_19970,N_17311,N_17273);
xor U19971 (N_19971,N_17496,N_16584);
and U19972 (N_19972,N_15793,N_15199);
nor U19973 (N_19973,N_17234,N_17422);
and U19974 (N_19974,N_15370,N_15375);
xnor U19975 (N_19975,N_15147,N_15568);
nand U19976 (N_19976,N_15706,N_17086);
or U19977 (N_19977,N_15468,N_16113);
and U19978 (N_19978,N_15485,N_16123);
nor U19979 (N_19979,N_15519,N_15987);
and U19980 (N_19980,N_16416,N_17468);
nand U19981 (N_19981,N_15864,N_15260);
or U19982 (N_19982,N_15704,N_16829);
and U19983 (N_19983,N_17083,N_16196);
or U19984 (N_19984,N_16997,N_16502);
nand U19985 (N_19985,N_15686,N_17296);
nor U19986 (N_19986,N_15843,N_17204);
nor U19987 (N_19987,N_15498,N_17149);
nor U19988 (N_19988,N_16109,N_17074);
or U19989 (N_19989,N_15491,N_15927);
xor U19990 (N_19990,N_16461,N_15858);
nor U19991 (N_19991,N_16858,N_17063);
nand U19992 (N_19992,N_16986,N_17112);
and U19993 (N_19993,N_16914,N_16265);
nor U19994 (N_19994,N_15603,N_17166);
nand U19995 (N_19995,N_16157,N_16090);
nor U19996 (N_19996,N_16995,N_17430);
xnor U19997 (N_19997,N_15107,N_16151);
or U19998 (N_19998,N_17119,N_16657);
nand U19999 (N_19999,N_17470,N_15123);
and U20000 (N_20000,N_19203,N_19234);
or U20001 (N_20001,N_19171,N_18303);
and U20002 (N_20002,N_19660,N_19609);
nand U20003 (N_20003,N_18580,N_19284);
or U20004 (N_20004,N_17569,N_19427);
xnor U20005 (N_20005,N_19201,N_18215);
nand U20006 (N_20006,N_19839,N_18375);
and U20007 (N_20007,N_19340,N_19191);
nand U20008 (N_20008,N_17893,N_17649);
xor U20009 (N_20009,N_18717,N_17756);
nor U20010 (N_20010,N_17629,N_18689);
or U20011 (N_20011,N_18780,N_18735);
or U20012 (N_20012,N_19827,N_18739);
or U20013 (N_20013,N_18946,N_18449);
nand U20014 (N_20014,N_19920,N_19715);
and U20015 (N_20015,N_19644,N_17774);
xor U20016 (N_20016,N_18013,N_18980);
nor U20017 (N_20017,N_18579,N_19147);
nor U20018 (N_20018,N_18820,N_19941);
or U20019 (N_20019,N_17980,N_17910);
nor U20020 (N_20020,N_17913,N_18070);
nor U20021 (N_20021,N_18959,N_17578);
xor U20022 (N_20022,N_18646,N_19413);
xnor U20023 (N_20023,N_18655,N_19455);
nor U20024 (N_20024,N_18041,N_18268);
xnor U20025 (N_20025,N_19145,N_19030);
or U20026 (N_20026,N_17834,N_19823);
and U20027 (N_20027,N_19865,N_18397);
xor U20028 (N_20028,N_19007,N_19228);
nand U20029 (N_20029,N_18290,N_18388);
nor U20030 (N_20030,N_17722,N_19965);
xor U20031 (N_20031,N_17602,N_19175);
nor U20032 (N_20032,N_19209,N_18373);
nor U20033 (N_20033,N_18639,N_19277);
nand U20034 (N_20034,N_18866,N_19112);
and U20035 (N_20035,N_18836,N_18441);
and U20036 (N_20036,N_17786,N_19970);
nand U20037 (N_20037,N_19775,N_18434);
nand U20038 (N_20038,N_18887,N_17622);
and U20039 (N_20039,N_19747,N_17995);
or U20040 (N_20040,N_19326,N_18052);
xnor U20041 (N_20041,N_19074,N_19297);
or U20042 (N_20042,N_19799,N_18599);
or U20043 (N_20043,N_18368,N_18092);
xnor U20044 (N_20044,N_19647,N_19801);
and U20045 (N_20045,N_17587,N_18586);
nand U20046 (N_20046,N_18164,N_18109);
nor U20047 (N_20047,N_17997,N_19378);
nand U20048 (N_20048,N_18988,N_19534);
xor U20049 (N_20049,N_18690,N_19946);
nor U20050 (N_20050,N_17585,N_17753);
nand U20051 (N_20051,N_18423,N_17627);
or U20052 (N_20052,N_17646,N_19515);
nor U20053 (N_20053,N_19876,N_19046);
and U20054 (N_20054,N_18912,N_19936);
and U20055 (N_20055,N_19282,N_18653);
nand U20056 (N_20056,N_17767,N_19097);
xnor U20057 (N_20057,N_18036,N_19873);
or U20058 (N_20058,N_19295,N_18654);
nor U20059 (N_20059,N_17556,N_19280);
nor U20060 (N_20060,N_17965,N_18117);
xnor U20061 (N_20061,N_19505,N_18517);
nor U20062 (N_20062,N_19819,N_18594);
nand U20063 (N_20063,N_19858,N_18811);
xnor U20064 (N_20064,N_17683,N_17591);
or U20065 (N_20065,N_19196,N_17616);
or U20066 (N_20066,N_17581,N_17594);
and U20067 (N_20067,N_18411,N_17668);
nand U20068 (N_20068,N_19997,N_19657);
and U20069 (N_20069,N_17961,N_19052);
or U20070 (N_20070,N_18663,N_19208);
nand U20071 (N_20071,N_17524,N_17750);
nand U20072 (N_20072,N_18455,N_19829);
nor U20073 (N_20073,N_19600,N_17917);
xor U20074 (N_20074,N_18754,N_18084);
or U20075 (N_20075,N_18349,N_19539);
nand U20076 (N_20076,N_19456,N_17692);
nand U20077 (N_20077,N_18393,N_18079);
and U20078 (N_20078,N_18855,N_17680);
nor U20079 (N_20079,N_18583,N_18021);
xor U20080 (N_20080,N_17988,N_19069);
or U20081 (N_20081,N_19878,N_19899);
nand U20082 (N_20082,N_19065,N_18243);
and U20083 (N_20083,N_18775,N_18899);
nor U20084 (N_20084,N_19963,N_18022);
nor U20085 (N_20085,N_19494,N_19240);
nand U20086 (N_20086,N_19791,N_19077);
nand U20087 (N_20087,N_18757,N_18809);
nor U20088 (N_20088,N_18324,N_18687);
or U20089 (N_20089,N_18996,N_18045);
nor U20090 (N_20090,N_18240,N_17542);
nand U20091 (N_20091,N_19532,N_19583);
nor U20092 (N_20092,N_19003,N_18982);
and U20093 (N_20093,N_17533,N_18512);
nor U20094 (N_20094,N_17638,N_19479);
xnor U20095 (N_20095,N_19258,N_19501);
xor U20096 (N_20096,N_19137,N_19437);
nor U20097 (N_20097,N_19931,N_18313);
xnor U20098 (N_20098,N_17945,N_19108);
and U20099 (N_20099,N_18112,N_19638);
nand U20100 (N_20100,N_18204,N_17943);
and U20101 (N_20101,N_17900,N_18800);
nand U20102 (N_20102,N_19754,N_18029);
xnor U20103 (N_20103,N_18573,N_17985);
nand U20104 (N_20104,N_19588,N_19338);
nand U20105 (N_20105,N_18130,N_18718);
xor U20106 (N_20106,N_19076,N_18776);
nand U20107 (N_20107,N_18475,N_17747);
nor U20108 (N_20108,N_17857,N_19058);
nor U20109 (N_20109,N_19336,N_19418);
nand U20110 (N_20110,N_18258,N_19803);
nor U20111 (N_20111,N_18154,N_19227);
xor U20112 (N_20112,N_19188,N_18424);
xnor U20113 (N_20113,N_19808,N_19582);
nor U20114 (N_20114,N_19810,N_19511);
and U20115 (N_20115,N_18960,N_18330);
nor U20116 (N_20116,N_18315,N_19843);
or U20117 (N_20117,N_18616,N_18014);
nand U20118 (N_20118,N_19700,N_18557);
or U20119 (N_20119,N_18385,N_17553);
or U20120 (N_20120,N_18951,N_17953);
xnor U20121 (N_20121,N_17826,N_19606);
nor U20122 (N_20122,N_19006,N_18514);
xor U20123 (N_20123,N_19397,N_19910);
and U20124 (N_20124,N_19812,N_17992);
nand U20125 (N_20125,N_17711,N_18958);
nor U20126 (N_20126,N_19620,N_18543);
nor U20127 (N_20127,N_19449,N_18762);
and U20128 (N_20128,N_17755,N_19376);
and U20129 (N_20129,N_19921,N_19541);
or U20130 (N_20130,N_19204,N_17510);
nand U20131 (N_20131,N_18012,N_18291);
nand U20132 (N_20132,N_19919,N_17549);
and U20133 (N_20133,N_18668,N_18231);
nor U20134 (N_20134,N_18892,N_18948);
or U20135 (N_20135,N_19636,N_17687);
nor U20136 (N_20136,N_18788,N_18321);
nand U20137 (N_20137,N_18636,N_18519);
xor U20138 (N_20138,N_19496,N_18587);
xnor U20139 (N_20139,N_18875,N_17665);
and U20140 (N_20140,N_18394,N_18938);
nor U20141 (N_20141,N_17563,N_19684);
nand U20142 (N_20142,N_19205,N_19372);
or U20143 (N_20143,N_18419,N_17684);
or U20144 (N_20144,N_18572,N_19522);
xor U20145 (N_20145,N_18310,N_18001);
nand U20146 (N_20146,N_19633,N_19691);
or U20147 (N_20147,N_19635,N_19781);
or U20148 (N_20148,N_17671,N_18561);
nor U20149 (N_20149,N_18340,N_19559);
xnor U20150 (N_20150,N_19987,N_18031);
and U20151 (N_20151,N_17879,N_18083);
nand U20152 (N_20152,N_18241,N_19009);
nor U20153 (N_20153,N_18223,N_18500);
and U20154 (N_20154,N_18382,N_18848);
nand U20155 (N_20155,N_19624,N_18984);
and U20156 (N_20156,N_18674,N_18644);
xor U20157 (N_20157,N_17850,N_19415);
or U20158 (N_20158,N_19663,N_19168);
xor U20159 (N_20159,N_18074,N_19520);
xor U20160 (N_20160,N_18128,N_19063);
nand U20161 (N_20161,N_18658,N_19883);
nand U20162 (N_20162,N_19802,N_18023);
and U20163 (N_20163,N_18358,N_19669);
or U20164 (N_20164,N_18546,N_19879);
nand U20165 (N_20165,N_19288,N_18795);
and U20166 (N_20166,N_17866,N_18915);
nand U20167 (N_20167,N_19521,N_18244);
and U20168 (N_20168,N_19637,N_19080);
nand U20169 (N_20169,N_17650,N_18486);
xnor U20170 (N_20170,N_19184,N_19574);
or U20171 (N_20171,N_18277,N_19032);
nand U20172 (N_20172,N_19840,N_18198);
nor U20173 (N_20173,N_18945,N_19938);
xor U20174 (N_20174,N_17895,N_19821);
nor U20175 (N_20175,N_18095,N_18671);
nor U20176 (N_20176,N_19547,N_17534);
xor U20177 (N_20177,N_17944,N_18008);
or U20178 (N_20178,N_19962,N_19194);
nand U20179 (N_20179,N_17809,N_19044);
xnor U20180 (N_20180,N_18961,N_19426);
or U20181 (N_20181,N_19986,N_19526);
nand U20182 (N_20182,N_19897,N_19922);
and U20183 (N_20183,N_18501,N_17908);
nand U20184 (N_20184,N_19849,N_19272);
or U20185 (N_20185,N_17874,N_17801);
nor U20186 (N_20186,N_17823,N_18220);
and U20187 (N_20187,N_19323,N_17807);
and U20188 (N_20188,N_19318,N_18759);
or U20189 (N_20189,N_19434,N_19560);
xnor U20190 (N_20190,N_19837,N_19422);
nor U20191 (N_20191,N_19195,N_18905);
nor U20192 (N_20192,N_18421,N_17623);
and U20193 (N_20193,N_18534,N_18177);
and U20194 (N_20194,N_18794,N_17564);
nor U20195 (N_20195,N_17886,N_19694);
xor U20196 (N_20196,N_19414,N_18347);
nand U20197 (N_20197,N_17509,N_19214);
and U20198 (N_20198,N_19450,N_17825);
xor U20199 (N_20199,N_17969,N_18480);
nand U20200 (N_20200,N_19551,N_18098);
nand U20201 (N_20201,N_18907,N_17625);
or U20202 (N_20202,N_17941,N_19890);
and U20203 (N_20203,N_18798,N_18054);
or U20204 (N_20204,N_17718,N_19010);
or U20205 (N_20205,N_17588,N_18765);
xnor U20206 (N_20206,N_18737,N_18554);
and U20207 (N_20207,N_19000,N_17685);
nor U20208 (N_20208,N_18099,N_19088);
xnor U20209 (N_20209,N_19474,N_19748);
and U20210 (N_20210,N_18357,N_18166);
and U20211 (N_20211,N_19590,N_19085);
nand U20212 (N_20212,N_18962,N_17951);
or U20213 (N_20213,N_19761,N_17847);
and U20214 (N_20214,N_19924,N_18100);
and U20215 (N_20215,N_18222,N_17604);
and U20216 (N_20216,N_18513,N_18863);
and U20217 (N_20217,N_18416,N_18481);
and U20218 (N_20218,N_18366,N_19223);
nand U20219 (N_20219,N_19374,N_18474);
nor U20220 (N_20220,N_18523,N_19724);
nor U20221 (N_20221,N_17781,N_19176);
nand U20222 (N_20222,N_18560,N_18448);
nor U20223 (N_20223,N_17572,N_18401);
nor U20224 (N_20224,N_19550,N_19460);
nand U20225 (N_20225,N_18977,N_18131);
and U20226 (N_20226,N_19210,N_19442);
nand U20227 (N_20227,N_18856,N_18732);
and U20228 (N_20228,N_19239,N_19777);
nor U20229 (N_20229,N_19867,N_17610);
nor U20230 (N_20230,N_19676,N_18123);
nand U20231 (N_20231,N_19198,N_19916);
or U20232 (N_20232,N_19463,N_18547);
nor U20233 (N_20233,N_19001,N_17603);
xnor U20234 (N_20234,N_19101,N_19394);
nand U20235 (N_20235,N_18115,N_18767);
nand U20236 (N_20236,N_17614,N_18816);
nor U20237 (N_20237,N_18544,N_17700);
nand U20238 (N_20238,N_18017,N_19653);
nand U20239 (N_20239,N_18778,N_19996);
nand U20240 (N_20240,N_18077,N_18069);
or U20241 (N_20241,N_19904,N_18728);
nor U20242 (N_20242,N_17624,N_17837);
or U20243 (N_20243,N_18018,N_19587);
nand U20244 (N_20244,N_17651,N_19557);
nor U20245 (N_20245,N_18921,N_17762);
nand U20246 (N_20246,N_19264,N_17738);
nand U20247 (N_20247,N_19093,N_19351);
nand U20248 (N_20248,N_19285,N_19842);
or U20249 (N_20249,N_19682,N_18659);
or U20250 (N_20250,N_19267,N_19433);
nand U20251 (N_20251,N_18155,N_17729);
nor U20252 (N_20252,N_19154,N_19537);
nor U20253 (N_20253,N_18807,N_19266);
nand U20254 (N_20254,N_19646,N_18588);
nand U20255 (N_20255,N_19424,N_18693);
or U20256 (N_20256,N_17559,N_18539);
nand U20257 (N_20257,N_18632,N_18064);
xnor U20258 (N_20258,N_18242,N_17686);
xnor U20259 (N_20259,N_19478,N_17708);
nand U20260 (N_20260,N_18652,N_17719);
and U20261 (N_20261,N_19788,N_19752);
and U20262 (N_20262,N_19298,N_18265);
and U20263 (N_20263,N_19882,N_19612);
xnor U20264 (N_20264,N_19991,N_19807);
nor U20265 (N_20265,N_19739,N_19571);
nor U20266 (N_20266,N_18857,N_19610);
nor U20267 (N_20267,N_19177,N_19385);
xnor U20268 (N_20268,N_18461,N_19130);
xnor U20269 (N_20269,N_19432,N_19743);
or U20270 (N_20270,N_17731,N_17820);
xnor U20271 (N_20271,N_19110,N_18338);
and U20272 (N_20272,N_18348,N_19850);
nand U20273 (N_20273,N_18483,N_18217);
xor U20274 (N_20274,N_19832,N_18159);
xor U20275 (N_20275,N_19325,N_18578);
or U20276 (N_20276,N_18950,N_18575);
or U20277 (N_20277,N_18142,N_18730);
or U20278 (N_20278,N_19746,N_17503);
and U20279 (N_20279,N_18153,N_17643);
or U20280 (N_20280,N_18633,N_18374);
xnor U20281 (N_20281,N_19341,N_18495);
and U20282 (N_20282,N_18426,N_17896);
and U20283 (N_20283,N_18367,N_19072);
nor U20284 (N_20284,N_18510,N_17771);
xnor U20285 (N_20285,N_19309,N_19441);
nor U20286 (N_20286,N_19666,N_18829);
nand U20287 (N_20287,N_19430,N_17570);
or U20288 (N_20288,N_17675,N_19079);
xor U20289 (N_20289,N_17979,N_18630);
nor U20290 (N_20290,N_19236,N_19985);
or U20291 (N_20291,N_18034,N_17792);
xnor U20292 (N_20292,N_19680,N_18381);
and U20293 (N_20293,N_18953,N_19678);
nand U20294 (N_20294,N_19891,N_18515);
or U20295 (N_20295,N_19507,N_19186);
nor U20296 (N_20296,N_18797,N_18695);
nand U20297 (N_20297,N_18876,N_19102);
nor U20298 (N_20298,N_17696,N_19768);
xor U20299 (N_20299,N_19081,N_19868);
nand U20300 (N_20300,N_19824,N_19956);
nor U20301 (N_20301,N_19770,N_17609);
and U20302 (N_20302,N_19874,N_19984);
nand U20303 (N_20303,N_18226,N_18460);
and U20304 (N_20304,N_19671,N_18882);
nand U20305 (N_20305,N_18102,N_19139);
nor U20306 (N_20306,N_18238,N_18346);
and U20307 (N_20307,N_19595,N_19448);
nand U20308 (N_20308,N_19216,N_18939);
nor U20309 (N_20309,N_17906,N_17612);
and U20310 (N_20310,N_17827,N_18667);
nand U20311 (N_20311,N_18647,N_18505);
or U20312 (N_20312,N_19159,N_19524);
nor U20313 (N_20313,N_17661,N_17778);
nand U20314 (N_20314,N_17514,N_18075);
nand U20315 (N_20315,N_18201,N_18997);
nand U20316 (N_20316,N_19673,N_19136);
xnor U20317 (N_20317,N_17543,N_19912);
nand U20318 (N_20318,N_18145,N_19632);
xor U20319 (N_20319,N_18901,N_18987);
nor U20320 (N_20320,N_19974,N_19654);
and U20321 (N_20321,N_17950,N_19623);
or U20322 (N_20322,N_18817,N_18040);
xnor U20323 (N_20323,N_17764,N_17601);
nand U20324 (N_20324,N_18600,N_17811);
and U20325 (N_20325,N_19569,N_19969);
or U20326 (N_20326,N_19625,N_17615);
and U20327 (N_20327,N_17983,N_18047);
xor U20328 (N_20328,N_18378,N_19324);
nor U20329 (N_20329,N_18685,N_19271);
or U20330 (N_20330,N_18278,N_18431);
and U20331 (N_20331,N_17586,N_18429);
or U20332 (N_20332,N_18071,N_19469);
xor U20333 (N_20333,N_19482,N_17517);
xnor U20334 (N_20334,N_18974,N_19199);
nor U20335 (N_20335,N_19627,N_19012);
nand U20336 (N_20336,N_18518,N_19056);
nor U20337 (N_20337,N_18136,N_17880);
or U20338 (N_20338,N_17676,N_18914);
xor U20339 (N_20339,N_19529,N_19034);
or U20340 (N_20340,N_17853,N_19446);
and U20341 (N_20341,N_19814,N_19202);
xnor U20342 (N_20342,N_18604,N_18403);
or U20343 (N_20343,N_19993,N_19047);
or U20344 (N_20344,N_19121,N_19779);
or U20345 (N_20345,N_19668,N_19545);
nand U20346 (N_20346,N_18398,N_18279);
nor U20347 (N_20347,N_18878,N_19525);
xor U20348 (N_20348,N_18504,N_17999);
or U20349 (N_20349,N_18952,N_18802);
and U20350 (N_20350,N_17710,N_19585);
or U20351 (N_20351,N_19117,N_17911);
nand U20352 (N_20352,N_17653,N_19346);
xnor U20353 (N_20353,N_19975,N_19407);
or U20354 (N_20354,N_19160,N_18967);
xor U20355 (N_20355,N_19115,N_18272);
xnor U20356 (N_20356,N_19445,N_18189);
xnor U20357 (N_20357,N_19572,N_18463);
or U20358 (N_20358,N_18993,N_18799);
nand U20359 (N_20359,N_18063,N_18631);
nand U20360 (N_20360,N_19020,N_19608);
and U20361 (N_20361,N_19417,N_18005);
or U20362 (N_20362,N_18270,N_19384);
xor U20363 (N_20363,N_19322,N_17730);
xnor U20364 (N_20364,N_17751,N_18839);
or U20365 (N_20365,N_17785,N_17986);
nand U20366 (N_20366,N_19253,N_18511);
xor U20367 (N_20367,N_18981,N_19262);
nor U20368 (N_20368,N_19717,N_19804);
xnor U20369 (N_20369,N_18453,N_17923);
and U20370 (N_20370,N_19294,N_19365);
nand U20371 (N_20371,N_19690,N_19465);
nand U20372 (N_20372,N_19190,N_18758);
and U20373 (N_20373,N_19584,N_19562);
and U20374 (N_20374,N_18004,N_18733);
and U20375 (N_20375,N_19734,N_19983);
nand U20376 (N_20376,N_18976,N_19287);
or U20377 (N_20377,N_19650,N_19800);
and U20378 (N_20378,N_18328,N_17991);
or U20379 (N_20379,N_18789,N_19630);
or U20380 (N_20380,N_18091,N_19075);
nor U20381 (N_20381,N_18471,N_19982);
and U20382 (N_20382,N_18492,N_18050);
and U20383 (N_20383,N_17737,N_19042);
nor U20384 (N_20384,N_19316,N_18752);
or U20385 (N_20385,N_17987,N_19221);
or U20386 (N_20386,N_17800,N_17916);
nand U20387 (N_20387,N_19548,N_19999);
nor U20388 (N_20388,N_18576,N_18716);
or U20389 (N_20389,N_19392,N_18094);
nand U20390 (N_20390,N_19181,N_18979);
and U20391 (N_20391,N_18656,N_19499);
nand U20392 (N_20392,N_18942,N_19943);
and U20393 (N_20393,N_19157,N_17688);
nand U20394 (N_20394,N_19447,N_19039);
and U20395 (N_20395,N_19254,N_18773);
or U20396 (N_20396,N_19213,N_18985);
nand U20397 (N_20397,N_19018,N_18266);
or U20398 (N_20398,N_19207,N_18086);
or U20399 (N_20399,N_19131,N_17791);
nand U20400 (N_20400,N_18288,N_19581);
or U20401 (N_20401,N_18184,N_19495);
and U20402 (N_20402,N_18305,N_19652);
and U20403 (N_20403,N_19579,N_19165);
nand U20404 (N_20404,N_18540,N_17597);
and U20405 (N_20405,N_19492,N_19621);
xnor U20406 (N_20406,N_19290,N_18582);
xnor U20407 (N_20407,N_19846,N_19396);
nor U20408 (N_20408,N_18456,N_19146);
nand U20409 (N_20409,N_18396,N_19477);
nor U20410 (N_20410,N_19771,N_18710);
and U20411 (N_20411,N_18812,N_19915);
nand U20412 (N_20412,N_18476,N_19733);
and U20413 (N_20413,N_19774,N_19320);
nor U20414 (N_20414,N_19352,N_17735);
or U20415 (N_20415,N_19778,N_17626);
xor U20416 (N_20416,N_19235,N_19906);
or U20417 (N_20417,N_19566,N_17842);
or U20418 (N_20418,N_18726,N_19467);
or U20419 (N_20419,N_19293,N_19838);
nor U20420 (N_20420,N_19642,N_18617);
or U20421 (N_20421,N_18181,N_19513);
or U20422 (N_20422,N_18193,N_17899);
nor U20423 (N_20423,N_19613,N_18384);
nor U20424 (N_20424,N_18746,N_19593);
nand U20425 (N_20425,N_18529,N_19831);
and U20426 (N_20426,N_18833,N_19930);
xnor U20427 (N_20427,N_18408,N_18202);
and U20428 (N_20428,N_18769,N_18623);
and U20429 (N_20429,N_17981,N_19751);
or U20430 (N_20430,N_17838,N_19935);
xor U20431 (N_20431,N_17511,N_19366);
nand U20432 (N_20432,N_18601,N_18885);
nand U20433 (N_20433,N_19933,N_19783);
xnor U20434 (N_20434,N_19119,N_18944);
nand U20435 (N_20435,N_18312,N_18565);
xnor U20436 (N_20436,N_18286,N_18254);
nand U20437 (N_20437,N_17971,N_18485);
or U20438 (N_20438,N_17724,N_18405);
xor U20439 (N_20439,N_19518,N_18584);
and U20440 (N_20440,N_19502,N_18611);
nand U20441 (N_20441,N_18669,N_17887);
and U20442 (N_20442,N_18719,N_19078);
and U20443 (N_20443,N_18249,N_19345);
nor U20444 (N_20444,N_17829,N_19408);
or U20445 (N_20445,N_19714,N_19880);
or U20446 (N_20446,N_18299,N_18256);
xnor U20447 (N_20447,N_18057,N_19311);
nor U20448 (N_20448,N_17743,N_19315);
or U20449 (N_20449,N_19556,N_19404);
xor U20450 (N_20450,N_18119,N_19973);
nand U20451 (N_20451,N_18770,N_18538);
and U20452 (N_20452,N_18457,N_18059);
or U20453 (N_20453,N_19674,N_18972);
or U20454 (N_20454,N_19640,N_19805);
xor U20455 (N_20455,N_17960,N_19382);
nor U20456 (N_20456,N_19022,N_18629);
nor U20457 (N_20457,N_17841,N_19765);
nand U20458 (N_20458,N_18725,N_18747);
nor U20459 (N_20459,N_18068,N_18955);
nor U20460 (N_20460,N_19677,N_19535);
nand U20461 (N_20461,N_18097,N_19737);
nor U20462 (N_20462,N_19604,N_19709);
or U20463 (N_20463,N_19084,N_19319);
and U20464 (N_20464,N_18415,N_18487);
and U20465 (N_20465,N_17888,N_19243);
xor U20466 (N_20466,N_18918,N_19538);
nor U20467 (N_20467,N_18285,N_17773);
nand U20468 (N_20468,N_18933,N_17975);
or U20469 (N_20469,N_18847,N_18870);
nand U20470 (N_20470,N_17790,N_17545);
and U20471 (N_20471,N_18503,N_18280);
nand U20472 (N_20472,N_19634,N_19332);
and U20473 (N_20473,N_17717,N_18462);
xnor U20474 (N_20474,N_17740,N_19237);
and U20475 (N_20475,N_19163,N_19905);
nor U20476 (N_20476,N_18205,N_18566);
xor U20477 (N_20477,N_19189,N_18026);
nand U20478 (N_20478,N_18530,N_18006);
or U20479 (N_20479,N_17930,N_17600);
or U20480 (N_20480,N_18383,N_18211);
nor U20481 (N_20481,N_17577,N_19813);
nand U20482 (N_20482,N_19051,N_19158);
nor U20483 (N_20483,N_18339,N_18821);
nor U20484 (N_20484,N_18978,N_17844);
nand U20485 (N_20485,N_18407,N_19344);
and U20486 (N_20486,N_19054,N_17636);
nand U20487 (N_20487,N_17652,N_19488);
nor U20488 (N_20488,N_19387,N_18046);
xnor U20489 (N_20489,N_18174,N_18402);
xnor U20490 (N_20490,N_18909,N_19749);
nand U20491 (N_20491,N_19383,N_19252);
nor U20492 (N_20492,N_17836,N_17561);
nand U20493 (N_20493,N_18729,N_19002);
or U20494 (N_20494,N_18236,N_19485);
nand U20495 (N_20495,N_18574,N_17904);
nor U20496 (N_20496,N_19528,N_19211);
xor U20497 (N_20497,N_19615,N_19589);
and U20498 (N_20498,N_19833,N_17878);
and U20499 (N_20499,N_18986,N_18218);
and U20500 (N_20500,N_18311,N_19607);
or U20501 (N_20501,N_19542,N_19603);
xor U20502 (N_20502,N_19767,N_18764);
nand U20503 (N_20503,N_19444,N_18742);
or U20504 (N_20504,N_18734,N_17905);
xor U20505 (N_20505,N_17967,N_18562);
nor U20506 (N_20506,N_19098,N_19464);
nor U20507 (N_20507,N_17647,N_18925);
nand U20508 (N_20508,N_17972,N_17933);
nand U20509 (N_20509,N_19742,N_18176);
nand U20510 (N_20510,N_19307,N_18323);
nor U20511 (N_20511,N_17537,N_18300);
and U20512 (N_20512,N_18536,N_19857);
nand U20513 (N_20513,N_18427,N_17544);
nor U20514 (N_20514,N_18372,N_19247);
xor U20515 (N_20515,N_17963,N_17558);
and U20516 (N_20516,N_18998,N_18360);
or U20517 (N_20517,N_18308,N_19178);
nand U20518 (N_20518,N_19575,N_18451);
xor U20519 (N_20519,N_18637,N_19955);
or U20520 (N_20520,N_19570,N_18105);
or U20521 (N_20521,N_17794,N_19103);
or U20522 (N_20522,N_18845,N_17984);
and U20523 (N_20523,N_19462,N_17645);
or U20524 (N_20524,N_19061,N_18420);
and U20525 (N_20525,N_18125,N_18852);
xnor U20526 (N_20526,N_19543,N_18889);
or U20527 (N_20527,N_19573,N_18930);
or U20528 (N_20528,N_18607,N_17787);
nand U20529 (N_20529,N_19889,N_18806);
xor U20530 (N_20530,N_18369,N_19645);
nand U20531 (N_20531,N_18060,N_18361);
nor U20532 (N_20532,N_19330,N_18715);
nor U20533 (N_20533,N_18395,N_18399);
and U20534 (N_20534,N_18787,N_17681);
and U20535 (N_20535,N_17552,N_19491);
and U20536 (N_20536,N_19967,N_17697);
or U20537 (N_20537,N_18609,N_18531);
xnor U20538 (N_20538,N_19519,N_17765);
and U20539 (N_20539,N_19500,N_19489);
or U20540 (N_20540,N_18731,N_17690);
nor U20541 (N_20541,N_19419,N_19784);
nor U20542 (N_20542,N_17940,N_18167);
nand U20543 (N_20543,N_19504,N_17573);
and U20544 (N_20544,N_18188,N_18853);
or U20545 (N_20545,N_18147,N_17956);
xor U20546 (N_20546,N_19818,N_18203);
xor U20547 (N_20547,N_19877,N_19333);
xnor U20548 (N_20548,N_18350,N_19468);
and U20549 (N_20549,N_18065,N_18871);
or U20550 (N_20550,N_17968,N_18877);
and U20551 (N_20551,N_18883,N_17901);
xor U20552 (N_20552,N_19859,N_17958);
or U20553 (N_20553,N_19483,N_19134);
or U20554 (N_20554,N_18854,N_19552);
nand U20555 (N_20555,N_18927,N_19934);
nand U20556 (N_20556,N_19286,N_19918);
nand U20557 (N_20557,N_19454,N_18180);
xor U20558 (N_20558,N_18454,N_18537);
nor U20559 (N_20559,N_18225,N_19256);
and U20560 (N_20560,N_17978,N_18319);
nor U20561 (N_20561,N_19370,N_18376);
and U20562 (N_20562,N_18559,N_19672);
nand U20563 (N_20563,N_19536,N_19992);
xor U20564 (N_20564,N_19452,N_19817);
xor U20565 (N_20565,N_19830,N_18468);
or U20566 (N_20566,N_18072,N_17877);
and U20567 (N_20567,N_17780,N_17760);
xnor U20568 (N_20568,N_18183,N_18651);
xor U20569 (N_20569,N_19728,N_18466);
and U20570 (N_20570,N_19692,N_18009);
and U20571 (N_20571,N_19192,N_19113);
nand U20572 (N_20572,N_19949,N_19968);
or U20573 (N_20573,N_19423,N_18263);
nand U20574 (N_20574,N_18790,N_18498);
or U20575 (N_20575,N_17890,N_19954);
nand U20576 (N_20576,N_18516,N_18963);
xnor U20577 (N_20577,N_18813,N_18294);
nor U20578 (N_20578,N_19231,N_19531);
and U20579 (N_20579,N_18801,N_19281);
nor U20580 (N_20580,N_18553,N_19816);
nor U20581 (N_20581,N_19241,N_18150);
or U20582 (N_20582,N_18973,N_19291);
nor U20583 (N_20583,N_18721,N_18199);
or U20584 (N_20584,N_18257,N_19390);
nor U20585 (N_20585,N_18822,N_18895);
xor U20586 (N_20586,N_19605,N_19353);
xor U20587 (N_20587,N_18470,N_18843);
and U20588 (N_20588,N_19435,N_19185);
nor U20589 (N_20589,N_19563,N_18133);
nor U20590 (N_20590,N_19270,N_18289);
xnor U20591 (N_20591,N_19095,N_18262);
xor U20592 (N_20592,N_19755,N_17725);
xnor U20593 (N_20593,N_19710,N_19699);
and U20594 (N_20594,N_18135,N_19038);
or U20595 (N_20595,N_18120,N_19031);
or U20596 (N_20596,N_19436,N_17793);
nand U20597 (N_20597,N_19440,N_17693);
nor U20598 (N_20598,N_17957,N_18774);
and U20599 (N_20599,N_18433,N_18569);
or U20600 (N_20600,N_18684,N_19402);
xor U20601 (N_20601,N_17889,N_18413);
nor U20602 (N_20602,N_18867,N_19082);
or U20603 (N_20603,N_19308,N_19594);
xor U20604 (N_20604,N_19212,N_18618);
or U20605 (N_20605,N_18160,N_18615);
and U20606 (N_20606,N_19327,N_18038);
and U20607 (N_20607,N_18784,N_19299);
xnor U20608 (N_20608,N_18824,N_17699);
xor U20609 (N_20609,N_19675,N_17550);
xnor U20610 (N_20610,N_19510,N_19126);
xnor U20611 (N_20611,N_19391,N_17810);
nor U20612 (N_20612,N_18314,N_19123);
and U20613 (N_20613,N_18763,N_19611);
or U20614 (N_20614,N_18612,N_18904);
or U20615 (N_20615,N_19166,N_19443);
nor U20616 (N_20616,N_19225,N_18956);
xor U20617 (N_20617,N_17639,N_19696);
xor U20618 (N_20618,N_17962,N_17855);
nand U20619 (N_20619,N_17560,N_19180);
nor U20620 (N_20620,N_19866,N_19957);
or U20621 (N_20621,N_17954,N_18702);
and U20622 (N_20622,N_18129,N_18840);
xnor U20623 (N_20623,N_18329,N_18722);
nor U20624 (N_20624,N_19116,N_17575);
nor U20625 (N_20625,N_18245,N_19961);
xor U20626 (N_20626,N_19041,N_19798);
xnor U20627 (N_20627,N_19527,N_18436);
nand U20628 (N_20628,N_18542,N_17659);
and U20629 (N_20629,N_18828,N_19664);
or U20630 (N_20630,N_19568,N_19355);
and U20631 (N_20631,N_18452,N_19648);
and U20632 (N_20632,N_19649,N_18228);
xor U20633 (N_20633,N_17734,N_17644);
xnor U20634 (N_20634,N_19120,N_18714);
and U20635 (N_20635,N_17802,N_17824);
and U20636 (N_20636,N_17507,N_17635);
and U20637 (N_20637,N_19722,N_19040);
nor U20638 (N_20638,N_18661,N_18425);
nand U20639 (N_20639,N_18049,N_17947);
nor U20640 (N_20640,N_17654,N_19481);
nor U20641 (N_20641,N_17830,N_19265);
nor U20642 (N_20642,N_18808,N_17536);
and U20643 (N_20643,N_18276,N_17746);
and U20644 (N_20644,N_18335,N_18971);
nor U20645 (N_20645,N_18248,N_19111);
nor U20646 (N_20646,N_19892,N_18171);
nand U20647 (N_20647,N_17831,N_17634);
xor U20648 (N_20648,N_18247,N_18192);
nor U20649 (N_20649,N_18620,N_18825);
xnor U20650 (N_20650,N_19451,N_19925);
or U20651 (N_20651,N_18649,N_18499);
nor U20652 (N_20652,N_18107,N_17512);
nand U20653 (N_20653,N_18896,N_19721);
or U20654 (N_20654,N_19245,N_19836);
nor U20655 (N_20655,N_19016,N_17694);
xor U20656 (N_20656,N_19903,N_18766);
and U20657 (N_20657,N_18657,N_19388);
nor U20658 (N_20658,N_18983,N_18191);
or U20659 (N_20659,N_18437,N_18085);
or U20660 (N_20660,N_19275,N_19894);
xor U20661 (N_20661,N_18819,N_18108);
xor U20662 (N_20662,N_19300,N_19458);
nand U20663 (N_20663,N_17858,N_19428);
or U20664 (N_20664,N_18010,N_18469);
or U20665 (N_20665,N_18744,N_18745);
nor U20666 (N_20666,N_19246,N_18298);
xnor U20667 (N_20667,N_18624,N_18989);
and U20668 (N_20668,N_18309,N_18482);
nor U20669 (N_20669,N_19151,N_18343);
xnor U20670 (N_20670,N_18114,N_18134);
nand U20671 (N_20671,N_19853,N_17522);
nor U20672 (N_20672,N_18545,N_18628);
xnor U20673 (N_20673,N_18634,N_18326);
nor U20674 (N_20674,N_17535,N_17921);
and U20675 (N_20675,N_17518,N_18796);
or U20676 (N_20676,N_18337,N_19193);
nand U20677 (N_20677,N_19851,N_18081);
or U20678 (N_20678,N_17727,N_19049);
and U20679 (N_20679,N_18214,N_18621);
or U20680 (N_20680,N_18027,N_18642);
or U20681 (N_20681,N_17589,N_17851);
and U20682 (N_20682,N_17974,N_18686);
nor U20683 (N_20683,N_18703,N_19218);
nand U20684 (N_20684,N_19347,N_17582);
nand U20685 (N_20685,N_18292,N_19662);
and U20686 (N_20686,N_18532,N_17523);
nand U20687 (N_20687,N_18409,N_18841);
and U20688 (N_20688,N_18080,N_19773);
xnor U20689 (N_20689,N_19944,N_18356);
xor U20690 (N_20690,N_17712,N_18489);
nand U20691 (N_20691,N_18391,N_17804);
nor U20692 (N_20692,N_17928,N_18858);
nor U20693 (N_20693,N_18253,N_19226);
or U20694 (N_20694,N_19546,N_17799);
nand U20695 (N_20695,N_19144,N_18352);
xnor U20696 (N_20696,N_17777,N_17715);
or U20697 (N_20697,N_18527,N_17633);
or U20698 (N_20698,N_17657,N_18528);
or U20699 (N_20699,N_18148,N_17935);
nand U20700 (N_20700,N_19472,N_19641);
nor U20701 (N_20701,N_17796,N_19170);
and U20702 (N_20702,N_17732,N_18488);
nand U20703 (N_20703,N_18152,N_19782);
xnor U20704 (N_20704,N_19224,N_19689);
or U20705 (N_20705,N_18761,N_19071);
and U20706 (N_20706,N_18318,N_19790);
nand U20707 (N_20707,N_19337,N_18704);
nor U20708 (N_20708,N_18246,N_18886);
nor U20709 (N_20709,N_17867,N_17562);
nand U20710 (N_20710,N_17752,N_19289);
nor U20711 (N_20711,N_19911,N_19685);
nand U20712 (N_20712,N_19329,N_18786);
nand U20713 (N_20713,N_18417,N_18182);
or U20714 (N_20714,N_17605,N_18713);
xor U20715 (N_20715,N_18900,N_19787);
and U20716 (N_20716,N_19011,N_17798);
xnor U20717 (N_20717,N_19244,N_19399);
nand U20718 (N_20718,N_19735,N_18791);
xor U20719 (N_20719,N_18753,N_19174);
and U20720 (N_20720,N_17598,N_17872);
nor U20721 (N_20721,N_17973,N_18011);
and U20722 (N_20722,N_19484,N_18779);
and U20723 (N_20723,N_18902,N_17839);
nand U20724 (N_20724,N_18273,N_19416);
xor U20725 (N_20725,N_17754,N_18506);
or U20726 (N_20726,N_19769,N_19533);
and U20727 (N_20727,N_17501,N_19182);
nand U20728 (N_20728,N_19037,N_17897);
or U20729 (N_20729,N_19960,N_18835);
nor U20730 (N_20730,N_17812,N_18304);
and U20731 (N_20731,N_19909,N_17705);
and U20732 (N_20732,N_19856,N_18336);
or U20733 (N_20733,N_17660,N_18558);
and U20734 (N_20734,N_19048,N_18535);
xnor U20735 (N_20735,N_17849,N_18297);
nand U20736 (N_20736,N_19806,N_17936);
or U20737 (N_20737,N_18302,N_18838);
nand U20738 (N_20738,N_19561,N_19549);
and U20739 (N_20739,N_19861,N_18570);
or U20740 (N_20740,N_18496,N_18943);
nand U20741 (N_20741,N_18024,N_17818);
nand U20742 (N_20742,N_19261,N_19470);
or U20743 (N_20743,N_18043,N_19403);
or U20744 (N_20744,N_19756,N_19506);
nor U20745 (N_20745,N_19888,N_19498);
and U20746 (N_20746,N_18947,N_19864);
or U20747 (N_20747,N_18931,N_19707);
xnor U20748 (N_20748,N_18389,N_18709);
or U20749 (N_20749,N_18364,N_18216);
nand U20750 (N_20750,N_19901,N_18665);
and U20751 (N_20751,N_18884,N_18724);
nand U20752 (N_20752,N_17758,N_17845);
xor U20753 (N_20753,N_17527,N_19055);
and U20754 (N_20754,N_19150,N_17576);
xnor U20755 (N_20755,N_18868,N_19401);
xnor U20756 (N_20756,N_19971,N_19053);
nor U20757 (N_20757,N_18768,N_19731);
or U20758 (N_20758,N_19643,N_19617);
xor U20759 (N_20759,N_18414,N_18645);
nor U20760 (N_20760,N_17832,N_19626);
nand U20761 (N_20761,N_19045,N_17881);
nor U20762 (N_20762,N_17806,N_17797);
and U20763 (N_20763,N_19004,N_18342);
nand U20764 (N_20764,N_18039,N_18333);
and U20765 (N_20765,N_19628,N_18048);
xor U20766 (N_20766,N_19425,N_18445);
or U20767 (N_20767,N_19486,N_18640);
xnor U20768 (N_20768,N_17779,N_18662);
nor U20769 (N_20769,N_17977,N_17606);
xor U20770 (N_20770,N_17689,N_18711);
nor U20771 (N_20771,N_18834,N_19599);
xnor U20772 (N_20772,N_19251,N_17990);
and U20773 (N_20773,N_19369,N_19953);
nor U20774 (N_20774,N_17915,N_19667);
nor U20775 (N_20775,N_19913,N_17541);
and U20776 (N_20776,N_17515,N_18844);
nor U20777 (N_20777,N_19860,N_18675);
or U20778 (N_20778,N_17863,N_17679);
and U20779 (N_20779,N_19328,N_17775);
nor U20780 (N_20780,N_17882,N_19597);
nand U20781 (N_20781,N_17768,N_18194);
or U20782 (N_20782,N_18316,N_17784);
nand U20783 (N_20783,N_19278,N_17593);
or U20784 (N_20784,N_18275,N_17621);
or U20785 (N_20785,N_19242,N_19757);
xnor U20786 (N_20786,N_17898,N_19907);
xnor U20787 (N_20787,N_17749,N_18941);
xnor U20788 (N_20788,N_17815,N_18598);
or U20789 (N_20789,N_17664,N_19023);
nor U20790 (N_20790,N_18861,N_19100);
and U20791 (N_20791,N_19555,N_19105);
or U20792 (N_20792,N_19279,N_18556);
nor U20793 (N_20793,N_19148,N_18705);
nor U20794 (N_20794,N_19222,N_19206);
or U20795 (N_20795,N_19708,N_19025);
nand U20796 (N_20796,N_17667,N_17828);
nor U20797 (N_20797,N_19567,N_19005);
and U20798 (N_20798,N_18044,N_18911);
xnor U20799 (N_20799,N_19043,N_18341);
xnor U20800 (N_20800,N_18581,N_18179);
and U20801 (N_20801,N_18992,N_19143);
nor U20802 (N_20802,N_19980,N_17516);
xnor U20803 (N_20803,N_18926,N_19792);
nor U20804 (N_20804,N_18917,N_17903);
and U20805 (N_20805,N_19162,N_17506);
and U20806 (N_20806,N_19033,N_19386);
xnor U20807 (N_20807,N_19273,N_18502);
and U20808 (N_20808,N_19848,N_17909);
or U20809 (N_20809,N_18030,N_19035);
nand U20810 (N_20810,N_17894,N_17757);
nand U20811 (N_20811,N_17822,N_18968);
or U20812 (N_20812,N_18567,N_18032);
nor U20813 (N_20813,N_18025,N_18227);
nor U20814 (N_20814,N_19586,N_17723);
and U20815 (N_20815,N_19884,N_18406);
or U20816 (N_20816,N_18287,N_17942);
xor U20817 (N_20817,N_19220,N_17728);
xnor U20818 (N_20818,N_18224,N_18234);
nand U20819 (N_20819,N_18771,N_19310);
or U20820 (N_20820,N_18804,N_19780);
nand U20821 (N_20821,N_19389,N_19854);
and U20822 (N_20822,N_19260,N_19947);
or U20823 (N_20823,N_18679,N_18697);
or U20824 (N_20824,N_19706,N_19681);
nand U20825 (N_20825,N_18593,N_19317);
xor U20826 (N_20826,N_18432,N_18688);
xnor U20827 (N_20827,N_19106,N_19380);
nor U20828 (N_20828,N_18003,N_17608);
and U20829 (N_20829,N_18660,N_18137);
xor U20830 (N_20830,N_19248,N_17931);
xor U20831 (N_20831,N_19367,N_17949);
or U20832 (N_20832,N_17502,N_18533);
and U20833 (N_20833,N_18410,N_18212);
nand U20834 (N_20834,N_19845,N_19013);
and U20835 (N_20835,N_19713,N_19128);
or U20836 (N_20836,N_18923,N_19429);
xor U20837 (N_20837,N_18261,N_17782);
nand U20838 (N_20838,N_19670,N_19565);
or U20839 (N_20839,N_19753,N_18066);
or U20840 (N_20840,N_18121,N_19927);
nand U20841 (N_20841,N_19269,N_18400);
and U20842 (N_20842,N_18862,N_17613);
nor U20843 (N_20843,N_19133,N_19368);
or U20844 (N_20844,N_19475,N_19683);
nor U20845 (N_20845,N_18736,N_18664);
and U20846 (N_20846,N_17803,N_18864);
xor U20847 (N_20847,N_18274,N_18803);
nand U20848 (N_20848,N_19411,N_18890);
nor U20849 (N_20849,N_19950,N_17776);
nor U20850 (N_20850,N_19091,N_17769);
nor U20851 (N_20851,N_19972,N_17856);
xor U20852 (N_20852,N_18879,N_17547);
nand U20853 (N_20853,N_18444,N_19118);
nand U20854 (N_20854,N_18701,N_17907);
and U20855 (N_20855,N_19558,N_18293);
xnor U20856 (N_20856,N_19978,N_19057);
xor U20857 (N_20857,N_19940,N_18966);
nand U20858 (N_20858,N_18842,N_17574);
xor U20859 (N_20859,N_17920,N_19335);
or U20860 (N_20860,N_19981,N_19886);
or U20861 (N_20861,N_18015,N_17970);
and U20862 (N_20862,N_19863,N_19109);
xnor U20863 (N_20863,N_17892,N_17805);
and U20864 (N_20864,N_19200,N_19598);
xnor U20865 (N_20865,N_17584,N_18740);
and U20866 (N_20866,N_18712,N_19990);
and U20867 (N_20867,N_18723,N_17736);
nor U20868 (N_20868,N_19512,N_18033);
nand U20869 (N_20869,N_18317,N_18781);
and U20870 (N_20870,N_19629,N_17555);
or U20871 (N_20871,N_19375,N_19759);
and U20872 (N_20872,N_19169,N_17583);
xnor U20873 (N_20873,N_19233,N_17865);
nand U20874 (N_20874,N_18990,N_18677);
or U20875 (N_20875,N_18439,N_19362);
xor U20876 (N_20876,N_19296,N_17937);
nor U20877 (N_20877,N_19702,N_18999);
and U20878 (N_20878,N_19926,N_18296);
nand U20879 (N_20879,N_19809,N_18355);
nor U20880 (N_20880,N_19420,N_19720);
xor U20881 (N_20881,N_19871,N_19409);
nand U20882 (N_20882,N_17551,N_19885);
nand U20883 (N_20883,N_18549,N_19008);
xnor U20884 (N_20884,N_18118,N_17870);
or U20885 (N_20885,N_18748,N_17673);
and U20886 (N_20886,N_18541,N_18673);
nor U20887 (N_20887,N_17532,N_19862);
nor U20888 (N_20888,N_19517,N_18269);
nor U20889 (N_20889,N_17672,N_19847);
xor U20890 (N_20890,N_18823,N_18363);
nor U20891 (N_20891,N_19219,N_19466);
and U20892 (N_20892,N_19197,N_19099);
xnor U20893 (N_20893,N_19738,N_18446);
xnor U20894 (N_20894,N_18073,N_17628);
and U20895 (N_20895,N_17707,N_19697);
xnor U20896 (N_20896,N_19073,N_18681);
nand U20897 (N_20897,N_17617,N_17925);
nor U20898 (N_20898,N_19135,N_17833);
xor U20899 (N_20899,N_18035,N_19658);
or U20900 (N_20900,N_18459,N_19132);
nand U20901 (N_20901,N_18334,N_18161);
or U20902 (N_20902,N_18386,N_18390);
nor U20903 (N_20903,N_18332,N_19686);
or U20904 (N_20904,N_18111,N_18260);
nor U20905 (N_20905,N_19744,N_19977);
xnor U20906 (N_20906,N_18613,N_18846);
or U20907 (N_20907,N_19917,N_17619);
xnor U20908 (N_20908,N_17580,N_19263);
nor U20909 (N_20909,N_19869,N_19381);
nand U20910 (N_20910,N_19622,N_17666);
nor U20911 (N_20911,N_19173,N_18141);
or U20912 (N_20912,N_17948,N_18850);
nor U20913 (N_20913,N_18162,N_17701);
nor U20914 (N_20914,N_19364,N_18144);
xnor U20915 (N_20915,N_17912,N_19343);
nand U20916 (N_20916,N_19453,N_17546);
xnor U20917 (N_20917,N_17808,N_18307);
or U20918 (N_20918,N_18590,N_19576);
and U20919 (N_20919,N_17964,N_17565);
nor U20920 (N_20920,N_18196,N_18259);
nor U20921 (N_20921,N_18826,N_18320);
xor U20922 (N_20922,N_19083,N_19966);
or U20923 (N_20923,N_19406,N_19094);
xnor U20924 (N_20924,N_19359,N_18916);
and U20925 (N_20925,N_18106,N_19480);
or U20926 (N_20926,N_18815,N_17982);
nand U20927 (N_20927,N_19793,N_18187);
nand U20928 (N_20928,N_18707,N_17658);
and U20929 (N_20929,N_18699,N_19070);
and U20930 (N_20930,N_19014,N_17713);
or U20931 (N_20931,N_19564,N_18555);
and U20932 (N_20932,N_18638,N_19473);
nor U20933 (N_20933,N_19421,N_17620);
nor U20934 (N_20934,N_19902,N_18377);
or U20935 (N_20935,N_18362,N_18200);
xor U20936 (N_20936,N_19503,N_19152);
or U20937 (N_20937,N_19716,N_19772);
nor U20938 (N_20938,N_19230,N_19619);
nor U20939 (N_20939,N_18888,N_18219);
nand U20940 (N_20940,N_19026,N_18772);
xnor U20941 (N_20941,N_19596,N_18650);
and U20942 (N_20942,N_17934,N_17611);
xnor U20943 (N_20943,N_18920,N_19736);
nand U20944 (N_20944,N_19929,N_18233);
xnor U20945 (N_20945,N_18969,N_19350);
nor U20946 (N_20946,N_19107,N_18970);
and U20947 (N_20947,N_19951,N_19896);
nor U20948 (N_20948,N_18306,N_19740);
xor U20949 (N_20949,N_18509,N_18881);
or U20950 (N_20950,N_18478,N_17529);
xnor U20951 (N_20951,N_18464,N_19687);
and U20952 (N_20952,N_19540,N_18146);
xor U20953 (N_20953,N_19639,N_17530);
nor U20954 (N_20954,N_18430,N_18206);
xor U20955 (N_20955,N_18874,N_19952);
or U20956 (N_20956,N_18093,N_18156);
nand U20957 (N_20957,N_17505,N_19789);
xor U20958 (N_20958,N_17656,N_17869);
nor U20959 (N_20959,N_18957,N_18597);
xor U20960 (N_20960,N_18016,N_18619);
xnor U20961 (N_20961,N_19577,N_19601);
nor U20962 (N_20962,N_17883,N_18255);
or U20963 (N_20963,N_18271,N_19487);
and U20964 (N_20964,N_18353,N_19125);
nand U20965 (N_20965,N_18484,N_18438);
xnor U20966 (N_20966,N_17789,N_19412);
and U20967 (N_20967,N_19741,N_17618);
xor U20968 (N_20968,N_18104,N_17976);
nor U20969 (N_20969,N_19321,N_18564);
xnor U20970 (N_20970,N_19834,N_18477);
xnor U20971 (N_20971,N_17655,N_19398);
nor U20972 (N_20972,N_18053,N_17520);
or U20973 (N_20973,N_17678,N_18096);
or U20974 (N_20974,N_18682,N_19766);
and U20975 (N_20975,N_18380,N_18467);
nand U20976 (N_20976,N_19651,N_17996);
nor U20977 (N_20977,N_18055,N_17709);
or U20978 (N_20978,N_18595,N_18458);
and U20979 (N_20979,N_17631,N_18042);
or U20980 (N_20980,N_19104,N_17766);
nand U20981 (N_20981,N_19457,N_18964);
or U20982 (N_20982,N_19250,N_19393);
nand U20983 (N_20983,N_17952,N_17548);
xor U20984 (N_20984,N_17873,N_19232);
nor U20985 (N_20985,N_18061,N_19718);
nor U20986 (N_20986,N_19908,N_18101);
or U20987 (N_20987,N_17519,N_18903);
nor U20988 (N_20988,N_18552,N_18490);
or U20989 (N_20989,N_19283,N_19820);
nand U20990 (N_20990,N_17677,N_19758);
nor U20991 (N_20991,N_17783,N_19363);
or U20992 (N_20992,N_17927,N_19872);
or U20993 (N_20993,N_18975,N_17557);
nand U20994 (N_20994,N_19760,N_17748);
nand U20995 (N_20995,N_18832,N_18232);
nand U20996 (N_20996,N_19060,N_19089);
nor U20997 (N_20997,N_17741,N_19828);
or U20998 (N_20998,N_18698,N_17795);
and U20999 (N_20999,N_17998,N_18720);
xnor U21000 (N_21000,N_18282,N_19656);
xnor U21001 (N_21001,N_19688,N_18058);
xnor U21002 (N_21002,N_17938,N_18007);
nand U21003 (N_21003,N_17642,N_18602);
xnor U21004 (N_21004,N_19187,N_18170);
nand U21005 (N_21005,N_18351,N_18472);
and U21006 (N_21006,N_19655,N_18221);
or U21007 (N_21007,N_19988,N_19096);
nand U21008 (N_21008,N_19377,N_18949);
nor U21009 (N_21009,N_18158,N_19086);
nor U21010 (N_21010,N_18422,N_19249);
or U21011 (N_21011,N_18894,N_19124);
xnor U21012 (N_21012,N_18830,N_18264);
nor U21013 (N_21013,N_19028,N_18869);
nand U21014 (N_21014,N_19811,N_18062);
nand U21015 (N_21015,N_19062,N_17902);
xor U21016 (N_21016,N_18810,N_19268);
nand U21017 (N_21017,N_19493,N_19217);
nand U21018 (N_21018,N_19841,N_18195);
nand U21019 (N_21019,N_18851,N_19024);
xor U21020 (N_21020,N_17924,N_18919);
nand U21021 (N_21021,N_19914,N_17568);
and U21022 (N_21022,N_19090,N_18087);
or U21023 (N_21023,N_18213,N_18526);
nand U21024 (N_21024,N_18491,N_17698);
xnor U21025 (N_21025,N_17571,N_19127);
or U21026 (N_21026,N_18370,N_18522);
nand U21027 (N_21027,N_19122,N_18139);
nand U21028 (N_21028,N_19155,N_18497);
and U21029 (N_21029,N_18563,N_18127);
and U21030 (N_21030,N_19183,N_18589);
or U21031 (N_21031,N_19238,N_18865);
xnor U21032 (N_21032,N_19698,N_18792);
and U21033 (N_21033,N_18283,N_18670);
xor U21034 (N_21034,N_19334,N_17939);
nor U21035 (N_21035,N_17932,N_17868);
nand U21036 (N_21036,N_19762,N_19019);
nand U21037 (N_21037,N_18435,N_19544);
nand U21038 (N_21038,N_19354,N_19149);
xnor U21039 (N_21039,N_19726,N_19431);
nor U21040 (N_21040,N_17663,N_18138);
xnor U21041 (N_21041,N_18250,N_18365);
and U21042 (N_21042,N_17521,N_18928);
or U21043 (N_21043,N_17528,N_18507);
xnor U21044 (N_21044,N_17596,N_17989);
xor U21045 (N_21045,N_17885,N_18122);
xnor U21046 (N_21046,N_17674,N_19461);
nor U21047 (N_21047,N_18749,N_19797);
xor U21048 (N_21048,N_19964,N_19614);
and U21049 (N_21049,N_18173,N_19661);
xor U21050 (N_21050,N_18521,N_18622);
and U21051 (N_21051,N_19306,N_17554);
or U21052 (N_21052,N_17640,N_17691);
xnor U21053 (N_21053,N_18680,N_17704);
nor U21054 (N_21054,N_18140,N_19825);
xnor U21055 (N_21055,N_18548,N_19928);
or U21056 (N_21056,N_18281,N_19989);
nand U21057 (N_21057,N_18157,N_18922);
or U21058 (N_21058,N_19618,N_17813);
and U21059 (N_21059,N_18239,N_17599);
or U21060 (N_21060,N_18585,N_18151);
nor U21061 (N_21061,N_19029,N_18908);
or U21062 (N_21062,N_18124,N_18929);
nand U21063 (N_21063,N_19497,N_18755);
and U21064 (N_21064,N_17670,N_17531);
nor U21065 (N_21065,N_18603,N_19471);
and U21066 (N_21066,N_18190,N_19021);
or U21067 (N_21067,N_18301,N_19301);
xor U21068 (N_21068,N_18172,N_18175);
and U21069 (N_21069,N_19602,N_19017);
nand U21070 (N_21070,N_18113,N_18473);
xor U21071 (N_21071,N_19745,N_18910);
nand U21072 (N_21072,N_19855,N_17994);
or U21073 (N_21073,N_19942,N_18344);
xnor U21074 (N_21074,N_17566,N_18209);
nor U21075 (N_21075,N_19592,N_19360);
or U21076 (N_21076,N_18325,N_17540);
and U21077 (N_21077,N_18936,N_19255);
xor U21078 (N_21078,N_19712,N_17770);
xor U21079 (N_21079,N_18252,N_19339);
and U21080 (N_21080,N_18132,N_17641);
xor U21081 (N_21081,N_19129,N_17814);
nand U21082 (N_21082,N_17843,N_19937);
nor U21083 (N_21083,N_18738,N_17744);
nor U21084 (N_21084,N_19959,N_19580);
or U21085 (N_21085,N_18551,N_18777);
or U21086 (N_21086,N_19172,N_17819);
nor U21087 (N_21087,N_19725,N_18322);
or U21088 (N_21088,N_18508,N_19898);
xnor U21089 (N_21089,N_18683,N_19379);
nor U21090 (N_21090,N_17772,N_18056);
nand U21091 (N_21091,N_17567,N_19142);
nand U21092 (N_21092,N_17761,N_19750);
nor U21093 (N_21093,N_17630,N_19729);
nand U21094 (N_21094,N_18608,N_19348);
or U21095 (N_21095,N_17955,N_18088);
nor U21096 (N_21096,N_19067,N_18078);
nor U21097 (N_21097,N_17846,N_18708);
and U21098 (N_21098,N_18116,N_19900);
xor U21099 (N_21099,N_18524,N_18359);
and U21100 (N_21100,N_17835,N_19215);
xnor U21101 (N_21101,N_19349,N_18404);
nor U21102 (N_21102,N_17525,N_19312);
nor U21103 (N_21103,N_17538,N_18849);
nand U21104 (N_21104,N_19578,N_19292);
nor U21105 (N_21105,N_18873,N_18331);
nor U21106 (N_21106,N_17763,N_18082);
or U21107 (N_21107,N_17821,N_18741);
or U21108 (N_21108,N_18465,N_18185);
xor U21109 (N_21109,N_18913,N_19361);
nor U21110 (N_21110,N_19776,N_17788);
nor U21111 (N_21111,N_18692,N_17852);
nand U21112 (N_21112,N_17508,N_19167);
xnor U21113 (N_21113,N_19844,N_17500);
xnor U21114 (N_21114,N_19050,N_18891);
and U21115 (N_21115,N_19796,N_18610);
or U21116 (N_21116,N_19958,N_18635);
nand U21117 (N_21117,N_18793,N_17742);
nand U21118 (N_21118,N_17632,N_18251);
and U21119 (N_21119,N_19723,N_17848);
and U21120 (N_21120,N_17662,N_19785);
and U21121 (N_21121,N_17922,N_19302);
or U21122 (N_21122,N_19161,N_18782);
xor U21123 (N_21123,N_18000,N_18934);
nand U21124 (N_21124,N_18089,N_18897);
and U21125 (N_21125,N_18295,N_18028);
nand U21126 (N_21126,N_17864,N_19732);
nand U21127 (N_21127,N_18591,N_17682);
nor U21128 (N_21128,N_18625,N_17871);
and U21129 (N_21129,N_17504,N_18443);
xor U21130 (N_21130,N_18706,N_19068);
or U21131 (N_21131,N_17592,N_18020);
or U21132 (N_21132,N_18924,N_18872);
or U21133 (N_21133,N_17817,N_19509);
nand U21134 (N_21134,N_18076,N_17884);
and U21135 (N_21135,N_18727,N_19893);
nor U21136 (N_21136,N_18940,N_19704);
and U21137 (N_21137,N_19730,N_18592);
nor U21138 (N_21138,N_18994,N_18230);
xnor U21139 (N_21139,N_18371,N_17648);
nor U21140 (N_21140,N_17745,N_19276);
xor U21141 (N_21141,N_18019,N_19764);
or U21142 (N_21142,N_19719,N_19976);
nor U21143 (N_21143,N_18387,N_19727);
xnor U21144 (N_21144,N_18418,N_19794);
and U21145 (N_21145,N_18090,N_19229);
and U21146 (N_21146,N_19554,N_18691);
xnor U21147 (N_21147,N_19138,N_19490);
nand U21148 (N_21148,N_18831,N_18143);
or U21149 (N_21149,N_18229,N_17959);
and U21150 (N_21150,N_17854,N_19304);
or U21151 (N_21151,N_19356,N_19945);
xnor U21152 (N_21152,N_19027,N_19140);
xnor U21153 (N_21153,N_18110,N_19679);
or U21154 (N_21154,N_18379,N_18207);
nor U21155 (N_21155,N_19795,N_18991);
or U21156 (N_21156,N_18935,N_18169);
or U21157 (N_21157,N_19631,N_18678);
nand U21158 (N_21158,N_18392,N_17840);
and U21159 (N_21159,N_18676,N_18954);
nand U21160 (N_21160,N_19476,N_17875);
nor U21161 (N_21161,N_18568,N_18641);
nand U21162 (N_21162,N_19373,N_19342);
nor U21163 (N_21163,N_19705,N_19357);
xnor U21164 (N_21164,N_19895,N_17966);
xor U21165 (N_21165,N_19852,N_19695);
xnor U21166 (N_21166,N_18627,N_17929);
xor U21167 (N_21167,N_18002,N_19156);
xor U21168 (N_21168,N_18893,N_18345);
nor U21169 (N_21169,N_19274,N_18208);
and U21170 (N_21170,N_18428,N_17695);
and U21171 (N_21171,N_18666,N_18165);
nand U21172 (N_21172,N_18284,N_17702);
or U21173 (N_21173,N_19395,N_17914);
nand U21174 (N_21174,N_18103,N_17595);
or U21175 (N_21175,N_19665,N_18571);
xnor U21176 (N_21176,N_18493,N_19153);
nand U21177 (N_21177,N_19508,N_19438);
and U21178 (N_21178,N_19516,N_19331);
nand U21179 (N_21179,N_18937,N_18785);
and U21180 (N_21180,N_18447,N_19870);
and U21181 (N_21181,N_17513,N_17721);
and U21182 (N_21182,N_18648,N_18932);
or U21183 (N_21183,N_19314,N_19887);
nand U21184 (N_21184,N_18440,N_18479);
nor U21185 (N_21185,N_19523,N_19659);
or U21186 (N_21186,N_18178,N_17918);
nor U21187 (N_21187,N_19939,N_19303);
or U21188 (N_21188,N_17919,N_18237);
and U21189 (N_21189,N_18814,N_19015);
and U21190 (N_21190,N_19141,N_19405);
and U21191 (N_21191,N_19616,N_19711);
and U21192 (N_21192,N_18494,N_18550);
xnor U21193 (N_21193,N_19371,N_17862);
xnor U21194 (N_21194,N_17720,N_19064);
nor U21195 (N_21195,N_18700,N_19179);
and U21196 (N_21196,N_17993,N_19835);
nor U21197 (N_21197,N_19530,N_19164);
or U21198 (N_21198,N_18525,N_19826);
xor U21199 (N_21199,N_19114,N_18859);
nand U21200 (N_21200,N_18412,N_18750);
nand U21201 (N_21201,N_19553,N_17816);
nand U21202 (N_21202,N_19994,N_18354);
nor U21203 (N_21203,N_17733,N_17579);
nand U21204 (N_21204,N_17716,N_18860);
or U21205 (N_21205,N_19257,N_18805);
nor U21206 (N_21206,N_19763,N_17637);
xor U21207 (N_21207,N_19786,N_19358);
nor U21208 (N_21208,N_19066,N_19439);
and U21209 (N_21209,N_18267,N_18965);
or U21210 (N_21210,N_18067,N_17590);
nor U21211 (N_21211,N_18051,N_19822);
nor U21212 (N_21212,N_17861,N_19087);
and U21213 (N_21213,N_17926,N_18837);
nor U21214 (N_21214,N_18743,N_18168);
xnor U21215 (N_21215,N_19410,N_18606);
nand U21216 (N_21216,N_19815,N_18827);
and U21217 (N_21217,N_18163,N_19591);
xor U21218 (N_21218,N_19998,N_17607);
or U21219 (N_21219,N_19259,N_19703);
and U21220 (N_21220,N_18880,N_18327);
and U21221 (N_21221,N_18751,N_19313);
nand U21222 (N_21222,N_19932,N_17860);
xor U21223 (N_21223,N_18149,N_19400);
xnor U21224 (N_21224,N_17714,N_19923);
or U21225 (N_21225,N_18037,N_18614);
nor U21226 (N_21226,N_18783,N_18235);
or U21227 (N_21227,N_18995,N_18210);
nand U21228 (N_21228,N_17876,N_17739);
xnor U21229 (N_21229,N_18643,N_18694);
nand U21230 (N_21230,N_17891,N_19514);
or U21231 (N_21231,N_19305,N_18818);
nor U21232 (N_21232,N_19092,N_18626);
or U21233 (N_21233,N_18126,N_18760);
or U21234 (N_21234,N_17526,N_19459);
nor U21235 (N_21235,N_19693,N_18442);
or U21236 (N_21236,N_18596,N_18672);
nand U21237 (N_21237,N_18906,N_17726);
nand U21238 (N_21238,N_19875,N_19036);
or U21239 (N_21239,N_17703,N_18577);
nor U21240 (N_21240,N_19979,N_19881);
and U21241 (N_21241,N_17539,N_18450);
nor U21242 (N_21242,N_17706,N_18605);
or U21243 (N_21243,N_17759,N_17859);
xnor U21244 (N_21244,N_19995,N_17669);
and U21245 (N_21245,N_18696,N_18756);
or U21246 (N_21246,N_18197,N_17946);
and U21247 (N_21247,N_18186,N_19948);
nor U21248 (N_21248,N_18898,N_19701);
xnor U21249 (N_21249,N_19059,N_18520);
xor U21250 (N_21250,N_17810,N_17793);
or U21251 (N_21251,N_19417,N_18877);
nor U21252 (N_21252,N_17889,N_19191);
and U21253 (N_21253,N_17666,N_18572);
xnor U21254 (N_21254,N_19690,N_19020);
or U21255 (N_21255,N_18292,N_18907);
and U21256 (N_21256,N_19203,N_19130);
or U21257 (N_21257,N_18398,N_17766);
and U21258 (N_21258,N_18880,N_18019);
and U21259 (N_21259,N_19068,N_17836);
or U21260 (N_21260,N_17881,N_19808);
or U21261 (N_21261,N_19304,N_17699);
nand U21262 (N_21262,N_19472,N_19675);
and U21263 (N_21263,N_18065,N_17911);
xnor U21264 (N_21264,N_19961,N_19657);
or U21265 (N_21265,N_19306,N_19287);
xnor U21266 (N_21266,N_18320,N_19130);
and U21267 (N_21267,N_18567,N_19166);
and U21268 (N_21268,N_19004,N_18142);
and U21269 (N_21269,N_19483,N_17566);
nand U21270 (N_21270,N_18111,N_17732);
and U21271 (N_21271,N_19045,N_18156);
xor U21272 (N_21272,N_19339,N_17614);
or U21273 (N_21273,N_17820,N_18297);
and U21274 (N_21274,N_19165,N_19203);
or U21275 (N_21275,N_17756,N_19760);
or U21276 (N_21276,N_19136,N_19481);
or U21277 (N_21277,N_19926,N_19637);
or U21278 (N_21278,N_19728,N_19214);
xnor U21279 (N_21279,N_19452,N_17910);
nor U21280 (N_21280,N_19107,N_19678);
nand U21281 (N_21281,N_19171,N_19153);
nand U21282 (N_21282,N_19100,N_18033);
or U21283 (N_21283,N_19810,N_17558);
or U21284 (N_21284,N_18906,N_18442);
xnor U21285 (N_21285,N_18989,N_18048);
xnor U21286 (N_21286,N_19045,N_19068);
xnor U21287 (N_21287,N_19226,N_18242);
nor U21288 (N_21288,N_17609,N_17608);
xnor U21289 (N_21289,N_18489,N_18536);
or U21290 (N_21290,N_19222,N_19143);
nand U21291 (N_21291,N_19153,N_17629);
or U21292 (N_21292,N_18706,N_18389);
nor U21293 (N_21293,N_18019,N_19073);
xnor U21294 (N_21294,N_18675,N_19604);
nor U21295 (N_21295,N_17547,N_17521);
xnor U21296 (N_21296,N_18866,N_19053);
nor U21297 (N_21297,N_17588,N_17651);
nor U21298 (N_21298,N_19544,N_17799);
xnor U21299 (N_21299,N_17644,N_17729);
and U21300 (N_21300,N_18202,N_18432);
xnor U21301 (N_21301,N_18995,N_17642);
nand U21302 (N_21302,N_17595,N_18390);
xnor U21303 (N_21303,N_18677,N_19850);
nor U21304 (N_21304,N_19850,N_18446);
or U21305 (N_21305,N_18392,N_18877);
or U21306 (N_21306,N_17843,N_19417);
and U21307 (N_21307,N_17680,N_19081);
nor U21308 (N_21308,N_18336,N_18233);
nor U21309 (N_21309,N_18606,N_17653);
nor U21310 (N_21310,N_18185,N_17811);
nand U21311 (N_21311,N_19133,N_19094);
or U21312 (N_21312,N_17632,N_17711);
xor U21313 (N_21313,N_18617,N_17909);
nand U21314 (N_21314,N_18183,N_19929);
xnor U21315 (N_21315,N_19190,N_17540);
nor U21316 (N_21316,N_19788,N_19500);
nand U21317 (N_21317,N_18530,N_17640);
nor U21318 (N_21318,N_18058,N_18410);
and U21319 (N_21319,N_17560,N_19371);
and U21320 (N_21320,N_19078,N_18561);
nand U21321 (N_21321,N_18551,N_18909);
nor U21322 (N_21322,N_19255,N_18948);
nand U21323 (N_21323,N_19690,N_18223);
and U21324 (N_21324,N_18346,N_19456);
and U21325 (N_21325,N_18260,N_18727);
and U21326 (N_21326,N_17535,N_19716);
xor U21327 (N_21327,N_18750,N_19858);
nand U21328 (N_21328,N_19976,N_18342);
and U21329 (N_21329,N_19239,N_17831);
nand U21330 (N_21330,N_17550,N_18986);
and U21331 (N_21331,N_19634,N_19734);
and U21332 (N_21332,N_19330,N_19976);
xor U21333 (N_21333,N_19659,N_19386);
and U21334 (N_21334,N_18450,N_19766);
xor U21335 (N_21335,N_19695,N_18391);
or U21336 (N_21336,N_19492,N_18485);
xor U21337 (N_21337,N_19574,N_18047);
or U21338 (N_21338,N_19000,N_17825);
or U21339 (N_21339,N_18743,N_17684);
or U21340 (N_21340,N_19390,N_18048);
nand U21341 (N_21341,N_19419,N_17582);
or U21342 (N_21342,N_17622,N_19467);
or U21343 (N_21343,N_18892,N_18604);
nand U21344 (N_21344,N_18259,N_17683);
nand U21345 (N_21345,N_19771,N_17691);
nand U21346 (N_21346,N_18623,N_19497);
or U21347 (N_21347,N_19106,N_18604);
and U21348 (N_21348,N_19671,N_19071);
and U21349 (N_21349,N_18660,N_18890);
xor U21350 (N_21350,N_18894,N_19295);
or U21351 (N_21351,N_19149,N_18661);
nand U21352 (N_21352,N_17873,N_18560);
nand U21353 (N_21353,N_18393,N_18209);
nand U21354 (N_21354,N_18440,N_19916);
nor U21355 (N_21355,N_19508,N_19860);
nand U21356 (N_21356,N_18580,N_19375);
or U21357 (N_21357,N_19292,N_18054);
or U21358 (N_21358,N_17701,N_18158);
and U21359 (N_21359,N_18763,N_19340);
xor U21360 (N_21360,N_19896,N_19027);
and U21361 (N_21361,N_18391,N_17570);
or U21362 (N_21362,N_17521,N_19289);
nor U21363 (N_21363,N_19891,N_17848);
nor U21364 (N_21364,N_19307,N_18448);
nand U21365 (N_21365,N_18119,N_18336);
or U21366 (N_21366,N_18324,N_19808);
and U21367 (N_21367,N_18834,N_19474);
or U21368 (N_21368,N_18605,N_19137);
nand U21369 (N_21369,N_18542,N_19212);
or U21370 (N_21370,N_18770,N_18191);
nand U21371 (N_21371,N_19134,N_18117);
and U21372 (N_21372,N_18307,N_18247);
or U21373 (N_21373,N_18485,N_19962);
or U21374 (N_21374,N_18115,N_17547);
nor U21375 (N_21375,N_18777,N_18682);
and U21376 (N_21376,N_18601,N_18148);
or U21377 (N_21377,N_18403,N_18321);
and U21378 (N_21378,N_18027,N_17939);
nor U21379 (N_21379,N_19307,N_18238);
nor U21380 (N_21380,N_17841,N_19691);
or U21381 (N_21381,N_18729,N_17634);
nor U21382 (N_21382,N_19258,N_19163);
xor U21383 (N_21383,N_19615,N_19282);
nor U21384 (N_21384,N_18249,N_18481);
and U21385 (N_21385,N_17638,N_17528);
nor U21386 (N_21386,N_19987,N_19696);
or U21387 (N_21387,N_19796,N_18009);
and U21388 (N_21388,N_17688,N_19209);
or U21389 (N_21389,N_17815,N_18457);
and U21390 (N_21390,N_17513,N_19094);
and U21391 (N_21391,N_18426,N_17771);
nand U21392 (N_21392,N_18523,N_19235);
nor U21393 (N_21393,N_18331,N_18040);
xnor U21394 (N_21394,N_18628,N_19970);
or U21395 (N_21395,N_19712,N_19249);
or U21396 (N_21396,N_19905,N_18099);
nor U21397 (N_21397,N_19680,N_19193);
and U21398 (N_21398,N_18916,N_19543);
nand U21399 (N_21399,N_17988,N_18090);
and U21400 (N_21400,N_18676,N_19448);
and U21401 (N_21401,N_18163,N_18908);
xnor U21402 (N_21402,N_18655,N_17835);
nor U21403 (N_21403,N_19814,N_18063);
and U21404 (N_21404,N_19990,N_18967);
nand U21405 (N_21405,N_18930,N_19046);
nor U21406 (N_21406,N_19598,N_18705);
and U21407 (N_21407,N_18955,N_18292);
xnor U21408 (N_21408,N_18064,N_18422);
nor U21409 (N_21409,N_17774,N_18890);
and U21410 (N_21410,N_18492,N_17712);
and U21411 (N_21411,N_17842,N_19805);
xor U21412 (N_21412,N_17790,N_18127);
and U21413 (N_21413,N_19352,N_18683);
nor U21414 (N_21414,N_18735,N_19154);
and U21415 (N_21415,N_18684,N_17975);
nor U21416 (N_21416,N_19536,N_19349);
xor U21417 (N_21417,N_18192,N_18789);
xor U21418 (N_21418,N_19503,N_17835);
nor U21419 (N_21419,N_19332,N_19092);
or U21420 (N_21420,N_19700,N_19915);
or U21421 (N_21421,N_19354,N_17795);
nand U21422 (N_21422,N_19082,N_18450);
nor U21423 (N_21423,N_19567,N_19782);
nand U21424 (N_21424,N_18308,N_17684);
nand U21425 (N_21425,N_19427,N_18209);
nor U21426 (N_21426,N_18968,N_17902);
nor U21427 (N_21427,N_18736,N_18014);
and U21428 (N_21428,N_18931,N_19728);
nand U21429 (N_21429,N_17707,N_19332);
nor U21430 (N_21430,N_18807,N_17675);
or U21431 (N_21431,N_18594,N_19835);
nand U21432 (N_21432,N_18766,N_17848);
or U21433 (N_21433,N_19415,N_18794);
nor U21434 (N_21434,N_18405,N_18531);
xor U21435 (N_21435,N_19109,N_17690);
xnor U21436 (N_21436,N_18554,N_19854);
xnor U21437 (N_21437,N_19744,N_17950);
or U21438 (N_21438,N_19772,N_18671);
and U21439 (N_21439,N_18438,N_19183);
nor U21440 (N_21440,N_17976,N_17975);
xnor U21441 (N_21441,N_18259,N_18728);
xor U21442 (N_21442,N_18589,N_18290);
nand U21443 (N_21443,N_19929,N_19741);
or U21444 (N_21444,N_19877,N_17612);
xnor U21445 (N_21445,N_18242,N_17503);
or U21446 (N_21446,N_18062,N_19744);
nor U21447 (N_21447,N_18251,N_18970);
nor U21448 (N_21448,N_17811,N_17781);
xor U21449 (N_21449,N_18730,N_18621);
and U21450 (N_21450,N_19111,N_18856);
nand U21451 (N_21451,N_19124,N_19056);
xor U21452 (N_21452,N_19290,N_19364);
or U21453 (N_21453,N_18671,N_19753);
xnor U21454 (N_21454,N_18545,N_19682);
and U21455 (N_21455,N_18735,N_19481);
and U21456 (N_21456,N_19729,N_19858);
nor U21457 (N_21457,N_17645,N_17524);
nor U21458 (N_21458,N_18790,N_18973);
or U21459 (N_21459,N_19788,N_17937);
and U21460 (N_21460,N_18996,N_18758);
and U21461 (N_21461,N_19586,N_19923);
nand U21462 (N_21462,N_18849,N_19173);
xnor U21463 (N_21463,N_18339,N_18365);
nor U21464 (N_21464,N_19200,N_19210);
nand U21465 (N_21465,N_17707,N_18833);
nor U21466 (N_21466,N_18895,N_19347);
nand U21467 (N_21467,N_19850,N_19920);
and U21468 (N_21468,N_19116,N_19230);
nand U21469 (N_21469,N_19592,N_17668);
nor U21470 (N_21470,N_18023,N_19615);
and U21471 (N_21471,N_18529,N_18208);
xnor U21472 (N_21472,N_18098,N_18060);
nand U21473 (N_21473,N_19386,N_18499);
and U21474 (N_21474,N_19095,N_19485);
or U21475 (N_21475,N_17933,N_18594);
nor U21476 (N_21476,N_18596,N_18739);
nand U21477 (N_21477,N_18297,N_17670);
and U21478 (N_21478,N_19346,N_18382);
xnor U21479 (N_21479,N_19018,N_18259);
nand U21480 (N_21480,N_19605,N_19576);
or U21481 (N_21481,N_18731,N_17868);
xor U21482 (N_21482,N_19023,N_18994);
and U21483 (N_21483,N_19075,N_18023);
nand U21484 (N_21484,N_19774,N_19876);
xnor U21485 (N_21485,N_19879,N_18322);
or U21486 (N_21486,N_18509,N_18919);
xnor U21487 (N_21487,N_19093,N_19553);
or U21488 (N_21488,N_19891,N_19818);
nor U21489 (N_21489,N_19212,N_17875);
nand U21490 (N_21490,N_19508,N_18958);
nor U21491 (N_21491,N_19263,N_19410);
nand U21492 (N_21492,N_18841,N_17889);
xnor U21493 (N_21493,N_19416,N_19676);
nand U21494 (N_21494,N_19840,N_19734);
xor U21495 (N_21495,N_17768,N_19774);
nor U21496 (N_21496,N_18142,N_19894);
nor U21497 (N_21497,N_19919,N_19324);
nor U21498 (N_21498,N_19388,N_19010);
xnor U21499 (N_21499,N_17677,N_19572);
and U21500 (N_21500,N_18569,N_17941);
nor U21501 (N_21501,N_19332,N_19820);
or U21502 (N_21502,N_17768,N_19028);
nand U21503 (N_21503,N_19857,N_19072);
and U21504 (N_21504,N_19204,N_17754);
xor U21505 (N_21505,N_17615,N_18748);
and U21506 (N_21506,N_17912,N_18272);
xnor U21507 (N_21507,N_19512,N_17728);
or U21508 (N_21508,N_18128,N_19235);
nor U21509 (N_21509,N_18650,N_18024);
or U21510 (N_21510,N_19262,N_18210);
nor U21511 (N_21511,N_19208,N_18584);
nand U21512 (N_21512,N_19629,N_18541);
or U21513 (N_21513,N_18963,N_19444);
and U21514 (N_21514,N_18297,N_19855);
or U21515 (N_21515,N_19759,N_19048);
nor U21516 (N_21516,N_19556,N_18988);
nor U21517 (N_21517,N_19507,N_18576);
or U21518 (N_21518,N_19442,N_19740);
nor U21519 (N_21519,N_18072,N_19246);
nand U21520 (N_21520,N_18493,N_19400);
xor U21521 (N_21521,N_18283,N_19651);
nor U21522 (N_21522,N_18067,N_19663);
or U21523 (N_21523,N_17706,N_18594);
nor U21524 (N_21524,N_18623,N_18829);
nand U21525 (N_21525,N_18514,N_18090);
or U21526 (N_21526,N_18522,N_18226);
and U21527 (N_21527,N_19933,N_19878);
or U21528 (N_21528,N_17606,N_17730);
or U21529 (N_21529,N_19664,N_19197);
nor U21530 (N_21530,N_17787,N_18210);
and U21531 (N_21531,N_18344,N_18017);
xnor U21532 (N_21532,N_17513,N_19237);
nand U21533 (N_21533,N_18742,N_17559);
xor U21534 (N_21534,N_17911,N_17671);
and U21535 (N_21535,N_18106,N_18471);
or U21536 (N_21536,N_18777,N_19578);
nor U21537 (N_21537,N_17824,N_19482);
or U21538 (N_21538,N_18960,N_18930);
xnor U21539 (N_21539,N_18289,N_19930);
and U21540 (N_21540,N_19897,N_19574);
and U21541 (N_21541,N_17546,N_18373);
or U21542 (N_21542,N_18639,N_18363);
xor U21543 (N_21543,N_18679,N_17800);
nand U21544 (N_21544,N_18876,N_17716);
nor U21545 (N_21545,N_19785,N_19673);
and U21546 (N_21546,N_18933,N_19161);
or U21547 (N_21547,N_19801,N_18251);
xor U21548 (N_21548,N_18707,N_19301);
or U21549 (N_21549,N_18149,N_19421);
and U21550 (N_21550,N_19450,N_19882);
xor U21551 (N_21551,N_17697,N_18668);
and U21552 (N_21552,N_18519,N_18488);
or U21553 (N_21553,N_19535,N_18541);
nor U21554 (N_21554,N_19706,N_18379);
xor U21555 (N_21555,N_19892,N_17718);
nand U21556 (N_21556,N_19846,N_18436);
or U21557 (N_21557,N_19609,N_19918);
nor U21558 (N_21558,N_18987,N_19171);
and U21559 (N_21559,N_18540,N_18672);
or U21560 (N_21560,N_17693,N_19698);
nor U21561 (N_21561,N_19768,N_19099);
or U21562 (N_21562,N_18094,N_17732);
nor U21563 (N_21563,N_17581,N_17896);
and U21564 (N_21564,N_19116,N_18373);
and U21565 (N_21565,N_18735,N_17645);
and U21566 (N_21566,N_19989,N_18103);
or U21567 (N_21567,N_18320,N_19032);
xor U21568 (N_21568,N_18471,N_18059);
and U21569 (N_21569,N_18758,N_17589);
xor U21570 (N_21570,N_18539,N_19009);
or U21571 (N_21571,N_17578,N_19389);
nand U21572 (N_21572,N_19633,N_19544);
nand U21573 (N_21573,N_17708,N_17733);
and U21574 (N_21574,N_18427,N_19525);
nand U21575 (N_21575,N_19963,N_19789);
and U21576 (N_21576,N_19160,N_18594);
nor U21577 (N_21577,N_17736,N_19257);
nand U21578 (N_21578,N_18606,N_18531);
or U21579 (N_21579,N_18440,N_19299);
nand U21580 (N_21580,N_18489,N_18530);
or U21581 (N_21581,N_18147,N_18221);
or U21582 (N_21582,N_19001,N_17564);
nor U21583 (N_21583,N_18898,N_19161);
and U21584 (N_21584,N_19072,N_19303);
or U21585 (N_21585,N_17898,N_19025);
nor U21586 (N_21586,N_19348,N_19874);
nor U21587 (N_21587,N_17740,N_18815);
nor U21588 (N_21588,N_18878,N_19377);
nand U21589 (N_21589,N_18945,N_19629);
and U21590 (N_21590,N_17788,N_18249);
xor U21591 (N_21591,N_18898,N_18084);
and U21592 (N_21592,N_19607,N_18126);
nand U21593 (N_21593,N_18292,N_17964);
xnor U21594 (N_21594,N_19768,N_19538);
nor U21595 (N_21595,N_18792,N_19911);
nand U21596 (N_21596,N_18975,N_19997);
nand U21597 (N_21597,N_18384,N_18540);
xor U21598 (N_21598,N_17840,N_19442);
nand U21599 (N_21599,N_17715,N_18144);
and U21600 (N_21600,N_17843,N_19814);
nand U21601 (N_21601,N_18196,N_18962);
nand U21602 (N_21602,N_19602,N_18716);
and U21603 (N_21603,N_18926,N_18511);
nor U21604 (N_21604,N_18650,N_18437);
or U21605 (N_21605,N_17550,N_18720);
and U21606 (N_21606,N_18649,N_18439);
nor U21607 (N_21607,N_19119,N_17832);
xnor U21608 (N_21608,N_18695,N_19080);
or U21609 (N_21609,N_18339,N_17944);
xor U21610 (N_21610,N_17541,N_19304);
and U21611 (N_21611,N_17940,N_19901);
xor U21612 (N_21612,N_18428,N_18650);
xnor U21613 (N_21613,N_18615,N_18745);
nor U21614 (N_21614,N_19893,N_19766);
nand U21615 (N_21615,N_17553,N_19654);
and U21616 (N_21616,N_18885,N_19386);
and U21617 (N_21617,N_17764,N_18156);
xor U21618 (N_21618,N_19983,N_18184);
xor U21619 (N_21619,N_17640,N_18544);
nand U21620 (N_21620,N_18207,N_19333);
nand U21621 (N_21621,N_19449,N_18465);
and U21622 (N_21622,N_17691,N_19905);
xnor U21623 (N_21623,N_18445,N_19761);
nor U21624 (N_21624,N_18341,N_19913);
nand U21625 (N_21625,N_19172,N_19361);
xnor U21626 (N_21626,N_18922,N_18409);
and U21627 (N_21627,N_18994,N_19391);
nor U21628 (N_21628,N_19964,N_18279);
and U21629 (N_21629,N_18708,N_18774);
or U21630 (N_21630,N_18179,N_17518);
nor U21631 (N_21631,N_19725,N_19709);
or U21632 (N_21632,N_19054,N_18947);
and U21633 (N_21633,N_17885,N_18860);
or U21634 (N_21634,N_18208,N_18353);
or U21635 (N_21635,N_18847,N_17975);
xor U21636 (N_21636,N_19755,N_18763);
xor U21637 (N_21637,N_17872,N_17593);
nor U21638 (N_21638,N_19825,N_17741);
nand U21639 (N_21639,N_18648,N_18999);
and U21640 (N_21640,N_19127,N_19865);
nand U21641 (N_21641,N_19880,N_18414);
xor U21642 (N_21642,N_18480,N_17844);
or U21643 (N_21643,N_18558,N_18022);
xnor U21644 (N_21644,N_19959,N_18867);
xnor U21645 (N_21645,N_19567,N_19296);
nor U21646 (N_21646,N_18911,N_18377);
nor U21647 (N_21647,N_17593,N_19651);
xnor U21648 (N_21648,N_18652,N_19318);
and U21649 (N_21649,N_17784,N_19046);
nor U21650 (N_21650,N_18275,N_17989);
or U21651 (N_21651,N_19504,N_17881);
xor U21652 (N_21652,N_18847,N_19088);
nand U21653 (N_21653,N_19921,N_18697);
and U21654 (N_21654,N_19761,N_19060);
nand U21655 (N_21655,N_18055,N_18184);
or U21656 (N_21656,N_18717,N_18316);
xor U21657 (N_21657,N_18498,N_18293);
nand U21658 (N_21658,N_18719,N_19618);
or U21659 (N_21659,N_18146,N_18687);
xnor U21660 (N_21660,N_19438,N_17969);
or U21661 (N_21661,N_19378,N_19349);
nand U21662 (N_21662,N_18580,N_19061);
xor U21663 (N_21663,N_19959,N_19139);
nor U21664 (N_21664,N_17639,N_19703);
or U21665 (N_21665,N_18022,N_18959);
xnor U21666 (N_21666,N_17831,N_19600);
xnor U21667 (N_21667,N_17595,N_19013);
or U21668 (N_21668,N_18826,N_17790);
or U21669 (N_21669,N_17877,N_18415);
and U21670 (N_21670,N_19780,N_18594);
nor U21671 (N_21671,N_19306,N_18967);
or U21672 (N_21672,N_17901,N_18638);
xnor U21673 (N_21673,N_18053,N_19672);
or U21674 (N_21674,N_19269,N_19589);
nand U21675 (N_21675,N_19997,N_18458);
xor U21676 (N_21676,N_19847,N_19757);
xor U21677 (N_21677,N_19486,N_18712);
nand U21678 (N_21678,N_19011,N_19335);
or U21679 (N_21679,N_18254,N_18595);
and U21680 (N_21680,N_18799,N_19822);
or U21681 (N_21681,N_18252,N_17797);
and U21682 (N_21682,N_19178,N_17880);
nand U21683 (N_21683,N_18995,N_18744);
and U21684 (N_21684,N_18001,N_18036);
nor U21685 (N_21685,N_17715,N_17925);
nor U21686 (N_21686,N_17644,N_18101);
nor U21687 (N_21687,N_19389,N_17505);
or U21688 (N_21688,N_18847,N_18143);
or U21689 (N_21689,N_18187,N_19388);
or U21690 (N_21690,N_18195,N_18828);
nor U21691 (N_21691,N_18386,N_18342);
or U21692 (N_21692,N_18530,N_18364);
nand U21693 (N_21693,N_19242,N_18288);
nand U21694 (N_21694,N_19141,N_17734);
xor U21695 (N_21695,N_17947,N_19403);
or U21696 (N_21696,N_18528,N_18186);
xnor U21697 (N_21697,N_18413,N_19257);
and U21698 (N_21698,N_19313,N_18495);
or U21699 (N_21699,N_17878,N_18260);
xor U21700 (N_21700,N_18589,N_17982);
nand U21701 (N_21701,N_18026,N_18506);
nor U21702 (N_21702,N_19060,N_19795);
nor U21703 (N_21703,N_17678,N_17694);
and U21704 (N_21704,N_18165,N_17574);
nand U21705 (N_21705,N_17823,N_19733);
xnor U21706 (N_21706,N_17956,N_18001);
xor U21707 (N_21707,N_19844,N_18457);
nor U21708 (N_21708,N_18946,N_17593);
nor U21709 (N_21709,N_19938,N_19581);
and U21710 (N_21710,N_17921,N_18605);
xnor U21711 (N_21711,N_19565,N_18615);
or U21712 (N_21712,N_19974,N_18871);
nand U21713 (N_21713,N_19373,N_18284);
nor U21714 (N_21714,N_19512,N_19101);
nand U21715 (N_21715,N_19319,N_18170);
and U21716 (N_21716,N_18446,N_19884);
xor U21717 (N_21717,N_19433,N_19171);
xor U21718 (N_21718,N_18601,N_18670);
nor U21719 (N_21719,N_18194,N_18761);
nor U21720 (N_21720,N_18021,N_17822);
xor U21721 (N_21721,N_18835,N_18176);
nand U21722 (N_21722,N_18977,N_18834);
or U21723 (N_21723,N_19076,N_19454);
nand U21724 (N_21724,N_19664,N_18611);
or U21725 (N_21725,N_19127,N_17899);
or U21726 (N_21726,N_19738,N_18175);
or U21727 (N_21727,N_18516,N_19527);
and U21728 (N_21728,N_18352,N_19079);
or U21729 (N_21729,N_17790,N_18070);
or U21730 (N_21730,N_19723,N_19828);
nand U21731 (N_21731,N_19728,N_18918);
nor U21732 (N_21732,N_17695,N_19700);
nand U21733 (N_21733,N_17827,N_19086);
and U21734 (N_21734,N_19619,N_18486);
xnor U21735 (N_21735,N_18418,N_19018);
xnor U21736 (N_21736,N_19673,N_17836);
or U21737 (N_21737,N_19702,N_19810);
nand U21738 (N_21738,N_18148,N_17733);
nor U21739 (N_21739,N_19167,N_18526);
nor U21740 (N_21740,N_19965,N_19814);
xor U21741 (N_21741,N_18794,N_18089);
xor U21742 (N_21742,N_17643,N_18717);
and U21743 (N_21743,N_18621,N_18122);
nor U21744 (N_21744,N_19759,N_18695);
and U21745 (N_21745,N_18657,N_19411);
nand U21746 (N_21746,N_19034,N_17755);
nand U21747 (N_21747,N_19054,N_19830);
xnor U21748 (N_21748,N_17999,N_19003);
nand U21749 (N_21749,N_18337,N_19068);
and U21750 (N_21750,N_19534,N_19021);
nor U21751 (N_21751,N_19709,N_19658);
nor U21752 (N_21752,N_19969,N_18432);
nand U21753 (N_21753,N_19265,N_19950);
nor U21754 (N_21754,N_17540,N_19330);
nor U21755 (N_21755,N_19549,N_17565);
xnor U21756 (N_21756,N_17869,N_19272);
nand U21757 (N_21757,N_18534,N_19389);
nand U21758 (N_21758,N_18116,N_18768);
nand U21759 (N_21759,N_19755,N_18138);
nand U21760 (N_21760,N_18835,N_19403);
and U21761 (N_21761,N_18536,N_17798);
and U21762 (N_21762,N_18409,N_19709);
nand U21763 (N_21763,N_18391,N_18628);
and U21764 (N_21764,N_17913,N_17544);
nand U21765 (N_21765,N_19842,N_17634);
xor U21766 (N_21766,N_17605,N_17679);
nand U21767 (N_21767,N_18048,N_18506);
and U21768 (N_21768,N_17572,N_19550);
xnor U21769 (N_21769,N_19549,N_18507);
and U21770 (N_21770,N_18409,N_19165);
xnor U21771 (N_21771,N_18151,N_18459);
and U21772 (N_21772,N_18492,N_19366);
nor U21773 (N_21773,N_18841,N_17703);
xnor U21774 (N_21774,N_18179,N_19883);
or U21775 (N_21775,N_17671,N_19336);
or U21776 (N_21776,N_19260,N_18904);
xnor U21777 (N_21777,N_18671,N_17696);
or U21778 (N_21778,N_17958,N_17674);
xor U21779 (N_21779,N_18645,N_18399);
nand U21780 (N_21780,N_18210,N_19757);
nand U21781 (N_21781,N_19490,N_18169);
and U21782 (N_21782,N_18587,N_18541);
xor U21783 (N_21783,N_18915,N_19143);
nor U21784 (N_21784,N_19745,N_18125);
or U21785 (N_21785,N_19761,N_19677);
and U21786 (N_21786,N_19456,N_18787);
xor U21787 (N_21787,N_17669,N_19520);
xor U21788 (N_21788,N_19454,N_19474);
or U21789 (N_21789,N_17603,N_18267);
nor U21790 (N_21790,N_17722,N_18407);
nor U21791 (N_21791,N_18685,N_18185);
nand U21792 (N_21792,N_19659,N_18808);
xnor U21793 (N_21793,N_18825,N_18097);
xor U21794 (N_21794,N_17597,N_19468);
nand U21795 (N_21795,N_18575,N_18122);
or U21796 (N_21796,N_18069,N_17928);
nor U21797 (N_21797,N_19194,N_17806);
or U21798 (N_21798,N_18062,N_19399);
nand U21799 (N_21799,N_19379,N_17511);
nand U21800 (N_21800,N_19022,N_18312);
and U21801 (N_21801,N_18799,N_19740);
xnor U21802 (N_21802,N_19210,N_19273);
nand U21803 (N_21803,N_18800,N_19051);
and U21804 (N_21804,N_18138,N_19358);
nand U21805 (N_21805,N_17931,N_18403);
and U21806 (N_21806,N_19171,N_17586);
nor U21807 (N_21807,N_18218,N_18561);
and U21808 (N_21808,N_19726,N_19108);
xor U21809 (N_21809,N_18443,N_18448);
nor U21810 (N_21810,N_19656,N_18356);
and U21811 (N_21811,N_19339,N_19083);
xnor U21812 (N_21812,N_18764,N_18437);
xor U21813 (N_21813,N_18635,N_19959);
nor U21814 (N_21814,N_17764,N_19775);
nor U21815 (N_21815,N_19955,N_18164);
nand U21816 (N_21816,N_18918,N_18904);
or U21817 (N_21817,N_18431,N_18270);
nand U21818 (N_21818,N_18961,N_19014);
and U21819 (N_21819,N_17970,N_18231);
nor U21820 (N_21820,N_18877,N_18041);
or U21821 (N_21821,N_19749,N_19940);
and U21822 (N_21822,N_17709,N_19464);
and U21823 (N_21823,N_18727,N_18263);
or U21824 (N_21824,N_18217,N_18571);
nand U21825 (N_21825,N_17636,N_19826);
and U21826 (N_21826,N_19895,N_19419);
and U21827 (N_21827,N_19036,N_19821);
xor U21828 (N_21828,N_19441,N_18118);
nand U21829 (N_21829,N_18874,N_18802);
xor U21830 (N_21830,N_18071,N_19008);
and U21831 (N_21831,N_18829,N_19458);
or U21832 (N_21832,N_19959,N_19650);
nor U21833 (N_21833,N_19069,N_17685);
xnor U21834 (N_21834,N_18900,N_19853);
xnor U21835 (N_21835,N_19193,N_17847);
nand U21836 (N_21836,N_19233,N_18623);
nand U21837 (N_21837,N_18452,N_19762);
or U21838 (N_21838,N_17872,N_18525);
nor U21839 (N_21839,N_17621,N_19973);
nand U21840 (N_21840,N_18035,N_19230);
nor U21841 (N_21841,N_19168,N_19420);
nand U21842 (N_21842,N_19741,N_18655);
xnor U21843 (N_21843,N_18769,N_19512);
nand U21844 (N_21844,N_18315,N_19273);
and U21845 (N_21845,N_19979,N_18451);
nand U21846 (N_21846,N_18482,N_17633);
or U21847 (N_21847,N_17541,N_18913);
xor U21848 (N_21848,N_19926,N_19984);
nand U21849 (N_21849,N_19245,N_18313);
nand U21850 (N_21850,N_19252,N_18212);
nand U21851 (N_21851,N_17581,N_18058);
nor U21852 (N_21852,N_19200,N_18119);
and U21853 (N_21853,N_18128,N_19565);
nor U21854 (N_21854,N_18509,N_19398);
xnor U21855 (N_21855,N_19497,N_19826);
or U21856 (N_21856,N_19175,N_19031);
and U21857 (N_21857,N_19251,N_19358);
nor U21858 (N_21858,N_17770,N_18295);
xor U21859 (N_21859,N_18295,N_19078);
xor U21860 (N_21860,N_17702,N_19956);
xnor U21861 (N_21861,N_17659,N_18903);
and U21862 (N_21862,N_19017,N_18801);
or U21863 (N_21863,N_18954,N_19195);
and U21864 (N_21864,N_18256,N_18473);
and U21865 (N_21865,N_19528,N_19869);
nand U21866 (N_21866,N_18905,N_17556);
nand U21867 (N_21867,N_18128,N_18871);
xnor U21868 (N_21868,N_18650,N_19685);
xor U21869 (N_21869,N_17617,N_17972);
or U21870 (N_21870,N_18275,N_19918);
xnor U21871 (N_21871,N_19995,N_19622);
or U21872 (N_21872,N_18563,N_18144);
nor U21873 (N_21873,N_18894,N_18547);
and U21874 (N_21874,N_19617,N_19017);
xor U21875 (N_21875,N_19543,N_18024);
nor U21876 (N_21876,N_19286,N_18892);
xnor U21877 (N_21877,N_17734,N_19297);
and U21878 (N_21878,N_19363,N_18725);
xor U21879 (N_21879,N_19060,N_19818);
and U21880 (N_21880,N_17636,N_18992);
nand U21881 (N_21881,N_18231,N_19008);
nor U21882 (N_21882,N_19336,N_18937);
and U21883 (N_21883,N_17803,N_18609);
or U21884 (N_21884,N_17780,N_17886);
or U21885 (N_21885,N_19775,N_19219);
xnor U21886 (N_21886,N_17960,N_19661);
nor U21887 (N_21887,N_19666,N_18281);
or U21888 (N_21888,N_19862,N_19953);
xor U21889 (N_21889,N_19959,N_19288);
nand U21890 (N_21890,N_18035,N_17694);
nand U21891 (N_21891,N_18005,N_18275);
and U21892 (N_21892,N_19652,N_17755);
nor U21893 (N_21893,N_19997,N_17670);
xor U21894 (N_21894,N_17543,N_19940);
and U21895 (N_21895,N_19975,N_17701);
or U21896 (N_21896,N_19374,N_18974);
nor U21897 (N_21897,N_18101,N_19666);
nor U21898 (N_21898,N_17771,N_17977);
or U21899 (N_21899,N_19487,N_18384);
nor U21900 (N_21900,N_19558,N_19873);
or U21901 (N_21901,N_19994,N_19609);
or U21902 (N_21902,N_19971,N_18531);
xnor U21903 (N_21903,N_17995,N_18797);
nand U21904 (N_21904,N_19895,N_18100);
xnor U21905 (N_21905,N_18278,N_18448);
nor U21906 (N_21906,N_18345,N_18450);
nand U21907 (N_21907,N_18654,N_17889);
xnor U21908 (N_21908,N_19443,N_19220);
xor U21909 (N_21909,N_18422,N_17685);
nor U21910 (N_21910,N_19948,N_19820);
xnor U21911 (N_21911,N_18485,N_17990);
xor U21912 (N_21912,N_18035,N_18421);
xor U21913 (N_21913,N_19087,N_18889);
or U21914 (N_21914,N_18182,N_19178);
xor U21915 (N_21915,N_19769,N_19798);
and U21916 (N_21916,N_19324,N_18866);
xnor U21917 (N_21917,N_18594,N_18896);
and U21918 (N_21918,N_18737,N_19301);
nand U21919 (N_21919,N_17926,N_19908);
xor U21920 (N_21920,N_18465,N_17903);
nor U21921 (N_21921,N_19893,N_19044);
or U21922 (N_21922,N_18036,N_19072);
nand U21923 (N_21923,N_18614,N_19902);
nor U21924 (N_21924,N_18804,N_19547);
or U21925 (N_21925,N_18691,N_17735);
xor U21926 (N_21926,N_18002,N_19340);
nor U21927 (N_21927,N_18942,N_18807);
nor U21928 (N_21928,N_19470,N_18397);
xor U21929 (N_21929,N_19336,N_17736);
or U21930 (N_21930,N_18853,N_19711);
nor U21931 (N_21931,N_19815,N_17629);
nor U21932 (N_21932,N_19453,N_19092);
nand U21933 (N_21933,N_19662,N_18385);
nor U21934 (N_21934,N_19962,N_18004);
and U21935 (N_21935,N_19586,N_19618);
nor U21936 (N_21936,N_19121,N_19520);
xor U21937 (N_21937,N_19047,N_19285);
and U21938 (N_21938,N_17532,N_19732);
nor U21939 (N_21939,N_18698,N_19743);
or U21940 (N_21940,N_17898,N_18401);
nor U21941 (N_21941,N_17798,N_18342);
nor U21942 (N_21942,N_19088,N_19906);
nor U21943 (N_21943,N_19999,N_19153);
nor U21944 (N_21944,N_17903,N_18978);
xnor U21945 (N_21945,N_19022,N_18829);
or U21946 (N_21946,N_19162,N_18081);
or U21947 (N_21947,N_19686,N_18582);
or U21948 (N_21948,N_17758,N_17674);
xor U21949 (N_21949,N_18927,N_19158);
xnor U21950 (N_21950,N_17875,N_17829);
nor U21951 (N_21951,N_19338,N_17940);
xnor U21952 (N_21952,N_18657,N_18840);
nor U21953 (N_21953,N_17739,N_17874);
nor U21954 (N_21954,N_17784,N_18537);
nor U21955 (N_21955,N_18084,N_19106);
nor U21956 (N_21956,N_18504,N_18680);
nand U21957 (N_21957,N_17733,N_18572);
nand U21958 (N_21958,N_17662,N_19329);
nand U21959 (N_21959,N_18511,N_19750);
or U21960 (N_21960,N_17894,N_19591);
and U21961 (N_21961,N_19111,N_18031);
and U21962 (N_21962,N_19674,N_18448);
and U21963 (N_21963,N_19478,N_17680);
or U21964 (N_21964,N_19033,N_19183);
nor U21965 (N_21965,N_19653,N_18577);
and U21966 (N_21966,N_19948,N_18492);
or U21967 (N_21967,N_18891,N_18561);
nand U21968 (N_21968,N_18364,N_17937);
xor U21969 (N_21969,N_19099,N_19793);
xor U21970 (N_21970,N_18453,N_19789);
nor U21971 (N_21971,N_18632,N_18687);
and U21972 (N_21972,N_18242,N_18048);
xor U21973 (N_21973,N_18988,N_18332);
nand U21974 (N_21974,N_19338,N_19144);
and U21975 (N_21975,N_19773,N_18134);
or U21976 (N_21976,N_18128,N_19242);
nor U21977 (N_21977,N_19696,N_18685);
xnor U21978 (N_21978,N_19429,N_19331);
or U21979 (N_21979,N_19430,N_19195);
xnor U21980 (N_21980,N_18092,N_17801);
nor U21981 (N_21981,N_18682,N_18407);
xnor U21982 (N_21982,N_19143,N_18423);
xnor U21983 (N_21983,N_18100,N_19106);
nand U21984 (N_21984,N_19248,N_19856);
nor U21985 (N_21985,N_18713,N_19398);
xor U21986 (N_21986,N_18158,N_18737);
xnor U21987 (N_21987,N_18087,N_18305);
nor U21988 (N_21988,N_17539,N_19388);
and U21989 (N_21989,N_19016,N_18255);
xor U21990 (N_21990,N_19176,N_17696);
and U21991 (N_21991,N_18754,N_19035);
nor U21992 (N_21992,N_19796,N_17547);
nand U21993 (N_21993,N_19712,N_17624);
nor U21994 (N_21994,N_19806,N_18054);
nor U21995 (N_21995,N_17759,N_18369);
or U21996 (N_21996,N_19970,N_19766);
and U21997 (N_21997,N_18754,N_19803);
or U21998 (N_21998,N_18220,N_19848);
or U21999 (N_21999,N_18349,N_17551);
nand U22000 (N_22000,N_19201,N_18592);
nand U22001 (N_22001,N_18169,N_18571);
xnor U22002 (N_22002,N_19644,N_17818);
nor U22003 (N_22003,N_18151,N_19661);
or U22004 (N_22004,N_19609,N_18462);
nand U22005 (N_22005,N_18431,N_19493);
nand U22006 (N_22006,N_19294,N_18768);
or U22007 (N_22007,N_18164,N_19598);
xnor U22008 (N_22008,N_19063,N_18526);
nor U22009 (N_22009,N_19089,N_19710);
or U22010 (N_22010,N_18174,N_17503);
and U22011 (N_22011,N_18080,N_18703);
and U22012 (N_22012,N_19637,N_18695);
nor U22013 (N_22013,N_19309,N_19752);
and U22014 (N_22014,N_18657,N_17762);
or U22015 (N_22015,N_18007,N_18544);
nor U22016 (N_22016,N_19035,N_18337);
nor U22017 (N_22017,N_19288,N_19335);
xor U22018 (N_22018,N_18665,N_19315);
nor U22019 (N_22019,N_19922,N_17870);
and U22020 (N_22020,N_18032,N_19099);
and U22021 (N_22021,N_18360,N_18142);
and U22022 (N_22022,N_18725,N_19422);
xnor U22023 (N_22023,N_17978,N_18400);
xor U22024 (N_22024,N_18773,N_19136);
nand U22025 (N_22025,N_18107,N_19946);
nor U22026 (N_22026,N_19943,N_18753);
xnor U22027 (N_22027,N_18635,N_19651);
or U22028 (N_22028,N_19690,N_19480);
or U22029 (N_22029,N_19755,N_18959);
nand U22030 (N_22030,N_19119,N_18365);
nor U22031 (N_22031,N_19815,N_18512);
nand U22032 (N_22032,N_19292,N_19389);
xnor U22033 (N_22033,N_19634,N_19065);
nand U22034 (N_22034,N_18385,N_19813);
nor U22035 (N_22035,N_18246,N_18159);
nor U22036 (N_22036,N_18751,N_19863);
nor U22037 (N_22037,N_19635,N_17920);
and U22038 (N_22038,N_18928,N_17553);
and U22039 (N_22039,N_18458,N_19371);
and U22040 (N_22040,N_18158,N_18445);
or U22041 (N_22041,N_19247,N_17766);
xnor U22042 (N_22042,N_19816,N_18503);
xor U22043 (N_22043,N_18600,N_17709);
or U22044 (N_22044,N_18823,N_18977);
nand U22045 (N_22045,N_19781,N_17504);
nor U22046 (N_22046,N_18768,N_19262);
nor U22047 (N_22047,N_18383,N_19170);
xnor U22048 (N_22048,N_18329,N_19938);
and U22049 (N_22049,N_19577,N_18418);
and U22050 (N_22050,N_19159,N_19004);
xor U22051 (N_22051,N_19113,N_18364);
and U22052 (N_22052,N_19914,N_17654);
nand U22053 (N_22053,N_19540,N_19779);
nor U22054 (N_22054,N_19545,N_18610);
nor U22055 (N_22055,N_18593,N_19983);
nand U22056 (N_22056,N_17599,N_18687);
or U22057 (N_22057,N_19892,N_18788);
xor U22058 (N_22058,N_17931,N_18361);
and U22059 (N_22059,N_18081,N_17933);
and U22060 (N_22060,N_19232,N_17731);
or U22061 (N_22061,N_18260,N_19849);
or U22062 (N_22062,N_19667,N_19458);
nand U22063 (N_22063,N_19595,N_19183);
or U22064 (N_22064,N_19411,N_19784);
nand U22065 (N_22065,N_18928,N_18152);
or U22066 (N_22066,N_19067,N_17990);
xnor U22067 (N_22067,N_17981,N_19977);
and U22068 (N_22068,N_18501,N_17691);
xnor U22069 (N_22069,N_19049,N_19163);
nor U22070 (N_22070,N_18920,N_19544);
and U22071 (N_22071,N_18318,N_18334);
xor U22072 (N_22072,N_18125,N_18095);
and U22073 (N_22073,N_18725,N_18917);
nand U22074 (N_22074,N_18241,N_18305);
xnor U22075 (N_22075,N_19786,N_17791);
nand U22076 (N_22076,N_17636,N_19337);
and U22077 (N_22077,N_19028,N_19928);
or U22078 (N_22078,N_18073,N_17686);
nand U22079 (N_22079,N_18778,N_19806);
and U22080 (N_22080,N_19765,N_17752);
nand U22081 (N_22081,N_18481,N_17953);
or U22082 (N_22082,N_19165,N_17850);
nor U22083 (N_22083,N_18486,N_19508);
nor U22084 (N_22084,N_18102,N_18597);
and U22085 (N_22085,N_18376,N_18255);
xor U22086 (N_22086,N_19348,N_18247);
and U22087 (N_22087,N_18214,N_18636);
nand U22088 (N_22088,N_19103,N_19292);
xnor U22089 (N_22089,N_18340,N_17812);
nor U22090 (N_22090,N_18860,N_19165);
nor U22091 (N_22091,N_19091,N_18777);
nand U22092 (N_22092,N_17972,N_18499);
or U22093 (N_22093,N_18861,N_19060);
or U22094 (N_22094,N_17630,N_17504);
xnor U22095 (N_22095,N_19989,N_19270);
and U22096 (N_22096,N_17646,N_17797);
nand U22097 (N_22097,N_17840,N_17728);
or U22098 (N_22098,N_18534,N_19773);
nand U22099 (N_22099,N_18758,N_19545);
or U22100 (N_22100,N_17662,N_19650);
nand U22101 (N_22101,N_19424,N_19471);
nand U22102 (N_22102,N_18891,N_19799);
and U22103 (N_22103,N_19188,N_18899);
nor U22104 (N_22104,N_18115,N_17769);
nor U22105 (N_22105,N_18469,N_19758);
nand U22106 (N_22106,N_19150,N_19046);
or U22107 (N_22107,N_17580,N_19898);
xnor U22108 (N_22108,N_19208,N_18990);
or U22109 (N_22109,N_19093,N_19418);
xor U22110 (N_22110,N_18945,N_17858);
or U22111 (N_22111,N_19300,N_17602);
nand U22112 (N_22112,N_17820,N_19195);
xnor U22113 (N_22113,N_18395,N_19017);
nand U22114 (N_22114,N_18183,N_19008);
or U22115 (N_22115,N_18325,N_18935);
or U22116 (N_22116,N_18055,N_19182);
or U22117 (N_22117,N_17698,N_18184);
nand U22118 (N_22118,N_17925,N_19478);
nand U22119 (N_22119,N_19571,N_18546);
or U22120 (N_22120,N_19232,N_17916);
nand U22121 (N_22121,N_18450,N_18610);
nor U22122 (N_22122,N_18252,N_18299);
or U22123 (N_22123,N_18262,N_18167);
nor U22124 (N_22124,N_18071,N_19848);
xor U22125 (N_22125,N_19514,N_18304);
nand U22126 (N_22126,N_19154,N_18379);
and U22127 (N_22127,N_17656,N_18648);
and U22128 (N_22128,N_17511,N_17880);
nor U22129 (N_22129,N_17958,N_18910);
or U22130 (N_22130,N_18496,N_19896);
xor U22131 (N_22131,N_19591,N_18978);
xor U22132 (N_22132,N_18578,N_19459);
nor U22133 (N_22133,N_17943,N_18953);
and U22134 (N_22134,N_19329,N_19383);
nand U22135 (N_22135,N_19151,N_19042);
xor U22136 (N_22136,N_19928,N_17538);
nand U22137 (N_22137,N_17986,N_17806);
or U22138 (N_22138,N_18538,N_18192);
xnor U22139 (N_22139,N_18239,N_18662);
and U22140 (N_22140,N_19081,N_17757);
xor U22141 (N_22141,N_17540,N_18736);
nand U22142 (N_22142,N_19006,N_17779);
or U22143 (N_22143,N_18500,N_19216);
nor U22144 (N_22144,N_18252,N_17877);
and U22145 (N_22145,N_18087,N_17957);
or U22146 (N_22146,N_19970,N_17810);
and U22147 (N_22147,N_19229,N_18755);
nand U22148 (N_22148,N_18505,N_18634);
xor U22149 (N_22149,N_19327,N_18672);
nand U22150 (N_22150,N_17722,N_17930);
xnor U22151 (N_22151,N_18794,N_18271);
and U22152 (N_22152,N_19418,N_17919);
xor U22153 (N_22153,N_19251,N_19175);
or U22154 (N_22154,N_17818,N_19647);
and U22155 (N_22155,N_17626,N_17669);
and U22156 (N_22156,N_18069,N_18986);
xor U22157 (N_22157,N_18363,N_18527);
xor U22158 (N_22158,N_19260,N_19677);
and U22159 (N_22159,N_19512,N_17893);
nand U22160 (N_22160,N_18584,N_18320);
and U22161 (N_22161,N_18733,N_18551);
or U22162 (N_22162,N_19136,N_18784);
and U22163 (N_22163,N_19979,N_18890);
nor U22164 (N_22164,N_19821,N_19356);
xor U22165 (N_22165,N_18724,N_19291);
and U22166 (N_22166,N_19604,N_18360);
and U22167 (N_22167,N_19878,N_18528);
nor U22168 (N_22168,N_19972,N_18357);
nor U22169 (N_22169,N_17825,N_19754);
xor U22170 (N_22170,N_19452,N_19555);
xnor U22171 (N_22171,N_18160,N_18617);
and U22172 (N_22172,N_19379,N_19629);
nand U22173 (N_22173,N_19195,N_18201);
nor U22174 (N_22174,N_17762,N_19020);
nor U22175 (N_22175,N_18887,N_17838);
xor U22176 (N_22176,N_19848,N_19960);
nor U22177 (N_22177,N_17929,N_19995);
xor U22178 (N_22178,N_17847,N_18674);
or U22179 (N_22179,N_19526,N_17563);
or U22180 (N_22180,N_19814,N_18940);
nor U22181 (N_22181,N_18454,N_17780);
and U22182 (N_22182,N_18577,N_18171);
nand U22183 (N_22183,N_19476,N_17723);
nand U22184 (N_22184,N_18985,N_18101);
and U22185 (N_22185,N_18516,N_18187);
nand U22186 (N_22186,N_17597,N_17866);
nand U22187 (N_22187,N_18659,N_19850);
and U22188 (N_22188,N_17702,N_18185);
or U22189 (N_22189,N_18028,N_19977);
and U22190 (N_22190,N_19888,N_19531);
nand U22191 (N_22191,N_18675,N_19296);
nor U22192 (N_22192,N_19645,N_18313);
xor U22193 (N_22193,N_17757,N_18208);
or U22194 (N_22194,N_18571,N_18026);
nor U22195 (N_22195,N_19574,N_19411);
xor U22196 (N_22196,N_19301,N_18836);
or U22197 (N_22197,N_19566,N_18448);
or U22198 (N_22198,N_17831,N_19819);
or U22199 (N_22199,N_19316,N_18021);
nand U22200 (N_22200,N_18728,N_19828);
and U22201 (N_22201,N_18639,N_19340);
nand U22202 (N_22202,N_19373,N_18761);
and U22203 (N_22203,N_19846,N_19658);
nor U22204 (N_22204,N_19182,N_19656);
nor U22205 (N_22205,N_19509,N_19077);
nor U22206 (N_22206,N_19645,N_19865);
xor U22207 (N_22207,N_19639,N_18778);
or U22208 (N_22208,N_18751,N_18278);
or U22209 (N_22209,N_19788,N_17551);
xnor U22210 (N_22210,N_18498,N_19586);
xnor U22211 (N_22211,N_18842,N_19412);
or U22212 (N_22212,N_18270,N_17950);
xor U22213 (N_22213,N_19457,N_17512);
nor U22214 (N_22214,N_18389,N_19405);
nand U22215 (N_22215,N_18284,N_18776);
or U22216 (N_22216,N_19618,N_19040);
nor U22217 (N_22217,N_18325,N_17570);
or U22218 (N_22218,N_19245,N_17531);
nand U22219 (N_22219,N_19080,N_19389);
nand U22220 (N_22220,N_18249,N_18491);
or U22221 (N_22221,N_17935,N_18295);
and U22222 (N_22222,N_18794,N_19793);
nand U22223 (N_22223,N_18479,N_19342);
nand U22224 (N_22224,N_18527,N_18312);
or U22225 (N_22225,N_19678,N_18431);
and U22226 (N_22226,N_17575,N_19487);
and U22227 (N_22227,N_19372,N_19163);
xnor U22228 (N_22228,N_18344,N_18314);
nor U22229 (N_22229,N_19898,N_17918);
and U22230 (N_22230,N_18479,N_19118);
xor U22231 (N_22231,N_19078,N_18127);
xor U22232 (N_22232,N_17635,N_18114);
nor U22233 (N_22233,N_17902,N_18796);
nand U22234 (N_22234,N_19852,N_18669);
or U22235 (N_22235,N_19447,N_19037);
or U22236 (N_22236,N_19257,N_19521);
or U22237 (N_22237,N_18311,N_17962);
or U22238 (N_22238,N_18892,N_18363);
and U22239 (N_22239,N_18910,N_19278);
nand U22240 (N_22240,N_18007,N_18186);
xnor U22241 (N_22241,N_19696,N_18815);
or U22242 (N_22242,N_19553,N_19173);
and U22243 (N_22243,N_18191,N_17904);
nor U22244 (N_22244,N_17519,N_19225);
and U22245 (N_22245,N_18318,N_18324);
nand U22246 (N_22246,N_18022,N_18099);
and U22247 (N_22247,N_18337,N_18748);
and U22248 (N_22248,N_18795,N_17879);
xnor U22249 (N_22249,N_18612,N_17598);
or U22250 (N_22250,N_18958,N_18727);
or U22251 (N_22251,N_18306,N_18698);
nor U22252 (N_22252,N_19606,N_18742);
nand U22253 (N_22253,N_17620,N_18632);
nand U22254 (N_22254,N_18824,N_17574);
xnor U22255 (N_22255,N_18267,N_19694);
nor U22256 (N_22256,N_18882,N_19586);
nand U22257 (N_22257,N_17508,N_18700);
xnor U22258 (N_22258,N_18549,N_17502);
nand U22259 (N_22259,N_19149,N_17796);
or U22260 (N_22260,N_19624,N_19662);
xor U22261 (N_22261,N_18342,N_19669);
or U22262 (N_22262,N_18860,N_18513);
or U22263 (N_22263,N_19611,N_17882);
nor U22264 (N_22264,N_19410,N_19617);
xnor U22265 (N_22265,N_19207,N_17730);
nor U22266 (N_22266,N_18615,N_19243);
xnor U22267 (N_22267,N_18021,N_18868);
nand U22268 (N_22268,N_19901,N_17884);
nor U22269 (N_22269,N_19035,N_19466);
or U22270 (N_22270,N_19267,N_18018);
or U22271 (N_22271,N_18038,N_19662);
nor U22272 (N_22272,N_19156,N_19024);
nand U22273 (N_22273,N_19438,N_19343);
nand U22274 (N_22274,N_18886,N_17526);
or U22275 (N_22275,N_19313,N_19168);
nor U22276 (N_22276,N_19129,N_18106);
xor U22277 (N_22277,N_19403,N_17570);
nand U22278 (N_22278,N_19369,N_19640);
or U22279 (N_22279,N_17614,N_18612);
xor U22280 (N_22280,N_18926,N_17695);
nand U22281 (N_22281,N_17809,N_19873);
and U22282 (N_22282,N_18688,N_17554);
xor U22283 (N_22283,N_17753,N_18215);
xor U22284 (N_22284,N_17741,N_17652);
nor U22285 (N_22285,N_19054,N_17902);
and U22286 (N_22286,N_19921,N_19720);
and U22287 (N_22287,N_18852,N_18781);
or U22288 (N_22288,N_17975,N_19112);
or U22289 (N_22289,N_19531,N_17635);
nor U22290 (N_22290,N_18140,N_19424);
xor U22291 (N_22291,N_17800,N_18114);
or U22292 (N_22292,N_18710,N_17870);
nor U22293 (N_22293,N_19440,N_19132);
nand U22294 (N_22294,N_18818,N_18071);
and U22295 (N_22295,N_19657,N_18182);
and U22296 (N_22296,N_18037,N_17818);
or U22297 (N_22297,N_19799,N_19523);
and U22298 (N_22298,N_18202,N_17752);
nor U22299 (N_22299,N_19309,N_18989);
nor U22300 (N_22300,N_19206,N_18284);
xnor U22301 (N_22301,N_19732,N_17623);
nor U22302 (N_22302,N_17865,N_17514);
xor U22303 (N_22303,N_18589,N_18324);
and U22304 (N_22304,N_18871,N_17913);
or U22305 (N_22305,N_19280,N_17661);
nand U22306 (N_22306,N_18604,N_19510);
nand U22307 (N_22307,N_19060,N_19253);
and U22308 (N_22308,N_19090,N_17686);
or U22309 (N_22309,N_19527,N_18195);
or U22310 (N_22310,N_19201,N_19655);
and U22311 (N_22311,N_19266,N_18676);
nand U22312 (N_22312,N_18632,N_18274);
xnor U22313 (N_22313,N_18275,N_17815);
nand U22314 (N_22314,N_18009,N_18389);
xnor U22315 (N_22315,N_18487,N_18591);
xor U22316 (N_22316,N_19856,N_19130);
xor U22317 (N_22317,N_18377,N_19272);
or U22318 (N_22318,N_18856,N_19609);
and U22319 (N_22319,N_19295,N_19030);
and U22320 (N_22320,N_18367,N_19253);
or U22321 (N_22321,N_19940,N_18814);
and U22322 (N_22322,N_19283,N_19995);
and U22323 (N_22323,N_17711,N_19052);
or U22324 (N_22324,N_18069,N_18198);
xor U22325 (N_22325,N_18850,N_19074);
nor U22326 (N_22326,N_19024,N_19493);
and U22327 (N_22327,N_18398,N_19579);
nand U22328 (N_22328,N_19511,N_19798);
nor U22329 (N_22329,N_19325,N_19621);
or U22330 (N_22330,N_18606,N_19232);
nor U22331 (N_22331,N_19604,N_19363);
xor U22332 (N_22332,N_19557,N_19850);
and U22333 (N_22333,N_19555,N_17599);
xnor U22334 (N_22334,N_18369,N_17512);
and U22335 (N_22335,N_19339,N_18514);
and U22336 (N_22336,N_17987,N_17950);
nor U22337 (N_22337,N_18964,N_19104);
and U22338 (N_22338,N_18215,N_17919);
and U22339 (N_22339,N_18196,N_17742);
nor U22340 (N_22340,N_18683,N_18275);
nor U22341 (N_22341,N_19397,N_18537);
nor U22342 (N_22342,N_19794,N_19544);
or U22343 (N_22343,N_18221,N_19350);
nor U22344 (N_22344,N_17735,N_19201);
and U22345 (N_22345,N_19168,N_19961);
xor U22346 (N_22346,N_18459,N_18427);
or U22347 (N_22347,N_18313,N_19757);
xnor U22348 (N_22348,N_19697,N_18356);
nor U22349 (N_22349,N_17527,N_19271);
nand U22350 (N_22350,N_18053,N_18819);
or U22351 (N_22351,N_18108,N_17927);
nand U22352 (N_22352,N_18482,N_17925);
or U22353 (N_22353,N_18345,N_19719);
xnor U22354 (N_22354,N_19975,N_17789);
nor U22355 (N_22355,N_19787,N_17762);
or U22356 (N_22356,N_19764,N_19440);
nor U22357 (N_22357,N_19232,N_18418);
or U22358 (N_22358,N_18723,N_18077);
nor U22359 (N_22359,N_19547,N_19933);
nor U22360 (N_22360,N_18238,N_18113);
and U22361 (N_22361,N_18152,N_18977);
nor U22362 (N_22362,N_18834,N_19266);
nand U22363 (N_22363,N_19855,N_18906);
or U22364 (N_22364,N_19594,N_17744);
nand U22365 (N_22365,N_18584,N_18354);
or U22366 (N_22366,N_18122,N_19083);
nand U22367 (N_22367,N_17908,N_18071);
nand U22368 (N_22368,N_19651,N_18046);
nand U22369 (N_22369,N_18552,N_18730);
nand U22370 (N_22370,N_19340,N_19535);
and U22371 (N_22371,N_19898,N_18377);
nand U22372 (N_22372,N_18515,N_19743);
xnor U22373 (N_22373,N_18128,N_19048);
nor U22374 (N_22374,N_19824,N_19512);
nand U22375 (N_22375,N_18717,N_17625);
nor U22376 (N_22376,N_18116,N_17706);
and U22377 (N_22377,N_18319,N_18310);
nand U22378 (N_22378,N_19756,N_19642);
xor U22379 (N_22379,N_18191,N_17969);
nand U22380 (N_22380,N_19474,N_18057);
or U22381 (N_22381,N_18333,N_17720);
and U22382 (N_22382,N_19947,N_18863);
nand U22383 (N_22383,N_18781,N_18533);
xnor U22384 (N_22384,N_18092,N_19654);
xnor U22385 (N_22385,N_19234,N_19921);
and U22386 (N_22386,N_17948,N_19984);
xor U22387 (N_22387,N_17835,N_19933);
and U22388 (N_22388,N_17949,N_19235);
or U22389 (N_22389,N_19113,N_18450);
nor U22390 (N_22390,N_19125,N_18480);
and U22391 (N_22391,N_17605,N_19606);
xor U22392 (N_22392,N_17882,N_18061);
xnor U22393 (N_22393,N_18436,N_18819);
xor U22394 (N_22394,N_19299,N_19304);
or U22395 (N_22395,N_18952,N_19554);
and U22396 (N_22396,N_19122,N_17850);
nand U22397 (N_22397,N_19782,N_19640);
nand U22398 (N_22398,N_17502,N_19907);
nand U22399 (N_22399,N_18826,N_18434);
or U22400 (N_22400,N_19955,N_18139);
nand U22401 (N_22401,N_18184,N_19658);
nor U22402 (N_22402,N_18623,N_18703);
xnor U22403 (N_22403,N_18373,N_18624);
nand U22404 (N_22404,N_17707,N_18590);
or U22405 (N_22405,N_18213,N_17984);
and U22406 (N_22406,N_19511,N_18356);
or U22407 (N_22407,N_17610,N_18851);
nor U22408 (N_22408,N_18921,N_17684);
nor U22409 (N_22409,N_17799,N_19494);
xnor U22410 (N_22410,N_19389,N_19342);
or U22411 (N_22411,N_19331,N_19648);
and U22412 (N_22412,N_19698,N_18387);
nor U22413 (N_22413,N_18575,N_17636);
nand U22414 (N_22414,N_18697,N_19052);
nand U22415 (N_22415,N_18436,N_18867);
xor U22416 (N_22416,N_19541,N_19822);
or U22417 (N_22417,N_18425,N_17912);
nand U22418 (N_22418,N_18746,N_19539);
or U22419 (N_22419,N_19527,N_19629);
nor U22420 (N_22420,N_19582,N_18109);
nor U22421 (N_22421,N_18107,N_19715);
or U22422 (N_22422,N_18592,N_17949);
xor U22423 (N_22423,N_17804,N_18122);
nor U22424 (N_22424,N_18010,N_19163);
or U22425 (N_22425,N_19205,N_19937);
or U22426 (N_22426,N_18403,N_18889);
nor U22427 (N_22427,N_18493,N_18416);
and U22428 (N_22428,N_19802,N_18694);
nor U22429 (N_22429,N_17967,N_18877);
nor U22430 (N_22430,N_18741,N_19124);
nor U22431 (N_22431,N_17872,N_18323);
xor U22432 (N_22432,N_19473,N_18596);
nor U22433 (N_22433,N_19098,N_18732);
xor U22434 (N_22434,N_19179,N_18020);
and U22435 (N_22435,N_19350,N_18987);
and U22436 (N_22436,N_18641,N_18075);
xnor U22437 (N_22437,N_19756,N_19667);
and U22438 (N_22438,N_18292,N_19215);
nand U22439 (N_22439,N_19022,N_18397);
or U22440 (N_22440,N_18154,N_18081);
nand U22441 (N_22441,N_19739,N_19229);
nand U22442 (N_22442,N_19585,N_19642);
or U22443 (N_22443,N_18018,N_17512);
xor U22444 (N_22444,N_18466,N_18523);
or U22445 (N_22445,N_18417,N_18315);
and U22446 (N_22446,N_17617,N_19502);
nor U22447 (N_22447,N_19940,N_19982);
and U22448 (N_22448,N_17820,N_18990);
xor U22449 (N_22449,N_19191,N_17805);
xnor U22450 (N_22450,N_19889,N_17581);
xnor U22451 (N_22451,N_19470,N_18855);
and U22452 (N_22452,N_18732,N_19331);
xnor U22453 (N_22453,N_19449,N_19593);
and U22454 (N_22454,N_19007,N_18741);
and U22455 (N_22455,N_19938,N_19299);
or U22456 (N_22456,N_18684,N_19085);
and U22457 (N_22457,N_17866,N_18531);
xnor U22458 (N_22458,N_19235,N_18720);
xor U22459 (N_22459,N_19592,N_17616);
xor U22460 (N_22460,N_19385,N_18507);
nor U22461 (N_22461,N_17514,N_17510);
xor U22462 (N_22462,N_18523,N_18219);
and U22463 (N_22463,N_19545,N_19308);
nor U22464 (N_22464,N_17785,N_19927);
nand U22465 (N_22465,N_19391,N_18242);
and U22466 (N_22466,N_18406,N_18747);
nor U22467 (N_22467,N_18288,N_19292);
xnor U22468 (N_22468,N_18402,N_19643);
nand U22469 (N_22469,N_19857,N_19598);
nand U22470 (N_22470,N_19573,N_19180);
xnor U22471 (N_22471,N_18041,N_19061);
nand U22472 (N_22472,N_18393,N_18504);
or U22473 (N_22473,N_19938,N_18050);
xnor U22474 (N_22474,N_18225,N_19766);
nor U22475 (N_22475,N_18817,N_18969);
and U22476 (N_22476,N_19983,N_18823);
or U22477 (N_22477,N_18298,N_19465);
and U22478 (N_22478,N_18848,N_17726);
and U22479 (N_22479,N_17952,N_18580);
nand U22480 (N_22480,N_17982,N_18779);
and U22481 (N_22481,N_19373,N_17637);
nand U22482 (N_22482,N_19911,N_18926);
and U22483 (N_22483,N_19395,N_19163);
xnor U22484 (N_22484,N_17707,N_18059);
xnor U22485 (N_22485,N_17928,N_19651);
and U22486 (N_22486,N_19815,N_19718);
xnor U22487 (N_22487,N_19556,N_19708);
nand U22488 (N_22488,N_18363,N_19491);
nand U22489 (N_22489,N_17937,N_19016);
or U22490 (N_22490,N_19978,N_19581);
or U22491 (N_22491,N_18292,N_18924);
xnor U22492 (N_22492,N_19478,N_18806);
xor U22493 (N_22493,N_19203,N_18687);
or U22494 (N_22494,N_18428,N_18345);
xnor U22495 (N_22495,N_17869,N_18375);
nor U22496 (N_22496,N_17943,N_18741);
xnor U22497 (N_22497,N_18160,N_18223);
xnor U22498 (N_22498,N_18516,N_18769);
and U22499 (N_22499,N_17718,N_18268);
nor U22500 (N_22500,N_20564,N_20569);
or U22501 (N_22501,N_21694,N_20893);
nand U22502 (N_22502,N_21649,N_21098);
nand U22503 (N_22503,N_22166,N_21191);
xor U22504 (N_22504,N_21943,N_21260);
xnor U22505 (N_22505,N_20237,N_21642);
nand U22506 (N_22506,N_21176,N_21501);
and U22507 (N_22507,N_22429,N_20779);
nor U22508 (N_22508,N_22030,N_20395);
nand U22509 (N_22509,N_20203,N_20012);
xor U22510 (N_22510,N_20407,N_20960);
nor U22511 (N_22511,N_21392,N_21491);
nor U22512 (N_22512,N_21937,N_21285);
xor U22513 (N_22513,N_20947,N_21825);
xnor U22514 (N_22514,N_21907,N_21883);
xor U22515 (N_22515,N_20558,N_22387);
xor U22516 (N_22516,N_21856,N_20673);
xnor U22517 (N_22517,N_21933,N_21964);
xnor U22518 (N_22518,N_20145,N_21543);
nor U22519 (N_22519,N_20210,N_22255);
and U22520 (N_22520,N_22238,N_20944);
nand U22521 (N_22521,N_20552,N_21468);
xnor U22522 (N_22522,N_22055,N_21999);
nand U22523 (N_22523,N_20497,N_20521);
nand U22524 (N_22524,N_20928,N_21798);
or U22525 (N_22525,N_20406,N_21521);
nor U22526 (N_22526,N_21261,N_22232);
nor U22527 (N_22527,N_21023,N_20638);
nand U22528 (N_22528,N_20584,N_20883);
and U22529 (N_22529,N_22186,N_22019);
and U22530 (N_22530,N_22367,N_20230);
nor U22531 (N_22531,N_20095,N_21060);
nand U22532 (N_22532,N_20362,N_20810);
nor U22533 (N_22533,N_21225,N_20926);
and U22534 (N_22534,N_21834,N_22118);
nor U22535 (N_22535,N_20402,N_22452);
and U22536 (N_22536,N_20380,N_21074);
or U22537 (N_22537,N_21743,N_22462);
xnor U22538 (N_22538,N_21925,N_21840);
and U22539 (N_22539,N_22069,N_20666);
nor U22540 (N_22540,N_22406,N_22280);
or U22541 (N_22541,N_21659,N_20118);
nor U22542 (N_22542,N_20057,N_21788);
and U22543 (N_22543,N_22291,N_22135);
nor U22544 (N_22544,N_20489,N_20382);
nand U22545 (N_22545,N_20387,N_22359);
nand U22546 (N_22546,N_21742,N_22008);
xor U22547 (N_22547,N_21799,N_21529);
or U22548 (N_22548,N_20847,N_20371);
nor U22549 (N_22549,N_20176,N_21820);
xnor U22550 (N_22550,N_21349,N_20021);
or U22551 (N_22551,N_21057,N_20843);
or U22552 (N_22552,N_20591,N_22259);
nor U22553 (N_22553,N_20300,N_21668);
xor U22554 (N_22554,N_20878,N_20703);
nor U22555 (N_22555,N_21487,N_20601);
or U22556 (N_22556,N_21751,N_20864);
nor U22557 (N_22557,N_21371,N_21830);
or U22558 (N_22558,N_21072,N_21711);
xnor U22559 (N_22559,N_21888,N_21294);
nor U22560 (N_22560,N_20888,N_20296);
nor U22561 (N_22561,N_22349,N_21372);
xnor U22562 (N_22562,N_20716,N_21105);
nand U22563 (N_22563,N_21973,N_20180);
nand U22564 (N_22564,N_21004,N_21877);
xor U22565 (N_22565,N_20797,N_20913);
and U22566 (N_22566,N_21413,N_21827);
nor U22567 (N_22567,N_20045,N_20634);
nand U22568 (N_22568,N_20904,N_21727);
or U22569 (N_22569,N_22327,N_21208);
xor U22570 (N_22570,N_22424,N_20124);
nor U22571 (N_22571,N_21740,N_20690);
nor U22572 (N_22572,N_21996,N_20549);
or U22573 (N_22573,N_20494,N_20148);
nand U22574 (N_22574,N_20799,N_20835);
nor U22575 (N_22575,N_21013,N_22453);
and U22576 (N_22576,N_21734,N_20289);
and U22577 (N_22577,N_22112,N_21787);
or U22578 (N_22578,N_22231,N_20929);
nor U22579 (N_22579,N_21815,N_21499);
nand U22580 (N_22580,N_21420,N_21324);
xor U22581 (N_22581,N_22218,N_22431);
and U22582 (N_22582,N_21351,N_20675);
and U22583 (N_22583,N_22066,N_20108);
nor U22584 (N_22584,N_22265,N_21424);
and U22585 (N_22585,N_20714,N_20891);
xor U22586 (N_22586,N_21164,N_21234);
nand U22587 (N_22587,N_21236,N_21990);
nor U22588 (N_22588,N_21494,N_21924);
nor U22589 (N_22589,N_21120,N_22119);
and U22590 (N_22590,N_20292,N_22063);
or U22591 (N_22591,N_20639,N_21247);
or U22592 (N_22592,N_20383,N_21240);
xnor U22593 (N_22593,N_20824,N_20499);
nand U22594 (N_22594,N_21812,N_21969);
or U22595 (N_22595,N_21053,N_21362);
or U22596 (N_22596,N_20557,N_20597);
nand U22597 (N_22597,N_21549,N_20577);
and U22598 (N_22598,N_21334,N_21216);
and U22599 (N_22599,N_20072,N_20876);
or U22600 (N_22600,N_21376,N_20811);
and U22601 (N_22601,N_20945,N_20694);
nand U22602 (N_22602,N_21921,N_22448);
and U22603 (N_22603,N_20850,N_22078);
or U22604 (N_22604,N_20887,N_20043);
nor U22605 (N_22605,N_21874,N_20092);
xnor U22606 (N_22606,N_21608,N_21142);
nand U22607 (N_22607,N_22077,N_20132);
nor U22608 (N_22608,N_20486,N_22148);
xor U22609 (N_22609,N_20711,N_20082);
nor U22610 (N_22610,N_21878,N_20604);
nand U22611 (N_22611,N_20539,N_21124);
or U22612 (N_22612,N_21960,N_22403);
xor U22613 (N_22613,N_20069,N_21656);
and U22614 (N_22614,N_20837,N_21381);
nand U22615 (N_22615,N_20135,N_21148);
nor U22616 (N_22616,N_21012,N_22330);
nor U22617 (N_22617,N_22152,N_21702);
and U22618 (N_22618,N_20063,N_20479);
xnor U22619 (N_22619,N_20324,N_21889);
nand U22620 (N_22620,N_20962,N_20918);
and U22621 (N_22621,N_21310,N_21335);
nand U22622 (N_22622,N_20940,N_21522);
or U22623 (N_22623,N_20017,N_20855);
nor U22624 (N_22624,N_20463,N_20753);
xnor U22625 (N_22625,N_22415,N_21390);
nand U22626 (N_22626,N_21532,N_20544);
and U22627 (N_22627,N_20979,N_21613);
nor U22628 (N_22628,N_21443,N_20275);
nor U22629 (N_22629,N_21988,N_21410);
or U22630 (N_22630,N_21461,N_22147);
or U22631 (N_22631,N_20568,N_21192);
and U22632 (N_22632,N_21810,N_21764);
and U22633 (N_22633,N_20050,N_21205);
nor U22634 (N_22634,N_21253,N_21576);
or U22635 (N_22635,N_20080,N_22056);
and U22636 (N_22636,N_22292,N_20542);
or U22637 (N_22637,N_21375,N_21651);
and U22638 (N_22638,N_21186,N_21887);
and U22639 (N_22639,N_21816,N_21384);
or U22640 (N_22640,N_22230,N_22303);
nor U22641 (N_22641,N_20496,N_21959);
xnor U22642 (N_22642,N_20846,N_20867);
xnor U22643 (N_22643,N_21564,N_20248);
nor U22644 (N_22644,N_21055,N_20239);
nand U22645 (N_22645,N_20309,N_20337);
and U22646 (N_22646,N_21238,N_21592);
nor U22647 (N_22647,N_21724,N_21805);
or U22648 (N_22648,N_21370,N_22458);
and U22649 (N_22649,N_22136,N_20485);
xor U22650 (N_22650,N_20646,N_21559);
and U22651 (N_22651,N_20439,N_20559);
and U22652 (N_22652,N_20922,N_21533);
xor U22653 (N_22653,N_22005,N_20038);
or U22654 (N_22654,N_22053,N_22271);
nand U22655 (N_22655,N_20720,N_21955);
or U22656 (N_22656,N_21493,N_21583);
nand U22657 (N_22657,N_20896,N_20375);
and U22658 (N_22658,N_20351,N_21223);
nand U22659 (N_22659,N_21962,N_21604);
xor U22660 (N_22660,N_20437,N_20713);
nand U22661 (N_22661,N_22102,N_22194);
nor U22662 (N_22662,N_21006,N_20515);
xnor U22663 (N_22663,N_20458,N_22495);
and U22664 (N_22664,N_22241,N_20882);
or U22665 (N_22665,N_20002,N_20413);
nor U22666 (N_22666,N_21752,N_20097);
nand U22667 (N_22667,N_21919,N_21337);
nand U22668 (N_22668,N_20778,N_22295);
xor U22669 (N_22669,N_20995,N_22414);
nand U22670 (N_22670,N_20781,N_21645);
xor U22671 (N_22671,N_22164,N_20519);
nand U22672 (N_22672,N_20774,N_21516);
nand U22673 (N_22673,N_22215,N_22060);
and U22674 (N_22674,N_20999,N_20310);
nand U22675 (N_22675,N_22162,N_21895);
and U22676 (N_22676,N_20526,N_21986);
nor U22677 (N_22677,N_22183,N_21712);
nor U22678 (N_22678,N_21116,N_20516);
and U22679 (N_22679,N_21056,N_22489);
nand U22680 (N_22680,N_20614,N_21052);
or U22681 (N_22681,N_21311,N_20366);
xnor U22682 (N_22682,N_20379,N_21101);
nand U22683 (N_22683,N_21399,N_21942);
nor U22684 (N_22684,N_21002,N_20302);
xor U22685 (N_22685,N_21927,N_20948);
nand U22686 (N_22686,N_21437,N_21910);
nand U22687 (N_22687,N_20386,N_20806);
or U22688 (N_22688,N_22443,N_21150);
and U22689 (N_22689,N_21330,N_21859);
and U22690 (N_22690,N_21553,N_20532);
nand U22691 (N_22691,N_20500,N_20360);
nor U22692 (N_22692,N_21081,N_20621);
and U22693 (N_22693,N_20652,N_20589);
nor U22694 (N_22694,N_22480,N_21278);
and U22695 (N_22695,N_21356,N_21771);
xor U22696 (N_22696,N_21763,N_20662);
nand U22697 (N_22697,N_20122,N_20640);
and U22698 (N_22698,N_21347,N_21119);
and U22699 (N_22699,N_21400,N_20868);
nand U22700 (N_22700,N_22320,N_21230);
nand U22701 (N_22701,N_22317,N_22377);
and U22702 (N_22702,N_21936,N_21784);
xor U22703 (N_22703,N_21721,N_22089);
or U22704 (N_22704,N_22070,N_22007);
nor U22705 (N_22705,N_21599,N_20553);
and U22706 (N_22706,N_21503,N_20411);
and U22707 (N_22707,N_20051,N_21976);
xnor U22708 (N_22708,N_22342,N_20465);
xor U22709 (N_22709,N_21630,N_22234);
or U22710 (N_22710,N_20821,N_21157);
nor U22711 (N_22711,N_20503,N_22014);
nor U22712 (N_22712,N_20256,N_21030);
nand U22713 (N_22713,N_22246,N_21881);
nand U22714 (N_22714,N_22251,N_20443);
or U22715 (N_22715,N_20538,N_20003);
or U22716 (N_22716,N_20985,N_21359);
xor U22717 (N_22717,N_21684,N_21644);
or U22718 (N_22718,N_20091,N_21961);
or U22719 (N_22719,N_21587,N_22306);
or U22720 (N_22720,N_20055,N_20919);
xor U22721 (N_22721,N_20715,N_21950);
xor U22722 (N_22722,N_20508,N_21147);
or U22723 (N_22723,N_21235,N_21786);
nand U22724 (N_22724,N_20692,N_20088);
or U22725 (N_22725,N_21560,N_20326);
or U22726 (N_22726,N_20206,N_21031);
and U22727 (N_22727,N_20481,N_20912);
nor U22728 (N_22728,N_21884,N_22028);
xor U22729 (N_22729,N_20520,N_21980);
xor U22730 (N_22730,N_21113,N_20814);
xnor U22731 (N_22731,N_21502,N_21891);
xor U22732 (N_22732,N_20684,N_21690);
or U22733 (N_22733,N_22297,N_21646);
nor U22734 (N_22734,N_20087,N_20341);
nor U22735 (N_22735,N_20936,N_21952);
nor U22736 (N_22736,N_20669,N_20727);
nor U22737 (N_22737,N_22451,N_20661);
nor U22738 (N_22738,N_21212,N_21233);
nor U22739 (N_22739,N_21534,N_22412);
and U22740 (N_22740,N_20113,N_20450);
xor U22741 (N_22741,N_22076,N_21361);
xor U22742 (N_22742,N_21893,N_21574);
xor U22743 (N_22743,N_22485,N_22180);
nand U22744 (N_22744,N_20178,N_21360);
nor U22745 (N_22745,N_21258,N_21303);
nand U22746 (N_22746,N_21920,N_22460);
and U22747 (N_22747,N_21094,N_20061);
xor U22748 (N_22748,N_21352,N_20253);
nand U22749 (N_22749,N_20712,N_20548);
xor U22750 (N_22750,N_20677,N_21829);
or U22751 (N_22751,N_22204,N_22219);
nor U22752 (N_22752,N_20531,N_20839);
or U22753 (N_22753,N_21290,N_21090);
xor U22754 (N_22754,N_20647,N_21875);
nand U22755 (N_22755,N_20361,N_21046);
nor U22756 (N_22756,N_22446,N_22022);
or U22757 (N_22757,N_22105,N_20160);
xnor U22758 (N_22758,N_21578,N_20653);
nor U22759 (N_22759,N_20342,N_21536);
nand U22760 (N_22760,N_22108,N_20518);
and U22761 (N_22761,N_20136,N_20472);
xnor U22762 (N_22762,N_21415,N_20348);
nor U22763 (N_22763,N_20244,N_22093);
or U22764 (N_22764,N_20773,N_20699);
xor U22765 (N_22765,N_20630,N_20191);
nand U22766 (N_22766,N_22399,N_21364);
xor U22767 (N_22767,N_21386,N_20075);
xor U22768 (N_22768,N_21251,N_21044);
and U22769 (N_22769,N_21153,N_20863);
and U22770 (N_22770,N_20881,N_20332);
xnor U22771 (N_22771,N_20410,N_20164);
or U22772 (N_22772,N_20809,N_21558);
nand U22773 (N_22773,N_21062,N_21267);
xor U22774 (N_22774,N_21729,N_20298);
nor U22775 (N_22775,N_22375,N_21231);
nor U22776 (N_22776,N_20202,N_21140);
or U22777 (N_22777,N_20171,N_22341);
or U22778 (N_22778,N_20798,N_22097);
nor U22779 (N_22779,N_20425,N_22339);
and U22780 (N_22780,N_22328,N_20197);
xnor U22781 (N_22781,N_20331,N_21042);
xor U22782 (N_22782,N_20620,N_22213);
and U22783 (N_22783,N_20031,N_20776);
xnor U22784 (N_22784,N_20844,N_20534);
nor U22785 (N_22785,N_20751,N_22103);
nor U22786 (N_22786,N_21145,N_20231);
nand U22787 (N_22787,N_20689,N_21527);
nor U22788 (N_22788,N_22045,N_22473);
nand U22789 (N_22789,N_22338,N_21713);
xor U22790 (N_22790,N_20916,N_22035);
nor U22791 (N_22791,N_21897,N_20259);
and U22792 (N_22792,N_21286,N_20190);
xnor U22793 (N_22793,N_20085,N_21391);
xnor U22794 (N_22794,N_20047,N_20528);
and U22795 (N_22795,N_20096,N_21279);
or U22796 (N_22796,N_22171,N_20364);
xnor U22797 (N_22797,N_21658,N_22463);
nor U22798 (N_22798,N_20530,N_20943);
nand U22799 (N_22799,N_21928,N_22475);
xnor U22800 (N_22800,N_21281,N_22132);
nor U22801 (N_22801,N_21026,N_21158);
nor U22802 (N_22802,N_22252,N_20129);
xor U22803 (N_22803,N_22457,N_21282);
or U22804 (N_22804,N_20414,N_20890);
xor U22805 (N_22805,N_21500,N_21802);
nand U22806 (N_22806,N_20812,N_21911);
xnor U22807 (N_22807,N_21607,N_20949);
nand U22808 (N_22808,N_20766,N_22018);
xor U22809 (N_22809,N_21638,N_20885);
and U22810 (N_22810,N_21814,N_22113);
xor U22811 (N_22811,N_20902,N_22382);
and U22812 (N_22812,N_22017,N_20232);
or U22813 (N_22813,N_22236,N_20571);
nor U22814 (N_22814,N_22484,N_20053);
nor U22815 (N_22815,N_22046,N_21600);
xnor U22816 (N_22816,N_20734,N_20724);
or U22817 (N_22817,N_20409,N_21535);
nand U22818 (N_22818,N_21862,N_21836);
nand U22819 (N_22819,N_20250,N_20344);
and U22820 (N_22820,N_21102,N_22188);
nor U22821 (N_22821,N_20400,N_20158);
nand U22822 (N_22822,N_21214,N_20596);
nand U22823 (N_22823,N_22174,N_20242);
xnor U22824 (N_22824,N_21997,N_21720);
xnor U22825 (N_22825,N_22197,N_20385);
nand U22826 (N_22826,N_22117,N_21709);
nand U22827 (N_22827,N_21038,N_22243);
xnor U22828 (N_22828,N_21027,N_21354);
xnor U22829 (N_22829,N_22343,N_20700);
or U22830 (N_22830,N_21904,N_21259);
xnor U22831 (N_22831,N_20915,N_22104);
nand U22832 (N_22832,N_22409,N_22413);
xnor U22833 (N_22833,N_21641,N_20709);
nand U22834 (N_22834,N_21710,N_21524);
nand U22835 (N_22835,N_22184,N_20551);
nand U22836 (N_22836,N_22356,N_20560);
nor U22837 (N_22837,N_22223,N_21946);
nand U22838 (N_22838,N_22193,N_20303);
and U22839 (N_22839,N_21367,N_20541);
nand U22840 (N_22840,N_22209,N_22207);
nand U22841 (N_22841,N_21470,N_21803);
nand U22842 (N_22842,N_22052,N_21588);
or U22843 (N_22843,N_20270,N_20431);
nand U22844 (N_22844,N_20907,N_20745);
and U22845 (N_22845,N_20886,N_20350);
nand U22846 (N_22846,N_21099,N_20029);
nor U22847 (N_22847,N_21109,N_21531);
xor U22848 (N_22848,N_21213,N_20079);
or U22849 (N_22849,N_22471,N_20009);
nand U22850 (N_22850,N_21923,N_20010);
or U22851 (N_22851,N_20512,N_20037);
xor U22852 (N_22852,N_20358,N_20968);
nor U22853 (N_22853,N_21477,N_21898);
nand U22854 (N_22854,N_21566,N_20735);
xnor U22855 (N_22855,N_20627,N_20126);
and U22856 (N_22856,N_20991,N_20609);
nand U22857 (N_22857,N_22160,N_20782);
or U22858 (N_22858,N_20290,N_22404);
and U22859 (N_22859,N_22386,N_22405);
or U22860 (N_22860,N_20856,N_22274);
nand U22861 (N_22861,N_20717,N_21466);
or U22862 (N_22862,N_21636,N_20187);
nand U22863 (N_22863,N_21725,N_20613);
nand U22864 (N_22864,N_20804,N_21079);
nand U22865 (N_22865,N_20156,N_20914);
nor U22866 (N_22866,N_21767,N_22192);
xnor U22867 (N_22867,N_20872,N_20624);
xnor U22868 (N_22868,N_20338,N_22438);
xor U22869 (N_22869,N_21979,N_22440);
nor U22870 (N_22870,N_22456,N_22477);
or U22871 (N_22871,N_22228,N_20033);
or U22872 (N_22872,N_21779,N_20134);
or U22873 (N_22873,N_20827,N_20723);
nor U22874 (N_22874,N_22325,N_22368);
or U22875 (N_22875,N_21210,N_20792);
and U22876 (N_22876,N_22101,N_21273);
or U22877 (N_22877,N_22167,N_20737);
and U22878 (N_22878,N_21823,N_21695);
and U22879 (N_22879,N_22275,N_20658);
nand U22880 (N_22880,N_21673,N_22313);
xor U22881 (N_22881,N_20246,N_20208);
nor U22882 (N_22882,N_20989,N_20123);
or U22883 (N_22883,N_20107,N_22235);
or U22884 (N_22884,N_20306,N_20174);
and U22885 (N_22885,N_21271,N_21992);
xor U22886 (N_22886,N_20073,N_20076);
nand U22887 (N_22887,N_21506,N_21488);
and U22888 (N_22888,N_21169,N_22114);
nor U22889 (N_22889,N_21945,N_20217);
or U22890 (N_22890,N_21317,N_22289);
nor U22891 (N_22891,N_20655,N_20098);
nor U22892 (N_22892,N_21083,N_20852);
nand U22893 (N_22893,N_22000,N_21341);
and U22894 (N_22894,N_21783,N_21831);
or U22895 (N_22895,N_21333,N_22276);
or U22896 (N_22896,N_20946,N_20314);
nor U22897 (N_22897,N_21139,N_21043);
xnor U22898 (N_22898,N_22237,N_22131);
nor U22899 (N_22899,N_20488,N_21086);
nor U22900 (N_22900,N_20034,N_22085);
or U22901 (N_22901,N_22314,N_20606);
and U22902 (N_22902,N_22165,N_21318);
nor U22903 (N_22903,N_22491,N_20649);
xor U22904 (N_22904,N_20874,N_21616);
xnor U22905 (N_22905,N_21793,N_20796);
xnor U22906 (N_22906,N_21185,N_21513);
nor U22907 (N_22907,N_21272,N_21672);
xnor U22908 (N_22908,N_21387,N_20861);
nor U22909 (N_22909,N_21379,N_20265);
nor U22910 (N_22910,N_20903,N_22425);
nand U22911 (N_22911,N_21439,N_20956);
xor U22912 (N_22912,N_20335,N_20408);
xnor U22913 (N_22913,N_22227,N_22421);
nor U22914 (N_22914,N_20697,N_21196);
or U22915 (N_22915,N_20163,N_20143);
and U22916 (N_22916,N_20533,N_21481);
or U22917 (N_22917,N_20719,N_20795);
and U22918 (N_22918,N_20923,N_22138);
nor U22919 (N_22919,N_22374,N_21402);
or U22920 (N_22920,N_22240,N_21288);
xnor U22921 (N_22921,N_21965,N_22109);
xor U22922 (N_22922,N_21570,N_20433);
and U22923 (N_22923,N_21161,N_21657);
xnor U22924 (N_22924,N_21675,N_22476);
xnor U22925 (N_22925,N_20865,N_22376);
and U22926 (N_22926,N_22470,N_21325);
nand U22927 (N_22927,N_21870,N_20958);
and U22928 (N_22928,N_22268,N_22288);
nor U22929 (N_22929,N_21476,N_20670);
and U22930 (N_22930,N_21598,N_21873);
xnor U22931 (N_22931,N_20832,N_20755);
and U22932 (N_22932,N_20039,N_20628);
xor U22933 (N_22933,N_21112,N_21422);
nor U22934 (N_22934,N_21671,N_20869);
nor U22935 (N_22935,N_22278,N_22407);
nor U22936 (N_22936,N_20605,N_20278);
xor U22937 (N_22937,N_20336,N_21908);
and U22938 (N_22938,N_20345,N_20554);
and U22939 (N_22939,N_22277,N_20580);
or U22940 (N_22940,N_20367,N_21498);
nand U22941 (N_22941,N_22329,N_20315);
nand U22942 (N_22942,N_20974,N_20860);
nor U22943 (N_22943,N_21841,N_21033);
xor U22944 (N_22944,N_21425,N_20468);
xor U22945 (N_22945,N_22099,N_21653);
or U22946 (N_22946,N_20941,N_20304);
nand U22947 (N_22947,N_20254,N_22107);
nand U22948 (N_22948,N_22263,N_21482);
xor U22949 (N_22949,N_21572,N_20742);
or U22950 (N_22950,N_22319,N_20939);
xnor U22951 (N_22951,N_20920,N_21121);
xnor U22952 (N_22952,N_22003,N_22144);
xnor U22953 (N_22953,N_21619,N_21606);
nor U22954 (N_22954,N_20957,N_21135);
or U22955 (N_22955,N_20642,N_22189);
xor U22956 (N_22956,N_20093,N_20060);
and U22957 (N_22957,N_21530,N_20299);
and U22958 (N_22958,N_20545,N_21663);
and U22959 (N_22959,N_22190,N_21329);
and U22960 (N_22960,N_20285,N_22366);
nand U22961 (N_22961,N_22157,N_21448);
nand U22962 (N_22962,N_21547,N_22392);
or U22963 (N_22963,N_21843,N_20808);
or U22964 (N_22964,N_21155,N_20822);
nand U22965 (N_22965,N_20866,N_21844);
nand U22966 (N_22966,N_22242,N_22151);
xnor U22967 (N_22967,N_20787,N_21762);
or U22968 (N_22968,N_21050,N_21523);
nor U22969 (N_22969,N_21546,N_22027);
nand U22970 (N_22970,N_21339,N_20721);
and U22971 (N_22971,N_22042,N_20783);
and U22972 (N_22972,N_21741,N_20255);
xnor U22973 (N_22973,N_20722,N_21239);
xnor U22974 (N_22974,N_20264,N_20477);
nor U22975 (N_22975,N_20139,N_21154);
xor U22976 (N_22976,N_22363,N_20436);
xor U22977 (N_22977,N_20225,N_20894);
nand U22978 (N_22978,N_20698,N_21706);
xor U22979 (N_22979,N_20970,N_20743);
nand U22980 (N_22980,N_20441,N_21757);
xor U22981 (N_22981,N_22058,N_22185);
xnor U22982 (N_22982,N_21863,N_21190);
or U22983 (N_22983,N_21331,N_21819);
or U22984 (N_22984,N_22331,N_21609);
and U22985 (N_22985,N_20058,N_22423);
or U22986 (N_22986,N_21899,N_20801);
or U22987 (N_22987,N_21755,N_20018);
and U22988 (N_22988,N_20911,N_22133);
nand U22989 (N_22989,N_20328,N_20462);
and U22990 (N_22990,N_20566,N_20325);
nor U22991 (N_22991,N_21595,N_21126);
xor U22992 (N_22992,N_20507,N_20600);
nand U22993 (N_22993,N_21772,N_21489);
nor U22994 (N_22994,N_20384,N_20937);
nor U22995 (N_22995,N_21037,N_21602);
or U22996 (N_22996,N_20444,N_20347);
or U22997 (N_22997,N_20416,N_20040);
xor U22998 (N_22998,N_20980,N_20857);
or U22999 (N_22999,N_21842,N_21545);
and U23000 (N_23000,N_21686,N_20167);
or U23001 (N_23001,N_21623,N_21474);
and U23002 (N_23002,N_21526,N_22318);
nor U23003 (N_23003,N_20168,N_22285);
nor U23004 (N_23004,N_20192,N_20682);
nor U23005 (N_23005,N_21504,N_20502);
or U23006 (N_23006,N_21207,N_20301);
nand U23007 (N_23007,N_21308,N_20466);
xnor U23008 (N_23008,N_20042,N_20322);
nand U23009 (N_23009,N_22094,N_20186);
nand U23010 (N_23010,N_20990,N_20678);
or U23011 (N_23011,N_20987,N_21839);
or U23012 (N_23012,N_22437,N_21754);
xnor U23013 (N_23013,N_22015,N_22469);
nand U23014 (N_23014,N_20982,N_22095);
or U23015 (N_23015,N_20119,N_21297);
nand U23016 (N_23016,N_22398,N_21024);
xor U23017 (N_23017,N_21346,N_21882);
xnor U23018 (N_23018,N_20710,N_20449);
and U23019 (N_23019,N_21737,N_22264);
nand U23020 (N_23020,N_20701,N_21590);
and U23021 (N_23021,N_21794,N_20008);
or U23022 (N_23022,N_20595,N_20219);
nand U23023 (N_23023,N_22370,N_20998);
or U23024 (N_23024,N_22287,N_21010);
or U23025 (N_23025,N_20924,N_20452);
nor U23026 (N_23026,N_21744,N_22400);
xor U23027 (N_23027,N_21005,N_20448);
nand U23028 (N_23028,N_21226,N_21639);
xor U23029 (N_23029,N_22323,N_22447);
nor U23030 (N_23030,N_20525,N_21224);
nor U23031 (N_23031,N_22355,N_20853);
xor U23032 (N_23032,N_21035,N_21987);
xnor U23033 (N_23033,N_20736,N_20378);
nand U23034 (N_23034,N_21229,N_20327);
nor U23035 (N_23035,N_21975,N_21565);
and U23036 (N_23036,N_21797,N_20199);
nor U23037 (N_23037,N_21756,N_20077);
nor U23038 (N_23038,N_21872,N_21640);
or U23039 (N_23039,N_21483,N_22153);
xor U23040 (N_23040,N_20594,N_20959);
xor U23041 (N_23041,N_21464,N_22454);
or U23042 (N_23042,N_22140,N_21861);
and U23043 (N_23043,N_21032,N_20704);
and U23044 (N_23044,N_20426,N_20975);
nand U23045 (N_23045,N_22439,N_20140);
and U23046 (N_23046,N_21465,N_20313);
and U23047 (N_23047,N_20262,N_22442);
nor U23048 (N_23048,N_20536,N_21123);
nor U23049 (N_23049,N_21193,N_20992);
and U23050 (N_23050,N_21342,N_22004);
nand U23051 (N_23051,N_21427,N_21938);
and U23052 (N_23052,N_21934,N_21248);
xnor U23053 (N_23053,N_21785,N_20157);
and U23054 (N_23054,N_20146,N_21373);
nor U23055 (N_23055,N_20487,N_21562);
nand U23056 (N_23056,N_21188,N_21745);
xnor U23057 (N_23057,N_21423,N_20818);
nand U23058 (N_23058,N_21774,N_20794);
xnor U23059 (N_23059,N_21255,N_20251);
xnor U23060 (N_23060,N_21141,N_20906);
xor U23061 (N_23061,N_22023,N_22357);
nor U23062 (N_23062,N_21088,N_21254);
and U23063 (N_23063,N_20048,N_20065);
xor U23064 (N_23064,N_21633,N_20741);
and U23065 (N_23065,N_20373,N_21518);
nand U23066 (N_23066,N_22365,N_21838);
and U23067 (N_23067,N_20688,N_22298);
or U23068 (N_23068,N_20330,N_20593);
nor U23069 (N_23069,N_21118,N_21896);
and U23070 (N_23070,N_21731,N_20537);
or U23071 (N_23071,N_20370,N_22472);
and U23072 (N_23072,N_20862,N_20052);
nor U23073 (N_23073,N_21567,N_20917);
nor U23074 (N_23074,N_21256,N_22072);
nand U23075 (N_23075,N_20765,N_20284);
or U23076 (N_23076,N_22041,N_21129);
nor U23077 (N_23077,N_20898,N_20873);
xnor U23078 (N_23078,N_21749,N_21879);
and U23079 (N_23079,N_20165,N_20169);
or U23080 (N_23080,N_22483,N_20603);
or U23081 (N_23081,N_20834,N_21584);
and U23082 (N_23082,N_22364,N_21707);
xnor U23083 (N_23083,N_21575,N_20826);
nand U23084 (N_23084,N_21432,N_20976);
and U23085 (N_23085,N_20112,N_21165);
xnor U23086 (N_23086,N_21683,N_20391);
nand U23087 (N_23087,N_21315,N_21107);
nor U23088 (N_23088,N_21374,N_20474);
nor U23089 (N_23089,N_20195,N_21430);
nor U23090 (N_23090,N_20667,N_20086);
xnor U23091 (N_23091,N_22344,N_22106);
xnor U23092 (N_23092,N_20993,N_20066);
nor U23093 (N_23093,N_20626,N_21485);
xor U23094 (N_23094,N_20768,N_22128);
nand U23095 (N_23095,N_21963,N_20368);
or U23096 (N_23096,N_21699,N_21219);
nor U23097 (N_23097,N_21681,N_21726);
and U23098 (N_23098,N_22261,N_20705);
nand U23099 (N_23099,N_22461,N_20308);
or U23100 (N_23100,N_20691,N_21156);
xor U23101 (N_23101,N_22206,N_20064);
or U23102 (N_23102,N_20359,N_20966);
and U23103 (N_23103,N_21837,N_21472);
nand U23104 (N_23104,N_21396,N_21625);
nand U23105 (N_23105,N_20590,N_22191);
nor U23106 (N_23106,N_22009,N_20813);
nor U23107 (N_23107,N_22432,N_20622);
nand U23108 (N_23108,N_21528,N_20293);
nand U23109 (N_23109,N_20725,N_21092);
or U23110 (N_23110,N_20319,N_21067);
nor U23111 (N_23111,N_21269,N_21867);
and U23112 (N_23112,N_20739,N_21939);
nand U23113 (N_23113,N_21495,N_21821);
and U23114 (N_23114,N_21070,N_21103);
and U23115 (N_23115,N_20438,N_20049);
nand U23116 (N_23116,N_20931,N_21036);
or U23117 (N_23117,N_20687,N_20563);
and U23118 (N_23118,N_22420,N_21344);
xnor U23119 (N_23119,N_20374,N_21462);
nand U23120 (N_23120,N_20889,N_21296);
xnor U23121 (N_23121,N_20241,N_20851);
nor U23122 (N_23122,N_20562,N_21589);
or U23123 (N_23123,N_21049,N_21554);
and U23124 (N_23124,N_21688,N_21781);
and U23125 (N_23125,N_22086,N_21394);
or U23126 (N_23126,N_21974,N_20027);
nand U23127 (N_23127,N_20573,N_20501);
xnor U23128 (N_23128,N_21304,N_21892);
and U23129 (N_23129,N_20786,N_20258);
or U23130 (N_23130,N_20556,N_20352);
nand U23131 (N_23131,N_21249,N_21520);
nand U23132 (N_23132,N_22333,N_20247);
nand U23133 (N_23133,N_20137,N_20988);
xnor U23134 (N_23134,N_21989,N_21063);
and U23135 (N_23135,N_20476,N_21201);
nand U23136 (N_23136,N_20650,N_21612);
or U23137 (N_23137,N_20243,N_21890);
and U23138 (N_23138,N_22426,N_21411);
and U23139 (N_23139,N_21971,N_22120);
and U23140 (N_23140,N_20224,N_20493);
nand U23141 (N_23141,N_20446,N_20651);
or U23142 (N_23142,N_21250,N_21434);
xor U23143 (N_23143,N_20637,N_22422);
xnor U23144 (N_23144,N_21539,N_20579);
and U23145 (N_23145,N_22212,N_20996);
nor U23146 (N_23146,N_20421,N_20471);
and U23147 (N_23147,N_21017,N_20680);
or U23148 (N_23148,N_21242,N_22247);
or U23149 (N_23149,N_21932,N_20757);
xor U23150 (N_23150,N_22396,N_21680);
and U23151 (N_23151,N_20166,N_21041);
xor U23152 (N_23152,N_21421,N_21982);
nand U23153 (N_23153,N_20204,N_20625);
xnor U23154 (N_23154,N_21790,N_20015);
xor U23155 (N_23155,N_22002,N_21097);
nand U23156 (N_23156,N_20656,N_20900);
and U23157 (N_23157,N_20505,N_20540);
nor U23158 (N_23158,N_21077,N_21136);
nor U23159 (N_23159,N_20070,N_22272);
or U23160 (N_23160,N_21401,N_20311);
or U23161 (N_23161,N_20294,N_22294);
xor U23162 (N_23162,N_21232,N_20041);
nand U23163 (N_23163,N_21438,N_21601);
nor U23164 (N_23164,N_20731,N_20777);
xor U23165 (N_23165,N_21813,N_20179);
xnor U23166 (N_23166,N_22308,N_21138);
xor U23167 (N_23167,N_20422,N_22048);
nand U23168 (N_23168,N_22125,N_20355);
nor U23169 (N_23169,N_20756,N_21894);
or U23170 (N_23170,N_21323,N_20184);
nand U23171 (N_23171,N_21778,N_22282);
or U23172 (N_23172,N_20921,N_20418);
and U23173 (N_23173,N_22059,N_22065);
xnor U23174 (N_23174,N_20235,N_21277);
or U23175 (N_23175,N_21029,N_21579);
nand U23176 (N_23176,N_21674,N_22044);
nor U23177 (N_23177,N_21983,N_20480);
nor U23178 (N_23178,N_20028,N_22096);
or U23179 (N_23179,N_22351,N_21807);
and U23180 (N_23180,N_21085,N_21419);
or U23181 (N_23181,N_20961,N_22467);
and U23182 (N_23182,N_22175,N_20173);
and U23183 (N_23183,N_20234,N_21106);
nand U23184 (N_23184,N_21620,N_22435);
xnor U23185 (N_23185,N_21700,N_21603);
and U23186 (N_23186,N_20583,N_20020);
or U23187 (N_23187,N_22079,N_20356);
xor U23188 (N_23188,N_21022,N_20201);
and U23189 (N_23189,N_21782,N_20749);
nor U23190 (N_23190,N_22428,N_21716);
nand U23191 (N_23191,N_21679,N_22337);
nor U23192 (N_23192,N_22441,N_20397);
or U23193 (N_23193,N_20576,N_21066);
xor U23194 (N_23194,N_21299,N_20196);
nand U23195 (N_23195,N_22111,N_20305);
nor U23196 (N_23196,N_22177,N_20429);
and U23197 (N_23197,N_21824,N_21048);
nor U23198 (N_23198,N_20588,N_21114);
nand U23199 (N_23199,N_20427,N_20513);
nand U23200 (N_23200,N_22169,N_20645);
xor U23201 (N_23201,N_21199,N_22182);
and U23202 (N_23202,N_20524,N_21395);
nand U23203 (N_23203,N_20428,N_20430);
and U23204 (N_23204,N_21198,N_21735);
or U23205 (N_23205,N_21635,N_20104);
xor U23206 (N_23206,N_20644,N_22321);
nand U23207 (N_23207,N_20641,N_22203);
nor U23208 (N_23208,N_20267,N_21828);
nand U23209 (N_23209,N_21733,N_20840);
xor U23210 (N_23210,N_20269,N_21622);
or U23211 (N_23211,N_21768,N_20120);
and U23212 (N_23212,N_21200,N_20130);
or U23213 (N_23213,N_21167,N_21850);
or U23214 (N_23214,N_21447,N_21322);
and U23215 (N_23215,N_20389,N_21718);
and U23216 (N_23216,N_20464,N_20623);
nand U23217 (N_23217,N_21064,N_21326);
and U23218 (N_23218,N_20829,N_20676);
nor U23219 (N_23219,N_21093,N_21096);
xor U23220 (N_23220,N_21615,N_21473);
nor U23221 (N_23221,N_21669,N_21866);
nor U23222 (N_23222,N_21458,N_21087);
nand U23223 (N_23223,N_20598,N_21698);
and U23224 (N_23224,N_22024,N_21478);
xnor U23225 (N_23225,N_22124,N_21610);
xor U23226 (N_23226,N_21252,N_22322);
nand U23227 (N_23227,N_22156,N_20599);
nor U23228 (N_23228,N_20245,N_22340);
nor U23229 (N_23229,N_22081,N_20222);
nor U23230 (N_23230,N_21509,N_22211);
nand U23231 (N_23231,N_20484,N_22418);
xnor U23232 (N_23232,N_22498,N_20074);
nor U23233 (N_23233,N_20405,N_20657);
xor U23234 (N_23234,N_20668,N_20965);
and U23235 (N_23235,N_21389,N_20504);
nor U23236 (N_23236,N_21885,N_20111);
nand U23237 (N_23237,N_20006,N_22179);
and U23238 (N_23238,N_20788,N_21418);
xnor U23239 (N_23239,N_20365,N_22496);
nor U23240 (N_23240,N_21054,N_20101);
and U23241 (N_23241,N_21941,N_21775);
or U23242 (N_23242,N_22464,N_20509);
xor U23243 (N_23243,N_21860,N_20933);
xor U23244 (N_23244,N_20215,N_21306);
xnor U23245 (N_23245,N_21557,N_21951);
or U23246 (N_23246,N_21480,N_21905);
nand U23247 (N_23247,N_21492,N_20106);
and U23248 (N_23248,N_20570,N_22239);
or U23249 (N_23249,N_20686,N_21991);
and U23250 (N_23250,N_21738,N_20266);
xor U23251 (N_23251,N_21868,N_21977);
nor U23252 (N_23252,N_20470,N_21314);
nor U23253 (N_23253,N_20261,N_20078);
nor U23254 (N_23254,N_20007,N_22142);
nand U23255 (N_23255,N_20775,N_21701);
and U23256 (N_23256,N_21691,N_21369);
or U23257 (N_23257,N_22408,N_22301);
xor U23258 (N_23258,N_20013,N_21345);
nand U23259 (N_23259,N_21507,N_21298);
nand U23260 (N_23260,N_22379,N_20218);
nor U23261 (N_23261,N_22312,N_20572);
or U23262 (N_23262,N_20228,N_20396);
nand U23263 (N_23263,N_21903,N_22244);
nand U23264 (N_23264,N_22378,N_21581);
nor U23265 (N_23265,N_21146,N_21409);
nand U23266 (N_23266,N_21170,N_21542);
or U23267 (N_23267,N_21160,N_21479);
xor U23268 (N_23268,N_21954,N_20744);
xnor U23269 (N_23269,N_22233,N_21222);
xor U23270 (N_23270,N_21456,N_21175);
and U23271 (N_23271,N_21496,N_20527);
xor U23272 (N_23272,N_22490,N_20321);
nand U23273 (N_23273,N_20895,N_21747);
nand U23274 (N_23274,N_21593,N_22013);
nor U23275 (N_23275,N_20575,N_22217);
xor U23276 (N_23276,N_20648,N_20942);
xor U23277 (N_23277,N_21944,N_20025);
nor U23278 (N_23278,N_22205,N_20257);
xnor U23279 (N_23279,N_20935,N_21984);
xor U23280 (N_23280,N_22090,N_21568);
or U23281 (N_23281,N_20263,N_21336);
or U23282 (N_23282,N_20227,N_21704);
and U23283 (N_23283,N_20859,N_21451);
nor U23284 (N_23284,N_20754,N_20784);
and U23285 (N_23285,N_21321,N_22220);
nor U23286 (N_23286,N_21217,N_22249);
nand U23287 (N_23287,N_21956,N_20412);
or U23288 (N_23288,N_21275,N_22390);
or U23289 (N_23289,N_22032,N_21241);
xnor U23290 (N_23290,N_22488,N_21817);
xnor U23291 (N_23291,N_20769,N_21913);
xnor U23292 (N_23292,N_21993,N_21748);
xnor U23293 (N_23293,N_21227,N_21416);
xor U23294 (N_23294,N_22129,N_20728);
or U23295 (N_23295,N_21808,N_21510);
or U23296 (N_23296,N_21505,N_21343);
nor U23297 (N_23297,N_20297,N_20340);
and U23298 (N_23298,N_21685,N_22139);
and U23299 (N_23299,N_22150,N_20155);
xnor U23300 (N_23300,N_20000,N_21655);
nor U23301 (N_23301,N_21243,N_20116);
nand U23302 (N_23302,N_20268,N_21039);
nor U23303 (N_23303,N_20807,N_20683);
xnor U23304 (N_23304,N_21110,N_22293);
nand U23305 (N_23305,N_20803,N_20702);
nand U23306 (N_23306,N_22402,N_21291);
xor U23307 (N_23307,N_22444,N_20535);
nand U23308 (N_23308,N_20718,N_20938);
nand U23309 (N_23309,N_20802,N_21467);
nand U23310 (N_23310,N_20044,N_21871);
and U23311 (N_23311,N_21075,N_22143);
nor U23312 (N_23312,N_21460,N_22345);
xor U23313 (N_23313,N_22088,N_20978);
or U23314 (N_23314,N_20457,N_22474);
nand U23315 (N_23315,N_21003,N_20440);
xnor U23316 (N_23316,N_22163,N_20550);
xnor U23317 (N_23317,N_22348,N_21596);
nor U23318 (N_23318,N_22481,N_22199);
or U23319 (N_23319,N_20213,N_22468);
xnor U23320 (N_23320,N_20291,N_20211);
and U23321 (N_23321,N_21922,N_20329);
nand U23322 (N_23322,N_22334,N_21811);
or U23323 (N_23323,N_21457,N_20973);
xor U23324 (N_23324,N_20295,N_21365);
and U23325 (N_23325,N_22497,N_20081);
and U23326 (N_23326,N_22250,N_22361);
or U23327 (N_23327,N_21071,N_20696);
or U23328 (N_23328,N_22026,N_22029);
nor U23329 (N_23329,N_21183,N_21902);
and U23330 (N_23330,N_22091,N_22449);
nand U23331 (N_23331,N_20260,N_20343);
nor U23332 (N_23332,N_20732,N_22168);
and U23333 (N_23333,N_21915,N_20607);
xor U23334 (N_23334,N_21569,N_20287);
and U23335 (N_23335,N_21202,N_22279);
nor U23336 (N_23336,N_21463,N_21571);
nor U23337 (N_23337,N_21011,N_20023);
or U23338 (N_23338,N_22459,N_20877);
nor U23339 (N_23339,N_21929,N_21059);
nand U23340 (N_23340,N_20403,N_21393);
or U23341 (N_23341,N_21152,N_21433);
nand U23342 (N_23342,N_20185,N_21732);
or U23343 (N_23343,N_21953,N_21388);
nor U23344 (N_23344,N_20016,N_20610);
and U23345 (N_23345,N_22149,N_21426);
and U23346 (N_23346,N_21900,N_20830);
nor U23347 (N_23347,N_21994,N_21517);
and U23348 (N_23348,N_22384,N_20659);
and U23349 (N_23349,N_20475,N_22115);
nor U23350 (N_23350,N_21776,N_20805);
xor U23351 (N_23351,N_21358,N_20963);
nand U23352 (N_23352,N_20793,N_22176);
or U23353 (N_23353,N_20899,N_21412);
and U23354 (N_23354,N_21730,N_20277);
and U23355 (N_23355,N_21414,N_22311);
nand U23356 (N_23356,N_22417,N_21293);
nor U23357 (N_23357,N_21265,N_20334);
and U23358 (N_23358,N_20631,N_21450);
or U23359 (N_23359,N_20177,N_22134);
xor U23360 (N_23360,N_21151,N_20880);
nand U23361 (N_23361,N_20459,N_20392);
xor U23362 (N_23362,N_22146,N_22074);
nand U23363 (N_23363,N_21264,N_21215);
xor U23364 (N_23364,N_21541,N_22229);
and U23365 (N_23365,N_20665,N_20401);
nand U23366 (N_23366,N_22332,N_20162);
nand U23367 (N_23367,N_20849,N_21289);
nor U23368 (N_23368,N_22290,N_22395);
xnor U23369 (N_23369,N_20771,N_22100);
or U23370 (N_23370,N_21228,N_20517);
xnor U23371 (N_23371,N_21930,N_21280);
nand U23372 (N_23372,N_21328,N_21173);
nor U23373 (N_23373,N_22383,N_20131);
nand U23374 (N_23374,N_20510,N_20791);
xor U23375 (N_23375,N_21512,N_20498);
or U23376 (N_23376,N_20848,N_22302);
or U23377 (N_23377,N_21985,N_21676);
or U23378 (N_23378,N_21664,N_21914);
nand U23379 (N_23379,N_21750,N_21687);
xnor U23380 (N_23380,N_21132,N_21363);
or U23381 (N_23381,N_20932,N_21538);
or U23382 (N_23382,N_22001,N_21431);
or U23383 (N_23383,N_21305,N_22393);
nor U23384 (N_23384,N_20019,N_22073);
xor U23385 (N_23385,N_21637,N_22075);
nor U23386 (N_23386,N_20442,N_20281);
or U23387 (N_23387,N_21846,N_21621);
and U23388 (N_23388,N_22307,N_21760);
xnor U23389 (N_23389,N_21667,N_21007);
nor U23390 (N_23390,N_21935,N_20194);
xor U23391 (N_23391,N_20207,N_21591);
nand U23392 (N_23392,N_21551,N_20357);
nand U23393 (N_23393,N_20909,N_21715);
xor U23394 (N_23394,N_20511,N_21015);
or U23395 (N_23395,N_20884,N_22187);
nand U23396 (N_23396,N_21051,N_22487);
and U23397 (N_23397,N_20994,N_22427);
nand U23398 (N_23398,N_21455,N_22178);
xor U23399 (N_23399,N_20307,N_21398);
or U23400 (N_23400,N_21332,N_21436);
xor U23401 (N_23401,N_22299,N_20240);
nand U23402 (N_23402,N_20740,N_22122);
and U23403 (N_23403,N_20608,N_22127);
or U23404 (N_23404,N_21624,N_22083);
nor U23405 (N_23405,N_22016,N_20758);
nor U23406 (N_23406,N_21268,N_22200);
or U23407 (N_23407,N_21182,N_20478);
or U23408 (N_23408,N_21926,N_22369);
or U23409 (N_23409,N_22482,N_22296);
nor U23410 (N_23410,N_21660,N_20964);
or U23411 (N_23411,N_20567,N_21940);
nand U23412 (N_23412,N_21832,N_20671);
and U23413 (N_23413,N_22305,N_20223);
or U23414 (N_23414,N_20823,N_21561);
xor U23415 (N_23415,N_20879,N_21319);
or U23416 (N_23416,N_22047,N_21221);
nor U23417 (N_23417,N_20035,N_21723);
nor U23418 (N_23418,N_21693,N_20875);
nand U23419 (N_23419,N_21100,N_20934);
and U23420 (N_23420,N_22436,N_20323);
or U23421 (N_23421,N_20618,N_20114);
nor U23422 (N_23422,N_21550,N_21149);
and U23423 (N_23423,N_20482,N_21970);
xnor U23424 (N_23424,N_22465,N_22039);
nand U23425 (N_23425,N_20394,N_21435);
xnor U23426 (N_23426,N_21058,N_21631);
nand U23427 (N_23427,N_20761,N_21108);
or U23428 (N_23428,N_22304,N_20908);
nand U23429 (N_23429,N_21034,N_20543);
nor U23430 (N_23430,N_22283,N_20312);
and U23431 (N_23431,N_22155,N_21773);
or U23432 (N_23432,N_21708,N_21257);
xor U23433 (N_23433,N_21791,N_21471);
xor U23434 (N_23434,N_20616,N_20685);
xor U23435 (N_23435,N_21858,N_21525);
xnor U23436 (N_23436,N_21909,N_21826);
and U23437 (N_23437,N_20490,N_20205);
and U23438 (N_23438,N_21736,N_22388);
nor U23439 (N_23439,N_20062,N_21245);
nor U23440 (N_23440,N_22499,N_20271);
or U23441 (N_23441,N_20790,N_21876);
or U23442 (N_23442,N_20660,N_21537);
or U23443 (N_23443,N_20059,N_20451);
nor U23444 (N_23444,N_21452,N_22269);
nor U23445 (N_23445,N_21018,N_21302);
xor U23446 (N_23446,N_20354,N_21274);
and U23447 (N_23447,N_21845,N_21203);
nand U23448 (N_23448,N_21133,N_21128);
and U23449 (N_23449,N_22057,N_20726);
or U23450 (N_23450,N_20363,N_22154);
nand U23451 (N_23451,N_20453,N_22346);
nor U23452 (N_23452,N_20815,N_20455);
xnor U23453 (N_23453,N_21417,N_20117);
or U23454 (N_23454,N_21643,N_21144);
xor U23455 (N_23455,N_21901,N_22494);
nor U23456 (N_23456,N_21348,N_21065);
or U23457 (N_23457,N_21327,N_20495);
nor U23458 (N_23458,N_22137,N_22195);
xor U23459 (N_23459,N_20672,N_21618);
nand U23460 (N_23460,N_22038,N_21309);
nor U23461 (N_23461,N_22245,N_21301);
xnor U23462 (N_23462,N_21078,N_21580);
nand U23463 (N_23463,N_21886,N_22221);
or U23464 (N_23464,N_20252,N_20030);
nor U23465 (N_23465,N_21670,N_21801);
or U23466 (N_23466,N_21804,N_21758);
or U23467 (N_23467,N_21445,N_21195);
nand U23468 (N_23468,N_20522,N_21405);
nand U23469 (N_23469,N_22450,N_21692);
or U23470 (N_23470,N_21340,N_21353);
nand U23471 (N_23471,N_21069,N_22479);
and U23472 (N_23472,N_21068,N_20611);
nor U23473 (N_23473,N_20212,N_22084);
xor U23474 (N_23474,N_20617,N_20997);
nand U23475 (N_23475,N_21122,N_22385);
nand U23476 (N_23476,N_21127,N_21552);
nand U23477 (N_23477,N_22034,N_22080);
or U23478 (N_23478,N_20154,N_22410);
or U23479 (N_23479,N_21276,N_21429);
nand U23480 (N_23480,N_21947,N_20738);
and U23481 (N_23481,N_21573,N_20730);
and U23482 (N_23482,N_21244,N_20434);
and U23483 (N_23483,N_21851,N_20390);
or U23484 (N_23484,N_20046,N_21211);
or U23485 (N_23485,N_20460,N_21047);
nand U23486 (N_23486,N_20981,N_21366);
nor U23487 (N_23487,N_22141,N_22126);
or U23488 (N_23488,N_21313,N_20333);
or U23489 (N_23489,N_20209,N_22037);
xnor U23490 (N_23490,N_21174,N_21172);
and U23491 (N_23491,N_20759,N_20133);
nand U23492 (N_23492,N_20679,N_21849);
or U23493 (N_23493,N_20967,N_21981);
nor U23494 (N_23494,N_20280,N_21582);
xor U23495 (N_23495,N_21917,N_21021);
nand U23496 (N_23496,N_21703,N_21444);
xnor U23497 (N_23497,N_21350,N_22284);
or U23498 (N_23498,N_21722,N_20102);
nand U23499 (N_23499,N_21194,N_21338);
or U23500 (N_23500,N_20897,N_20972);
nor U23501 (N_23501,N_21131,N_22416);
or U23502 (N_23502,N_21091,N_22208);
and U23503 (N_23503,N_21407,N_20417);
and U23504 (N_23504,N_21084,N_22262);
xor U23505 (N_23505,N_20664,N_22445);
nor U23506 (N_23506,N_20121,N_22493);
nor U23507 (N_23507,N_22224,N_21020);
and U23508 (N_23508,N_22158,N_21008);
and U23509 (N_23509,N_20249,N_22478);
nor U23510 (N_23510,N_20767,N_20149);
or U23511 (N_23511,N_21795,N_21662);
xor U23512 (N_23512,N_22326,N_20969);
or U23513 (N_23513,N_20785,N_20153);
nor U23514 (N_23514,N_21800,N_21514);
and U23515 (N_23515,N_20585,N_21220);
xnor U23516 (N_23516,N_21854,N_20024);
or U23517 (N_23517,N_22121,N_21143);
and U23518 (N_23518,N_21014,N_22315);
xor U23519 (N_23519,N_21300,N_21406);
nor U23520 (N_23520,N_21237,N_21931);
xor U23521 (N_23521,N_20905,N_20110);
xnor U23522 (N_23522,N_21728,N_20986);
or U23523 (N_23523,N_21181,N_20141);
and U23524 (N_23524,N_21469,N_21864);
nand U23525 (N_23525,N_20339,N_21204);
or U23526 (N_23526,N_21869,N_22040);
or U23527 (N_23527,N_20615,N_21661);
and U23528 (N_23528,N_20103,N_21459);
xnor U23529 (N_23529,N_21796,N_20561);
xnor U23530 (N_23530,N_22248,N_22159);
or U23531 (N_23531,N_20952,N_21104);
nand U23532 (N_23532,N_20927,N_20152);
xor U23533 (N_23533,N_20910,N_20125);
nor U23534 (N_23534,N_20483,N_21995);
xnor U23535 (N_23535,N_20193,N_22098);
and U23536 (N_23536,N_20094,N_20750);
or U23537 (N_23537,N_20004,N_21833);
nand U23538 (N_23538,N_21918,N_21766);
xor U23539 (N_23539,N_20346,N_20635);
xnor U23540 (N_23540,N_21865,N_21490);
xnor U23541 (N_23541,N_21544,N_21912);
and U23542 (N_23542,N_20369,N_20214);
and U23543 (N_23543,N_20925,N_21577);
or U23544 (N_23544,N_21777,N_21045);
and U23545 (N_23545,N_21307,N_20032);
or U23546 (N_23546,N_20188,N_21082);
xnor U23547 (N_23547,N_20183,N_20770);
and U23548 (N_23548,N_22286,N_21719);
or U23549 (N_23549,N_22010,N_21292);
nand U23550 (N_23550,N_22064,N_22266);
and U23551 (N_23551,N_20233,N_21449);
or U23552 (N_23552,N_21403,N_20447);
or U23553 (N_23553,N_21028,N_20388);
nor U23554 (N_23554,N_20831,N_20272);
nor U23555 (N_23555,N_20279,N_20636);
and U23556 (N_23556,N_20420,N_20419);
or U23557 (N_23557,N_20693,N_21770);
nor U23558 (N_23558,N_20067,N_22049);
xor U23559 (N_23559,N_21761,N_20707);
or U23560 (N_23560,N_21948,N_20026);
and U23561 (N_23561,N_21263,N_21454);
or U23562 (N_23562,N_20415,N_21654);
xnor U23563 (N_23563,N_20099,N_20318);
nor U23564 (N_23564,N_20587,N_21397);
nor U23565 (N_23565,N_20316,N_20372);
or U23566 (N_23566,N_20381,N_21677);
or U23567 (N_23567,N_20011,N_22145);
and U23568 (N_23568,N_21594,N_21040);
and U23569 (N_23569,N_20816,N_22214);
nor U23570 (N_23570,N_22394,N_22216);
nand U23571 (N_23571,N_21629,N_20555);
xnor U23572 (N_23572,N_20216,N_21189);
or U23573 (N_23573,N_21597,N_22335);
xnor U23574 (N_23574,N_21442,N_21001);
or U23575 (N_23575,N_21632,N_21025);
xnor U23576 (N_23576,N_21958,N_21486);
xnor U23577 (N_23577,N_21076,N_21689);
or U23578 (N_23578,N_20674,N_20983);
xnor U23579 (N_23579,N_22181,N_20054);
and U23580 (N_23580,N_22021,N_21666);
xnor U23581 (N_23581,N_21792,N_21382);
nor U23582 (N_23582,N_20175,N_21968);
nand U23583 (N_23583,N_20456,N_22466);
and U23584 (N_23584,N_21166,N_20858);
xor U23585 (N_23585,N_20491,N_21705);
or U23586 (N_23586,N_20353,N_20147);
or U23587 (N_23587,N_22198,N_20772);
or U23588 (N_23588,N_22358,N_21972);
nand U23589 (N_23589,N_22006,N_22067);
nor U23590 (N_23590,N_21295,N_22350);
nand U23591 (N_23591,N_21385,N_21080);
and U23592 (N_23592,N_21853,N_21746);
and U23593 (N_23593,N_21246,N_20836);
nand U23594 (N_23594,N_20036,N_21073);
nand U23595 (N_23595,N_22381,N_20629);
and U23596 (N_23596,N_21089,N_20871);
nor U23597 (N_23597,N_20746,N_20161);
nor U23598 (N_23598,N_20930,N_21163);
and U23599 (N_23599,N_20056,N_20001);
xor U23600 (N_23600,N_20586,N_21266);
or U23601 (N_23601,N_21180,N_21316);
nor U23602 (N_23602,N_21125,N_22161);
nand U23603 (N_23603,N_20142,N_21508);
nand U23604 (N_23604,N_22430,N_20633);
and U23605 (N_23605,N_20632,N_21847);
nand U23606 (N_23606,N_20288,N_22362);
or U23607 (N_23607,N_22281,N_21822);
and U23608 (N_23608,N_22201,N_22486);
or U23609 (N_23609,N_21806,N_20445);
xnor U23610 (N_23610,N_22062,N_21855);
and U23611 (N_23611,N_20951,N_20105);
nand U23612 (N_23612,N_20529,N_22433);
nor U23613 (N_23613,N_21611,N_20547);
or U23614 (N_23614,N_21130,N_22391);
nand U23615 (N_23615,N_22380,N_21515);
xnor U23616 (N_23616,N_20473,N_20901);
nand U23617 (N_23617,N_20435,N_22434);
and U23618 (N_23618,N_21179,N_22225);
and U23619 (N_23619,N_20763,N_20565);
nor U23620 (N_23620,N_22061,N_21284);
nand U23621 (N_23621,N_20424,N_20127);
xor U23622 (N_23622,N_20838,N_21428);
xnor U23623 (N_23623,N_20523,N_21115);
and U23624 (N_23624,N_22226,N_21016);
and U23625 (N_23625,N_20221,N_22110);
nand U23626 (N_23626,N_21678,N_20182);
nand U23627 (N_23627,N_22254,N_22353);
nand U23628 (N_23628,N_22043,N_22210);
nand U23629 (N_23629,N_21441,N_22025);
and U23630 (N_23630,N_21262,N_21880);
nor U23631 (N_23631,N_22316,N_21453);
and U23632 (N_23632,N_22020,N_21617);
nor U23633 (N_23633,N_20144,N_20841);
nor U23634 (N_23634,N_20971,N_21162);
and U23635 (N_23635,N_21563,N_21978);
xor U23636 (N_23636,N_22455,N_21697);
and U23637 (N_23637,N_20954,N_20014);
and U23638 (N_23638,N_22419,N_22123);
or U23639 (N_23639,N_21916,N_22373);
nand U23640 (N_23640,N_20833,N_20828);
xnor U23641 (N_23641,N_21647,N_22371);
xnor U23642 (N_23642,N_22087,N_20376);
xnor U23643 (N_23643,N_20708,N_21484);
and U23644 (N_23644,N_21765,N_20109);
xnor U23645 (N_23645,N_20578,N_21665);
nand U23646 (N_23646,N_21739,N_21168);
or U23647 (N_23647,N_21627,N_20612);
xor U23648 (N_23648,N_20151,N_20733);
nand U23649 (N_23649,N_20602,N_21134);
nand U23650 (N_23650,N_22170,N_21998);
or U23651 (N_23651,N_20825,N_20398);
nor U23652 (N_23652,N_20800,N_21714);
xnor U23653 (N_23653,N_22258,N_21061);
nor U23654 (N_23654,N_20984,N_21383);
xnor U23655 (N_23655,N_21548,N_21408);
nand U23656 (N_23656,N_22033,N_20349);
and U23657 (N_23657,N_21966,N_21270);
nand U23658 (N_23658,N_20198,N_20663);
or U23659 (N_23659,N_20432,N_20729);
and U23660 (N_23660,N_21650,N_22324);
or U23661 (N_23661,N_22309,N_21682);
nor U23662 (N_23662,N_21769,N_20170);
xor U23663 (N_23663,N_21857,N_20286);
xnor U23664 (N_23664,N_21380,N_22347);
nor U23665 (N_23665,N_20071,N_20150);
nand U23666 (N_23666,N_20317,N_20747);
nand U23667 (N_23667,N_21178,N_20780);
xor U23668 (N_23668,N_21634,N_21187);
nor U23669 (N_23669,N_20654,N_20220);
nand U23670 (N_23670,N_22267,N_20695);
xnor U23671 (N_23671,N_21759,N_22492);
xnor U23672 (N_23672,N_20229,N_20404);
xor U23673 (N_23673,N_21949,N_22389);
nand U23674 (N_23674,N_21378,N_20892);
or U23675 (N_23675,N_22354,N_21184);
nor U23676 (N_23676,N_21809,N_22253);
nand U23677 (N_23677,N_21614,N_22310);
nor U23678 (N_23678,N_22270,N_20546);
xnor U23679 (N_23679,N_22256,N_20005);
nor U23680 (N_23680,N_21218,N_22036);
and U23681 (N_23681,N_20619,N_20273);
and U23682 (N_23682,N_21320,N_20454);
nor U23683 (N_23683,N_22068,N_21848);
xor U23684 (N_23684,N_22411,N_20870);
or U23685 (N_23685,N_21626,N_20706);
nor U23686 (N_23686,N_20236,N_20181);
and U23687 (N_23687,N_20950,N_21835);
and U23688 (N_23688,N_21019,N_20789);
nand U23689 (N_23689,N_20592,N_20226);
nor U23690 (N_23690,N_21111,N_20238);
and U23691 (N_23691,N_20953,N_21906);
xnor U23692 (N_23692,N_22050,N_20752);
nor U23693 (N_23693,N_21177,N_21095);
and U23694 (N_23694,N_20068,N_21586);
nor U23695 (N_23695,N_21519,N_21652);
xnor U23696 (N_23696,N_20022,N_20764);
nor U23697 (N_23697,N_21511,N_20100);
nand U23698 (N_23698,N_22116,N_22196);
and U23699 (N_23699,N_21628,N_20469);
and U23700 (N_23700,N_20819,N_20393);
xor U23701 (N_23701,N_20467,N_21497);
or U23702 (N_23702,N_22397,N_22300);
xnor U23703 (N_23703,N_22401,N_22222);
nor U23704 (N_23704,N_22011,N_21696);
or U23705 (N_23705,N_20574,N_22012);
nand U23706 (N_23706,N_20276,N_20274);
and U23707 (N_23707,N_21556,N_20089);
nand U23708 (N_23708,N_20115,N_20283);
or U23709 (N_23709,N_20581,N_21789);
or U23710 (N_23710,N_21440,N_20320);
xor U23711 (N_23711,N_22202,N_21209);
xor U23712 (N_23712,N_21818,N_21368);
xor U23713 (N_23713,N_21137,N_20643);
xor U23714 (N_23714,N_21648,N_21540);
xnor U23715 (N_23715,N_22173,N_20172);
and U23716 (N_23716,N_21009,N_20842);
and U23717 (N_23717,N_20845,N_22054);
and U23718 (N_23718,N_22172,N_21206);
nor U23719 (N_23719,N_22372,N_21753);
and U23720 (N_23720,N_20492,N_20681);
xor U23721 (N_23721,N_20817,N_21585);
nor U23722 (N_23722,N_21171,N_21312);
nor U23723 (N_23723,N_20138,N_20159);
and U23724 (N_23724,N_20423,N_20977);
and U23725 (N_23725,N_20854,N_20083);
nor U23726 (N_23726,N_21159,N_21957);
or U23727 (N_23727,N_20084,N_21555);
xnor U23728 (N_23728,N_22273,N_21197);
or U23729 (N_23729,N_20820,N_21000);
or U23730 (N_23730,N_22092,N_20582);
nand U23731 (N_23731,N_20200,N_22360);
and U23732 (N_23732,N_21283,N_21605);
nor U23733 (N_23733,N_20760,N_22260);
nand U23734 (N_23734,N_22071,N_20955);
or U23735 (N_23735,N_21967,N_21117);
nand U23736 (N_23736,N_21717,N_20461);
nor U23737 (N_23737,N_20090,N_22082);
or U23738 (N_23738,N_22031,N_21404);
nor U23739 (N_23739,N_20128,N_21780);
nor U23740 (N_23740,N_20282,N_21287);
or U23741 (N_23741,N_20514,N_21377);
and U23742 (N_23742,N_20748,N_21852);
and U23743 (N_23743,N_20399,N_22130);
nor U23744 (N_23744,N_21355,N_21475);
xor U23745 (N_23745,N_22051,N_20506);
xor U23746 (N_23746,N_20762,N_22352);
nand U23747 (N_23747,N_20189,N_21357);
nand U23748 (N_23748,N_21446,N_22336);
nor U23749 (N_23749,N_20377,N_22257);
and U23750 (N_23750,N_22068,N_21732);
xnor U23751 (N_23751,N_21718,N_22300);
nor U23752 (N_23752,N_21572,N_21264);
or U23753 (N_23753,N_22481,N_20816);
and U23754 (N_23754,N_21157,N_20020);
xor U23755 (N_23755,N_21371,N_21043);
nor U23756 (N_23756,N_21785,N_20646);
xnor U23757 (N_23757,N_20217,N_20201);
or U23758 (N_23758,N_22118,N_22207);
nor U23759 (N_23759,N_21864,N_21182);
nor U23760 (N_23760,N_22052,N_22296);
xor U23761 (N_23761,N_21552,N_21141);
and U23762 (N_23762,N_21621,N_21116);
nand U23763 (N_23763,N_20869,N_20365);
nand U23764 (N_23764,N_20228,N_22063);
and U23765 (N_23765,N_21522,N_20326);
nor U23766 (N_23766,N_20765,N_21975);
nand U23767 (N_23767,N_20807,N_20902);
xnor U23768 (N_23768,N_21733,N_22254);
xor U23769 (N_23769,N_21126,N_21390);
or U23770 (N_23770,N_21378,N_22264);
nand U23771 (N_23771,N_20084,N_21915);
or U23772 (N_23772,N_20017,N_20939);
nor U23773 (N_23773,N_22362,N_21686);
xnor U23774 (N_23774,N_21509,N_21662);
nor U23775 (N_23775,N_21686,N_20522);
xnor U23776 (N_23776,N_20037,N_20073);
xnor U23777 (N_23777,N_21405,N_22408);
or U23778 (N_23778,N_21410,N_20675);
nor U23779 (N_23779,N_20234,N_21007);
or U23780 (N_23780,N_21235,N_22017);
nor U23781 (N_23781,N_22072,N_21511);
or U23782 (N_23782,N_21836,N_21451);
nor U23783 (N_23783,N_21422,N_20431);
nand U23784 (N_23784,N_22170,N_21983);
nor U23785 (N_23785,N_20763,N_21034);
and U23786 (N_23786,N_21421,N_20432);
xnor U23787 (N_23787,N_21756,N_21041);
nor U23788 (N_23788,N_22461,N_20738);
or U23789 (N_23789,N_21289,N_21321);
and U23790 (N_23790,N_21175,N_20101);
or U23791 (N_23791,N_22423,N_22365);
and U23792 (N_23792,N_20219,N_21068);
nor U23793 (N_23793,N_21919,N_21634);
nand U23794 (N_23794,N_21425,N_21245);
or U23795 (N_23795,N_20014,N_20323);
xor U23796 (N_23796,N_21216,N_20046);
and U23797 (N_23797,N_21848,N_20596);
xor U23798 (N_23798,N_20542,N_22102);
xor U23799 (N_23799,N_21624,N_21316);
xnor U23800 (N_23800,N_20459,N_20272);
or U23801 (N_23801,N_21133,N_20757);
and U23802 (N_23802,N_20449,N_22499);
or U23803 (N_23803,N_22276,N_20961);
and U23804 (N_23804,N_20418,N_20223);
xnor U23805 (N_23805,N_22181,N_21650);
xor U23806 (N_23806,N_21752,N_21247);
nor U23807 (N_23807,N_22446,N_21723);
nor U23808 (N_23808,N_20278,N_21926);
nor U23809 (N_23809,N_21481,N_21499);
xnor U23810 (N_23810,N_20767,N_20502);
nor U23811 (N_23811,N_22311,N_21832);
xor U23812 (N_23812,N_20792,N_21096);
xor U23813 (N_23813,N_21355,N_22019);
nor U23814 (N_23814,N_21169,N_20368);
nand U23815 (N_23815,N_20436,N_21521);
and U23816 (N_23816,N_21458,N_22263);
xor U23817 (N_23817,N_21247,N_20691);
or U23818 (N_23818,N_20766,N_21989);
nand U23819 (N_23819,N_22097,N_22286);
and U23820 (N_23820,N_21236,N_21595);
or U23821 (N_23821,N_21893,N_22447);
or U23822 (N_23822,N_21669,N_22210);
or U23823 (N_23823,N_20354,N_20183);
or U23824 (N_23824,N_20185,N_21155);
xor U23825 (N_23825,N_20900,N_21329);
nor U23826 (N_23826,N_20004,N_20404);
nand U23827 (N_23827,N_20237,N_22381);
and U23828 (N_23828,N_20103,N_21696);
and U23829 (N_23829,N_22248,N_20205);
or U23830 (N_23830,N_20341,N_22103);
and U23831 (N_23831,N_22431,N_21529);
nor U23832 (N_23832,N_22107,N_20386);
and U23833 (N_23833,N_22125,N_21707);
nor U23834 (N_23834,N_21251,N_22053);
and U23835 (N_23835,N_21209,N_20058);
nor U23836 (N_23836,N_21811,N_21158);
or U23837 (N_23837,N_21138,N_21042);
and U23838 (N_23838,N_22239,N_21507);
xnor U23839 (N_23839,N_20950,N_21695);
nor U23840 (N_23840,N_20460,N_21836);
nor U23841 (N_23841,N_22098,N_22131);
nor U23842 (N_23842,N_22349,N_21892);
xor U23843 (N_23843,N_21511,N_20688);
xnor U23844 (N_23844,N_21663,N_21458);
or U23845 (N_23845,N_20246,N_20381);
or U23846 (N_23846,N_20768,N_20972);
xnor U23847 (N_23847,N_21784,N_22052);
xor U23848 (N_23848,N_21911,N_20502);
nor U23849 (N_23849,N_22211,N_21790);
nor U23850 (N_23850,N_20921,N_21017);
or U23851 (N_23851,N_20113,N_21024);
and U23852 (N_23852,N_20505,N_20046);
and U23853 (N_23853,N_21575,N_20146);
xnor U23854 (N_23854,N_20337,N_20914);
nand U23855 (N_23855,N_21078,N_20916);
and U23856 (N_23856,N_21122,N_21677);
nand U23857 (N_23857,N_20914,N_21386);
nor U23858 (N_23858,N_20974,N_20670);
xor U23859 (N_23859,N_21173,N_21197);
or U23860 (N_23860,N_20134,N_20985);
nand U23861 (N_23861,N_21658,N_20606);
nor U23862 (N_23862,N_20405,N_20204);
and U23863 (N_23863,N_20484,N_22400);
or U23864 (N_23864,N_20207,N_21264);
xor U23865 (N_23865,N_20525,N_21526);
or U23866 (N_23866,N_22067,N_20698);
xnor U23867 (N_23867,N_21847,N_21872);
or U23868 (N_23868,N_21444,N_22149);
or U23869 (N_23869,N_21180,N_22396);
and U23870 (N_23870,N_22254,N_20841);
and U23871 (N_23871,N_20465,N_21473);
xnor U23872 (N_23872,N_21192,N_21140);
or U23873 (N_23873,N_20166,N_20299);
nor U23874 (N_23874,N_21454,N_21926);
or U23875 (N_23875,N_21801,N_20337);
or U23876 (N_23876,N_20220,N_20313);
nor U23877 (N_23877,N_21319,N_20488);
or U23878 (N_23878,N_21875,N_21731);
or U23879 (N_23879,N_20104,N_21748);
nor U23880 (N_23880,N_21613,N_21791);
xnor U23881 (N_23881,N_20752,N_22064);
xor U23882 (N_23882,N_21084,N_20761);
and U23883 (N_23883,N_20059,N_21045);
or U23884 (N_23884,N_22366,N_21171);
xor U23885 (N_23885,N_20303,N_21291);
nor U23886 (N_23886,N_20118,N_20300);
or U23887 (N_23887,N_21589,N_21416);
and U23888 (N_23888,N_20880,N_21901);
nor U23889 (N_23889,N_21739,N_20153);
or U23890 (N_23890,N_22390,N_21076);
nand U23891 (N_23891,N_20824,N_21870);
and U23892 (N_23892,N_20405,N_22180);
nor U23893 (N_23893,N_20175,N_21616);
and U23894 (N_23894,N_20584,N_21948);
xor U23895 (N_23895,N_20927,N_20265);
or U23896 (N_23896,N_20165,N_21437);
nand U23897 (N_23897,N_22323,N_21932);
or U23898 (N_23898,N_20469,N_21005);
nor U23899 (N_23899,N_21834,N_22212);
nor U23900 (N_23900,N_20372,N_21003);
xor U23901 (N_23901,N_21696,N_21929);
xnor U23902 (N_23902,N_20706,N_21370);
and U23903 (N_23903,N_20729,N_21440);
and U23904 (N_23904,N_21060,N_21603);
xnor U23905 (N_23905,N_21938,N_21548);
and U23906 (N_23906,N_20715,N_20445);
and U23907 (N_23907,N_21481,N_20085);
nand U23908 (N_23908,N_20159,N_21195);
and U23909 (N_23909,N_21520,N_20657);
nand U23910 (N_23910,N_21619,N_21909);
nand U23911 (N_23911,N_20987,N_20451);
or U23912 (N_23912,N_20956,N_22042);
nor U23913 (N_23913,N_20088,N_20298);
nand U23914 (N_23914,N_20382,N_20914);
nor U23915 (N_23915,N_20054,N_22331);
xnor U23916 (N_23916,N_21954,N_21132);
nand U23917 (N_23917,N_20659,N_20564);
nand U23918 (N_23918,N_20088,N_22238);
and U23919 (N_23919,N_21769,N_22159);
xnor U23920 (N_23920,N_20671,N_21528);
or U23921 (N_23921,N_21217,N_20662);
nand U23922 (N_23922,N_21418,N_22267);
and U23923 (N_23923,N_21904,N_20296);
and U23924 (N_23924,N_21244,N_20064);
and U23925 (N_23925,N_21692,N_20404);
nand U23926 (N_23926,N_21819,N_21114);
and U23927 (N_23927,N_21359,N_21686);
or U23928 (N_23928,N_20865,N_22187);
and U23929 (N_23929,N_21570,N_22284);
nor U23930 (N_23930,N_21806,N_21091);
or U23931 (N_23931,N_20074,N_20221);
nand U23932 (N_23932,N_20068,N_20025);
and U23933 (N_23933,N_21704,N_21543);
and U23934 (N_23934,N_20100,N_21599);
nor U23935 (N_23935,N_21774,N_22408);
nand U23936 (N_23936,N_20748,N_21821);
and U23937 (N_23937,N_21169,N_22166);
nand U23938 (N_23938,N_20831,N_22479);
and U23939 (N_23939,N_21173,N_22260);
nor U23940 (N_23940,N_21688,N_21233);
and U23941 (N_23941,N_21220,N_21597);
xnor U23942 (N_23942,N_21474,N_21926);
and U23943 (N_23943,N_22467,N_21591);
nand U23944 (N_23944,N_20429,N_22497);
nand U23945 (N_23945,N_21972,N_22021);
nor U23946 (N_23946,N_20344,N_21743);
xor U23947 (N_23947,N_22388,N_21880);
and U23948 (N_23948,N_20930,N_21839);
and U23949 (N_23949,N_22148,N_22127);
and U23950 (N_23950,N_20618,N_22167);
nor U23951 (N_23951,N_21079,N_22278);
nand U23952 (N_23952,N_22311,N_22144);
nor U23953 (N_23953,N_22016,N_20074);
and U23954 (N_23954,N_21634,N_21969);
nand U23955 (N_23955,N_20934,N_21267);
and U23956 (N_23956,N_21143,N_20023);
nand U23957 (N_23957,N_21891,N_20554);
nor U23958 (N_23958,N_20656,N_21683);
and U23959 (N_23959,N_21335,N_21797);
and U23960 (N_23960,N_21888,N_21846);
and U23961 (N_23961,N_21121,N_21611);
and U23962 (N_23962,N_22051,N_21796);
nor U23963 (N_23963,N_20741,N_22128);
nor U23964 (N_23964,N_21441,N_21354);
nor U23965 (N_23965,N_21409,N_20627);
xnor U23966 (N_23966,N_21635,N_22213);
and U23967 (N_23967,N_20502,N_21374);
nand U23968 (N_23968,N_21213,N_20296);
nand U23969 (N_23969,N_21881,N_20779);
nand U23970 (N_23970,N_22297,N_21122);
nor U23971 (N_23971,N_21957,N_21836);
and U23972 (N_23972,N_20746,N_20920);
xor U23973 (N_23973,N_22114,N_21799);
and U23974 (N_23974,N_21430,N_21495);
or U23975 (N_23975,N_20844,N_21791);
xnor U23976 (N_23976,N_21427,N_21035);
or U23977 (N_23977,N_22053,N_21112);
nor U23978 (N_23978,N_22028,N_21483);
nand U23979 (N_23979,N_20331,N_20488);
nor U23980 (N_23980,N_20377,N_20797);
xor U23981 (N_23981,N_21615,N_20527);
xnor U23982 (N_23982,N_20071,N_21275);
and U23983 (N_23983,N_22086,N_22277);
nand U23984 (N_23984,N_21259,N_21102);
nor U23985 (N_23985,N_20341,N_20784);
or U23986 (N_23986,N_21444,N_21679);
nand U23987 (N_23987,N_20840,N_20163);
and U23988 (N_23988,N_20835,N_21704);
or U23989 (N_23989,N_21083,N_20587);
and U23990 (N_23990,N_20022,N_21287);
nor U23991 (N_23991,N_20821,N_20964);
nand U23992 (N_23992,N_22041,N_20791);
and U23993 (N_23993,N_20546,N_20293);
nand U23994 (N_23994,N_22190,N_21595);
nand U23995 (N_23995,N_21278,N_21949);
nor U23996 (N_23996,N_20522,N_20125);
or U23997 (N_23997,N_21892,N_21151);
nor U23998 (N_23998,N_21765,N_20718);
xor U23999 (N_23999,N_20215,N_20557);
or U24000 (N_24000,N_20483,N_21412);
nand U24001 (N_24001,N_20753,N_22467);
or U24002 (N_24002,N_20165,N_20331);
nand U24003 (N_24003,N_22223,N_20671);
nand U24004 (N_24004,N_20474,N_21210);
xor U24005 (N_24005,N_20729,N_21189);
nor U24006 (N_24006,N_21545,N_20940);
nand U24007 (N_24007,N_20624,N_20046);
nand U24008 (N_24008,N_21336,N_20901);
and U24009 (N_24009,N_20388,N_21332);
nand U24010 (N_24010,N_20594,N_20303);
or U24011 (N_24011,N_20943,N_22072);
xor U24012 (N_24012,N_21823,N_20450);
xnor U24013 (N_24013,N_21683,N_21266);
and U24014 (N_24014,N_21135,N_22272);
nand U24015 (N_24015,N_20945,N_22457);
xnor U24016 (N_24016,N_21416,N_20617);
or U24017 (N_24017,N_20229,N_21727);
nand U24018 (N_24018,N_20502,N_21218);
and U24019 (N_24019,N_21703,N_21192);
nand U24020 (N_24020,N_21302,N_20574);
xor U24021 (N_24021,N_21598,N_20922);
xor U24022 (N_24022,N_21308,N_20105);
nor U24023 (N_24023,N_22101,N_21673);
xnor U24024 (N_24024,N_20002,N_21481);
and U24025 (N_24025,N_20702,N_20271);
nor U24026 (N_24026,N_21701,N_22488);
nor U24027 (N_24027,N_20633,N_21557);
and U24028 (N_24028,N_21302,N_20291);
or U24029 (N_24029,N_20576,N_22498);
or U24030 (N_24030,N_20942,N_20663);
nand U24031 (N_24031,N_22121,N_21376);
or U24032 (N_24032,N_21179,N_21009);
and U24033 (N_24033,N_21701,N_20234);
nand U24034 (N_24034,N_21864,N_20498);
nand U24035 (N_24035,N_21175,N_21056);
or U24036 (N_24036,N_21744,N_20813);
or U24037 (N_24037,N_21619,N_20011);
nor U24038 (N_24038,N_21688,N_22156);
nand U24039 (N_24039,N_22403,N_20380);
nand U24040 (N_24040,N_22082,N_20118);
nand U24041 (N_24041,N_21968,N_21625);
or U24042 (N_24042,N_20405,N_20795);
or U24043 (N_24043,N_20304,N_22165);
and U24044 (N_24044,N_21336,N_22322);
nor U24045 (N_24045,N_20449,N_21629);
or U24046 (N_24046,N_21499,N_22341);
or U24047 (N_24047,N_22002,N_21449);
nand U24048 (N_24048,N_21465,N_21776);
xor U24049 (N_24049,N_21524,N_21617);
xnor U24050 (N_24050,N_20386,N_22495);
or U24051 (N_24051,N_21764,N_20151);
nand U24052 (N_24052,N_22016,N_21480);
and U24053 (N_24053,N_20540,N_21015);
and U24054 (N_24054,N_20935,N_22374);
nor U24055 (N_24055,N_21955,N_22054);
and U24056 (N_24056,N_20652,N_21246);
nor U24057 (N_24057,N_20025,N_21570);
xor U24058 (N_24058,N_20888,N_22279);
nand U24059 (N_24059,N_20561,N_21108);
xnor U24060 (N_24060,N_22257,N_21121);
xnor U24061 (N_24061,N_21180,N_22325);
and U24062 (N_24062,N_22376,N_20348);
and U24063 (N_24063,N_20028,N_21801);
or U24064 (N_24064,N_21981,N_20404);
nand U24065 (N_24065,N_20665,N_22350);
xnor U24066 (N_24066,N_21547,N_20683);
or U24067 (N_24067,N_21797,N_20264);
nor U24068 (N_24068,N_21074,N_20263);
or U24069 (N_24069,N_22174,N_20465);
xor U24070 (N_24070,N_21446,N_22192);
nand U24071 (N_24071,N_21282,N_22303);
nand U24072 (N_24072,N_21730,N_20095);
or U24073 (N_24073,N_22224,N_21337);
and U24074 (N_24074,N_20339,N_22014);
xnor U24075 (N_24075,N_21912,N_20005);
nor U24076 (N_24076,N_21555,N_22244);
xor U24077 (N_24077,N_22123,N_20057);
nor U24078 (N_24078,N_21110,N_22096);
or U24079 (N_24079,N_22332,N_22016);
or U24080 (N_24080,N_22161,N_21651);
xor U24081 (N_24081,N_21629,N_21789);
nand U24082 (N_24082,N_21498,N_20194);
nand U24083 (N_24083,N_21556,N_21061);
nor U24084 (N_24084,N_20480,N_21597);
or U24085 (N_24085,N_22121,N_21225);
nor U24086 (N_24086,N_20687,N_20442);
or U24087 (N_24087,N_21944,N_20619);
xor U24088 (N_24088,N_22059,N_20554);
xnor U24089 (N_24089,N_21571,N_22215);
or U24090 (N_24090,N_21246,N_22021);
xnor U24091 (N_24091,N_20864,N_20538);
nor U24092 (N_24092,N_21524,N_22422);
and U24093 (N_24093,N_21509,N_20053);
nor U24094 (N_24094,N_20173,N_22422);
xor U24095 (N_24095,N_21168,N_21489);
nor U24096 (N_24096,N_20676,N_20124);
nor U24097 (N_24097,N_20511,N_21799);
nor U24098 (N_24098,N_22480,N_20513);
xnor U24099 (N_24099,N_20462,N_20693);
xor U24100 (N_24100,N_20217,N_22158);
nor U24101 (N_24101,N_20980,N_20533);
and U24102 (N_24102,N_21358,N_20176);
nor U24103 (N_24103,N_21569,N_20396);
nor U24104 (N_24104,N_20313,N_22172);
nand U24105 (N_24105,N_21278,N_20623);
and U24106 (N_24106,N_20506,N_21664);
xnor U24107 (N_24107,N_20381,N_21919);
and U24108 (N_24108,N_21609,N_21407);
nand U24109 (N_24109,N_20803,N_21364);
nand U24110 (N_24110,N_22051,N_21997);
or U24111 (N_24111,N_21449,N_20292);
xnor U24112 (N_24112,N_21085,N_20649);
nor U24113 (N_24113,N_20976,N_21622);
nand U24114 (N_24114,N_22285,N_20635);
nand U24115 (N_24115,N_22468,N_21620);
and U24116 (N_24116,N_21228,N_20969);
xnor U24117 (N_24117,N_20326,N_20725);
xor U24118 (N_24118,N_21283,N_22230);
and U24119 (N_24119,N_20555,N_20175);
nand U24120 (N_24120,N_20135,N_21631);
and U24121 (N_24121,N_21538,N_21696);
nand U24122 (N_24122,N_20024,N_21477);
nand U24123 (N_24123,N_20487,N_20500);
nor U24124 (N_24124,N_20223,N_22006);
nand U24125 (N_24125,N_22481,N_21832);
and U24126 (N_24126,N_21597,N_20838);
xnor U24127 (N_24127,N_20302,N_20060);
xor U24128 (N_24128,N_20629,N_20446);
or U24129 (N_24129,N_21513,N_20269);
nand U24130 (N_24130,N_20693,N_21119);
xnor U24131 (N_24131,N_22045,N_21011);
xnor U24132 (N_24132,N_22349,N_20206);
and U24133 (N_24133,N_21034,N_20217);
and U24134 (N_24134,N_20148,N_22486);
xnor U24135 (N_24135,N_20484,N_22109);
xor U24136 (N_24136,N_21614,N_21242);
and U24137 (N_24137,N_20473,N_21639);
and U24138 (N_24138,N_21966,N_20808);
nor U24139 (N_24139,N_22283,N_20419);
or U24140 (N_24140,N_21981,N_21960);
or U24141 (N_24141,N_21121,N_21094);
and U24142 (N_24142,N_20136,N_20191);
or U24143 (N_24143,N_21105,N_20801);
nand U24144 (N_24144,N_20606,N_22363);
xor U24145 (N_24145,N_21328,N_21802);
nand U24146 (N_24146,N_21045,N_20649);
nand U24147 (N_24147,N_21062,N_21665);
nand U24148 (N_24148,N_21536,N_22308);
or U24149 (N_24149,N_20529,N_20070);
and U24150 (N_24150,N_20803,N_22346);
nor U24151 (N_24151,N_20935,N_20865);
xnor U24152 (N_24152,N_20791,N_22248);
xor U24153 (N_24153,N_20153,N_22315);
or U24154 (N_24154,N_20572,N_21128);
xor U24155 (N_24155,N_21986,N_21279);
nand U24156 (N_24156,N_21618,N_21622);
or U24157 (N_24157,N_20249,N_20209);
nand U24158 (N_24158,N_20099,N_20222);
or U24159 (N_24159,N_20849,N_22131);
xnor U24160 (N_24160,N_21775,N_22446);
xor U24161 (N_24161,N_21950,N_22224);
nand U24162 (N_24162,N_20116,N_21362);
xnor U24163 (N_24163,N_21672,N_21837);
or U24164 (N_24164,N_21849,N_22182);
or U24165 (N_24165,N_21313,N_21809);
nor U24166 (N_24166,N_20702,N_20618);
and U24167 (N_24167,N_21762,N_20301);
or U24168 (N_24168,N_20796,N_20040);
nand U24169 (N_24169,N_20766,N_21319);
or U24170 (N_24170,N_20351,N_20886);
xnor U24171 (N_24171,N_22089,N_20576);
xor U24172 (N_24172,N_21670,N_21863);
xnor U24173 (N_24173,N_21025,N_20906);
nand U24174 (N_24174,N_22288,N_21153);
xor U24175 (N_24175,N_21177,N_20148);
or U24176 (N_24176,N_21011,N_20842);
nand U24177 (N_24177,N_21290,N_20030);
and U24178 (N_24178,N_20138,N_20413);
xor U24179 (N_24179,N_20887,N_21067);
or U24180 (N_24180,N_20166,N_21675);
and U24181 (N_24181,N_20922,N_21151);
xnor U24182 (N_24182,N_20776,N_21280);
nor U24183 (N_24183,N_21257,N_21162);
and U24184 (N_24184,N_21774,N_20781);
and U24185 (N_24185,N_21171,N_20018);
xor U24186 (N_24186,N_21629,N_21160);
or U24187 (N_24187,N_21576,N_21951);
and U24188 (N_24188,N_20824,N_22207);
nand U24189 (N_24189,N_21528,N_21078);
and U24190 (N_24190,N_21210,N_21279);
nor U24191 (N_24191,N_21384,N_20953);
xnor U24192 (N_24192,N_20335,N_21757);
xor U24193 (N_24193,N_20871,N_20747);
nor U24194 (N_24194,N_20481,N_21132);
xor U24195 (N_24195,N_21648,N_20696);
xor U24196 (N_24196,N_22440,N_21412);
nor U24197 (N_24197,N_21480,N_22119);
and U24198 (N_24198,N_21180,N_22357);
nor U24199 (N_24199,N_22216,N_20197);
and U24200 (N_24200,N_21613,N_21556);
xnor U24201 (N_24201,N_21794,N_20366);
and U24202 (N_24202,N_20659,N_22112);
or U24203 (N_24203,N_21984,N_22444);
and U24204 (N_24204,N_21623,N_20874);
and U24205 (N_24205,N_21758,N_20045);
and U24206 (N_24206,N_20978,N_21865);
nor U24207 (N_24207,N_21798,N_21736);
and U24208 (N_24208,N_22101,N_21791);
xor U24209 (N_24209,N_22369,N_21837);
and U24210 (N_24210,N_22452,N_20502);
xor U24211 (N_24211,N_20311,N_22389);
xnor U24212 (N_24212,N_21003,N_22148);
nor U24213 (N_24213,N_21465,N_20426);
nor U24214 (N_24214,N_21408,N_21740);
and U24215 (N_24215,N_21677,N_20812);
or U24216 (N_24216,N_22224,N_21728);
nand U24217 (N_24217,N_21817,N_20384);
xor U24218 (N_24218,N_21270,N_22137);
nand U24219 (N_24219,N_20699,N_20154);
xor U24220 (N_24220,N_22134,N_20743);
nand U24221 (N_24221,N_21041,N_22116);
xnor U24222 (N_24222,N_21102,N_21576);
or U24223 (N_24223,N_22359,N_21792);
xnor U24224 (N_24224,N_20359,N_20350);
xnor U24225 (N_24225,N_21964,N_21710);
xor U24226 (N_24226,N_20006,N_21950);
nor U24227 (N_24227,N_20080,N_21184);
or U24228 (N_24228,N_22125,N_22166);
or U24229 (N_24229,N_20577,N_20666);
nor U24230 (N_24230,N_20354,N_22161);
nor U24231 (N_24231,N_22140,N_20104);
or U24232 (N_24232,N_21631,N_22309);
nand U24233 (N_24233,N_21691,N_21360);
nor U24234 (N_24234,N_22438,N_21955);
nor U24235 (N_24235,N_20699,N_21655);
xor U24236 (N_24236,N_22196,N_21623);
nand U24237 (N_24237,N_22449,N_22418);
nand U24238 (N_24238,N_20582,N_22141);
nand U24239 (N_24239,N_21000,N_22111);
and U24240 (N_24240,N_22460,N_21436);
nor U24241 (N_24241,N_21017,N_20384);
or U24242 (N_24242,N_22129,N_20384);
nor U24243 (N_24243,N_22102,N_20064);
nand U24244 (N_24244,N_22390,N_22004);
or U24245 (N_24245,N_20588,N_20439);
nand U24246 (N_24246,N_21597,N_20886);
nor U24247 (N_24247,N_20706,N_20218);
or U24248 (N_24248,N_20171,N_21220);
nand U24249 (N_24249,N_20731,N_20133);
or U24250 (N_24250,N_21573,N_21102);
or U24251 (N_24251,N_21309,N_21272);
and U24252 (N_24252,N_20208,N_21234);
nand U24253 (N_24253,N_20473,N_21902);
nor U24254 (N_24254,N_22332,N_22410);
nand U24255 (N_24255,N_21502,N_21587);
nand U24256 (N_24256,N_20353,N_20165);
nor U24257 (N_24257,N_20951,N_21669);
and U24258 (N_24258,N_20009,N_22259);
xnor U24259 (N_24259,N_20457,N_20588);
and U24260 (N_24260,N_22438,N_20220);
xnor U24261 (N_24261,N_22434,N_21937);
xnor U24262 (N_24262,N_20663,N_21023);
or U24263 (N_24263,N_20263,N_21109);
xor U24264 (N_24264,N_20948,N_21802);
or U24265 (N_24265,N_20695,N_21841);
and U24266 (N_24266,N_22373,N_21303);
or U24267 (N_24267,N_20502,N_22053);
or U24268 (N_24268,N_21678,N_22279);
nor U24269 (N_24269,N_21711,N_20386);
nand U24270 (N_24270,N_21614,N_21011);
nand U24271 (N_24271,N_21187,N_20513);
xor U24272 (N_24272,N_20052,N_20774);
nor U24273 (N_24273,N_20676,N_20820);
or U24274 (N_24274,N_21635,N_20060);
nand U24275 (N_24275,N_20307,N_20199);
nor U24276 (N_24276,N_20328,N_21314);
nand U24277 (N_24277,N_20584,N_20771);
and U24278 (N_24278,N_22229,N_21373);
and U24279 (N_24279,N_22159,N_20929);
nor U24280 (N_24280,N_20802,N_21491);
and U24281 (N_24281,N_21044,N_21027);
xnor U24282 (N_24282,N_21608,N_20852);
nand U24283 (N_24283,N_22221,N_21239);
nand U24284 (N_24284,N_22151,N_22282);
xor U24285 (N_24285,N_21292,N_21832);
nor U24286 (N_24286,N_21023,N_20589);
or U24287 (N_24287,N_21797,N_21110);
nand U24288 (N_24288,N_21288,N_20652);
nand U24289 (N_24289,N_21556,N_22318);
and U24290 (N_24290,N_21731,N_21570);
xor U24291 (N_24291,N_20060,N_20103);
or U24292 (N_24292,N_20435,N_21439);
nor U24293 (N_24293,N_20678,N_22321);
and U24294 (N_24294,N_22358,N_22077);
and U24295 (N_24295,N_20239,N_20198);
or U24296 (N_24296,N_22094,N_20981);
and U24297 (N_24297,N_20462,N_20853);
nor U24298 (N_24298,N_21426,N_21850);
xor U24299 (N_24299,N_20647,N_20179);
nor U24300 (N_24300,N_20282,N_21289);
and U24301 (N_24301,N_21703,N_21451);
xor U24302 (N_24302,N_21835,N_20414);
nor U24303 (N_24303,N_21929,N_22118);
xor U24304 (N_24304,N_22284,N_20039);
nand U24305 (N_24305,N_21596,N_20513);
nand U24306 (N_24306,N_21515,N_20832);
xor U24307 (N_24307,N_21097,N_20070);
or U24308 (N_24308,N_22412,N_20542);
and U24309 (N_24309,N_21729,N_21719);
nor U24310 (N_24310,N_20157,N_21639);
xnor U24311 (N_24311,N_21862,N_21867);
xnor U24312 (N_24312,N_20704,N_20022);
and U24313 (N_24313,N_20444,N_20468);
or U24314 (N_24314,N_21322,N_20151);
or U24315 (N_24315,N_21131,N_22260);
and U24316 (N_24316,N_20673,N_22091);
nor U24317 (N_24317,N_20800,N_20724);
nand U24318 (N_24318,N_21206,N_20878);
xor U24319 (N_24319,N_21182,N_22014);
and U24320 (N_24320,N_22400,N_21361);
and U24321 (N_24321,N_21033,N_22270);
and U24322 (N_24322,N_21403,N_21552);
xor U24323 (N_24323,N_21323,N_22074);
nor U24324 (N_24324,N_21525,N_21685);
xnor U24325 (N_24325,N_20414,N_21884);
or U24326 (N_24326,N_20396,N_21648);
and U24327 (N_24327,N_20679,N_21663);
and U24328 (N_24328,N_22329,N_20754);
xnor U24329 (N_24329,N_20366,N_21502);
xor U24330 (N_24330,N_22458,N_20049);
xnor U24331 (N_24331,N_20339,N_22084);
xnor U24332 (N_24332,N_20220,N_21878);
xor U24333 (N_24333,N_20481,N_21639);
nand U24334 (N_24334,N_20906,N_21758);
xor U24335 (N_24335,N_21521,N_21114);
xor U24336 (N_24336,N_21401,N_21823);
nor U24337 (N_24337,N_21322,N_20155);
xnor U24338 (N_24338,N_20129,N_20313);
or U24339 (N_24339,N_22165,N_21935);
nand U24340 (N_24340,N_20712,N_20332);
nand U24341 (N_24341,N_22478,N_20274);
xor U24342 (N_24342,N_20221,N_20940);
xor U24343 (N_24343,N_20831,N_20506);
nor U24344 (N_24344,N_20942,N_21873);
or U24345 (N_24345,N_22183,N_20636);
nand U24346 (N_24346,N_20325,N_21461);
xnor U24347 (N_24347,N_22494,N_20893);
or U24348 (N_24348,N_20575,N_20995);
and U24349 (N_24349,N_22497,N_22394);
xor U24350 (N_24350,N_20848,N_20153);
xnor U24351 (N_24351,N_21551,N_21637);
xor U24352 (N_24352,N_22005,N_21118);
nand U24353 (N_24353,N_20879,N_20159);
xor U24354 (N_24354,N_21525,N_20008);
nor U24355 (N_24355,N_21130,N_20479);
or U24356 (N_24356,N_21454,N_21382);
and U24357 (N_24357,N_22385,N_22375);
nand U24358 (N_24358,N_20989,N_21025);
nand U24359 (N_24359,N_20809,N_21528);
and U24360 (N_24360,N_22057,N_21690);
and U24361 (N_24361,N_21364,N_21582);
nand U24362 (N_24362,N_20943,N_21812);
nand U24363 (N_24363,N_20474,N_21262);
nand U24364 (N_24364,N_21532,N_20695);
or U24365 (N_24365,N_22215,N_20511);
or U24366 (N_24366,N_21294,N_21356);
and U24367 (N_24367,N_22474,N_22264);
nand U24368 (N_24368,N_21939,N_22497);
xor U24369 (N_24369,N_20124,N_22335);
or U24370 (N_24370,N_21015,N_20600);
nand U24371 (N_24371,N_20210,N_20789);
nor U24372 (N_24372,N_20348,N_20058);
nor U24373 (N_24373,N_20609,N_20682);
nand U24374 (N_24374,N_20716,N_20122);
xor U24375 (N_24375,N_22047,N_21014);
or U24376 (N_24376,N_22046,N_20579);
and U24377 (N_24377,N_21618,N_20267);
and U24378 (N_24378,N_20176,N_20559);
or U24379 (N_24379,N_20009,N_21796);
or U24380 (N_24380,N_22120,N_20430);
and U24381 (N_24381,N_20515,N_20594);
nand U24382 (N_24382,N_21873,N_21585);
nor U24383 (N_24383,N_20733,N_20852);
nand U24384 (N_24384,N_21870,N_21775);
nand U24385 (N_24385,N_20188,N_21452);
or U24386 (N_24386,N_21387,N_21767);
or U24387 (N_24387,N_22406,N_20952);
and U24388 (N_24388,N_20965,N_21761);
and U24389 (N_24389,N_20417,N_21610);
nor U24390 (N_24390,N_20669,N_20478);
nand U24391 (N_24391,N_22310,N_21893);
nand U24392 (N_24392,N_22364,N_21423);
or U24393 (N_24393,N_20483,N_22140);
nand U24394 (N_24394,N_22018,N_21110);
xor U24395 (N_24395,N_20392,N_21055);
and U24396 (N_24396,N_22475,N_21064);
and U24397 (N_24397,N_21184,N_20235);
nor U24398 (N_24398,N_20872,N_20095);
or U24399 (N_24399,N_21815,N_21072);
xnor U24400 (N_24400,N_20295,N_20314);
or U24401 (N_24401,N_21536,N_20724);
and U24402 (N_24402,N_20645,N_20105);
and U24403 (N_24403,N_20187,N_22173);
nand U24404 (N_24404,N_20488,N_21015);
and U24405 (N_24405,N_20322,N_22453);
xor U24406 (N_24406,N_20827,N_21408);
nor U24407 (N_24407,N_22298,N_21885);
xor U24408 (N_24408,N_21773,N_21672);
and U24409 (N_24409,N_21691,N_21519);
nand U24410 (N_24410,N_21875,N_22287);
and U24411 (N_24411,N_22219,N_20864);
or U24412 (N_24412,N_22305,N_20557);
nand U24413 (N_24413,N_22099,N_21686);
or U24414 (N_24414,N_21180,N_21840);
and U24415 (N_24415,N_21883,N_21632);
nor U24416 (N_24416,N_22211,N_20101);
or U24417 (N_24417,N_21165,N_20134);
or U24418 (N_24418,N_21694,N_20906);
or U24419 (N_24419,N_20433,N_20110);
and U24420 (N_24420,N_21679,N_20037);
or U24421 (N_24421,N_21456,N_20931);
nor U24422 (N_24422,N_20062,N_22100);
nand U24423 (N_24423,N_20803,N_21530);
nand U24424 (N_24424,N_21566,N_21444);
nand U24425 (N_24425,N_21811,N_22007);
and U24426 (N_24426,N_21708,N_20781);
nand U24427 (N_24427,N_21402,N_20831);
nor U24428 (N_24428,N_22018,N_21445);
nand U24429 (N_24429,N_21172,N_20051);
and U24430 (N_24430,N_21589,N_20678);
nor U24431 (N_24431,N_21860,N_21869);
nand U24432 (N_24432,N_22004,N_20049);
nor U24433 (N_24433,N_20002,N_20845);
and U24434 (N_24434,N_22291,N_20701);
nor U24435 (N_24435,N_21616,N_22398);
xor U24436 (N_24436,N_21418,N_20097);
xor U24437 (N_24437,N_20656,N_20291);
or U24438 (N_24438,N_21967,N_20352);
nand U24439 (N_24439,N_20667,N_21301);
xnor U24440 (N_24440,N_22271,N_20627);
and U24441 (N_24441,N_20008,N_21723);
nand U24442 (N_24442,N_21014,N_20979);
xnor U24443 (N_24443,N_20301,N_20461);
and U24444 (N_24444,N_21950,N_20203);
nor U24445 (N_24445,N_21748,N_21304);
or U24446 (N_24446,N_20274,N_21128);
xor U24447 (N_24447,N_20598,N_22226);
or U24448 (N_24448,N_21776,N_22048);
xor U24449 (N_24449,N_20564,N_21402);
nor U24450 (N_24450,N_20472,N_20683);
or U24451 (N_24451,N_20298,N_20737);
or U24452 (N_24452,N_22345,N_21935);
nand U24453 (N_24453,N_20817,N_21254);
nor U24454 (N_24454,N_20022,N_20924);
xor U24455 (N_24455,N_21112,N_21543);
xnor U24456 (N_24456,N_22237,N_22476);
and U24457 (N_24457,N_21091,N_20558);
or U24458 (N_24458,N_20658,N_21535);
and U24459 (N_24459,N_21939,N_22338);
and U24460 (N_24460,N_21890,N_20454);
nor U24461 (N_24461,N_20236,N_21286);
or U24462 (N_24462,N_20708,N_22051);
and U24463 (N_24463,N_22344,N_20392);
or U24464 (N_24464,N_22160,N_21082);
nand U24465 (N_24465,N_20450,N_20340);
or U24466 (N_24466,N_21118,N_21355);
or U24467 (N_24467,N_20499,N_21628);
and U24468 (N_24468,N_21758,N_20658);
xnor U24469 (N_24469,N_22273,N_20906);
and U24470 (N_24470,N_21299,N_21454);
and U24471 (N_24471,N_22093,N_21685);
nand U24472 (N_24472,N_22048,N_21777);
xnor U24473 (N_24473,N_21967,N_22436);
nor U24474 (N_24474,N_20987,N_20627);
nor U24475 (N_24475,N_21446,N_22095);
xor U24476 (N_24476,N_20633,N_21605);
or U24477 (N_24477,N_20499,N_21018);
and U24478 (N_24478,N_20943,N_22357);
or U24479 (N_24479,N_22242,N_22374);
or U24480 (N_24480,N_22114,N_20993);
nand U24481 (N_24481,N_20028,N_21892);
nand U24482 (N_24482,N_20813,N_22108);
nor U24483 (N_24483,N_21640,N_22178);
nor U24484 (N_24484,N_22450,N_20327);
nor U24485 (N_24485,N_22488,N_22460);
nor U24486 (N_24486,N_21473,N_22498);
nand U24487 (N_24487,N_22462,N_22115);
nor U24488 (N_24488,N_21615,N_21289);
nor U24489 (N_24489,N_20320,N_21035);
or U24490 (N_24490,N_20754,N_20690);
nor U24491 (N_24491,N_21362,N_22313);
xor U24492 (N_24492,N_21949,N_21190);
nor U24493 (N_24493,N_20801,N_22349);
and U24494 (N_24494,N_22166,N_21213);
and U24495 (N_24495,N_21182,N_20102);
and U24496 (N_24496,N_20867,N_20105);
and U24497 (N_24497,N_21878,N_20438);
and U24498 (N_24498,N_20767,N_20664);
nand U24499 (N_24499,N_20281,N_21892);
xnor U24500 (N_24500,N_20678,N_20286);
and U24501 (N_24501,N_21093,N_20486);
and U24502 (N_24502,N_20723,N_20199);
nor U24503 (N_24503,N_22047,N_20367);
nor U24504 (N_24504,N_21302,N_21541);
or U24505 (N_24505,N_21712,N_20958);
or U24506 (N_24506,N_21948,N_20018);
nor U24507 (N_24507,N_21211,N_21167);
nand U24508 (N_24508,N_20032,N_21155);
or U24509 (N_24509,N_20088,N_20812);
and U24510 (N_24510,N_21055,N_22045);
xor U24511 (N_24511,N_20296,N_22422);
nor U24512 (N_24512,N_20343,N_20814);
nor U24513 (N_24513,N_22192,N_20011);
or U24514 (N_24514,N_21793,N_20205);
xnor U24515 (N_24515,N_20621,N_22183);
or U24516 (N_24516,N_20771,N_20399);
nor U24517 (N_24517,N_21400,N_22453);
nand U24518 (N_24518,N_21269,N_21811);
nand U24519 (N_24519,N_21603,N_21483);
nand U24520 (N_24520,N_21982,N_21972);
or U24521 (N_24521,N_20106,N_20078);
and U24522 (N_24522,N_21327,N_21063);
nor U24523 (N_24523,N_20295,N_21876);
or U24524 (N_24524,N_21901,N_21170);
nor U24525 (N_24525,N_21810,N_20358);
nand U24526 (N_24526,N_21119,N_20306);
and U24527 (N_24527,N_21135,N_21499);
or U24528 (N_24528,N_21465,N_21294);
nand U24529 (N_24529,N_20706,N_20908);
nor U24530 (N_24530,N_21961,N_22209);
xnor U24531 (N_24531,N_20278,N_22012);
and U24532 (N_24532,N_22242,N_20739);
nand U24533 (N_24533,N_21513,N_22232);
xnor U24534 (N_24534,N_20396,N_21069);
and U24535 (N_24535,N_20969,N_21819);
nor U24536 (N_24536,N_20407,N_20502);
nand U24537 (N_24537,N_21888,N_20453);
nor U24538 (N_24538,N_21531,N_20159);
or U24539 (N_24539,N_22369,N_20254);
xnor U24540 (N_24540,N_22496,N_20104);
nor U24541 (N_24541,N_21944,N_20581);
nor U24542 (N_24542,N_20461,N_21063);
xnor U24543 (N_24543,N_21659,N_20927);
or U24544 (N_24544,N_22442,N_21746);
nor U24545 (N_24545,N_22474,N_20453);
xor U24546 (N_24546,N_20561,N_21479);
or U24547 (N_24547,N_21624,N_22354);
xnor U24548 (N_24548,N_20473,N_21959);
xor U24549 (N_24549,N_21971,N_20115);
xor U24550 (N_24550,N_20710,N_21203);
and U24551 (N_24551,N_20943,N_20233);
xor U24552 (N_24552,N_22421,N_21028);
xnor U24553 (N_24553,N_20818,N_22467);
nand U24554 (N_24554,N_20337,N_20940);
and U24555 (N_24555,N_20410,N_21657);
and U24556 (N_24556,N_20629,N_20445);
and U24557 (N_24557,N_21596,N_21752);
xor U24558 (N_24558,N_21712,N_21680);
xnor U24559 (N_24559,N_22318,N_21718);
xor U24560 (N_24560,N_21584,N_22042);
and U24561 (N_24561,N_22195,N_22145);
xnor U24562 (N_24562,N_22174,N_21839);
nand U24563 (N_24563,N_22243,N_20548);
nand U24564 (N_24564,N_21264,N_20094);
nand U24565 (N_24565,N_20719,N_22291);
and U24566 (N_24566,N_22186,N_22231);
nand U24567 (N_24567,N_20895,N_21501);
and U24568 (N_24568,N_20105,N_22222);
nor U24569 (N_24569,N_20246,N_21720);
nand U24570 (N_24570,N_21149,N_20468);
and U24571 (N_24571,N_22115,N_20092);
xnor U24572 (N_24572,N_20717,N_21384);
nor U24573 (N_24573,N_22100,N_20238);
nand U24574 (N_24574,N_22221,N_22128);
and U24575 (N_24575,N_20942,N_20474);
nor U24576 (N_24576,N_21913,N_21189);
or U24577 (N_24577,N_21487,N_20729);
nor U24578 (N_24578,N_21021,N_20296);
nand U24579 (N_24579,N_21207,N_21240);
nand U24580 (N_24580,N_21490,N_20483);
xnor U24581 (N_24581,N_21224,N_21962);
and U24582 (N_24582,N_21719,N_21570);
and U24583 (N_24583,N_22219,N_22159);
xor U24584 (N_24584,N_20397,N_21318);
and U24585 (N_24585,N_21930,N_22172);
xor U24586 (N_24586,N_20617,N_20912);
and U24587 (N_24587,N_20304,N_22270);
nand U24588 (N_24588,N_20088,N_20433);
nor U24589 (N_24589,N_21844,N_22185);
nand U24590 (N_24590,N_21141,N_21971);
nand U24591 (N_24591,N_20483,N_21449);
nor U24592 (N_24592,N_22415,N_22499);
xnor U24593 (N_24593,N_22410,N_21976);
nand U24594 (N_24594,N_21767,N_22497);
and U24595 (N_24595,N_22424,N_21090);
nand U24596 (N_24596,N_20395,N_22334);
and U24597 (N_24597,N_21311,N_20100);
xor U24598 (N_24598,N_21444,N_21973);
xor U24599 (N_24599,N_21815,N_21565);
nand U24600 (N_24600,N_22057,N_20235);
nand U24601 (N_24601,N_20029,N_21558);
or U24602 (N_24602,N_22011,N_20465);
nand U24603 (N_24603,N_21973,N_21237);
nor U24604 (N_24604,N_20666,N_21120);
and U24605 (N_24605,N_22483,N_21185);
or U24606 (N_24606,N_20735,N_20376);
nor U24607 (N_24607,N_21208,N_20270);
xnor U24608 (N_24608,N_20685,N_20925);
and U24609 (N_24609,N_21529,N_20346);
and U24610 (N_24610,N_22329,N_21925);
nand U24611 (N_24611,N_21857,N_20453);
nand U24612 (N_24612,N_21110,N_20495);
or U24613 (N_24613,N_20458,N_22468);
nand U24614 (N_24614,N_20670,N_21907);
xnor U24615 (N_24615,N_21174,N_20399);
or U24616 (N_24616,N_22361,N_21327);
and U24617 (N_24617,N_21000,N_20250);
nor U24618 (N_24618,N_20252,N_20321);
nand U24619 (N_24619,N_20520,N_21222);
or U24620 (N_24620,N_21182,N_21263);
xor U24621 (N_24621,N_20421,N_21662);
and U24622 (N_24622,N_20215,N_21058);
xnor U24623 (N_24623,N_20485,N_20735);
nand U24624 (N_24624,N_22124,N_20272);
and U24625 (N_24625,N_20190,N_20662);
nor U24626 (N_24626,N_20714,N_22205);
nor U24627 (N_24627,N_20972,N_20203);
nand U24628 (N_24628,N_21285,N_20827);
or U24629 (N_24629,N_20521,N_20626);
nand U24630 (N_24630,N_22119,N_20556);
xor U24631 (N_24631,N_20532,N_22159);
xnor U24632 (N_24632,N_22114,N_20411);
or U24633 (N_24633,N_21768,N_21917);
xnor U24634 (N_24634,N_22172,N_20527);
and U24635 (N_24635,N_20193,N_22443);
or U24636 (N_24636,N_21845,N_21232);
and U24637 (N_24637,N_20540,N_21597);
nand U24638 (N_24638,N_20301,N_21438);
nand U24639 (N_24639,N_20990,N_21601);
xor U24640 (N_24640,N_22346,N_20980);
xor U24641 (N_24641,N_21974,N_20749);
or U24642 (N_24642,N_20254,N_21323);
xor U24643 (N_24643,N_20084,N_21655);
or U24644 (N_24644,N_21453,N_22434);
nand U24645 (N_24645,N_21551,N_21480);
nand U24646 (N_24646,N_22026,N_21442);
and U24647 (N_24647,N_20606,N_21031);
nand U24648 (N_24648,N_20290,N_20631);
and U24649 (N_24649,N_21643,N_20254);
nand U24650 (N_24650,N_20047,N_20835);
xor U24651 (N_24651,N_21019,N_21584);
nor U24652 (N_24652,N_21687,N_20733);
or U24653 (N_24653,N_20875,N_22238);
nand U24654 (N_24654,N_21934,N_21905);
and U24655 (N_24655,N_21896,N_22218);
nor U24656 (N_24656,N_21124,N_21005);
xor U24657 (N_24657,N_20104,N_21131);
and U24658 (N_24658,N_22077,N_21531);
nand U24659 (N_24659,N_21679,N_20373);
nand U24660 (N_24660,N_22401,N_20756);
xnor U24661 (N_24661,N_22293,N_20046);
xor U24662 (N_24662,N_21324,N_20560);
and U24663 (N_24663,N_21767,N_20534);
xor U24664 (N_24664,N_20758,N_20033);
nand U24665 (N_24665,N_21052,N_20636);
nand U24666 (N_24666,N_21984,N_22197);
nand U24667 (N_24667,N_20800,N_20940);
nor U24668 (N_24668,N_21671,N_20333);
nor U24669 (N_24669,N_22433,N_21193);
and U24670 (N_24670,N_21651,N_21776);
or U24671 (N_24671,N_20322,N_20305);
xnor U24672 (N_24672,N_20943,N_20550);
xor U24673 (N_24673,N_22249,N_21680);
xor U24674 (N_24674,N_20303,N_20257);
nand U24675 (N_24675,N_20814,N_21693);
nand U24676 (N_24676,N_21101,N_21758);
or U24677 (N_24677,N_21599,N_22482);
or U24678 (N_24678,N_21110,N_21578);
nand U24679 (N_24679,N_20016,N_21006);
and U24680 (N_24680,N_20825,N_22409);
or U24681 (N_24681,N_21780,N_22438);
and U24682 (N_24682,N_20700,N_20370);
nand U24683 (N_24683,N_20844,N_20662);
or U24684 (N_24684,N_21974,N_21269);
or U24685 (N_24685,N_21154,N_20908);
nand U24686 (N_24686,N_20327,N_22241);
nand U24687 (N_24687,N_20106,N_21384);
or U24688 (N_24688,N_22362,N_21483);
nor U24689 (N_24689,N_21198,N_21337);
nand U24690 (N_24690,N_22149,N_20324);
nor U24691 (N_24691,N_20613,N_21440);
nor U24692 (N_24692,N_20790,N_20270);
xor U24693 (N_24693,N_20819,N_22404);
xor U24694 (N_24694,N_22226,N_20599);
or U24695 (N_24695,N_21352,N_21116);
xnor U24696 (N_24696,N_20239,N_21558);
and U24697 (N_24697,N_22115,N_22476);
or U24698 (N_24698,N_21544,N_20299);
nand U24699 (N_24699,N_21976,N_20878);
or U24700 (N_24700,N_21955,N_20721);
nor U24701 (N_24701,N_22227,N_20137);
xor U24702 (N_24702,N_20271,N_20317);
xnor U24703 (N_24703,N_22447,N_22448);
nor U24704 (N_24704,N_21675,N_22418);
or U24705 (N_24705,N_21638,N_20555);
or U24706 (N_24706,N_21813,N_21244);
or U24707 (N_24707,N_20230,N_20253);
xor U24708 (N_24708,N_21903,N_20078);
and U24709 (N_24709,N_20743,N_22411);
nand U24710 (N_24710,N_22057,N_20315);
and U24711 (N_24711,N_21131,N_20389);
xor U24712 (N_24712,N_20077,N_21713);
xnor U24713 (N_24713,N_21053,N_22320);
nand U24714 (N_24714,N_20234,N_21524);
or U24715 (N_24715,N_20951,N_20213);
or U24716 (N_24716,N_21904,N_21383);
xor U24717 (N_24717,N_22066,N_20913);
xor U24718 (N_24718,N_22070,N_20937);
nor U24719 (N_24719,N_20047,N_21186);
and U24720 (N_24720,N_20564,N_20798);
xnor U24721 (N_24721,N_22466,N_21943);
xnor U24722 (N_24722,N_21507,N_20705);
or U24723 (N_24723,N_20972,N_20487);
xor U24724 (N_24724,N_21838,N_20536);
and U24725 (N_24725,N_21724,N_21413);
xor U24726 (N_24726,N_21526,N_20809);
or U24727 (N_24727,N_21520,N_20760);
xor U24728 (N_24728,N_20209,N_20537);
nor U24729 (N_24729,N_20805,N_21743);
xor U24730 (N_24730,N_21732,N_21449);
and U24731 (N_24731,N_20134,N_20396);
xor U24732 (N_24732,N_20272,N_20999);
or U24733 (N_24733,N_21213,N_22476);
nand U24734 (N_24734,N_21911,N_21213);
and U24735 (N_24735,N_20902,N_21647);
or U24736 (N_24736,N_20338,N_20460);
or U24737 (N_24737,N_21320,N_21923);
and U24738 (N_24738,N_21487,N_21307);
or U24739 (N_24739,N_20198,N_20152);
nor U24740 (N_24740,N_21747,N_20094);
and U24741 (N_24741,N_22480,N_21102);
or U24742 (N_24742,N_21575,N_20906);
nor U24743 (N_24743,N_21316,N_20285);
nand U24744 (N_24744,N_21215,N_20600);
nor U24745 (N_24745,N_21912,N_21313);
or U24746 (N_24746,N_20430,N_21509);
nor U24747 (N_24747,N_21167,N_21721);
nand U24748 (N_24748,N_20671,N_22260);
nor U24749 (N_24749,N_21411,N_20063);
or U24750 (N_24750,N_20285,N_21624);
nor U24751 (N_24751,N_21154,N_20077);
and U24752 (N_24752,N_20280,N_21417);
nand U24753 (N_24753,N_21378,N_21924);
and U24754 (N_24754,N_20463,N_20806);
nand U24755 (N_24755,N_20017,N_21414);
or U24756 (N_24756,N_20598,N_20610);
or U24757 (N_24757,N_20835,N_21956);
xor U24758 (N_24758,N_21775,N_21318);
nand U24759 (N_24759,N_21973,N_21587);
or U24760 (N_24760,N_20413,N_21067);
xor U24761 (N_24761,N_21729,N_20415);
and U24762 (N_24762,N_22119,N_21008);
nor U24763 (N_24763,N_20180,N_21272);
nor U24764 (N_24764,N_22348,N_22166);
and U24765 (N_24765,N_21268,N_22347);
nand U24766 (N_24766,N_20221,N_21009);
nand U24767 (N_24767,N_20385,N_21650);
nor U24768 (N_24768,N_21069,N_21267);
nand U24769 (N_24769,N_21112,N_20278);
nand U24770 (N_24770,N_21394,N_20959);
nor U24771 (N_24771,N_21613,N_21936);
xnor U24772 (N_24772,N_21965,N_21910);
xor U24773 (N_24773,N_21460,N_21220);
or U24774 (N_24774,N_21796,N_20792);
and U24775 (N_24775,N_21164,N_20598);
xor U24776 (N_24776,N_21575,N_20833);
nand U24777 (N_24777,N_20716,N_21993);
and U24778 (N_24778,N_21615,N_22154);
xnor U24779 (N_24779,N_21289,N_21754);
nand U24780 (N_24780,N_20926,N_20873);
nand U24781 (N_24781,N_21928,N_21831);
xor U24782 (N_24782,N_20256,N_21207);
and U24783 (N_24783,N_20638,N_21000);
xor U24784 (N_24784,N_22468,N_21560);
nand U24785 (N_24785,N_22396,N_21529);
and U24786 (N_24786,N_21125,N_21010);
nand U24787 (N_24787,N_20463,N_20947);
or U24788 (N_24788,N_20579,N_21573);
or U24789 (N_24789,N_22308,N_20964);
or U24790 (N_24790,N_21804,N_22288);
nand U24791 (N_24791,N_22457,N_22232);
and U24792 (N_24792,N_22240,N_20560);
nand U24793 (N_24793,N_21624,N_20232);
xor U24794 (N_24794,N_20934,N_22332);
or U24795 (N_24795,N_22376,N_21679);
nand U24796 (N_24796,N_21760,N_21583);
nand U24797 (N_24797,N_20268,N_20304);
and U24798 (N_24798,N_22371,N_20079);
nand U24799 (N_24799,N_21045,N_22463);
xor U24800 (N_24800,N_20034,N_21509);
xnor U24801 (N_24801,N_21514,N_20505);
nand U24802 (N_24802,N_22387,N_20948);
nand U24803 (N_24803,N_22325,N_22198);
xnor U24804 (N_24804,N_22304,N_21988);
nand U24805 (N_24805,N_21348,N_20362);
nand U24806 (N_24806,N_21127,N_20576);
and U24807 (N_24807,N_22396,N_20131);
nand U24808 (N_24808,N_21213,N_21515);
and U24809 (N_24809,N_21052,N_20978);
nor U24810 (N_24810,N_20008,N_21270);
or U24811 (N_24811,N_21293,N_20237);
nor U24812 (N_24812,N_22097,N_21191);
nor U24813 (N_24813,N_22430,N_20296);
or U24814 (N_24814,N_20893,N_20818);
or U24815 (N_24815,N_21373,N_21399);
or U24816 (N_24816,N_21383,N_21972);
and U24817 (N_24817,N_20034,N_20751);
nor U24818 (N_24818,N_21443,N_20772);
nand U24819 (N_24819,N_21060,N_21567);
nor U24820 (N_24820,N_21335,N_21052);
and U24821 (N_24821,N_20515,N_21946);
nand U24822 (N_24822,N_20567,N_20704);
nand U24823 (N_24823,N_21039,N_20166);
or U24824 (N_24824,N_20370,N_20398);
or U24825 (N_24825,N_21617,N_21730);
xnor U24826 (N_24826,N_20464,N_21386);
nor U24827 (N_24827,N_20777,N_20641);
xnor U24828 (N_24828,N_20314,N_20036);
xnor U24829 (N_24829,N_21243,N_20901);
xor U24830 (N_24830,N_20189,N_21057);
nand U24831 (N_24831,N_22498,N_20892);
nor U24832 (N_24832,N_22413,N_21536);
nor U24833 (N_24833,N_20061,N_22041);
or U24834 (N_24834,N_20803,N_20442);
nor U24835 (N_24835,N_20298,N_21005);
nor U24836 (N_24836,N_21290,N_20814);
and U24837 (N_24837,N_20997,N_20319);
nor U24838 (N_24838,N_20635,N_22486);
nor U24839 (N_24839,N_21747,N_22299);
xor U24840 (N_24840,N_21363,N_21798);
xor U24841 (N_24841,N_21480,N_20447);
and U24842 (N_24842,N_20448,N_20893);
nand U24843 (N_24843,N_21186,N_21496);
nand U24844 (N_24844,N_20099,N_20111);
nand U24845 (N_24845,N_22269,N_22096);
and U24846 (N_24846,N_21107,N_21284);
nand U24847 (N_24847,N_21679,N_21297);
xnor U24848 (N_24848,N_22377,N_20368);
and U24849 (N_24849,N_20737,N_20640);
nand U24850 (N_24850,N_20078,N_22398);
xor U24851 (N_24851,N_20887,N_20061);
nor U24852 (N_24852,N_22487,N_20946);
xor U24853 (N_24853,N_20826,N_20318);
nand U24854 (N_24854,N_22333,N_21705);
or U24855 (N_24855,N_22292,N_22360);
nor U24856 (N_24856,N_22462,N_21033);
or U24857 (N_24857,N_22169,N_20803);
or U24858 (N_24858,N_20482,N_21598);
nand U24859 (N_24859,N_20175,N_20878);
xnor U24860 (N_24860,N_21757,N_21901);
or U24861 (N_24861,N_22468,N_20425);
or U24862 (N_24862,N_20849,N_20914);
xnor U24863 (N_24863,N_21056,N_21954);
and U24864 (N_24864,N_21003,N_22455);
xnor U24865 (N_24865,N_20684,N_22228);
and U24866 (N_24866,N_20256,N_20106);
and U24867 (N_24867,N_21334,N_21825);
xor U24868 (N_24868,N_20211,N_21494);
or U24869 (N_24869,N_21600,N_22300);
and U24870 (N_24870,N_21754,N_21575);
nand U24871 (N_24871,N_21959,N_21284);
nand U24872 (N_24872,N_22052,N_21950);
and U24873 (N_24873,N_21789,N_21188);
and U24874 (N_24874,N_20440,N_20430);
nor U24875 (N_24875,N_22088,N_21800);
or U24876 (N_24876,N_20657,N_21003);
nand U24877 (N_24877,N_21424,N_21998);
nor U24878 (N_24878,N_20812,N_20279);
xor U24879 (N_24879,N_21991,N_21304);
nor U24880 (N_24880,N_22017,N_21148);
or U24881 (N_24881,N_21368,N_21420);
xnor U24882 (N_24882,N_20780,N_22160);
xnor U24883 (N_24883,N_22031,N_21962);
and U24884 (N_24884,N_20049,N_20147);
xnor U24885 (N_24885,N_21823,N_20812);
nand U24886 (N_24886,N_21256,N_20050);
or U24887 (N_24887,N_20760,N_21909);
or U24888 (N_24888,N_20136,N_20946);
xor U24889 (N_24889,N_22249,N_20575);
and U24890 (N_24890,N_21318,N_21558);
xnor U24891 (N_24891,N_20724,N_22115);
or U24892 (N_24892,N_22179,N_21553);
and U24893 (N_24893,N_20119,N_21506);
and U24894 (N_24894,N_22467,N_22216);
nand U24895 (N_24895,N_20156,N_21597);
xnor U24896 (N_24896,N_21362,N_21119);
nor U24897 (N_24897,N_21132,N_20671);
xnor U24898 (N_24898,N_20204,N_21567);
or U24899 (N_24899,N_20540,N_21891);
nand U24900 (N_24900,N_21251,N_21433);
nor U24901 (N_24901,N_20824,N_21407);
and U24902 (N_24902,N_20858,N_20296);
nor U24903 (N_24903,N_21821,N_22475);
or U24904 (N_24904,N_21183,N_21067);
and U24905 (N_24905,N_22450,N_22308);
xor U24906 (N_24906,N_20575,N_21439);
nor U24907 (N_24907,N_20573,N_22441);
xnor U24908 (N_24908,N_21468,N_21079);
or U24909 (N_24909,N_22193,N_20089);
and U24910 (N_24910,N_22139,N_20096);
xnor U24911 (N_24911,N_22116,N_20630);
xnor U24912 (N_24912,N_21312,N_21245);
xnor U24913 (N_24913,N_20870,N_20620);
nor U24914 (N_24914,N_22404,N_20638);
or U24915 (N_24915,N_21561,N_21911);
or U24916 (N_24916,N_21711,N_22015);
and U24917 (N_24917,N_21695,N_20184);
xor U24918 (N_24918,N_22119,N_22017);
or U24919 (N_24919,N_20200,N_20886);
nor U24920 (N_24920,N_22045,N_20774);
or U24921 (N_24921,N_21308,N_22335);
and U24922 (N_24922,N_21989,N_20642);
nor U24923 (N_24923,N_20425,N_21539);
xor U24924 (N_24924,N_20847,N_20295);
xor U24925 (N_24925,N_20746,N_20740);
nor U24926 (N_24926,N_21840,N_21185);
or U24927 (N_24927,N_20252,N_21363);
and U24928 (N_24928,N_21086,N_21895);
xnor U24929 (N_24929,N_20925,N_20964);
nor U24930 (N_24930,N_20234,N_20559);
xnor U24931 (N_24931,N_22407,N_20008);
nor U24932 (N_24932,N_21168,N_21750);
nand U24933 (N_24933,N_20243,N_22372);
nand U24934 (N_24934,N_21508,N_22266);
or U24935 (N_24935,N_21253,N_22346);
or U24936 (N_24936,N_20636,N_20448);
xnor U24937 (N_24937,N_22314,N_22325);
nand U24938 (N_24938,N_20992,N_21276);
nand U24939 (N_24939,N_20080,N_20966);
nor U24940 (N_24940,N_20221,N_22388);
xnor U24941 (N_24941,N_22221,N_22214);
and U24942 (N_24942,N_21424,N_22490);
nor U24943 (N_24943,N_20371,N_20413);
and U24944 (N_24944,N_20684,N_20128);
xor U24945 (N_24945,N_21244,N_22373);
nand U24946 (N_24946,N_21797,N_21029);
and U24947 (N_24947,N_20625,N_20081);
nand U24948 (N_24948,N_22096,N_20515);
and U24949 (N_24949,N_21064,N_21508);
or U24950 (N_24950,N_20591,N_22099);
nand U24951 (N_24951,N_21448,N_21975);
xor U24952 (N_24952,N_21172,N_20129);
xor U24953 (N_24953,N_22066,N_21106);
or U24954 (N_24954,N_22354,N_21464);
or U24955 (N_24955,N_21222,N_20319);
and U24956 (N_24956,N_21934,N_21480);
nand U24957 (N_24957,N_20698,N_20892);
nor U24958 (N_24958,N_20445,N_20353);
nand U24959 (N_24959,N_21121,N_22060);
and U24960 (N_24960,N_20881,N_20055);
nor U24961 (N_24961,N_20171,N_20428);
and U24962 (N_24962,N_20165,N_21738);
nor U24963 (N_24963,N_20955,N_21845);
and U24964 (N_24964,N_20388,N_21022);
xor U24965 (N_24965,N_21096,N_21087);
or U24966 (N_24966,N_20183,N_21970);
and U24967 (N_24967,N_21998,N_20383);
nand U24968 (N_24968,N_21238,N_21424);
nand U24969 (N_24969,N_20984,N_21756);
nand U24970 (N_24970,N_20586,N_21386);
and U24971 (N_24971,N_20547,N_20053);
and U24972 (N_24972,N_21441,N_22167);
nor U24973 (N_24973,N_20093,N_20246);
nor U24974 (N_24974,N_22481,N_20806);
nor U24975 (N_24975,N_22430,N_21453);
or U24976 (N_24976,N_20977,N_21701);
xor U24977 (N_24977,N_22022,N_20398);
or U24978 (N_24978,N_22249,N_20124);
xnor U24979 (N_24979,N_21418,N_22305);
nand U24980 (N_24980,N_21731,N_21668);
and U24981 (N_24981,N_20847,N_20239);
or U24982 (N_24982,N_22080,N_21754);
nand U24983 (N_24983,N_21652,N_22155);
and U24984 (N_24984,N_22408,N_22285);
xnor U24985 (N_24985,N_20321,N_21839);
or U24986 (N_24986,N_21377,N_20227);
nand U24987 (N_24987,N_20673,N_20769);
nor U24988 (N_24988,N_20485,N_22096);
and U24989 (N_24989,N_20663,N_20528);
and U24990 (N_24990,N_22203,N_20587);
and U24991 (N_24991,N_21820,N_22366);
or U24992 (N_24992,N_20585,N_20897);
xor U24993 (N_24993,N_22479,N_20528);
xnor U24994 (N_24994,N_21305,N_22004);
xnor U24995 (N_24995,N_20389,N_20473);
and U24996 (N_24996,N_22402,N_21425);
xnor U24997 (N_24997,N_20795,N_22197);
xnor U24998 (N_24998,N_21010,N_20939);
xnor U24999 (N_24999,N_20055,N_20701);
nor UO_0 (O_0,N_24380,N_22973);
xor UO_1 (O_1,N_24096,N_22612);
or UO_2 (O_2,N_24200,N_24420);
nor UO_3 (O_3,N_23185,N_23349);
xnor UO_4 (O_4,N_24386,N_24730);
or UO_5 (O_5,N_24383,N_24019);
xnor UO_6 (O_6,N_23175,N_24795);
xnor UO_7 (O_7,N_24761,N_23042);
and UO_8 (O_8,N_24458,N_22515);
or UO_9 (O_9,N_24174,N_23062);
or UO_10 (O_10,N_23144,N_23098);
nand UO_11 (O_11,N_24493,N_23207);
nand UO_12 (O_12,N_23549,N_23463);
nor UO_13 (O_13,N_23842,N_24496);
or UO_14 (O_14,N_24506,N_24508);
and UO_15 (O_15,N_22746,N_23634);
nor UO_16 (O_16,N_23196,N_23419);
or UO_17 (O_17,N_23749,N_23069);
and UO_18 (O_18,N_24548,N_23688);
nand UO_19 (O_19,N_24712,N_22638);
and UO_20 (O_20,N_24707,N_23570);
nand UO_21 (O_21,N_24047,N_24612);
or UO_22 (O_22,N_23183,N_23600);
xor UO_23 (O_23,N_23981,N_23537);
or UO_24 (O_24,N_23929,N_24491);
nand UO_25 (O_25,N_24071,N_24819);
or UO_26 (O_26,N_24594,N_24361);
and UO_27 (O_27,N_24466,N_22866);
and UO_28 (O_28,N_24020,N_24518);
xnor UO_29 (O_29,N_24510,N_23885);
or UO_30 (O_30,N_24823,N_24624);
and UO_31 (O_31,N_24989,N_24043);
nand UO_32 (O_32,N_24341,N_23230);
nor UO_33 (O_33,N_24643,N_24093);
nor UO_34 (O_34,N_23064,N_24159);
or UO_35 (O_35,N_23732,N_22628);
xnor UO_36 (O_36,N_22917,N_23912);
or UO_37 (O_37,N_22908,N_24303);
and UO_38 (O_38,N_23123,N_22933);
or UO_39 (O_39,N_23642,N_22873);
nor UO_40 (O_40,N_22928,N_22969);
xnor UO_41 (O_41,N_23938,N_23339);
and UO_42 (O_42,N_23477,N_24562);
xor UO_43 (O_43,N_23414,N_23913);
nand UO_44 (O_44,N_24099,N_23375);
nand UO_45 (O_45,N_24297,N_24088);
or UO_46 (O_46,N_23485,N_24404);
and UO_47 (O_47,N_22957,N_23168);
nor UO_48 (O_48,N_23193,N_23934);
and UO_49 (O_49,N_22966,N_23776);
and UO_50 (O_50,N_24902,N_24275);
and UO_51 (O_51,N_23517,N_22899);
or UO_52 (O_52,N_22802,N_22841);
and UO_53 (O_53,N_24340,N_24324);
nand UO_54 (O_54,N_22632,N_22926);
or UO_55 (O_55,N_23927,N_24217);
or UO_56 (O_56,N_24193,N_22907);
nand UO_57 (O_57,N_24842,N_23143);
xor UO_58 (O_58,N_24015,N_23733);
nor UO_59 (O_59,N_22567,N_24391);
and UO_60 (O_60,N_23678,N_24641);
nand UO_61 (O_61,N_23614,N_24547);
nand UO_62 (O_62,N_24978,N_24794);
or UO_63 (O_63,N_23918,N_23280);
nor UO_64 (O_64,N_22674,N_24500);
nand UO_65 (O_65,N_23910,N_22843);
xor UO_66 (O_66,N_24938,N_22665);
or UO_67 (O_67,N_24559,N_23886);
nand UO_68 (O_68,N_23294,N_24481);
nor UO_69 (O_69,N_22975,N_24941);
nand UO_70 (O_70,N_24954,N_23790);
nor UO_71 (O_71,N_24589,N_22505);
and UO_72 (O_72,N_22934,N_23310);
or UO_73 (O_73,N_22876,N_23953);
or UO_74 (O_74,N_22924,N_24172);
or UO_75 (O_75,N_23229,N_23773);
or UO_76 (O_76,N_23216,N_23033);
nand UO_77 (O_77,N_24167,N_24091);
xnor UO_78 (O_78,N_24958,N_24209);
nand UO_79 (O_79,N_23114,N_23336);
nand UO_80 (O_80,N_24453,N_23148);
xor UO_81 (O_81,N_23353,N_23075);
xor UO_82 (O_82,N_24539,N_23383);
and UO_83 (O_83,N_22513,N_24266);
xnor UO_84 (O_84,N_23977,N_23119);
or UO_85 (O_85,N_23290,N_23514);
nor UO_86 (O_86,N_22660,N_24026);
nor UO_87 (O_87,N_24642,N_24044);
nand UO_88 (O_88,N_23510,N_23670);
or UO_89 (O_89,N_23701,N_23416);
and UO_90 (O_90,N_23051,N_22960);
or UO_91 (O_91,N_22525,N_24084);
nor UO_92 (O_92,N_24129,N_23071);
nand UO_93 (O_93,N_24435,N_23975);
or UO_94 (O_94,N_24146,N_24579);
or UO_95 (O_95,N_22722,N_23984);
nand UO_96 (O_96,N_23034,N_22870);
nand UO_97 (O_97,N_24219,N_22850);
nor UO_98 (O_98,N_24205,N_23863);
nand UO_99 (O_99,N_23129,N_22935);
or UO_100 (O_100,N_24462,N_23831);
and UO_101 (O_101,N_23364,N_22792);
xnor UO_102 (O_102,N_24742,N_23544);
nor UO_103 (O_103,N_24294,N_24975);
xnor UO_104 (O_104,N_24580,N_23063);
xor UO_105 (O_105,N_24316,N_23362);
and UO_106 (O_106,N_22998,N_24703);
and UO_107 (O_107,N_24583,N_23906);
xnor UO_108 (O_108,N_23415,N_24308);
nor UO_109 (O_109,N_22882,N_22982);
xor UO_110 (O_110,N_24764,N_22782);
nand UO_111 (O_111,N_23552,N_22629);
nor UO_112 (O_112,N_23425,N_24046);
or UO_113 (O_113,N_23645,N_24041);
or UO_114 (O_114,N_23759,N_23122);
nand UO_115 (O_115,N_23251,N_22885);
xnor UO_116 (O_116,N_23374,N_23291);
and UO_117 (O_117,N_22656,N_23440);
or UO_118 (O_118,N_22569,N_24149);
or UO_119 (O_119,N_24281,N_23734);
nand UO_120 (O_120,N_24609,N_24923);
and UO_121 (O_121,N_24603,N_24657);
or UO_122 (O_122,N_22653,N_24869);
nor UO_123 (O_123,N_24886,N_23870);
or UO_124 (O_124,N_24223,N_23516);
nand UO_125 (O_125,N_24858,N_23320);
or UO_126 (O_126,N_22589,N_23354);
nor UO_127 (O_127,N_24541,N_24976);
nand UO_128 (O_128,N_23292,N_24252);
xor UO_129 (O_129,N_22791,N_23556);
nor UO_130 (O_130,N_24996,N_24213);
or UO_131 (O_131,N_23028,N_24578);
nor UO_132 (O_132,N_24852,N_22657);
or UO_133 (O_133,N_23761,N_23533);
nand UO_134 (O_134,N_22565,N_24532);
or UO_135 (O_135,N_23055,N_24155);
nand UO_136 (O_136,N_24287,N_22783);
nand UO_137 (O_137,N_24323,N_24867);
or UO_138 (O_138,N_23579,N_24658);
nor UO_139 (O_139,N_22856,N_24639);
nand UO_140 (O_140,N_22826,N_22552);
nand UO_141 (O_141,N_23053,N_23306);
or UO_142 (O_142,N_24835,N_24924);
and UO_143 (O_143,N_23786,N_22750);
and UO_144 (O_144,N_24467,N_24182);
or UO_145 (O_145,N_23573,N_23277);
nand UO_146 (O_146,N_23894,N_24554);
or UO_147 (O_147,N_24606,N_23174);
nor UO_148 (O_148,N_22587,N_23565);
or UO_149 (O_149,N_23772,N_24895);
nor UO_150 (O_150,N_22737,N_22765);
nand UO_151 (O_151,N_24225,N_23213);
xor UO_152 (O_152,N_24948,N_22991);
nor UO_153 (O_153,N_23014,N_23311);
nor UO_154 (O_154,N_22706,N_24169);
xor UO_155 (O_155,N_24527,N_22667);
xnor UO_156 (O_156,N_23072,N_24107);
xor UO_157 (O_157,N_24878,N_23039);
and UO_158 (O_158,N_23828,N_23057);
and UO_159 (O_159,N_24906,N_23676);
xnor UO_160 (O_160,N_24273,N_24454);
nor UO_161 (O_161,N_24979,N_24911);
and UO_162 (O_162,N_23128,N_23723);
xor UO_163 (O_163,N_24064,N_23852);
or UO_164 (O_164,N_24232,N_23618);
xor UO_165 (O_165,N_23282,N_23647);
nor UO_166 (O_166,N_24338,N_23762);
and UO_167 (O_167,N_23352,N_23355);
or UO_168 (O_168,N_24009,N_22538);
nor UO_169 (O_169,N_22532,N_23684);
and UO_170 (O_170,N_23518,N_24802);
or UO_171 (O_171,N_22571,N_22760);
and UO_172 (O_172,N_24384,N_22644);
and UO_173 (O_173,N_24803,N_24899);
or UO_174 (O_174,N_23238,N_23750);
nand UO_175 (O_175,N_23536,N_23351);
nand UO_176 (O_176,N_22752,N_23638);
nor UO_177 (O_177,N_24249,N_23503);
and UO_178 (O_178,N_23234,N_23359);
nand UO_179 (O_179,N_23893,N_24673);
and UO_180 (O_180,N_23884,N_24409);
nand UO_181 (O_181,N_22568,N_24451);
or UO_182 (O_182,N_23704,N_22685);
xnor UO_183 (O_183,N_23276,N_24670);
nor UO_184 (O_184,N_23027,N_24950);
nand UO_185 (O_185,N_24744,N_24348);
or UO_186 (O_186,N_22600,N_23696);
or UO_187 (O_187,N_23837,N_23711);
nand UO_188 (O_188,N_23830,N_23209);
nand UO_189 (O_189,N_23316,N_24929);
xnor UO_190 (O_190,N_24908,N_22820);
nand UO_191 (O_191,N_23659,N_24021);
nor UO_192 (O_192,N_23961,N_22586);
and UO_193 (O_193,N_24962,N_23653);
xor UO_194 (O_194,N_23337,N_24874);
nand UO_195 (O_195,N_22661,N_24049);
or UO_196 (O_196,N_23641,N_24263);
or UO_197 (O_197,N_23655,N_23753);
and UO_198 (O_198,N_23236,N_24356);
or UO_199 (O_199,N_23222,N_23987);
xnor UO_200 (O_200,N_24739,N_24234);
nand UO_201 (O_201,N_24125,N_24299);
and UO_202 (O_202,N_23322,N_23758);
or UO_203 (O_203,N_23079,N_24664);
and UO_204 (O_204,N_22534,N_23748);
nor UO_205 (O_205,N_23275,N_22803);
or UO_206 (O_206,N_23454,N_22541);
nand UO_207 (O_207,N_23202,N_22812);
and UO_208 (O_208,N_24177,N_24346);
xnor UO_209 (O_209,N_24357,N_23259);
xnor UO_210 (O_210,N_23038,N_22972);
nand UO_211 (O_211,N_22593,N_24930);
and UO_212 (O_212,N_24659,N_23265);
xnor UO_213 (O_213,N_23443,N_23289);
nand UO_214 (O_214,N_23767,N_22902);
nand UO_215 (O_215,N_22700,N_22522);
or UO_216 (O_216,N_23747,N_23908);
nand UO_217 (O_217,N_23417,N_22786);
xor UO_218 (O_218,N_24914,N_23086);
or UO_219 (O_219,N_24716,N_23268);
nand UO_220 (O_220,N_23488,N_24077);
or UO_221 (O_221,N_23134,N_24244);
xor UO_222 (O_222,N_24521,N_22740);
nand UO_223 (O_223,N_23307,N_23065);
and UO_224 (O_224,N_23411,N_23077);
nor UO_225 (O_225,N_23288,N_23464);
and UO_226 (O_226,N_24050,N_22890);
or UO_227 (O_227,N_23471,N_22611);
or UO_228 (O_228,N_22971,N_22728);
nor UO_229 (O_229,N_24726,N_23789);
nand UO_230 (O_230,N_24184,N_22814);
xor UO_231 (O_231,N_23804,N_24873);
nand UO_232 (O_232,N_23505,N_23117);
or UO_233 (O_233,N_24880,N_22897);
nand UO_234 (O_234,N_23609,N_23922);
nor UO_235 (O_235,N_22805,N_23891);
and UO_236 (O_236,N_23935,N_23127);
xor UO_237 (O_237,N_24854,N_22609);
or UO_238 (O_238,N_22630,N_23816);
xor UO_239 (O_239,N_23170,N_23799);
nor UO_240 (O_240,N_23532,N_23626);
nand UO_241 (O_241,N_23694,N_23744);
xnor UO_242 (O_242,N_24157,N_24227);
or UO_243 (O_243,N_22811,N_23287);
nor UO_244 (O_244,N_23166,N_24315);
or UO_245 (O_245,N_22516,N_23864);
and UO_246 (O_246,N_24736,N_23757);
and UO_247 (O_247,N_23521,N_24571);
or UO_248 (O_248,N_23346,N_24469);
xor UO_249 (O_249,N_24052,N_24829);
xor UO_250 (O_250,N_24085,N_23598);
xnor UO_251 (O_251,N_22852,N_23142);
xor UO_252 (O_252,N_24588,N_24889);
and UO_253 (O_253,N_23001,N_22775);
or UO_254 (O_254,N_24745,N_24550);
or UO_255 (O_255,N_23644,N_23774);
nand UO_256 (O_256,N_24390,N_23372);
nor UO_257 (O_257,N_24023,N_23835);
nand UO_258 (O_258,N_23896,N_23500);
and UO_259 (O_259,N_22663,N_23137);
nor UO_260 (O_260,N_24337,N_23255);
and UO_261 (O_261,N_22868,N_23736);
or UO_262 (O_262,N_24845,N_24305);
or UO_263 (O_263,N_24198,N_24971);
nor UO_264 (O_264,N_22709,N_22925);
xnor UO_265 (O_265,N_23685,N_22634);
xor UO_266 (O_266,N_23487,N_22542);
nand UO_267 (O_267,N_22818,N_22861);
nand UO_268 (O_268,N_24524,N_23445);
xnor UO_269 (O_269,N_23082,N_23667);
xnor UO_270 (O_270,N_23361,N_24546);
or UO_271 (O_271,N_22635,N_24511);
and UO_272 (O_272,N_23943,N_22625);
or UO_273 (O_273,N_24953,N_23872);
xor UO_274 (O_274,N_23564,N_23652);
nand UO_275 (O_275,N_24598,N_24286);
xor UO_276 (O_276,N_23915,N_24313);
and UO_277 (O_277,N_24022,N_23857);
xnor UO_278 (O_278,N_24916,N_23365);
or UO_279 (O_279,N_24201,N_24214);
nand UO_280 (O_280,N_22622,N_24468);
nor UO_281 (O_281,N_23606,N_24464);
and UO_282 (O_282,N_24708,N_24277);
nor UO_283 (O_283,N_24743,N_23952);
nor UO_284 (O_284,N_24408,N_23782);
and UO_285 (O_285,N_23809,N_23406);
xnor UO_286 (O_286,N_23775,N_23687);
nand UO_287 (O_287,N_23635,N_23107);
or UO_288 (O_288,N_23865,N_22537);
nand UO_289 (O_289,N_23637,N_23706);
and UO_290 (O_290,N_23456,N_22647);
and UO_291 (O_291,N_23571,N_24661);
and UO_292 (O_292,N_23624,N_24188);
nand UO_293 (O_293,N_23597,N_23827);
and UO_294 (O_294,N_23887,N_24635);
nor UO_295 (O_295,N_23035,N_24495);
and UO_296 (O_296,N_23444,N_23283);
nor UO_297 (O_297,N_24522,N_23046);
nor UO_298 (O_298,N_24966,N_23451);
nand UO_299 (O_299,N_24977,N_23088);
nand UO_300 (O_300,N_23545,N_24434);
xnor UO_301 (O_301,N_24872,N_24355);
nor UO_302 (O_302,N_24582,N_23332);
and UO_303 (O_303,N_23165,N_24211);
or UO_304 (O_304,N_23883,N_24246);
or UO_305 (O_305,N_23955,N_22527);
nand UO_306 (O_306,N_22574,N_23699);
nor UO_307 (O_307,N_23373,N_24343);
and UO_308 (O_308,N_24885,N_23543);
nor UO_309 (O_309,N_23538,N_24358);
and UO_310 (O_310,N_22502,N_23431);
xnor UO_311 (O_311,N_23607,N_22977);
xnor UO_312 (O_312,N_24255,N_23794);
xnor UO_313 (O_313,N_23264,N_24699);
xor UO_314 (O_314,N_23680,N_24497);
or UO_315 (O_315,N_24126,N_24059);
nand UO_316 (O_316,N_22872,N_24893);
or UO_317 (O_317,N_23085,N_22954);
nor UO_318 (O_318,N_23056,N_23081);
nor UO_319 (O_319,N_23410,N_24967);
and UO_320 (O_320,N_24120,N_24186);
or UO_321 (O_321,N_22887,N_23483);
or UO_322 (O_322,N_23735,N_23920);
nor UO_323 (O_323,N_23327,N_24862);
and UO_324 (O_324,N_24793,N_23858);
or UO_325 (O_325,N_23878,N_22789);
nand UO_326 (O_326,N_24959,N_24002);
or UO_327 (O_327,N_22785,N_23386);
nor UO_328 (O_328,N_23660,N_24407);
nor UO_329 (O_329,N_24332,N_24145);
nand UO_330 (O_330,N_22579,N_22799);
nor UO_331 (O_331,N_23881,N_22504);
xnor UO_332 (O_332,N_23092,N_24759);
xor UO_333 (O_333,N_24711,N_24832);
nor UO_334 (O_334,N_22566,N_23221);
nand UO_335 (O_335,N_22672,N_24654);
xor UO_336 (O_336,N_23482,N_23492);
nand UO_337 (O_337,N_24668,N_23742);
nand UO_338 (O_338,N_23076,N_24768);
nor UO_339 (O_339,N_22506,N_23130);
nand UO_340 (O_340,N_22664,N_22863);
nor UO_341 (O_341,N_24124,N_23839);
nand UO_342 (O_342,N_24933,N_23161);
xnor UO_343 (O_343,N_24560,N_24203);
xnor UO_344 (O_344,N_23875,N_24551);
or UO_345 (O_345,N_23714,N_23700);
and UO_346 (O_346,N_23980,N_23525);
nor UO_347 (O_347,N_22543,N_23849);
nor UO_348 (O_348,N_24839,N_24636);
and UO_349 (O_349,N_24713,N_23147);
nor UO_350 (O_350,N_23966,N_22682);
xnor UO_351 (O_351,N_23720,N_24780);
nand UO_352 (O_352,N_24753,N_22596);
nand UO_353 (O_353,N_22573,N_24411);
or UO_354 (O_354,N_24498,N_23184);
nor UO_355 (O_355,N_22512,N_24304);
nand UO_356 (O_356,N_23401,N_24861);
or UO_357 (O_357,N_24786,N_23208);
nand UO_358 (O_358,N_23692,N_24375);
nand UO_359 (O_359,N_23133,N_23025);
or UO_360 (O_360,N_23965,N_22749);
and UO_361 (O_361,N_22712,N_24545);
nor UO_362 (O_362,N_24185,N_23523);
xnor UO_363 (O_363,N_22906,N_22619);
or UO_364 (O_364,N_22594,N_24100);
nor UO_365 (O_365,N_23709,N_24490);
nor UO_366 (O_366,N_24445,N_22742);
or UO_367 (O_367,N_22981,N_24108);
nand UO_368 (O_368,N_22913,N_24896);
and UO_369 (O_369,N_24265,N_23240);
nand UO_370 (O_370,N_22707,N_23555);
nand UO_371 (O_371,N_23993,N_22809);
nor UO_372 (O_372,N_23859,N_24827);
or UO_373 (O_373,N_22747,N_24489);
xor UO_374 (O_374,N_24302,N_23409);
xor UO_375 (O_375,N_22894,N_23377);
xnor UO_376 (O_376,N_24282,N_23160);
nand UO_377 (O_377,N_24161,N_22608);
nand UO_378 (O_378,N_24653,N_22881);
xor UO_379 (O_379,N_23806,N_24116);
nand UO_380 (O_380,N_24239,N_23737);
or UO_381 (O_381,N_22892,N_23413);
xnor UO_382 (O_382,N_23568,N_23020);
xnor UO_383 (O_383,N_24986,N_23198);
nor UO_384 (O_384,N_23338,N_24342);
and UO_385 (O_385,N_22561,N_24494);
or UO_386 (O_386,N_24817,N_24504);
or UO_387 (O_387,N_22732,N_22617);
and UO_388 (O_388,N_24306,N_22531);
and UO_389 (O_389,N_23496,N_23224);
or UO_390 (O_390,N_23560,N_24805);
xnor UO_391 (O_391,N_23101,N_24060);
and UO_392 (O_392,N_22918,N_24733);
and UO_393 (O_393,N_24620,N_22539);
nor UO_394 (O_394,N_24027,N_24311);
or UO_395 (O_395,N_24472,N_24318);
or UO_396 (O_396,N_24807,N_24425);
xor UO_397 (O_397,N_24056,N_23619);
nor UO_398 (O_398,N_24692,N_24741);
or UO_399 (O_399,N_24222,N_22948);
nor UO_400 (O_400,N_24112,N_23248);
or UO_401 (O_401,N_23163,N_24173);
nand UO_402 (O_402,N_22550,N_23601);
nand UO_403 (O_403,N_24396,N_23649);
xnor UO_404 (O_404,N_23381,N_24737);
and UO_405 (O_405,N_24290,N_23743);
xor UO_406 (O_406,N_23693,N_23094);
nand UO_407 (O_407,N_23330,N_22825);
nor UO_408 (O_408,N_23671,N_22845);
nor UO_409 (O_409,N_23475,N_24175);
nor UO_410 (O_410,N_24629,N_23719);
nor UO_411 (O_411,N_23242,N_22734);
or UO_412 (O_412,N_23682,N_23084);
xnor UO_413 (O_413,N_24563,N_24850);
nand UO_414 (O_414,N_23040,N_24105);
nand UO_415 (O_415,N_23557,N_24417);
nor UO_416 (O_416,N_23018,N_23580);
nand UO_417 (O_417,N_23003,N_23779);
or UO_418 (O_418,N_23422,N_23593);
nor UO_419 (O_419,N_23246,N_24725);
xor UO_420 (O_420,N_24421,N_23959);
and UO_421 (O_421,N_24492,N_23979);
xor UO_422 (O_422,N_22710,N_23149);
xnor UO_423 (O_423,N_23850,N_23746);
nand UO_424 (O_424,N_23590,N_23195);
nand UO_425 (O_425,N_24471,N_22570);
nor UO_426 (O_426,N_22901,N_24840);
nand UO_427 (O_427,N_23104,N_23326);
or UO_428 (O_428,N_23400,N_24879);
and UO_429 (O_429,N_24429,N_22668);
nand UO_430 (O_430,N_23029,N_22654);
xnor UO_431 (O_431,N_23215,N_24946);
nand UO_432 (O_432,N_22950,N_22697);
xor UO_433 (O_433,N_23793,N_24660);
nand UO_434 (O_434,N_23554,N_22875);
or UO_435 (O_435,N_24631,N_24680);
xor UO_436 (O_436,N_23895,N_24478);
nor UO_437 (O_437,N_24095,N_24011);
or UO_438 (O_438,N_24456,N_23845);
nand UO_439 (O_439,N_23928,N_22692);
xor UO_440 (O_440,N_23313,N_23394);
or UO_441 (O_441,N_24727,N_22683);
nand UO_442 (O_442,N_23718,N_24907);
nor UO_443 (O_443,N_24540,N_24766);
or UO_444 (O_444,N_24814,N_24663);
xnor UO_445 (O_445,N_22713,N_24686);
nor UO_446 (O_446,N_22738,N_23112);
and UO_447 (O_447,N_24892,N_24370);
xnor UO_448 (O_448,N_23620,N_24216);
and UO_449 (O_449,N_24798,N_24317);
nor UO_450 (O_450,N_23467,N_24974);
nand UO_451 (O_451,N_24076,N_24307);
nand UO_452 (O_452,N_23106,N_23465);
nand UO_453 (O_453,N_24600,N_24309);
nand UO_454 (O_454,N_24509,N_24119);
nand UO_455 (O_455,N_23992,N_24477);
and UO_456 (O_456,N_23628,N_22736);
nor UO_457 (O_457,N_22988,N_23506);
and UO_458 (O_458,N_24152,N_22762);
nor UO_459 (O_459,N_24993,N_22666);
nand UO_460 (O_460,N_23190,N_23486);
and UO_461 (O_461,N_24310,N_22944);
or UO_462 (O_462,N_24502,N_23279);
nand UO_463 (O_463,N_22912,N_24373);
and UO_464 (O_464,N_23562,N_23924);
xnor UO_465 (O_465,N_23838,N_23769);
xnor UO_466 (O_466,N_24666,N_23582);
and UO_467 (O_467,N_24517,N_24752);
or UO_468 (O_468,N_23797,N_22636);
nor UO_469 (O_469,N_23841,N_24553);
nor UO_470 (O_470,N_24256,N_23921);
or UO_471 (O_471,N_23548,N_24611);
and UO_472 (O_472,N_23293,N_23049);
or UO_473 (O_473,N_24593,N_23889);
xor UO_474 (O_474,N_24207,N_23227);
and UO_475 (O_475,N_24801,N_24784);
and UO_476 (O_476,N_24614,N_23468);
and UO_477 (O_477,N_24233,N_23946);
and UO_478 (O_478,N_22605,N_24877);
nor UO_479 (O_479,N_24109,N_23155);
or UO_480 (O_480,N_24732,N_22519);
or UO_481 (O_481,N_22637,N_22974);
nor UO_482 (O_482,N_22679,N_23446);
or UO_483 (O_483,N_22815,N_23803);
xor UO_484 (O_484,N_23851,N_23449);
and UO_485 (O_485,N_24296,N_22761);
nor UO_486 (O_486,N_23390,N_22914);
nor UO_487 (O_487,N_23572,N_23302);
or UO_488 (O_488,N_24197,N_23504);
and UO_489 (O_489,N_23387,N_24901);
and UO_490 (O_490,N_24176,N_24884);
xnor UO_491 (O_491,N_22951,N_23630);
and UO_492 (O_492,N_23203,N_24816);
xnor UO_493 (O_493,N_24072,N_24830);
and UO_494 (O_494,N_24229,N_23530);
or UO_495 (O_495,N_23998,N_22877);
nor UO_496 (O_496,N_24017,N_24824);
xnor UO_497 (O_497,N_24621,N_23668);
and UO_498 (O_498,N_24087,N_22693);
nor UO_499 (O_499,N_24718,N_24094);
nor UO_500 (O_500,N_23933,N_24678);
nand UO_501 (O_501,N_24164,N_24682);
and UO_502 (O_502,N_24051,N_23507);
nand UO_503 (O_503,N_22846,N_23581);
nor UO_504 (O_504,N_23541,N_23931);
nor UO_505 (O_505,N_23214,N_22575);
nor UO_506 (O_506,N_24283,N_23017);
nand UO_507 (O_507,N_22514,N_24040);
nand UO_508 (O_508,N_24860,N_24561);
nor UO_509 (O_509,N_23902,N_22669);
or UO_510 (O_510,N_22915,N_23960);
and UO_511 (O_511,N_22784,N_22857);
or UO_512 (O_512,N_22649,N_24697);
nor UO_513 (O_513,N_23531,N_24655);
or UO_514 (O_514,N_23724,N_24608);
nand UO_515 (O_515,N_23204,N_24577);
nand UO_516 (O_516,N_22743,N_24833);
nor UO_517 (O_517,N_23663,N_22819);
nor UO_518 (O_518,N_24062,N_24269);
and UO_519 (O_519,N_22959,N_23610);
nand UO_520 (O_520,N_24864,N_24143);
xnor UO_521 (O_521,N_23524,N_24783);
nand UO_522 (O_522,N_24134,N_23206);
or UO_523 (O_523,N_23967,N_24248);
xnor UO_524 (O_524,N_23340,N_24194);
nor UO_525 (O_525,N_22758,N_23253);
nor UO_526 (O_526,N_23932,N_23392);
or UO_527 (O_527,N_23066,N_24754);
nand UO_528 (O_528,N_24909,N_23191);
xnor UO_529 (O_529,N_22922,N_24382);
xnor UO_530 (O_530,N_23890,N_23223);
nand UO_531 (O_531,N_23599,N_24769);
or UO_532 (O_532,N_22955,N_23664);
nand UO_533 (O_533,N_24291,N_24934);
xor UO_534 (O_534,N_24117,N_22686);
and UO_535 (O_535,N_24415,N_23455);
nor UO_536 (O_536,N_22614,N_22874);
nand UO_537 (O_537,N_23651,N_24844);
xor UO_538 (O_538,N_24276,N_23771);
xor UO_539 (O_539,N_22938,N_24945);
or UO_540 (O_540,N_23423,N_22896);
or UO_541 (O_541,N_24330,N_24905);
and UO_542 (O_542,N_24627,N_22956);
or UO_543 (O_543,N_24368,N_24927);
or UO_544 (O_544,N_24110,N_22606);
or UO_545 (O_545,N_24778,N_24289);
xor UO_546 (O_546,N_24279,N_22919);
and UO_547 (O_547,N_22602,N_23131);
xor UO_548 (O_548,N_23172,N_22536);
nor UO_549 (O_549,N_24665,N_24645);
nor UO_550 (O_550,N_24092,N_24853);
xnor UO_551 (O_551,N_24166,N_22958);
nand UO_552 (O_552,N_23476,N_23271);
nand UO_553 (O_553,N_23811,N_24765);
xor UO_554 (O_554,N_23237,N_24325);
or UO_555 (O_555,N_23820,N_23379);
xor UO_556 (O_556,N_24714,N_24587);
and UO_557 (O_557,N_24347,N_22702);
and UO_558 (O_558,N_24328,N_23698);
and UO_559 (O_559,N_23939,N_24192);
and UO_560 (O_560,N_24689,N_23672);
xnor UO_561 (O_561,N_23019,N_24586);
nand UO_562 (O_562,N_23199,N_24988);
nor UO_563 (O_563,N_24972,N_24376);
xnor UO_564 (O_564,N_24849,N_24863);
nor UO_565 (O_565,N_23569,N_24104);
xor UO_566 (O_566,N_23800,N_23345);
or UO_567 (O_567,N_24038,N_24891);
xnor UO_568 (O_568,N_22952,N_24334);
nand UO_569 (O_569,N_23179,N_24843);
and UO_570 (O_570,N_22551,N_24617);
and UO_571 (O_571,N_23426,N_22766);
nor UO_572 (O_572,N_23988,N_22592);
or UO_573 (O_573,N_24841,N_22849);
nand UO_574 (O_574,N_24034,N_23944);
xnor UO_575 (O_575,N_24516,N_22962);
or UO_576 (O_576,N_23563,N_24082);
nor UO_577 (O_577,N_24156,N_23146);
xnor UO_578 (O_578,N_23515,N_24693);
nor UO_579 (O_579,N_24067,N_23489);
or UO_580 (O_580,N_22905,N_22931);
nor UO_581 (O_581,N_23257,N_24133);
nand UO_582 (O_582,N_23187,N_23868);
xnor UO_583 (O_583,N_24163,N_24018);
nand UO_584 (O_584,N_24327,N_23710);
and UO_585 (O_585,N_24097,N_23551);
or UO_586 (O_586,N_23182,N_23061);
xnor UO_587 (O_587,N_24231,N_23249);
nand UO_588 (O_588,N_22945,N_23550);
xnor UO_589 (O_589,N_23108,N_24208);
nor UO_590 (O_590,N_24704,N_23105);
nor UO_591 (O_591,N_23169,N_22595);
and UO_592 (O_592,N_24433,N_24118);
or UO_593 (O_593,N_24918,N_24969);
nand UO_594 (O_594,N_22544,N_24394);
xor UO_595 (O_595,N_23244,N_24048);
and UO_596 (O_596,N_24808,N_24771);
and UO_597 (O_597,N_23333,N_22853);
and UO_598 (O_598,N_22714,N_23836);
nor UO_599 (O_599,N_23435,N_24029);
xnor UO_600 (O_600,N_24656,N_24187);
nor UO_601 (O_601,N_23405,N_23380);
and UO_602 (O_602,N_24581,N_23903);
xnor UO_603 (O_603,N_23032,N_24443);
nor UO_604 (O_604,N_24364,N_22941);
xor UO_605 (O_605,N_24857,N_24651);
nor UO_606 (O_606,N_24961,N_22723);
nor UO_607 (O_607,N_23617,N_23115);
xor UO_608 (O_608,N_22961,N_23138);
nor UO_609 (O_609,N_23587,N_24724);
nor UO_610 (O_610,N_22858,N_23384);
nand UO_611 (O_611,N_23323,N_23427);
and UO_612 (O_612,N_23765,N_22524);
or UO_613 (O_613,N_22699,N_23300);
and UO_614 (O_614,N_23009,N_24865);
or UO_615 (O_615,N_24452,N_23805);
or UO_616 (O_616,N_24055,N_24999);
nand UO_617 (O_617,N_23194,N_24140);
or UO_618 (O_618,N_23589,N_23625);
or UO_619 (O_619,N_22548,N_24381);
and UO_620 (O_620,N_23739,N_23462);
xnor UO_621 (O_621,N_24951,N_24650);
xnor UO_622 (O_622,N_24288,N_22833);
nand UO_623 (O_623,N_23627,N_22745);
xnor UO_624 (O_624,N_23357,N_23690);
or UO_625 (O_625,N_24760,N_24010);
nand UO_626 (O_626,N_24649,N_24749);
and UO_627 (O_627,N_23861,N_24543);
nand UO_628 (O_628,N_24701,N_24212);
xor UO_629 (O_629,N_24881,N_23470);
xnor UO_630 (O_630,N_23823,N_22800);
xor UO_631 (O_631,N_24568,N_24128);
and UO_632 (O_632,N_23022,N_23360);
or UO_633 (O_633,N_22963,N_23783);
or UO_634 (O_634,N_24767,N_23245);
and UO_635 (O_635,N_24903,N_24810);
nand UO_636 (O_636,N_24735,N_23102);
nor UO_637 (O_637,N_23250,N_23983);
or UO_638 (O_638,N_23371,N_22585);
xnor UO_639 (O_639,N_23241,N_23755);
nand UO_640 (O_640,N_23233,N_22718);
nand UO_641 (O_641,N_24262,N_23499);
nand UO_642 (O_642,N_22643,N_23011);
nor UO_643 (O_643,N_23778,N_23643);
xnor UO_644 (O_644,N_23054,N_24813);
xor UO_645 (O_645,N_23262,N_24350);
and UO_646 (O_646,N_22824,N_24397);
or UO_647 (O_647,N_23989,N_24709);
nand UO_648 (O_648,N_22980,N_24405);
and UO_649 (O_649,N_23367,N_23583);
nand UO_650 (O_650,N_23254,N_23673);
nor UO_651 (O_651,N_23923,N_23197);
xor UO_652 (O_652,N_23512,N_23869);
nor UO_653 (O_653,N_24033,N_24915);
nand UO_654 (O_654,N_24403,N_24387);
or UO_655 (O_655,N_24257,N_24413);
nand UO_656 (O_656,N_22695,N_22999);
xor UO_657 (O_657,N_24779,N_24576);
xor UO_658 (O_658,N_22559,N_24788);
and UO_659 (O_659,N_23389,N_24025);
nor UO_660 (O_660,N_22779,N_23278);
nand UO_661 (O_661,N_22923,N_24499);
nand UO_662 (O_662,N_22965,N_24039);
or UO_663 (O_663,N_24834,N_23491);
nor UO_664 (O_664,N_23662,N_24601);
and UO_665 (O_665,N_22726,N_22970);
or UO_666 (O_666,N_24333,N_24189);
nor UO_667 (O_667,N_23519,N_24520);
and UO_668 (O_668,N_23150,N_23613);
nand UO_669 (O_669,N_24012,N_23898);
nand UO_670 (O_670,N_24301,N_23153);
nand UO_671 (O_671,N_22801,N_22648);
and UO_672 (O_672,N_23629,N_23576);
xor UO_673 (O_673,N_23498,N_24618);
nand UO_674 (O_674,N_23947,N_24254);
nand UO_675 (O_675,N_24781,N_24887);
xor UO_676 (O_676,N_24446,N_24322);
nor UO_677 (O_677,N_23024,N_24970);
nand UO_678 (O_678,N_24956,N_23534);
nor UO_679 (O_679,N_23260,N_24964);
nor UO_680 (O_680,N_23479,N_24998);
xor UO_681 (O_681,N_23754,N_24868);
nor UO_682 (O_682,N_24787,N_24549);
nand UO_683 (O_683,N_24121,N_24894);
and UO_684 (O_684,N_23526,N_23595);
nor UO_685 (O_685,N_24910,N_24013);
nor UO_686 (O_686,N_23829,N_24354);
and UO_687 (O_687,N_22620,N_23815);
and UO_688 (O_688,N_23691,N_24534);
xor UO_689 (O_689,N_24395,N_24782);
or UO_690 (O_690,N_23391,N_24684);
and UO_691 (O_691,N_23180,N_24599);
nor UO_692 (O_692,N_23269,N_23031);
xor UO_693 (O_693,N_24883,N_24103);
or UO_694 (O_694,N_22711,N_23796);
or UO_695 (O_695,N_23252,N_22626);
nand UO_696 (O_696,N_24345,N_24567);
xor UO_697 (O_697,N_22755,N_23996);
nand UO_698 (O_698,N_22871,N_24470);
xor UO_699 (O_699,N_22984,N_24785);
and UO_700 (O_700,N_23826,N_23157);
xnor UO_701 (O_701,N_24036,N_24921);
nor UO_702 (O_702,N_23452,N_22526);
xnor UO_703 (O_703,N_22721,N_24440);
nand UO_704 (O_704,N_22888,N_23273);
or UO_705 (O_705,N_23258,N_24035);
xor UO_706 (O_706,N_24272,N_23281);
and UO_707 (O_707,N_24379,N_24392);
or UO_708 (O_708,N_22893,N_22994);
nand UO_709 (O_709,N_23412,N_24775);
xnor UO_710 (O_710,N_22869,N_24702);
or UO_711 (O_711,N_23118,N_23535);
xor UO_712 (O_712,N_24218,N_22978);
nand UO_713 (O_713,N_24122,N_24698);
or UO_714 (O_714,N_23712,N_24685);
xor UO_715 (O_715,N_24757,N_22631);
and UO_716 (O_716,N_23393,N_24774);
and UO_717 (O_717,N_22741,N_23008);
nand UO_718 (O_718,N_22946,N_24267);
nand UO_719 (O_719,N_24943,N_24081);
nand UO_720 (O_720,N_22949,N_24130);
nor UO_721 (O_721,N_23824,N_23856);
nor UO_722 (O_722,N_24137,N_24821);
nand UO_723 (O_723,N_22684,N_22879);
nand UO_724 (O_724,N_22822,N_24530);
and UO_725 (O_725,N_24258,N_23100);
or UO_726 (O_726,N_24162,N_23074);
and UO_727 (O_727,N_23950,N_23867);
nor UO_728 (O_728,N_22744,N_24772);
nor UO_729 (O_729,N_23370,N_23819);
and UO_730 (O_730,N_24533,N_23015);
nand UO_731 (O_731,N_24637,N_23954);
xor UO_732 (O_732,N_23801,N_23695);
nor UO_733 (O_733,N_23304,N_24876);
nor UO_734 (O_734,N_22835,N_24339);
nor UO_735 (O_735,N_24042,N_24990);
xnor UO_736 (O_736,N_24461,N_22808);
xor UO_737 (O_737,N_22708,N_24806);
nand UO_738 (O_738,N_24920,N_22676);
or UO_739 (O_739,N_23080,N_22528);
nor UO_740 (O_740,N_22719,N_23763);
nand UO_741 (O_741,N_23448,N_23103);
nand UO_742 (O_742,N_24939,N_23752);
nor UO_743 (O_743,N_22681,N_23113);
or UO_744 (O_744,N_24240,N_24210);
xor UO_745 (O_745,N_23023,N_23408);
nor UO_746 (O_746,N_23052,N_22533);
or UO_747 (O_747,N_24628,N_24362);
xnor UO_748 (O_748,N_24555,N_23860);
or UO_749 (O_749,N_23200,N_24083);
nand UO_750 (O_750,N_22836,N_23559);
nor UO_751 (O_751,N_23437,N_24811);
xnor UO_752 (O_752,N_22832,N_24139);
xnor UO_753 (O_753,N_24585,N_24158);
or UO_754 (O_754,N_24569,N_24871);
nand UO_755 (O_755,N_22767,N_24992);
xnor UO_756 (O_756,N_22563,N_23026);
xnor UO_757 (O_757,N_24450,N_22986);
nand UO_758 (O_758,N_24416,N_24572);
nand UO_759 (O_759,N_23295,N_24280);
and UO_760 (O_760,N_22807,N_22652);
and UO_761 (O_761,N_22511,N_23716);
xor UO_762 (O_762,N_24630,N_22727);
nand UO_763 (O_763,N_22997,N_23447);
nor UO_764 (O_764,N_24994,N_23745);
nand UO_765 (O_765,N_24503,N_23808);
and UO_766 (O_766,N_24058,N_24075);
and UO_767 (O_767,N_22834,N_24412);
nand UO_768 (O_768,N_23740,N_22501);
nand UO_769 (O_769,N_24004,N_22547);
or UO_770 (O_770,N_24171,N_22549);
or UO_771 (O_771,N_23472,N_24809);
or UO_772 (O_772,N_23073,N_24037);
or UO_773 (O_773,N_24410,N_22508);
xor UO_774 (O_774,N_24168,N_22645);
nand UO_775 (O_775,N_23116,N_23154);
nand UO_776 (O_776,N_22806,N_22788);
or UO_777 (O_777,N_23272,N_24113);
xor UO_778 (O_778,N_23050,N_24828);
or UO_779 (O_779,N_24981,N_24619);
or UO_780 (O_780,N_24359,N_23574);
nand UO_781 (O_781,N_23239,N_22564);
or UO_782 (O_782,N_22725,N_23111);
xnor UO_783 (O_783,N_24270,N_23021);
xnor UO_784 (O_784,N_24913,N_22968);
nor UO_785 (O_785,N_23124,N_23368);
nand UO_786 (O_786,N_23926,N_23900);
nand UO_787 (O_787,N_24947,N_23679);
or UO_788 (O_788,N_23091,N_23460);
nand UO_789 (O_789,N_23683,N_23798);
or UO_790 (O_790,N_24138,N_23632);
nor UO_791 (O_791,N_24154,N_24447);
nand UO_792 (O_792,N_23439,N_24652);
nand UO_793 (O_793,N_23605,N_22895);
nor UO_794 (O_794,N_23136,N_24190);
xnor UO_795 (O_795,N_22936,N_23528);
nor UO_796 (O_796,N_24762,N_24388);
nand UO_797 (O_797,N_22909,N_23738);
xor UO_798 (O_798,N_24952,N_24773);
nor UO_799 (O_799,N_23925,N_23067);
and UO_800 (O_800,N_24264,N_22837);
or UO_801 (O_801,N_24066,N_23388);
or UO_802 (O_802,N_23527,N_23715);
or UO_803 (O_803,N_24196,N_22976);
nor UO_804 (O_804,N_23318,N_24519);
nand UO_805 (O_805,N_24369,N_22529);
xnor UO_806 (O_806,N_23843,N_24090);
xnor UO_807 (O_807,N_23232,N_24931);
xnor UO_808 (O_808,N_24102,N_23751);
and UO_809 (O_809,N_24320,N_23436);
xnor UO_810 (O_810,N_22964,N_24607);
nand UO_811 (O_811,N_23247,N_24465);
or UO_812 (O_812,N_22658,N_23567);
nand UO_813 (O_813,N_24061,N_22878);
or UO_814 (O_814,N_24336,N_22840);
xnor UO_815 (O_815,N_24633,N_23270);
nand UO_816 (O_816,N_24073,N_23167);
xor UO_817 (O_817,N_24089,N_22553);
nand UO_818 (O_818,N_22756,N_23139);
and UO_819 (O_819,N_24326,N_22523);
nand UO_820 (O_820,N_24750,N_24728);
nor UO_821 (O_821,N_23713,N_24285);
xnor UO_822 (O_822,N_22557,N_24250);
and UO_823 (O_823,N_24268,N_24991);
xor UO_824 (O_824,N_23369,N_23398);
or UO_825 (O_825,N_23004,N_23547);
nand UO_826 (O_826,N_22503,N_24584);
nand UO_827 (O_827,N_22680,N_22675);
nand UO_828 (O_828,N_24935,N_23243);
and UO_829 (O_829,N_22903,N_24922);
or UO_830 (O_830,N_22703,N_22610);
nor UO_831 (O_831,N_22599,N_23396);
and UO_832 (O_832,N_24398,N_23089);
nor UO_833 (O_833,N_23721,N_24748);
or UO_834 (O_834,N_23484,N_23309);
xnor UO_835 (O_835,N_24590,N_23844);
xor UO_836 (O_836,N_24738,N_23095);
nand UO_837 (O_837,N_24888,N_23726);
or UO_838 (O_838,N_24144,N_24444);
xnor UO_839 (O_839,N_23905,N_24001);
nor UO_840 (O_840,N_24602,N_23497);
and UO_841 (O_841,N_22854,N_24024);
nor UO_842 (O_842,N_22572,N_24312);
nand UO_843 (O_843,N_23833,N_22990);
or UO_844 (O_844,N_23834,N_24078);
and UO_845 (O_845,N_22796,N_22546);
nand UO_846 (O_846,N_24335,N_24797);
and UO_847 (O_847,N_24514,N_24353);
or UO_848 (O_848,N_23999,N_23177);
or UO_849 (O_849,N_23060,N_23561);
and UO_850 (O_850,N_23006,N_23513);
or UO_851 (O_851,N_22839,N_24482);
nor UO_852 (O_852,N_23577,N_23874);
and UO_853 (O_853,N_24366,N_23453);
nor UO_854 (O_854,N_23348,N_24937);
nor UO_855 (O_855,N_24419,N_23358);
nand UO_856 (O_856,N_23708,N_24393);
or UO_857 (O_857,N_24191,N_24000);
nor UO_858 (O_858,N_24178,N_23218);
nor UO_859 (O_859,N_22828,N_22646);
nand UO_860 (O_860,N_23399,N_23974);
and UO_861 (O_861,N_23016,N_23529);
nand UO_862 (O_862,N_22633,N_24720);
nor UO_863 (O_863,N_23325,N_23228);
and UO_864 (O_864,N_24488,N_23942);
nor UO_865 (O_865,N_24422,N_23586);
xor UO_866 (O_866,N_24148,N_22615);
nor UO_867 (O_867,N_23546,N_23892);
nand UO_868 (O_868,N_23780,N_24676);
xor UO_869 (O_869,N_23397,N_23854);
or UO_870 (O_870,N_22983,N_24791);
nand UO_871 (O_871,N_22754,N_22838);
nand UO_872 (O_872,N_23882,N_22810);
and UO_873 (O_873,N_24800,N_23877);
or UO_874 (O_874,N_22583,N_24792);
nand UO_875 (O_875,N_23433,N_24622);
or UO_876 (O_876,N_23159,N_24298);
and UO_877 (O_877,N_23985,N_22580);
nor UO_878 (O_878,N_23681,N_24057);
and UO_879 (O_879,N_23434,N_22555);
or UO_880 (O_880,N_23430,N_24501);
nand UO_881 (O_881,N_22886,N_23657);
and UO_882 (O_882,N_24674,N_23315);
and UO_883 (O_883,N_24687,N_24080);
xor UO_884 (O_884,N_22844,N_23441);
nand UO_885 (O_885,N_22916,N_24596);
and UO_886 (O_886,N_24897,N_24804);
nor UO_887 (O_887,N_23899,N_23731);
and UO_888 (O_888,N_23951,N_22509);
nand UO_889 (O_889,N_24556,N_24646);
and UO_890 (O_890,N_23217,N_22673);
or UO_891 (O_891,N_23677,N_22535);
xor UO_892 (O_892,N_22798,N_24826);
xor UO_893 (O_893,N_24181,N_24329);
xor UO_894 (O_894,N_23125,N_22987);
nor UO_895 (O_895,N_22671,N_22584);
and UO_896 (O_896,N_23909,N_24681);
or UO_897 (O_897,N_23817,N_24790);
nand UO_898 (O_898,N_22704,N_23982);
nor UO_899 (O_899,N_23420,N_24705);
nand UO_900 (O_900,N_23787,N_24777);
nand UO_901 (O_901,N_23297,N_22716);
xnor UO_902 (O_902,N_24968,N_22698);
xnor UO_903 (O_903,N_24944,N_24746);
or UO_904 (O_904,N_24150,N_22864);
nand UO_905 (O_905,N_22558,N_23666);
and UO_906 (O_906,N_24295,N_23722);
xor UO_907 (O_907,N_23299,N_24512);
and UO_908 (O_908,N_24431,N_24505);
xnor UO_909 (O_909,N_24526,N_23047);
nand UO_910 (O_910,N_24202,N_24677);
or UO_911 (O_911,N_24053,N_22943);
nor UO_912 (O_912,N_24151,N_23897);
or UO_913 (O_913,N_23509,N_23002);
and UO_914 (O_914,N_23424,N_24721);
and UO_915 (O_915,N_23822,N_22545);
xor UO_916 (O_916,N_24423,N_22624);
nand UO_917 (O_917,N_23639,N_22773);
or UO_918 (O_918,N_23044,N_24715);
or UO_919 (O_919,N_23225,N_24932);
nor UO_920 (O_920,N_24525,N_22768);
and UO_921 (O_921,N_23376,N_24822);
and UO_922 (O_922,N_22860,N_23914);
or UO_923 (O_923,N_22859,N_24439);
xor UO_924 (O_924,N_24430,N_24457);
and UO_925 (O_925,N_22604,N_22662);
or UO_926 (O_926,N_24251,N_24449);
nand UO_927 (O_927,N_23395,N_22889);
and UO_928 (O_928,N_24623,N_23459);
and UO_929 (O_929,N_23366,N_24063);
xnor UO_930 (O_930,N_23916,N_24101);
or UO_931 (O_931,N_22641,N_24983);
nor UO_932 (O_932,N_22518,N_22627);
or UO_933 (O_933,N_24605,N_23957);
or UO_934 (O_934,N_24960,N_23347);
nand UO_935 (O_935,N_23096,N_24575);
nor UO_936 (O_936,N_24963,N_22930);
or UO_937 (O_937,N_23911,N_24851);
nand UO_938 (O_938,N_23812,N_23948);
nor UO_939 (O_939,N_22989,N_24259);
and UO_940 (O_940,N_23070,N_24542);
nand UO_941 (O_941,N_24796,N_24006);
nor UO_942 (O_942,N_24751,N_24242);
and UO_943 (O_943,N_23592,N_23231);
nor UO_944 (O_944,N_23494,N_22678);
xor UO_945 (O_945,N_22910,N_22562);
and UO_946 (O_946,N_23930,N_24595);
xnor UO_947 (O_947,N_23970,N_23825);
nor UO_948 (O_948,N_24831,N_24875);
and UO_949 (O_949,N_22804,N_24957);
and UO_950 (O_950,N_24574,N_24424);
or UO_951 (O_951,N_22588,N_24127);
or UO_952 (O_952,N_22640,N_22797);
xor UO_953 (O_953,N_24591,N_23575);
or UO_954 (O_954,N_23045,N_24898);
xnor UO_955 (O_955,N_24179,N_22757);
and UO_956 (O_956,N_24566,N_24224);
or UO_957 (O_957,N_22937,N_23785);
xnor UO_958 (O_958,N_24473,N_23478);
nor UO_959 (O_959,N_23622,N_23152);
nor UO_960 (O_960,N_24284,N_24437);
and UO_961 (O_961,N_23363,N_23888);
and UO_962 (O_962,N_22687,N_24815);
xor UO_963 (O_963,N_23539,N_24274);
or UO_964 (O_964,N_24980,N_23284);
or UO_965 (O_965,N_24710,N_23594);
xnor UO_966 (O_966,N_22769,N_23697);
xor UO_967 (O_967,N_22821,N_23876);
xnor UO_968 (O_968,N_24045,N_23540);
xor UO_969 (O_969,N_22780,N_24882);
nand UO_970 (O_970,N_24890,N_22794);
nand UO_971 (O_971,N_22510,N_23429);
or UO_972 (O_972,N_24640,N_23235);
nor UO_973 (O_973,N_23588,N_24722);
or UO_974 (O_974,N_23991,N_24374);
and UO_975 (O_975,N_22751,N_24111);
nand UO_976 (O_976,N_24402,N_23604);
nand UO_977 (O_977,N_22597,N_23350);
xnor UO_978 (O_978,N_23378,N_24700);
nor UO_979 (O_979,N_24131,N_23591);
xor UO_980 (O_980,N_24293,N_23802);
xnor UO_981 (O_981,N_22947,N_23474);
xor UO_982 (O_982,N_24995,N_23616);
nand UO_983 (O_983,N_24160,N_22735);
nand UO_984 (O_984,N_24054,N_22603);
xnor UO_985 (O_985,N_24672,N_23904);
and UO_986 (O_986,N_23810,N_23956);
nand UO_987 (O_987,N_24838,N_23717);
and UO_988 (O_988,N_23404,N_23848);
nand UO_989 (O_989,N_24731,N_23331);
nand UO_990 (O_990,N_24086,N_24544);
or UO_991 (O_991,N_24228,N_24648);
or UO_992 (O_992,N_24719,N_24812);
and UO_993 (O_993,N_23917,N_23219);
or UO_994 (O_994,N_24949,N_23729);
nand UO_995 (O_995,N_23963,N_22607);
or UO_996 (O_996,N_24142,N_23458);
or UO_997 (O_997,N_22577,N_24300);
and UO_998 (O_998,N_24570,N_24235);
and UO_999 (O_999,N_23520,N_22776);
and UO_1000 (O_1000,N_22927,N_24638);
nand UO_1001 (O_1001,N_23226,N_22651);
nand UO_1002 (O_1002,N_24385,N_22781);
nand UO_1003 (O_1003,N_23969,N_22842);
nand UO_1004 (O_1004,N_23344,N_24626);
xor UO_1005 (O_1005,N_24706,N_23220);
and UO_1006 (O_1006,N_24789,N_22898);
and UO_1007 (O_1007,N_22690,N_24238);
xor UO_1008 (O_1008,N_23341,N_23493);
xnor UO_1009 (O_1009,N_23792,N_23990);
and UO_1010 (O_1010,N_23151,N_24558);
nor UO_1011 (O_1011,N_24592,N_23788);
or UO_1012 (O_1012,N_24432,N_23994);
xor UO_1013 (O_1013,N_23037,N_22764);
xnor UO_1014 (O_1014,N_23821,N_23090);
nand UO_1015 (O_1015,N_24688,N_24436);
nor UO_1016 (O_1016,N_24729,N_24459);
xor UO_1017 (O_1017,N_23402,N_23995);
or UO_1018 (O_1018,N_22521,N_23665);
xor UO_1019 (O_1019,N_23646,N_24400);
or UO_1020 (O_1020,N_23286,N_23186);
and UO_1021 (O_1021,N_23442,N_23314);
nor UO_1022 (O_1022,N_24351,N_22829);
or UO_1023 (O_1023,N_23135,N_24866);
or UO_1024 (O_1024,N_24220,N_24074);
nand UO_1025 (O_1025,N_22932,N_22953);
nand UO_1026 (O_1026,N_22696,N_23940);
nor UO_1027 (O_1027,N_24528,N_24241);
or UO_1028 (O_1028,N_24367,N_24675);
nand UO_1029 (O_1029,N_24904,N_22556);
or UO_1030 (O_1030,N_23005,N_22816);
nand UO_1031 (O_1031,N_22655,N_24377);
nand UO_1032 (O_1032,N_23880,N_22618);
and UO_1033 (O_1033,N_23490,N_22677);
or UO_1034 (O_1034,N_24615,N_23178);
nor UO_1035 (O_1035,N_22530,N_23511);
and UO_1036 (O_1036,N_24515,N_23558);
or UO_1037 (O_1037,N_24818,N_24253);
or UO_1038 (O_1038,N_24484,N_24442);
nor UO_1039 (O_1039,N_23173,N_22855);
nand UO_1040 (O_1040,N_24215,N_23968);
and UO_1041 (O_1041,N_22730,N_22880);
xor UO_1042 (O_1042,N_23171,N_23432);
nand UO_1043 (O_1043,N_22688,N_24441);
or UO_1044 (O_1044,N_23266,N_22985);
nand UO_1045 (O_1045,N_24438,N_23356);
nand UO_1046 (O_1046,N_23385,N_22771);
nor UO_1047 (O_1047,N_23784,N_24538);
nand UO_1048 (O_1048,N_24507,N_22670);
nor UO_1049 (O_1049,N_22817,N_22848);
xor UO_1050 (O_1050,N_24479,N_24755);
and UO_1051 (O_1051,N_23703,N_24070);
nand UO_1052 (O_1052,N_23192,N_24997);
nor UO_1053 (O_1053,N_24418,N_22920);
or UO_1054 (O_1054,N_23382,N_23596);
nand UO_1055 (O_1055,N_24597,N_22939);
xor UO_1056 (O_1056,N_23585,N_23608);
xor UO_1057 (O_1057,N_24221,N_23048);
xor UO_1058 (O_1058,N_24401,N_23301);
nor UO_1059 (O_1059,N_24016,N_22642);
or UO_1060 (O_1060,N_22731,N_22867);
and UO_1061 (O_1061,N_23741,N_24776);
nand UO_1062 (O_1062,N_24523,N_22623);
nand UO_1063 (O_1063,N_23964,N_22772);
xnor UO_1064 (O_1064,N_24372,N_24292);
nand UO_1065 (O_1065,N_23457,N_22720);
nor UO_1066 (O_1066,N_24669,N_23986);
or UO_1067 (O_1067,N_23879,N_24987);
nor UO_1068 (O_1068,N_24230,N_23466);
nor UO_1069 (O_1069,N_22891,N_23000);
nand UO_1070 (O_1070,N_24007,N_24448);
nand UO_1071 (O_1071,N_24153,N_24406);
or UO_1072 (O_1072,N_22770,N_23728);
nor UO_1073 (O_1073,N_23093,N_23068);
xnor UO_1074 (O_1074,N_23205,N_22865);
nand UO_1075 (O_1075,N_23030,N_23109);
and UO_1076 (O_1076,N_23636,N_24900);
xor UO_1077 (O_1077,N_23176,N_22813);
or UO_1078 (O_1078,N_23907,N_24610);
nor UO_1079 (O_1079,N_24114,N_24028);
nor UO_1080 (O_1080,N_24005,N_24734);
or UO_1081 (O_1081,N_23480,N_23777);
nand UO_1082 (O_1082,N_23832,N_23012);
or UO_1083 (O_1083,N_23707,N_22701);
or UO_1084 (O_1084,N_24331,N_23855);
or UO_1085 (O_1085,N_24389,N_22904);
nand UO_1086 (O_1086,N_22900,N_23312);
or UO_1087 (O_1087,N_23126,N_24557);
and UO_1088 (O_1088,N_23972,N_24147);
xor UO_1089 (O_1089,N_24799,N_23633);
or UO_1090 (O_1090,N_24848,N_24032);
nand UO_1091 (O_1091,N_22787,N_24531);
or UO_1092 (O_1092,N_22581,N_23781);
xnor UO_1093 (O_1093,N_22823,N_24261);
nor UO_1094 (O_1094,N_22705,N_24132);
nand UO_1095 (O_1095,N_23329,N_23481);
and UO_1096 (O_1096,N_23873,N_22940);
or UO_1097 (O_1097,N_24535,N_23705);
or UO_1098 (O_1098,N_23727,N_23162);
or UO_1099 (O_1099,N_23656,N_22883);
and UO_1100 (O_1100,N_23256,N_23962);
and UO_1101 (O_1101,N_23807,N_24030);
nand UO_1102 (O_1102,N_23110,N_23553);
or UO_1103 (O_1103,N_23334,N_23901);
nor UO_1104 (O_1104,N_23648,N_24536);
nand UO_1105 (O_1105,N_23603,N_24926);
and UO_1106 (O_1106,N_22576,N_24206);
or UO_1107 (O_1107,N_23407,N_23795);
or UO_1108 (O_1108,N_23097,N_23421);
xnor UO_1109 (O_1109,N_23997,N_23650);
or UO_1110 (O_1110,N_22979,N_23317);
nor UO_1111 (O_1111,N_24475,N_24260);
and UO_1112 (O_1112,N_23818,N_23342);
nand UO_1113 (O_1113,N_23267,N_24942);
or UO_1114 (O_1114,N_23654,N_22650);
nor UO_1115 (O_1115,N_23495,N_23760);
nor UO_1116 (O_1116,N_24691,N_22993);
xnor UO_1117 (O_1117,N_24696,N_24226);
xnor UO_1118 (O_1118,N_24690,N_22691);
or UO_1119 (O_1119,N_23189,N_22578);
xor UO_1120 (O_1120,N_24604,N_23866);
or UO_1121 (O_1121,N_23261,N_23611);
xnor UO_1122 (O_1122,N_24427,N_24414);
xor UO_1123 (O_1123,N_23689,N_24428);
and UO_1124 (O_1124,N_24564,N_23158);
nor UO_1125 (O_1125,N_23791,N_22520);
or UO_1126 (O_1126,N_23099,N_24271);
or UO_1127 (O_1127,N_24069,N_23730);
or UO_1128 (O_1128,N_22795,N_22763);
nand UO_1129 (O_1129,N_24625,N_24480);
nor UO_1130 (O_1130,N_22694,N_23263);
xor UO_1131 (O_1131,N_23631,N_24647);
nor UO_1132 (O_1132,N_24683,N_24837);
xor UO_1133 (O_1133,N_23847,N_24925);
xnor UO_1134 (O_1134,N_24068,N_24513);
xnor UO_1135 (O_1135,N_23764,N_22921);
and UO_1136 (O_1136,N_23303,N_22724);
nand UO_1137 (O_1137,N_23615,N_24667);
nor UO_1138 (O_1138,N_24552,N_23120);
xor UO_1139 (O_1139,N_22715,N_22942);
or UO_1140 (O_1140,N_22540,N_23501);
nand UO_1141 (O_1141,N_23036,N_24847);
nor UO_1142 (O_1142,N_24141,N_23661);
and UO_1143 (O_1143,N_23428,N_23438);
nand UO_1144 (O_1144,N_24723,N_23201);
nor UO_1145 (O_1145,N_24965,N_24079);
and UO_1146 (O_1146,N_24855,N_22554);
nor UO_1147 (O_1147,N_24694,N_22759);
xor UO_1148 (O_1148,N_23132,N_22639);
and UO_1149 (O_1149,N_24912,N_24483);
xnor UO_1150 (O_1150,N_22616,N_23298);
xor UO_1151 (O_1151,N_23328,N_23936);
xnor UO_1152 (O_1152,N_23308,N_24573);
nand UO_1153 (O_1153,N_24165,N_24098);
or UO_1154 (O_1154,N_22774,N_23941);
and UO_1155 (O_1155,N_22911,N_24717);
or UO_1156 (O_1156,N_24917,N_23814);
nor UO_1157 (O_1157,N_24314,N_23973);
and UO_1158 (O_1158,N_23210,N_22689);
and UO_1159 (O_1159,N_24632,N_23403);
xnor UO_1160 (O_1160,N_23058,N_23156);
or UO_1161 (O_1161,N_22862,N_24463);
or UO_1162 (O_1162,N_24662,N_23658);
xor UO_1163 (O_1163,N_23059,N_24135);
and UO_1164 (O_1164,N_23335,N_22517);
xnor UO_1165 (O_1165,N_23937,N_23041);
and UO_1166 (O_1166,N_22847,N_22967);
nand UO_1167 (O_1167,N_23578,N_24537);
and UO_1168 (O_1168,N_24486,N_23976);
or UO_1169 (O_1169,N_24679,N_24106);
or UO_1170 (O_1170,N_23602,N_24695);
and UO_1171 (O_1171,N_23686,N_22831);
nand UO_1172 (O_1172,N_23319,N_23285);
or UO_1173 (O_1173,N_24426,N_23756);
nand UO_1174 (O_1174,N_23945,N_22621);
nor UO_1175 (O_1175,N_24644,N_24859);
nand UO_1176 (O_1176,N_23702,N_22601);
and UO_1177 (O_1177,N_24740,N_23211);
nor UO_1178 (O_1178,N_24031,N_23121);
and UO_1179 (O_1179,N_24399,N_24487);
and UO_1180 (O_1180,N_24236,N_22729);
xnor UO_1181 (O_1181,N_24940,N_24003);
or UO_1182 (O_1182,N_24237,N_23584);
or UO_1183 (O_1183,N_22598,N_23164);
xnor UO_1184 (O_1184,N_23305,N_24136);
nor UO_1185 (O_1185,N_24616,N_24985);
nand UO_1186 (O_1186,N_23675,N_24008);
xnor UO_1187 (O_1187,N_22790,N_24870);
nand UO_1188 (O_1188,N_24836,N_24474);
and UO_1189 (O_1189,N_24371,N_22591);
and UO_1190 (O_1190,N_24955,N_24973);
nor UO_1191 (O_1191,N_22659,N_24247);
nor UO_1192 (O_1192,N_23674,N_23522);
and UO_1193 (O_1193,N_24195,N_24476);
or UO_1194 (O_1194,N_22827,N_23212);
xor UO_1195 (O_1195,N_22507,N_24485);
xnor UO_1196 (O_1196,N_22733,N_23473);
xnor UO_1197 (O_1197,N_23141,N_22992);
nand UO_1198 (O_1198,N_23078,N_22582);
nand UO_1199 (O_1199,N_23469,N_22753);
nand UO_1200 (O_1200,N_24065,N_24319);
nand UO_1201 (O_1201,N_23621,N_23725);
nand UO_1202 (O_1202,N_24378,N_24014);
and UO_1203 (O_1203,N_23043,N_24183);
and UO_1204 (O_1204,N_23853,N_24455);
nand UO_1205 (O_1205,N_24363,N_24634);
xor UO_1206 (O_1206,N_23566,N_24846);
and UO_1207 (O_1207,N_22777,N_23949);
nand UO_1208 (O_1208,N_23343,N_22590);
nor UO_1209 (O_1209,N_24919,N_24170);
xnor UO_1210 (O_1210,N_24825,N_24820);
xnor UO_1211 (O_1211,N_23083,N_23871);
or UO_1212 (O_1212,N_22500,N_23612);
nor UO_1213 (O_1213,N_24928,N_22717);
nor UO_1214 (O_1214,N_24460,N_24245);
nand UO_1215 (O_1215,N_24758,N_24278);
or UO_1216 (O_1216,N_23766,N_22996);
nand UO_1217 (O_1217,N_23958,N_23010);
xor UO_1218 (O_1218,N_22995,N_23296);
and UO_1219 (O_1219,N_23140,N_23846);
and UO_1220 (O_1220,N_22851,N_24763);
xor UO_1221 (O_1221,N_23978,N_24243);
nand UO_1222 (O_1222,N_23862,N_23450);
nand UO_1223 (O_1223,N_24204,N_24199);
or UO_1224 (O_1224,N_24123,N_22884);
and UO_1225 (O_1225,N_23640,N_23502);
nor UO_1226 (O_1226,N_22778,N_23145);
and UO_1227 (O_1227,N_22830,N_24671);
xnor UO_1228 (O_1228,N_22739,N_24529);
nand UO_1229 (O_1229,N_24565,N_23461);
xor UO_1230 (O_1230,N_24747,N_22613);
nand UO_1231 (O_1231,N_23669,N_23007);
and UO_1232 (O_1232,N_23013,N_22560);
and UO_1233 (O_1233,N_24613,N_24352);
xnor UO_1234 (O_1234,N_23813,N_23324);
or UO_1235 (O_1235,N_23770,N_22793);
or UO_1236 (O_1236,N_24984,N_23971);
xnor UO_1237 (O_1237,N_23274,N_24344);
xor UO_1238 (O_1238,N_23321,N_22929);
nor UO_1239 (O_1239,N_24856,N_24936);
nor UO_1240 (O_1240,N_24115,N_23768);
or UO_1241 (O_1241,N_23919,N_24321);
nand UO_1242 (O_1242,N_23181,N_24756);
nor UO_1243 (O_1243,N_23418,N_24770);
and UO_1244 (O_1244,N_24180,N_23840);
nand UO_1245 (O_1245,N_24982,N_24360);
nand UO_1246 (O_1246,N_23623,N_23087);
nand UO_1247 (O_1247,N_23542,N_23508);
nand UO_1248 (O_1248,N_24349,N_24365);
nand UO_1249 (O_1249,N_22748,N_23188);
or UO_1250 (O_1250,N_23098,N_24627);
nand UO_1251 (O_1251,N_22909,N_23706);
nor UO_1252 (O_1252,N_22697,N_23395);
xnor UO_1253 (O_1253,N_23561,N_24965);
nor UO_1254 (O_1254,N_24120,N_22839);
and UO_1255 (O_1255,N_23333,N_23784);
and UO_1256 (O_1256,N_24238,N_24727);
nor UO_1257 (O_1257,N_23848,N_23546);
xor UO_1258 (O_1258,N_24828,N_23562);
nand UO_1259 (O_1259,N_24631,N_24283);
nor UO_1260 (O_1260,N_23675,N_23454);
xnor UO_1261 (O_1261,N_24555,N_24288);
nor UO_1262 (O_1262,N_24173,N_23722);
and UO_1263 (O_1263,N_22526,N_22643);
or UO_1264 (O_1264,N_24934,N_23716);
nand UO_1265 (O_1265,N_24628,N_22860);
or UO_1266 (O_1266,N_24072,N_24236);
xor UO_1267 (O_1267,N_24783,N_24577);
nor UO_1268 (O_1268,N_24759,N_23367);
xor UO_1269 (O_1269,N_24090,N_24061);
nand UO_1270 (O_1270,N_22694,N_22963);
and UO_1271 (O_1271,N_22750,N_22662);
nor UO_1272 (O_1272,N_23906,N_22609);
nand UO_1273 (O_1273,N_22650,N_23536);
or UO_1274 (O_1274,N_24811,N_23682);
nand UO_1275 (O_1275,N_23095,N_22957);
or UO_1276 (O_1276,N_24140,N_24820);
and UO_1277 (O_1277,N_22636,N_22813);
nor UO_1278 (O_1278,N_24410,N_23579);
nor UO_1279 (O_1279,N_24545,N_24564);
nand UO_1280 (O_1280,N_24605,N_24550);
nand UO_1281 (O_1281,N_23063,N_24127);
or UO_1282 (O_1282,N_22968,N_24096);
nand UO_1283 (O_1283,N_23526,N_23049);
and UO_1284 (O_1284,N_24317,N_23123);
and UO_1285 (O_1285,N_24923,N_23952);
nand UO_1286 (O_1286,N_23074,N_24628);
and UO_1287 (O_1287,N_24944,N_22619);
or UO_1288 (O_1288,N_24246,N_23099);
nand UO_1289 (O_1289,N_22797,N_23953);
xnor UO_1290 (O_1290,N_24762,N_23418);
and UO_1291 (O_1291,N_23720,N_24625);
xor UO_1292 (O_1292,N_24352,N_24146);
xnor UO_1293 (O_1293,N_22915,N_24104);
or UO_1294 (O_1294,N_24591,N_23206);
or UO_1295 (O_1295,N_23678,N_23892);
nor UO_1296 (O_1296,N_23820,N_24104);
xnor UO_1297 (O_1297,N_23516,N_22910);
or UO_1298 (O_1298,N_23512,N_23098);
xor UO_1299 (O_1299,N_22813,N_22916);
xor UO_1300 (O_1300,N_23130,N_23437);
or UO_1301 (O_1301,N_23411,N_24305);
xor UO_1302 (O_1302,N_22594,N_24422);
nor UO_1303 (O_1303,N_24894,N_23927);
xnor UO_1304 (O_1304,N_24692,N_24446);
and UO_1305 (O_1305,N_24579,N_24893);
and UO_1306 (O_1306,N_23009,N_24580);
or UO_1307 (O_1307,N_23039,N_23866);
xor UO_1308 (O_1308,N_23825,N_24609);
and UO_1309 (O_1309,N_24875,N_24660);
nor UO_1310 (O_1310,N_22813,N_22634);
and UO_1311 (O_1311,N_24550,N_23821);
nand UO_1312 (O_1312,N_23522,N_24585);
nand UO_1313 (O_1313,N_24039,N_24452);
nand UO_1314 (O_1314,N_24116,N_23393);
or UO_1315 (O_1315,N_24354,N_24788);
and UO_1316 (O_1316,N_23141,N_24143);
or UO_1317 (O_1317,N_24488,N_24334);
or UO_1318 (O_1318,N_22927,N_24194);
or UO_1319 (O_1319,N_23875,N_24755);
nand UO_1320 (O_1320,N_24031,N_23573);
or UO_1321 (O_1321,N_23861,N_24491);
xor UO_1322 (O_1322,N_23391,N_24568);
nor UO_1323 (O_1323,N_24588,N_22629);
xor UO_1324 (O_1324,N_24081,N_23443);
or UO_1325 (O_1325,N_23868,N_23863);
xor UO_1326 (O_1326,N_24414,N_24552);
nand UO_1327 (O_1327,N_23433,N_24506);
xor UO_1328 (O_1328,N_24529,N_23986);
nor UO_1329 (O_1329,N_24457,N_22585);
nor UO_1330 (O_1330,N_23982,N_24395);
nand UO_1331 (O_1331,N_24006,N_23643);
nor UO_1332 (O_1332,N_22527,N_24559);
nand UO_1333 (O_1333,N_22792,N_24787);
nand UO_1334 (O_1334,N_24767,N_23985);
nor UO_1335 (O_1335,N_24903,N_23239);
or UO_1336 (O_1336,N_24189,N_23271);
and UO_1337 (O_1337,N_24103,N_24969);
or UO_1338 (O_1338,N_22521,N_23479);
xor UO_1339 (O_1339,N_23040,N_22556);
and UO_1340 (O_1340,N_24757,N_24153);
nor UO_1341 (O_1341,N_23270,N_23434);
or UO_1342 (O_1342,N_22723,N_24562);
and UO_1343 (O_1343,N_23043,N_22989);
nor UO_1344 (O_1344,N_23790,N_23085);
nor UO_1345 (O_1345,N_24074,N_24159);
xnor UO_1346 (O_1346,N_24267,N_23896);
xor UO_1347 (O_1347,N_23245,N_24803);
nor UO_1348 (O_1348,N_23535,N_22802);
or UO_1349 (O_1349,N_22856,N_23479);
and UO_1350 (O_1350,N_23210,N_23798);
xor UO_1351 (O_1351,N_24252,N_24045);
xor UO_1352 (O_1352,N_22703,N_24357);
nand UO_1353 (O_1353,N_23421,N_22848);
xnor UO_1354 (O_1354,N_22565,N_23792);
nor UO_1355 (O_1355,N_24567,N_24614);
nor UO_1356 (O_1356,N_23867,N_22691);
nand UO_1357 (O_1357,N_24047,N_23020);
or UO_1358 (O_1358,N_23950,N_22639);
nor UO_1359 (O_1359,N_24845,N_23818);
nor UO_1360 (O_1360,N_23156,N_23688);
or UO_1361 (O_1361,N_22951,N_24339);
and UO_1362 (O_1362,N_22689,N_23314);
xnor UO_1363 (O_1363,N_24171,N_24460);
nor UO_1364 (O_1364,N_23610,N_23611);
xnor UO_1365 (O_1365,N_23676,N_22625);
nand UO_1366 (O_1366,N_23945,N_23771);
xnor UO_1367 (O_1367,N_22668,N_23406);
or UO_1368 (O_1368,N_23366,N_23437);
nor UO_1369 (O_1369,N_23992,N_23896);
nand UO_1370 (O_1370,N_24424,N_22574);
and UO_1371 (O_1371,N_24871,N_24318);
nand UO_1372 (O_1372,N_22983,N_24278);
nor UO_1373 (O_1373,N_24587,N_22801);
or UO_1374 (O_1374,N_22920,N_23595);
xnor UO_1375 (O_1375,N_23233,N_22900);
and UO_1376 (O_1376,N_23052,N_23307);
xnor UO_1377 (O_1377,N_23010,N_24786);
nand UO_1378 (O_1378,N_24315,N_23014);
nor UO_1379 (O_1379,N_23445,N_23983);
nand UO_1380 (O_1380,N_24544,N_22549);
nor UO_1381 (O_1381,N_23500,N_24143);
or UO_1382 (O_1382,N_23898,N_23437);
or UO_1383 (O_1383,N_23129,N_23951);
nand UO_1384 (O_1384,N_24407,N_24307);
nand UO_1385 (O_1385,N_23876,N_24889);
nor UO_1386 (O_1386,N_23729,N_24389);
nand UO_1387 (O_1387,N_24182,N_22685);
xor UO_1388 (O_1388,N_24645,N_22903);
nor UO_1389 (O_1389,N_22948,N_23161);
xnor UO_1390 (O_1390,N_22551,N_24098);
xor UO_1391 (O_1391,N_23257,N_23634);
xor UO_1392 (O_1392,N_23298,N_24475);
xor UO_1393 (O_1393,N_24244,N_24948);
and UO_1394 (O_1394,N_24713,N_24960);
and UO_1395 (O_1395,N_24329,N_23276);
nor UO_1396 (O_1396,N_23430,N_24942);
nor UO_1397 (O_1397,N_24569,N_22685);
nand UO_1398 (O_1398,N_24794,N_24049);
nor UO_1399 (O_1399,N_22613,N_23083);
xor UO_1400 (O_1400,N_24955,N_24374);
xnor UO_1401 (O_1401,N_24512,N_23026);
nand UO_1402 (O_1402,N_23678,N_23968);
nor UO_1403 (O_1403,N_24334,N_23165);
xor UO_1404 (O_1404,N_23054,N_24318);
xnor UO_1405 (O_1405,N_24620,N_23648);
xor UO_1406 (O_1406,N_24084,N_24336);
nand UO_1407 (O_1407,N_22929,N_22798);
and UO_1408 (O_1408,N_23756,N_22719);
nand UO_1409 (O_1409,N_24466,N_23476);
or UO_1410 (O_1410,N_23124,N_23445);
or UO_1411 (O_1411,N_23501,N_23117);
and UO_1412 (O_1412,N_24997,N_24087);
nor UO_1413 (O_1413,N_23347,N_22523);
xnor UO_1414 (O_1414,N_23050,N_24731);
and UO_1415 (O_1415,N_24680,N_24819);
xnor UO_1416 (O_1416,N_24572,N_24290);
or UO_1417 (O_1417,N_23008,N_24722);
xor UO_1418 (O_1418,N_24977,N_23125);
and UO_1419 (O_1419,N_22535,N_23563);
xnor UO_1420 (O_1420,N_22670,N_23711);
or UO_1421 (O_1421,N_24497,N_23056);
nand UO_1422 (O_1422,N_23125,N_24325);
and UO_1423 (O_1423,N_24027,N_23539);
nor UO_1424 (O_1424,N_23876,N_22815);
or UO_1425 (O_1425,N_23232,N_23859);
nand UO_1426 (O_1426,N_24232,N_23385);
xor UO_1427 (O_1427,N_24432,N_22965);
or UO_1428 (O_1428,N_23759,N_23549);
nor UO_1429 (O_1429,N_23466,N_24949);
nor UO_1430 (O_1430,N_23820,N_23048);
nor UO_1431 (O_1431,N_23301,N_24490);
or UO_1432 (O_1432,N_24408,N_23724);
nand UO_1433 (O_1433,N_24337,N_23951);
or UO_1434 (O_1434,N_24393,N_23267);
nor UO_1435 (O_1435,N_24666,N_22545);
or UO_1436 (O_1436,N_23302,N_24069);
and UO_1437 (O_1437,N_23957,N_22989);
nor UO_1438 (O_1438,N_24197,N_22702);
or UO_1439 (O_1439,N_23892,N_23199);
nor UO_1440 (O_1440,N_24594,N_24807);
xnor UO_1441 (O_1441,N_23421,N_22615);
nor UO_1442 (O_1442,N_23852,N_22606);
and UO_1443 (O_1443,N_23542,N_23316);
nand UO_1444 (O_1444,N_23083,N_24870);
nor UO_1445 (O_1445,N_24073,N_23323);
or UO_1446 (O_1446,N_23084,N_23757);
nand UO_1447 (O_1447,N_23951,N_22932);
nor UO_1448 (O_1448,N_23412,N_23058);
nand UO_1449 (O_1449,N_22970,N_23197);
nor UO_1450 (O_1450,N_22683,N_22606);
or UO_1451 (O_1451,N_23931,N_22853);
nor UO_1452 (O_1452,N_23311,N_24499);
xor UO_1453 (O_1453,N_23764,N_23780);
or UO_1454 (O_1454,N_22721,N_24608);
nand UO_1455 (O_1455,N_24046,N_24296);
or UO_1456 (O_1456,N_22504,N_24329);
nand UO_1457 (O_1457,N_23916,N_23311);
and UO_1458 (O_1458,N_23656,N_24011);
nor UO_1459 (O_1459,N_23013,N_23951);
nor UO_1460 (O_1460,N_23335,N_23088);
or UO_1461 (O_1461,N_23883,N_23739);
nand UO_1462 (O_1462,N_23273,N_23601);
nor UO_1463 (O_1463,N_22606,N_22855);
and UO_1464 (O_1464,N_23379,N_23639);
and UO_1465 (O_1465,N_23980,N_23102);
nor UO_1466 (O_1466,N_22864,N_24817);
nor UO_1467 (O_1467,N_22763,N_24937);
nor UO_1468 (O_1468,N_22863,N_23259);
and UO_1469 (O_1469,N_24746,N_23551);
or UO_1470 (O_1470,N_22506,N_22593);
nand UO_1471 (O_1471,N_23552,N_23116);
or UO_1472 (O_1472,N_23710,N_23195);
xor UO_1473 (O_1473,N_22881,N_24241);
or UO_1474 (O_1474,N_24273,N_24855);
xnor UO_1475 (O_1475,N_23198,N_24139);
or UO_1476 (O_1476,N_23996,N_24973);
nor UO_1477 (O_1477,N_23475,N_24243);
and UO_1478 (O_1478,N_24506,N_23108);
nand UO_1479 (O_1479,N_24819,N_23439);
nand UO_1480 (O_1480,N_23375,N_24192);
or UO_1481 (O_1481,N_22709,N_24959);
or UO_1482 (O_1482,N_23775,N_23214);
nor UO_1483 (O_1483,N_24453,N_22923);
xnor UO_1484 (O_1484,N_24534,N_23886);
nand UO_1485 (O_1485,N_24726,N_24380);
or UO_1486 (O_1486,N_23255,N_24128);
nand UO_1487 (O_1487,N_22936,N_24198);
nand UO_1488 (O_1488,N_22864,N_24467);
and UO_1489 (O_1489,N_22979,N_24619);
nand UO_1490 (O_1490,N_22781,N_23845);
xnor UO_1491 (O_1491,N_24730,N_24432);
and UO_1492 (O_1492,N_23136,N_23065);
nor UO_1493 (O_1493,N_23557,N_24538);
or UO_1494 (O_1494,N_23898,N_24026);
xnor UO_1495 (O_1495,N_23793,N_24870);
or UO_1496 (O_1496,N_23938,N_22607);
nand UO_1497 (O_1497,N_22589,N_22733);
nand UO_1498 (O_1498,N_24747,N_24563);
nand UO_1499 (O_1499,N_24981,N_23515);
or UO_1500 (O_1500,N_22564,N_22737);
xor UO_1501 (O_1501,N_24812,N_24933);
or UO_1502 (O_1502,N_22684,N_24466);
and UO_1503 (O_1503,N_23128,N_24158);
and UO_1504 (O_1504,N_24089,N_23096);
nor UO_1505 (O_1505,N_22633,N_24988);
or UO_1506 (O_1506,N_24103,N_24838);
or UO_1507 (O_1507,N_24602,N_22752);
xor UO_1508 (O_1508,N_24434,N_24391);
or UO_1509 (O_1509,N_23910,N_24077);
nand UO_1510 (O_1510,N_24632,N_23882);
nor UO_1511 (O_1511,N_22867,N_23457);
and UO_1512 (O_1512,N_24983,N_22861);
or UO_1513 (O_1513,N_22573,N_24546);
nor UO_1514 (O_1514,N_23700,N_24017);
nor UO_1515 (O_1515,N_22956,N_23937);
xnor UO_1516 (O_1516,N_24076,N_24212);
nand UO_1517 (O_1517,N_22523,N_23304);
nor UO_1518 (O_1518,N_24150,N_24968);
nand UO_1519 (O_1519,N_24948,N_22591);
and UO_1520 (O_1520,N_24556,N_23804);
or UO_1521 (O_1521,N_22936,N_24340);
and UO_1522 (O_1522,N_24237,N_23636);
nor UO_1523 (O_1523,N_22835,N_23209);
or UO_1524 (O_1524,N_23846,N_24313);
nor UO_1525 (O_1525,N_22545,N_22584);
nand UO_1526 (O_1526,N_22652,N_23547);
nand UO_1527 (O_1527,N_22805,N_23180);
xnor UO_1528 (O_1528,N_24309,N_24441);
nand UO_1529 (O_1529,N_22839,N_23782);
nor UO_1530 (O_1530,N_24396,N_24653);
or UO_1531 (O_1531,N_24649,N_24755);
nor UO_1532 (O_1532,N_22832,N_24986);
and UO_1533 (O_1533,N_23370,N_24634);
xor UO_1534 (O_1534,N_22843,N_24161);
and UO_1535 (O_1535,N_23027,N_23598);
nand UO_1536 (O_1536,N_24653,N_24843);
nand UO_1537 (O_1537,N_22950,N_23607);
nand UO_1538 (O_1538,N_24042,N_24525);
and UO_1539 (O_1539,N_24074,N_24882);
and UO_1540 (O_1540,N_23859,N_23425);
and UO_1541 (O_1541,N_22652,N_22688);
xor UO_1542 (O_1542,N_23451,N_23639);
nor UO_1543 (O_1543,N_24829,N_22893);
xor UO_1544 (O_1544,N_24608,N_22801);
nor UO_1545 (O_1545,N_23868,N_22554);
nand UO_1546 (O_1546,N_24547,N_24811);
xnor UO_1547 (O_1547,N_23546,N_22618);
nor UO_1548 (O_1548,N_23027,N_24198);
and UO_1549 (O_1549,N_24190,N_24114);
or UO_1550 (O_1550,N_24800,N_23239);
nor UO_1551 (O_1551,N_22523,N_23069);
and UO_1552 (O_1552,N_22714,N_24488);
nand UO_1553 (O_1553,N_23061,N_22861);
or UO_1554 (O_1554,N_23960,N_24024);
or UO_1555 (O_1555,N_24014,N_24766);
nand UO_1556 (O_1556,N_23835,N_24427);
and UO_1557 (O_1557,N_24684,N_22666);
nand UO_1558 (O_1558,N_24980,N_23250);
and UO_1559 (O_1559,N_24779,N_22755);
and UO_1560 (O_1560,N_22604,N_24357);
nor UO_1561 (O_1561,N_23356,N_22867);
or UO_1562 (O_1562,N_24826,N_24424);
and UO_1563 (O_1563,N_24726,N_23141);
and UO_1564 (O_1564,N_22795,N_23794);
or UO_1565 (O_1565,N_23571,N_24501);
or UO_1566 (O_1566,N_24395,N_24119);
or UO_1567 (O_1567,N_24367,N_24578);
nor UO_1568 (O_1568,N_24540,N_24088);
nor UO_1569 (O_1569,N_24569,N_23626);
or UO_1570 (O_1570,N_23175,N_24198);
or UO_1571 (O_1571,N_23305,N_24194);
and UO_1572 (O_1572,N_22501,N_23647);
and UO_1573 (O_1573,N_23806,N_23647);
or UO_1574 (O_1574,N_24317,N_24926);
nand UO_1575 (O_1575,N_23007,N_24566);
and UO_1576 (O_1576,N_23648,N_22703);
and UO_1577 (O_1577,N_22601,N_23723);
xor UO_1578 (O_1578,N_24932,N_22716);
nor UO_1579 (O_1579,N_23600,N_22658);
xnor UO_1580 (O_1580,N_22852,N_23363);
nand UO_1581 (O_1581,N_24317,N_22862);
or UO_1582 (O_1582,N_24373,N_24513);
or UO_1583 (O_1583,N_24506,N_24723);
nand UO_1584 (O_1584,N_23721,N_23272);
or UO_1585 (O_1585,N_24313,N_23272);
and UO_1586 (O_1586,N_23556,N_22575);
xnor UO_1587 (O_1587,N_22514,N_24563);
xnor UO_1588 (O_1588,N_22588,N_23257);
xnor UO_1589 (O_1589,N_22548,N_23153);
nand UO_1590 (O_1590,N_24697,N_24014);
nand UO_1591 (O_1591,N_23444,N_23940);
nand UO_1592 (O_1592,N_22970,N_24904);
nand UO_1593 (O_1593,N_24087,N_23418);
xor UO_1594 (O_1594,N_22933,N_24899);
or UO_1595 (O_1595,N_23344,N_22780);
nand UO_1596 (O_1596,N_24873,N_22517);
nor UO_1597 (O_1597,N_23582,N_22926);
and UO_1598 (O_1598,N_24997,N_24560);
and UO_1599 (O_1599,N_23783,N_24803);
nand UO_1600 (O_1600,N_24151,N_24563);
xor UO_1601 (O_1601,N_23785,N_24537);
and UO_1602 (O_1602,N_24077,N_22812);
or UO_1603 (O_1603,N_23883,N_23452);
xor UO_1604 (O_1604,N_24385,N_23654);
nor UO_1605 (O_1605,N_24333,N_22952);
xnor UO_1606 (O_1606,N_23976,N_23083);
nor UO_1607 (O_1607,N_23628,N_23422);
nor UO_1608 (O_1608,N_22991,N_24188);
xnor UO_1609 (O_1609,N_22959,N_24133);
nor UO_1610 (O_1610,N_23101,N_24536);
nand UO_1611 (O_1611,N_23754,N_23209);
nor UO_1612 (O_1612,N_23488,N_22614);
and UO_1613 (O_1613,N_22693,N_24122);
nor UO_1614 (O_1614,N_23347,N_24901);
nor UO_1615 (O_1615,N_24965,N_23521);
and UO_1616 (O_1616,N_24147,N_23132);
xor UO_1617 (O_1617,N_24848,N_24539);
and UO_1618 (O_1618,N_22803,N_24293);
or UO_1619 (O_1619,N_23313,N_24178);
nand UO_1620 (O_1620,N_23755,N_23336);
xnor UO_1621 (O_1621,N_24049,N_24873);
nor UO_1622 (O_1622,N_22951,N_23084);
and UO_1623 (O_1623,N_23725,N_23434);
nor UO_1624 (O_1624,N_23728,N_23016);
and UO_1625 (O_1625,N_23323,N_24210);
nand UO_1626 (O_1626,N_24927,N_24074);
xnor UO_1627 (O_1627,N_22577,N_24475);
and UO_1628 (O_1628,N_24458,N_24761);
nor UO_1629 (O_1629,N_24793,N_24896);
nor UO_1630 (O_1630,N_23315,N_23853);
or UO_1631 (O_1631,N_23924,N_24797);
xnor UO_1632 (O_1632,N_24886,N_24377);
xnor UO_1633 (O_1633,N_23330,N_24673);
xor UO_1634 (O_1634,N_23532,N_22860);
or UO_1635 (O_1635,N_22617,N_23947);
and UO_1636 (O_1636,N_23968,N_24273);
nor UO_1637 (O_1637,N_22839,N_23052);
nand UO_1638 (O_1638,N_24149,N_23127);
nor UO_1639 (O_1639,N_24931,N_24278);
nor UO_1640 (O_1640,N_24555,N_22585);
nor UO_1641 (O_1641,N_23996,N_22776);
and UO_1642 (O_1642,N_22869,N_22729);
nand UO_1643 (O_1643,N_23040,N_24739);
nand UO_1644 (O_1644,N_22562,N_24421);
xor UO_1645 (O_1645,N_23397,N_23626);
and UO_1646 (O_1646,N_23622,N_24634);
or UO_1647 (O_1647,N_23884,N_23033);
and UO_1648 (O_1648,N_23368,N_23574);
xor UO_1649 (O_1649,N_23115,N_24386);
and UO_1650 (O_1650,N_24701,N_22624);
nand UO_1651 (O_1651,N_24954,N_23019);
and UO_1652 (O_1652,N_22916,N_24826);
or UO_1653 (O_1653,N_22709,N_23765);
nand UO_1654 (O_1654,N_23141,N_22787);
nand UO_1655 (O_1655,N_23402,N_24935);
nor UO_1656 (O_1656,N_24327,N_24083);
nand UO_1657 (O_1657,N_24596,N_24906);
xnor UO_1658 (O_1658,N_23554,N_24877);
and UO_1659 (O_1659,N_23235,N_23942);
nor UO_1660 (O_1660,N_24255,N_23704);
or UO_1661 (O_1661,N_23532,N_23841);
nand UO_1662 (O_1662,N_24098,N_24100);
and UO_1663 (O_1663,N_23735,N_23581);
nor UO_1664 (O_1664,N_23571,N_22926);
nand UO_1665 (O_1665,N_23299,N_24072);
xnor UO_1666 (O_1666,N_24855,N_24445);
and UO_1667 (O_1667,N_24338,N_24178);
or UO_1668 (O_1668,N_23222,N_23896);
nand UO_1669 (O_1669,N_22970,N_22568);
or UO_1670 (O_1670,N_23341,N_24371);
nor UO_1671 (O_1671,N_23020,N_23370);
nand UO_1672 (O_1672,N_23108,N_23418);
nand UO_1673 (O_1673,N_22969,N_23512);
or UO_1674 (O_1674,N_23310,N_24210);
nor UO_1675 (O_1675,N_24885,N_23027);
nand UO_1676 (O_1676,N_23042,N_24975);
and UO_1677 (O_1677,N_24308,N_22876);
or UO_1678 (O_1678,N_23751,N_22967);
nand UO_1679 (O_1679,N_24748,N_24876);
or UO_1680 (O_1680,N_23128,N_22844);
nand UO_1681 (O_1681,N_23141,N_23172);
and UO_1682 (O_1682,N_24455,N_24995);
nand UO_1683 (O_1683,N_23689,N_24187);
and UO_1684 (O_1684,N_23821,N_23659);
nand UO_1685 (O_1685,N_23399,N_23451);
nand UO_1686 (O_1686,N_23399,N_24687);
nand UO_1687 (O_1687,N_24165,N_23282);
or UO_1688 (O_1688,N_24814,N_24506);
or UO_1689 (O_1689,N_24479,N_24542);
or UO_1690 (O_1690,N_22615,N_23198);
and UO_1691 (O_1691,N_24093,N_23549);
nor UO_1692 (O_1692,N_23567,N_23241);
nand UO_1693 (O_1693,N_22591,N_24028);
xor UO_1694 (O_1694,N_24893,N_24838);
nand UO_1695 (O_1695,N_24283,N_23163);
nor UO_1696 (O_1696,N_23192,N_24498);
nor UO_1697 (O_1697,N_24219,N_24409);
and UO_1698 (O_1698,N_23075,N_22712);
xor UO_1699 (O_1699,N_24972,N_24768);
nand UO_1700 (O_1700,N_22522,N_24389);
and UO_1701 (O_1701,N_23252,N_24103);
and UO_1702 (O_1702,N_24748,N_22770);
xnor UO_1703 (O_1703,N_23622,N_23048);
xnor UO_1704 (O_1704,N_23707,N_22867);
nand UO_1705 (O_1705,N_24392,N_22914);
or UO_1706 (O_1706,N_24842,N_23395);
and UO_1707 (O_1707,N_24596,N_23616);
nand UO_1708 (O_1708,N_23382,N_24511);
nand UO_1709 (O_1709,N_23171,N_23580);
nand UO_1710 (O_1710,N_24142,N_22931);
xnor UO_1711 (O_1711,N_24801,N_24426);
or UO_1712 (O_1712,N_24461,N_23057);
or UO_1713 (O_1713,N_22842,N_24514);
xnor UO_1714 (O_1714,N_24331,N_24939);
xnor UO_1715 (O_1715,N_23309,N_23734);
nor UO_1716 (O_1716,N_23829,N_24933);
nand UO_1717 (O_1717,N_24868,N_23345);
nor UO_1718 (O_1718,N_24216,N_24988);
or UO_1719 (O_1719,N_23221,N_24963);
or UO_1720 (O_1720,N_23109,N_23456);
and UO_1721 (O_1721,N_23744,N_23789);
xnor UO_1722 (O_1722,N_23620,N_22802);
nor UO_1723 (O_1723,N_22738,N_23196);
and UO_1724 (O_1724,N_23759,N_22715);
and UO_1725 (O_1725,N_24414,N_22844);
and UO_1726 (O_1726,N_23662,N_23107);
or UO_1727 (O_1727,N_22654,N_24316);
nand UO_1728 (O_1728,N_23684,N_24723);
or UO_1729 (O_1729,N_22631,N_24864);
nand UO_1730 (O_1730,N_23867,N_22576);
nor UO_1731 (O_1731,N_22901,N_22676);
nand UO_1732 (O_1732,N_24655,N_24455);
or UO_1733 (O_1733,N_23894,N_24679);
nor UO_1734 (O_1734,N_24965,N_22725);
nor UO_1735 (O_1735,N_24515,N_23252);
or UO_1736 (O_1736,N_24233,N_23817);
and UO_1737 (O_1737,N_23485,N_24067);
nand UO_1738 (O_1738,N_23168,N_23229);
nor UO_1739 (O_1739,N_23595,N_24449);
xor UO_1740 (O_1740,N_22581,N_23441);
or UO_1741 (O_1741,N_22591,N_23979);
nand UO_1742 (O_1742,N_24315,N_23128);
xor UO_1743 (O_1743,N_24395,N_22626);
xor UO_1744 (O_1744,N_24833,N_24594);
xor UO_1745 (O_1745,N_23413,N_24080);
xnor UO_1746 (O_1746,N_23992,N_23670);
or UO_1747 (O_1747,N_24021,N_24125);
or UO_1748 (O_1748,N_24860,N_23730);
nor UO_1749 (O_1749,N_23154,N_24357);
xor UO_1750 (O_1750,N_23118,N_23494);
or UO_1751 (O_1751,N_22999,N_23533);
nor UO_1752 (O_1752,N_24653,N_24233);
or UO_1753 (O_1753,N_24397,N_22665);
and UO_1754 (O_1754,N_24338,N_24661);
xnor UO_1755 (O_1755,N_22642,N_22754);
and UO_1756 (O_1756,N_23716,N_24660);
nand UO_1757 (O_1757,N_24405,N_24231);
or UO_1758 (O_1758,N_23941,N_22988);
nand UO_1759 (O_1759,N_24225,N_23387);
and UO_1760 (O_1760,N_23461,N_23139);
and UO_1761 (O_1761,N_22606,N_23235);
and UO_1762 (O_1762,N_24679,N_23713);
nor UO_1763 (O_1763,N_22918,N_24070);
and UO_1764 (O_1764,N_24743,N_24494);
xnor UO_1765 (O_1765,N_24266,N_24520);
and UO_1766 (O_1766,N_22585,N_24324);
or UO_1767 (O_1767,N_22573,N_24552);
xnor UO_1768 (O_1768,N_24600,N_23525);
and UO_1769 (O_1769,N_22771,N_24231);
nand UO_1770 (O_1770,N_22871,N_23877);
or UO_1771 (O_1771,N_23726,N_24623);
xor UO_1772 (O_1772,N_24879,N_23632);
or UO_1773 (O_1773,N_24339,N_23416);
nand UO_1774 (O_1774,N_23311,N_24502);
xnor UO_1775 (O_1775,N_23401,N_23450);
xor UO_1776 (O_1776,N_24881,N_24061);
and UO_1777 (O_1777,N_24269,N_23636);
nand UO_1778 (O_1778,N_22729,N_24718);
nor UO_1779 (O_1779,N_24808,N_23682);
or UO_1780 (O_1780,N_23639,N_24528);
nor UO_1781 (O_1781,N_23370,N_23799);
and UO_1782 (O_1782,N_22665,N_23417);
nand UO_1783 (O_1783,N_23722,N_24226);
nor UO_1784 (O_1784,N_22837,N_24210);
or UO_1785 (O_1785,N_22666,N_24907);
and UO_1786 (O_1786,N_24489,N_23995);
nand UO_1787 (O_1787,N_24057,N_24397);
nor UO_1788 (O_1788,N_22871,N_24007);
and UO_1789 (O_1789,N_22538,N_24961);
xor UO_1790 (O_1790,N_23915,N_23366);
nor UO_1791 (O_1791,N_23311,N_22571);
xor UO_1792 (O_1792,N_23265,N_23517);
nor UO_1793 (O_1793,N_23159,N_24558);
xor UO_1794 (O_1794,N_24476,N_24829);
or UO_1795 (O_1795,N_22536,N_24872);
nand UO_1796 (O_1796,N_24835,N_24771);
nor UO_1797 (O_1797,N_22796,N_23397);
and UO_1798 (O_1798,N_23619,N_24690);
nand UO_1799 (O_1799,N_23650,N_24650);
and UO_1800 (O_1800,N_23094,N_23489);
and UO_1801 (O_1801,N_23588,N_23058);
or UO_1802 (O_1802,N_23544,N_24404);
or UO_1803 (O_1803,N_23817,N_23751);
nor UO_1804 (O_1804,N_23364,N_24342);
or UO_1805 (O_1805,N_23019,N_24841);
nand UO_1806 (O_1806,N_24279,N_24641);
and UO_1807 (O_1807,N_23148,N_24391);
nand UO_1808 (O_1808,N_24146,N_23705);
xor UO_1809 (O_1809,N_24663,N_23968);
or UO_1810 (O_1810,N_24256,N_22584);
nor UO_1811 (O_1811,N_24156,N_22608);
xor UO_1812 (O_1812,N_22670,N_23977);
or UO_1813 (O_1813,N_22970,N_23517);
nand UO_1814 (O_1814,N_23999,N_24594);
xnor UO_1815 (O_1815,N_24775,N_23447);
nand UO_1816 (O_1816,N_23165,N_23009);
and UO_1817 (O_1817,N_22681,N_23755);
nand UO_1818 (O_1818,N_23972,N_22702);
or UO_1819 (O_1819,N_24874,N_23516);
and UO_1820 (O_1820,N_23342,N_23992);
xnor UO_1821 (O_1821,N_23775,N_24020);
nand UO_1822 (O_1822,N_24264,N_22738);
nand UO_1823 (O_1823,N_24257,N_23401);
xnor UO_1824 (O_1824,N_23765,N_24919);
or UO_1825 (O_1825,N_24027,N_24402);
xnor UO_1826 (O_1826,N_22830,N_24657);
xnor UO_1827 (O_1827,N_22674,N_22640);
or UO_1828 (O_1828,N_22982,N_23073);
or UO_1829 (O_1829,N_24150,N_24398);
and UO_1830 (O_1830,N_23034,N_23883);
nor UO_1831 (O_1831,N_23213,N_24342);
or UO_1832 (O_1832,N_23183,N_24552);
nand UO_1833 (O_1833,N_23175,N_23128);
or UO_1834 (O_1834,N_23275,N_23607);
or UO_1835 (O_1835,N_23597,N_23696);
nor UO_1836 (O_1836,N_22683,N_22708);
xnor UO_1837 (O_1837,N_22611,N_24252);
and UO_1838 (O_1838,N_23555,N_22856);
and UO_1839 (O_1839,N_23090,N_23304);
nand UO_1840 (O_1840,N_22568,N_22597);
nand UO_1841 (O_1841,N_23474,N_22635);
xnor UO_1842 (O_1842,N_23306,N_24564);
or UO_1843 (O_1843,N_23670,N_23083);
xnor UO_1844 (O_1844,N_22905,N_24160);
nor UO_1845 (O_1845,N_22646,N_24535);
or UO_1846 (O_1846,N_22961,N_24919);
nand UO_1847 (O_1847,N_23172,N_22530);
nand UO_1848 (O_1848,N_23952,N_22744);
xor UO_1849 (O_1849,N_23664,N_22939);
nor UO_1850 (O_1850,N_23523,N_22720);
nand UO_1851 (O_1851,N_23163,N_24289);
xnor UO_1852 (O_1852,N_22840,N_23474);
nand UO_1853 (O_1853,N_22622,N_24923);
nor UO_1854 (O_1854,N_23099,N_24040);
xnor UO_1855 (O_1855,N_24184,N_23682);
and UO_1856 (O_1856,N_23566,N_22556);
nand UO_1857 (O_1857,N_22957,N_23462);
nand UO_1858 (O_1858,N_23228,N_24772);
xor UO_1859 (O_1859,N_24551,N_23214);
nor UO_1860 (O_1860,N_23437,N_23674);
nor UO_1861 (O_1861,N_24688,N_24180);
or UO_1862 (O_1862,N_23744,N_23443);
xnor UO_1863 (O_1863,N_24001,N_22627);
nand UO_1864 (O_1864,N_24892,N_24931);
and UO_1865 (O_1865,N_24379,N_22521);
and UO_1866 (O_1866,N_24477,N_24521);
or UO_1867 (O_1867,N_23416,N_24780);
nand UO_1868 (O_1868,N_24603,N_23531);
xnor UO_1869 (O_1869,N_23958,N_24002);
nand UO_1870 (O_1870,N_24635,N_24251);
and UO_1871 (O_1871,N_23949,N_24070);
xor UO_1872 (O_1872,N_23950,N_23580);
xor UO_1873 (O_1873,N_23425,N_24207);
nor UO_1874 (O_1874,N_24479,N_24870);
xnor UO_1875 (O_1875,N_24525,N_22743);
nand UO_1876 (O_1876,N_24556,N_23558);
and UO_1877 (O_1877,N_23054,N_24008);
xnor UO_1878 (O_1878,N_23202,N_22678);
nand UO_1879 (O_1879,N_24027,N_24294);
nor UO_1880 (O_1880,N_23895,N_23377);
nand UO_1881 (O_1881,N_24319,N_22536);
or UO_1882 (O_1882,N_22505,N_22672);
and UO_1883 (O_1883,N_22943,N_23641);
and UO_1884 (O_1884,N_23416,N_22893);
xnor UO_1885 (O_1885,N_23844,N_24588);
nor UO_1886 (O_1886,N_23666,N_23556);
nor UO_1887 (O_1887,N_23868,N_24992);
nor UO_1888 (O_1888,N_23860,N_23369);
and UO_1889 (O_1889,N_22721,N_24237);
and UO_1890 (O_1890,N_23767,N_23394);
or UO_1891 (O_1891,N_23101,N_22829);
xnor UO_1892 (O_1892,N_24461,N_24266);
nor UO_1893 (O_1893,N_24451,N_23197);
xnor UO_1894 (O_1894,N_23566,N_24358);
xnor UO_1895 (O_1895,N_23312,N_23420);
and UO_1896 (O_1896,N_22784,N_23370);
or UO_1897 (O_1897,N_22745,N_22778);
xnor UO_1898 (O_1898,N_23808,N_24691);
and UO_1899 (O_1899,N_24088,N_24119);
or UO_1900 (O_1900,N_24340,N_24238);
or UO_1901 (O_1901,N_22592,N_23082);
nand UO_1902 (O_1902,N_24629,N_22542);
or UO_1903 (O_1903,N_22759,N_24408);
xnor UO_1904 (O_1904,N_24539,N_22802);
and UO_1905 (O_1905,N_23777,N_22789);
nor UO_1906 (O_1906,N_23193,N_23550);
and UO_1907 (O_1907,N_23175,N_22984);
and UO_1908 (O_1908,N_23116,N_22563);
or UO_1909 (O_1909,N_22850,N_22944);
nand UO_1910 (O_1910,N_22690,N_22724);
nand UO_1911 (O_1911,N_23893,N_23396);
nor UO_1912 (O_1912,N_23484,N_24712);
nor UO_1913 (O_1913,N_22619,N_22773);
nor UO_1914 (O_1914,N_22806,N_23819);
and UO_1915 (O_1915,N_22961,N_23503);
nor UO_1916 (O_1916,N_23799,N_22894);
xor UO_1917 (O_1917,N_23827,N_24607);
nor UO_1918 (O_1918,N_24956,N_22754);
nand UO_1919 (O_1919,N_24329,N_23834);
xor UO_1920 (O_1920,N_22962,N_23041);
nor UO_1921 (O_1921,N_22541,N_23049);
nand UO_1922 (O_1922,N_22698,N_24472);
nand UO_1923 (O_1923,N_23975,N_24070);
xnor UO_1924 (O_1924,N_23551,N_23669);
nand UO_1925 (O_1925,N_24526,N_22637);
nor UO_1926 (O_1926,N_22619,N_24838);
nor UO_1927 (O_1927,N_24577,N_24251);
xor UO_1928 (O_1928,N_24549,N_24454);
xor UO_1929 (O_1929,N_24894,N_24165);
and UO_1930 (O_1930,N_22921,N_23619);
and UO_1931 (O_1931,N_24541,N_23514);
nand UO_1932 (O_1932,N_24211,N_24512);
nor UO_1933 (O_1933,N_23162,N_24745);
and UO_1934 (O_1934,N_23514,N_23139);
or UO_1935 (O_1935,N_24284,N_24111);
or UO_1936 (O_1936,N_23093,N_24929);
or UO_1937 (O_1937,N_24976,N_24475);
nand UO_1938 (O_1938,N_23348,N_22888);
or UO_1939 (O_1939,N_23857,N_24087);
xor UO_1940 (O_1940,N_23550,N_24484);
xnor UO_1941 (O_1941,N_24291,N_23832);
and UO_1942 (O_1942,N_22644,N_24870);
nor UO_1943 (O_1943,N_24983,N_23227);
nor UO_1944 (O_1944,N_24686,N_23207);
xor UO_1945 (O_1945,N_23043,N_24159);
nand UO_1946 (O_1946,N_24200,N_23780);
and UO_1947 (O_1947,N_22591,N_24405);
and UO_1948 (O_1948,N_24715,N_23367);
nand UO_1949 (O_1949,N_22804,N_24867);
xnor UO_1950 (O_1950,N_24887,N_24302);
and UO_1951 (O_1951,N_24757,N_22535);
or UO_1952 (O_1952,N_23476,N_24082);
or UO_1953 (O_1953,N_24051,N_24489);
nor UO_1954 (O_1954,N_24917,N_24641);
nand UO_1955 (O_1955,N_22859,N_24027);
and UO_1956 (O_1956,N_22879,N_24699);
nor UO_1957 (O_1957,N_23482,N_24642);
nor UO_1958 (O_1958,N_23944,N_22867);
or UO_1959 (O_1959,N_24087,N_24735);
xnor UO_1960 (O_1960,N_24217,N_23865);
xor UO_1961 (O_1961,N_24598,N_23290);
nand UO_1962 (O_1962,N_23690,N_22660);
xor UO_1963 (O_1963,N_24949,N_24407);
or UO_1964 (O_1964,N_24267,N_24611);
and UO_1965 (O_1965,N_23603,N_22852);
or UO_1966 (O_1966,N_24301,N_22778);
and UO_1967 (O_1967,N_23856,N_23945);
and UO_1968 (O_1968,N_23226,N_23236);
nor UO_1969 (O_1969,N_22987,N_24784);
or UO_1970 (O_1970,N_22553,N_24326);
xnor UO_1971 (O_1971,N_24070,N_22533);
or UO_1972 (O_1972,N_23115,N_22782);
nor UO_1973 (O_1973,N_23730,N_23056);
nor UO_1974 (O_1974,N_24302,N_23717);
xor UO_1975 (O_1975,N_22931,N_23400);
xor UO_1976 (O_1976,N_23583,N_24886);
nor UO_1977 (O_1977,N_23391,N_23094);
and UO_1978 (O_1978,N_23331,N_24358);
and UO_1979 (O_1979,N_23718,N_24731);
nand UO_1980 (O_1980,N_23217,N_23547);
and UO_1981 (O_1981,N_23899,N_24998);
nand UO_1982 (O_1982,N_23941,N_22771);
and UO_1983 (O_1983,N_22889,N_23968);
nor UO_1984 (O_1984,N_23252,N_22877);
or UO_1985 (O_1985,N_24504,N_24410);
nand UO_1986 (O_1986,N_24863,N_24916);
and UO_1987 (O_1987,N_24002,N_22732);
and UO_1988 (O_1988,N_22960,N_23054);
xor UO_1989 (O_1989,N_23286,N_23547);
and UO_1990 (O_1990,N_23877,N_22513);
and UO_1991 (O_1991,N_23043,N_23337);
nand UO_1992 (O_1992,N_24991,N_24608);
nand UO_1993 (O_1993,N_22670,N_24342);
or UO_1994 (O_1994,N_23184,N_22924);
or UO_1995 (O_1995,N_23082,N_23375);
nand UO_1996 (O_1996,N_22896,N_22710);
xnor UO_1997 (O_1997,N_22600,N_22995);
nor UO_1998 (O_1998,N_22937,N_23556);
or UO_1999 (O_1999,N_23390,N_23534);
and UO_2000 (O_2000,N_23936,N_23417);
nand UO_2001 (O_2001,N_22787,N_23711);
or UO_2002 (O_2002,N_24131,N_24125);
or UO_2003 (O_2003,N_22699,N_23227);
xor UO_2004 (O_2004,N_22642,N_24873);
or UO_2005 (O_2005,N_22784,N_24565);
nand UO_2006 (O_2006,N_23278,N_23851);
nand UO_2007 (O_2007,N_23765,N_22519);
and UO_2008 (O_2008,N_23610,N_22955);
xor UO_2009 (O_2009,N_24048,N_23076);
nand UO_2010 (O_2010,N_22891,N_24883);
nor UO_2011 (O_2011,N_24652,N_23168);
and UO_2012 (O_2012,N_24009,N_22633);
and UO_2013 (O_2013,N_22979,N_23992);
and UO_2014 (O_2014,N_23525,N_22885);
nor UO_2015 (O_2015,N_23817,N_23270);
or UO_2016 (O_2016,N_23391,N_22978);
or UO_2017 (O_2017,N_24393,N_22562);
xor UO_2018 (O_2018,N_22893,N_23825);
nand UO_2019 (O_2019,N_22688,N_24972);
nand UO_2020 (O_2020,N_23918,N_22725);
nand UO_2021 (O_2021,N_24440,N_23409);
nand UO_2022 (O_2022,N_23800,N_24967);
nor UO_2023 (O_2023,N_23562,N_23301);
or UO_2024 (O_2024,N_22742,N_23265);
xor UO_2025 (O_2025,N_24683,N_23713);
and UO_2026 (O_2026,N_24328,N_23430);
nand UO_2027 (O_2027,N_22979,N_22578);
and UO_2028 (O_2028,N_23163,N_24073);
nor UO_2029 (O_2029,N_24986,N_23299);
nor UO_2030 (O_2030,N_24466,N_23486);
or UO_2031 (O_2031,N_23925,N_24373);
or UO_2032 (O_2032,N_23387,N_23476);
xor UO_2033 (O_2033,N_22726,N_24919);
nor UO_2034 (O_2034,N_22698,N_23723);
xor UO_2035 (O_2035,N_23265,N_24779);
nor UO_2036 (O_2036,N_24072,N_23343);
nand UO_2037 (O_2037,N_24444,N_24819);
and UO_2038 (O_2038,N_24285,N_24338);
nor UO_2039 (O_2039,N_24655,N_22944);
and UO_2040 (O_2040,N_24810,N_24892);
nand UO_2041 (O_2041,N_22710,N_24415);
nor UO_2042 (O_2042,N_24724,N_24037);
and UO_2043 (O_2043,N_22841,N_24485);
and UO_2044 (O_2044,N_24542,N_22537);
nor UO_2045 (O_2045,N_24301,N_23294);
nand UO_2046 (O_2046,N_24847,N_24715);
and UO_2047 (O_2047,N_24790,N_23659);
xor UO_2048 (O_2048,N_22695,N_23275);
nor UO_2049 (O_2049,N_23414,N_23740);
nand UO_2050 (O_2050,N_23942,N_24270);
or UO_2051 (O_2051,N_23200,N_23749);
nor UO_2052 (O_2052,N_23732,N_22874);
xor UO_2053 (O_2053,N_23792,N_24496);
or UO_2054 (O_2054,N_24864,N_24238);
xnor UO_2055 (O_2055,N_24470,N_23996);
nand UO_2056 (O_2056,N_23273,N_22924);
or UO_2057 (O_2057,N_24035,N_22856);
xnor UO_2058 (O_2058,N_23424,N_24523);
nand UO_2059 (O_2059,N_24375,N_22848);
xnor UO_2060 (O_2060,N_24753,N_24279);
nor UO_2061 (O_2061,N_22668,N_23270);
nand UO_2062 (O_2062,N_24423,N_23201);
xor UO_2063 (O_2063,N_23808,N_24846);
and UO_2064 (O_2064,N_23553,N_23827);
nand UO_2065 (O_2065,N_23320,N_24728);
and UO_2066 (O_2066,N_22708,N_24267);
xnor UO_2067 (O_2067,N_24595,N_24532);
nand UO_2068 (O_2068,N_23715,N_23063);
nand UO_2069 (O_2069,N_24772,N_23206);
xnor UO_2070 (O_2070,N_24494,N_23121);
or UO_2071 (O_2071,N_22959,N_24651);
nor UO_2072 (O_2072,N_23253,N_23177);
nand UO_2073 (O_2073,N_23109,N_22548);
and UO_2074 (O_2074,N_22800,N_24919);
xor UO_2075 (O_2075,N_22830,N_23201);
or UO_2076 (O_2076,N_24999,N_23454);
or UO_2077 (O_2077,N_24265,N_24814);
xnor UO_2078 (O_2078,N_24173,N_24363);
or UO_2079 (O_2079,N_24376,N_24988);
nor UO_2080 (O_2080,N_24274,N_23141);
and UO_2081 (O_2081,N_22857,N_24515);
nand UO_2082 (O_2082,N_24726,N_24092);
nand UO_2083 (O_2083,N_23559,N_24083);
nor UO_2084 (O_2084,N_22836,N_23255);
and UO_2085 (O_2085,N_23658,N_24458);
and UO_2086 (O_2086,N_23855,N_23137);
nor UO_2087 (O_2087,N_23095,N_22925);
nand UO_2088 (O_2088,N_23504,N_23854);
nor UO_2089 (O_2089,N_22745,N_24358);
nor UO_2090 (O_2090,N_23260,N_22625);
nor UO_2091 (O_2091,N_23216,N_24669);
and UO_2092 (O_2092,N_23077,N_23460);
xnor UO_2093 (O_2093,N_24906,N_23307);
or UO_2094 (O_2094,N_22904,N_23774);
or UO_2095 (O_2095,N_23415,N_22635);
nor UO_2096 (O_2096,N_24769,N_23868);
or UO_2097 (O_2097,N_24012,N_24758);
or UO_2098 (O_2098,N_23483,N_22895);
xnor UO_2099 (O_2099,N_24698,N_23374);
nor UO_2100 (O_2100,N_24957,N_24390);
or UO_2101 (O_2101,N_23124,N_24131);
nor UO_2102 (O_2102,N_24493,N_22594);
xor UO_2103 (O_2103,N_23385,N_22664);
xnor UO_2104 (O_2104,N_24657,N_24164);
or UO_2105 (O_2105,N_24945,N_22832);
nor UO_2106 (O_2106,N_24817,N_23516);
nor UO_2107 (O_2107,N_23306,N_24313);
nor UO_2108 (O_2108,N_22538,N_23809);
nand UO_2109 (O_2109,N_24881,N_22955);
and UO_2110 (O_2110,N_23223,N_24315);
nand UO_2111 (O_2111,N_22599,N_23587);
nor UO_2112 (O_2112,N_22664,N_23216);
and UO_2113 (O_2113,N_24165,N_23071);
nand UO_2114 (O_2114,N_23134,N_22833);
nand UO_2115 (O_2115,N_23042,N_22914);
nor UO_2116 (O_2116,N_24726,N_22972);
nand UO_2117 (O_2117,N_24968,N_24644);
and UO_2118 (O_2118,N_22736,N_23713);
and UO_2119 (O_2119,N_22779,N_22804);
or UO_2120 (O_2120,N_23359,N_22593);
xnor UO_2121 (O_2121,N_24319,N_24359);
nand UO_2122 (O_2122,N_24885,N_24238);
and UO_2123 (O_2123,N_24432,N_22608);
nand UO_2124 (O_2124,N_23238,N_23923);
nor UO_2125 (O_2125,N_22596,N_23201);
nand UO_2126 (O_2126,N_24751,N_23117);
xor UO_2127 (O_2127,N_24504,N_23394);
and UO_2128 (O_2128,N_24010,N_24225);
xor UO_2129 (O_2129,N_24315,N_23966);
and UO_2130 (O_2130,N_22856,N_24668);
and UO_2131 (O_2131,N_24120,N_24526);
nor UO_2132 (O_2132,N_23302,N_23271);
or UO_2133 (O_2133,N_22948,N_23824);
and UO_2134 (O_2134,N_24802,N_24845);
nor UO_2135 (O_2135,N_22507,N_24586);
and UO_2136 (O_2136,N_23443,N_22964);
and UO_2137 (O_2137,N_24204,N_23777);
nor UO_2138 (O_2138,N_23001,N_23647);
and UO_2139 (O_2139,N_22825,N_23590);
and UO_2140 (O_2140,N_22531,N_24205);
xor UO_2141 (O_2141,N_24463,N_24866);
nor UO_2142 (O_2142,N_23149,N_23726);
nor UO_2143 (O_2143,N_23419,N_22750);
and UO_2144 (O_2144,N_24407,N_22598);
nand UO_2145 (O_2145,N_24265,N_24613);
xnor UO_2146 (O_2146,N_24835,N_23603);
nor UO_2147 (O_2147,N_24742,N_23101);
and UO_2148 (O_2148,N_24858,N_24705);
and UO_2149 (O_2149,N_22643,N_22745);
xor UO_2150 (O_2150,N_22919,N_24703);
or UO_2151 (O_2151,N_23679,N_24032);
nand UO_2152 (O_2152,N_23679,N_22904);
xnor UO_2153 (O_2153,N_23730,N_22676);
and UO_2154 (O_2154,N_22763,N_22586);
nand UO_2155 (O_2155,N_22659,N_24330);
xor UO_2156 (O_2156,N_22623,N_22982);
nand UO_2157 (O_2157,N_24980,N_23240);
xor UO_2158 (O_2158,N_23634,N_23105);
nor UO_2159 (O_2159,N_24830,N_23784);
nand UO_2160 (O_2160,N_23273,N_24330);
or UO_2161 (O_2161,N_24650,N_24652);
or UO_2162 (O_2162,N_24168,N_24567);
nand UO_2163 (O_2163,N_23911,N_23857);
or UO_2164 (O_2164,N_24918,N_23513);
xnor UO_2165 (O_2165,N_24265,N_23083);
nand UO_2166 (O_2166,N_24130,N_24227);
nor UO_2167 (O_2167,N_24604,N_24847);
nand UO_2168 (O_2168,N_24548,N_23563);
xor UO_2169 (O_2169,N_24991,N_24829);
and UO_2170 (O_2170,N_23370,N_24102);
or UO_2171 (O_2171,N_23293,N_23833);
xnor UO_2172 (O_2172,N_24550,N_23219);
xor UO_2173 (O_2173,N_23849,N_22962);
xor UO_2174 (O_2174,N_24253,N_22578);
nand UO_2175 (O_2175,N_23250,N_24584);
nor UO_2176 (O_2176,N_24223,N_24955);
nand UO_2177 (O_2177,N_24015,N_24452);
and UO_2178 (O_2178,N_22749,N_24612);
nor UO_2179 (O_2179,N_24615,N_22762);
xnor UO_2180 (O_2180,N_24289,N_24166);
nor UO_2181 (O_2181,N_22993,N_23386);
and UO_2182 (O_2182,N_23049,N_23811);
nor UO_2183 (O_2183,N_23828,N_24238);
and UO_2184 (O_2184,N_22654,N_22860);
nand UO_2185 (O_2185,N_23486,N_23020);
or UO_2186 (O_2186,N_23381,N_24743);
nor UO_2187 (O_2187,N_24750,N_23581);
xor UO_2188 (O_2188,N_23021,N_24901);
nor UO_2189 (O_2189,N_22989,N_23049);
xnor UO_2190 (O_2190,N_23936,N_22625);
nand UO_2191 (O_2191,N_23797,N_23945);
xor UO_2192 (O_2192,N_23114,N_23802);
or UO_2193 (O_2193,N_23647,N_22778);
xnor UO_2194 (O_2194,N_24966,N_24596);
nand UO_2195 (O_2195,N_24089,N_23977);
or UO_2196 (O_2196,N_22910,N_22602);
xnor UO_2197 (O_2197,N_23354,N_23248);
nand UO_2198 (O_2198,N_22751,N_22833);
nor UO_2199 (O_2199,N_23340,N_22980);
nor UO_2200 (O_2200,N_24375,N_24936);
and UO_2201 (O_2201,N_24087,N_23450);
nor UO_2202 (O_2202,N_23479,N_23253);
nand UO_2203 (O_2203,N_22584,N_23524);
nor UO_2204 (O_2204,N_22561,N_22688);
nor UO_2205 (O_2205,N_23859,N_23958);
and UO_2206 (O_2206,N_23069,N_24885);
xnor UO_2207 (O_2207,N_24541,N_22679);
or UO_2208 (O_2208,N_24625,N_24471);
nand UO_2209 (O_2209,N_23923,N_23973);
or UO_2210 (O_2210,N_23054,N_24591);
or UO_2211 (O_2211,N_24770,N_22714);
or UO_2212 (O_2212,N_23046,N_23457);
or UO_2213 (O_2213,N_22893,N_23166);
nand UO_2214 (O_2214,N_24684,N_23980);
xnor UO_2215 (O_2215,N_24892,N_23576);
xor UO_2216 (O_2216,N_23728,N_23363);
nor UO_2217 (O_2217,N_23292,N_24028);
xnor UO_2218 (O_2218,N_23839,N_22732);
nand UO_2219 (O_2219,N_23585,N_22731);
xnor UO_2220 (O_2220,N_23849,N_24938);
nor UO_2221 (O_2221,N_24910,N_22708);
xnor UO_2222 (O_2222,N_23939,N_24228);
or UO_2223 (O_2223,N_24160,N_23588);
xor UO_2224 (O_2224,N_23285,N_24529);
xnor UO_2225 (O_2225,N_24408,N_24745);
and UO_2226 (O_2226,N_24749,N_23030);
or UO_2227 (O_2227,N_23254,N_22933);
nor UO_2228 (O_2228,N_24896,N_24853);
nor UO_2229 (O_2229,N_23904,N_23760);
nand UO_2230 (O_2230,N_24144,N_22720);
or UO_2231 (O_2231,N_23411,N_23795);
nor UO_2232 (O_2232,N_24244,N_22744);
or UO_2233 (O_2233,N_24950,N_23908);
or UO_2234 (O_2234,N_24714,N_24457);
and UO_2235 (O_2235,N_23717,N_24289);
and UO_2236 (O_2236,N_24764,N_22519);
nand UO_2237 (O_2237,N_24786,N_23612);
and UO_2238 (O_2238,N_23459,N_24707);
nor UO_2239 (O_2239,N_24497,N_23575);
xor UO_2240 (O_2240,N_24023,N_23824);
or UO_2241 (O_2241,N_24634,N_23364);
nand UO_2242 (O_2242,N_24699,N_24275);
xnor UO_2243 (O_2243,N_23215,N_24507);
nand UO_2244 (O_2244,N_24964,N_23704);
and UO_2245 (O_2245,N_24979,N_23068);
nand UO_2246 (O_2246,N_24596,N_24260);
nand UO_2247 (O_2247,N_24524,N_24923);
nor UO_2248 (O_2248,N_22666,N_22603);
nand UO_2249 (O_2249,N_22777,N_24523);
xnor UO_2250 (O_2250,N_24916,N_24136);
xnor UO_2251 (O_2251,N_23491,N_24613);
and UO_2252 (O_2252,N_24313,N_23392);
nor UO_2253 (O_2253,N_24550,N_23342);
xor UO_2254 (O_2254,N_24581,N_24197);
nor UO_2255 (O_2255,N_24908,N_24647);
nand UO_2256 (O_2256,N_23223,N_24742);
and UO_2257 (O_2257,N_23748,N_23646);
nand UO_2258 (O_2258,N_23605,N_23241);
or UO_2259 (O_2259,N_24072,N_23798);
xnor UO_2260 (O_2260,N_22775,N_22904);
nand UO_2261 (O_2261,N_23776,N_22648);
nand UO_2262 (O_2262,N_24417,N_24992);
or UO_2263 (O_2263,N_24642,N_24289);
or UO_2264 (O_2264,N_24741,N_23601);
nor UO_2265 (O_2265,N_24195,N_24046);
xnor UO_2266 (O_2266,N_23295,N_22833);
or UO_2267 (O_2267,N_24869,N_24373);
xnor UO_2268 (O_2268,N_24823,N_22919);
and UO_2269 (O_2269,N_23862,N_23065);
or UO_2270 (O_2270,N_23628,N_24437);
nand UO_2271 (O_2271,N_23524,N_23299);
and UO_2272 (O_2272,N_24211,N_23919);
nand UO_2273 (O_2273,N_24787,N_24396);
and UO_2274 (O_2274,N_22633,N_24341);
nor UO_2275 (O_2275,N_23933,N_23215);
and UO_2276 (O_2276,N_24133,N_24904);
or UO_2277 (O_2277,N_23811,N_23833);
xnor UO_2278 (O_2278,N_23434,N_23405);
and UO_2279 (O_2279,N_24510,N_23292);
xor UO_2280 (O_2280,N_24883,N_24827);
or UO_2281 (O_2281,N_24744,N_23527);
nand UO_2282 (O_2282,N_24954,N_22662);
or UO_2283 (O_2283,N_23941,N_24720);
xor UO_2284 (O_2284,N_24135,N_23409);
nor UO_2285 (O_2285,N_24474,N_23284);
and UO_2286 (O_2286,N_23474,N_22904);
or UO_2287 (O_2287,N_23194,N_24241);
nand UO_2288 (O_2288,N_23509,N_23078);
nor UO_2289 (O_2289,N_24480,N_23499);
and UO_2290 (O_2290,N_23305,N_23921);
nor UO_2291 (O_2291,N_24991,N_24616);
xor UO_2292 (O_2292,N_24920,N_22682);
or UO_2293 (O_2293,N_23765,N_22809);
nand UO_2294 (O_2294,N_23002,N_23958);
or UO_2295 (O_2295,N_24433,N_24252);
and UO_2296 (O_2296,N_23127,N_23096);
nor UO_2297 (O_2297,N_23115,N_23301);
nor UO_2298 (O_2298,N_24668,N_22916);
and UO_2299 (O_2299,N_22572,N_24572);
and UO_2300 (O_2300,N_22903,N_24635);
nand UO_2301 (O_2301,N_24855,N_24007);
nor UO_2302 (O_2302,N_23990,N_22788);
nand UO_2303 (O_2303,N_24865,N_24924);
xnor UO_2304 (O_2304,N_24277,N_24482);
nor UO_2305 (O_2305,N_23204,N_24573);
or UO_2306 (O_2306,N_23626,N_24310);
or UO_2307 (O_2307,N_24930,N_24375);
or UO_2308 (O_2308,N_24517,N_24252);
xor UO_2309 (O_2309,N_24298,N_24653);
nand UO_2310 (O_2310,N_24614,N_24019);
or UO_2311 (O_2311,N_23220,N_23454);
xor UO_2312 (O_2312,N_23920,N_23126);
and UO_2313 (O_2313,N_24032,N_23873);
or UO_2314 (O_2314,N_24558,N_23049);
nand UO_2315 (O_2315,N_22629,N_23352);
or UO_2316 (O_2316,N_24514,N_24799);
xnor UO_2317 (O_2317,N_23390,N_24156);
xor UO_2318 (O_2318,N_24559,N_23375);
or UO_2319 (O_2319,N_22813,N_24001);
nor UO_2320 (O_2320,N_24369,N_22806);
or UO_2321 (O_2321,N_23285,N_22941);
xor UO_2322 (O_2322,N_22633,N_24524);
xnor UO_2323 (O_2323,N_24712,N_24406);
or UO_2324 (O_2324,N_23528,N_23162);
xor UO_2325 (O_2325,N_23045,N_24130);
nor UO_2326 (O_2326,N_23180,N_22514);
xnor UO_2327 (O_2327,N_22507,N_24021);
nor UO_2328 (O_2328,N_23309,N_23925);
and UO_2329 (O_2329,N_23944,N_24836);
nand UO_2330 (O_2330,N_23876,N_24099);
nor UO_2331 (O_2331,N_22743,N_24194);
xor UO_2332 (O_2332,N_22892,N_23326);
nor UO_2333 (O_2333,N_23936,N_23897);
nor UO_2334 (O_2334,N_24534,N_24843);
nand UO_2335 (O_2335,N_22951,N_23306);
or UO_2336 (O_2336,N_22907,N_24771);
xnor UO_2337 (O_2337,N_22545,N_23622);
nor UO_2338 (O_2338,N_24597,N_24675);
nor UO_2339 (O_2339,N_24078,N_22545);
or UO_2340 (O_2340,N_23643,N_24503);
xor UO_2341 (O_2341,N_23834,N_24065);
or UO_2342 (O_2342,N_22644,N_24263);
nor UO_2343 (O_2343,N_23683,N_23881);
nand UO_2344 (O_2344,N_23662,N_22944);
nand UO_2345 (O_2345,N_23262,N_22777);
nand UO_2346 (O_2346,N_22603,N_23048);
or UO_2347 (O_2347,N_24183,N_22850);
nand UO_2348 (O_2348,N_24499,N_24114);
nor UO_2349 (O_2349,N_23935,N_24093);
nand UO_2350 (O_2350,N_23638,N_24070);
nand UO_2351 (O_2351,N_24280,N_23084);
and UO_2352 (O_2352,N_23186,N_22755);
nor UO_2353 (O_2353,N_23737,N_23299);
and UO_2354 (O_2354,N_24443,N_24594);
nand UO_2355 (O_2355,N_24553,N_23712);
and UO_2356 (O_2356,N_24252,N_24565);
or UO_2357 (O_2357,N_24820,N_24391);
xor UO_2358 (O_2358,N_23628,N_22938);
nand UO_2359 (O_2359,N_24495,N_23914);
nand UO_2360 (O_2360,N_23949,N_22947);
xnor UO_2361 (O_2361,N_22655,N_23411);
xnor UO_2362 (O_2362,N_23394,N_22628);
nand UO_2363 (O_2363,N_22747,N_22774);
xnor UO_2364 (O_2364,N_23912,N_24145);
xor UO_2365 (O_2365,N_24429,N_23896);
xor UO_2366 (O_2366,N_24300,N_23424);
or UO_2367 (O_2367,N_23712,N_22655);
and UO_2368 (O_2368,N_24727,N_23116);
and UO_2369 (O_2369,N_23511,N_24282);
nand UO_2370 (O_2370,N_23775,N_24527);
xor UO_2371 (O_2371,N_24668,N_22688);
or UO_2372 (O_2372,N_24112,N_23088);
nor UO_2373 (O_2373,N_23144,N_24264);
xor UO_2374 (O_2374,N_23230,N_22751);
or UO_2375 (O_2375,N_24509,N_24708);
and UO_2376 (O_2376,N_24098,N_24338);
xor UO_2377 (O_2377,N_23637,N_23677);
or UO_2378 (O_2378,N_22668,N_22862);
or UO_2379 (O_2379,N_24033,N_24368);
and UO_2380 (O_2380,N_24267,N_23179);
and UO_2381 (O_2381,N_24317,N_23869);
xor UO_2382 (O_2382,N_23013,N_24496);
xnor UO_2383 (O_2383,N_23250,N_23996);
nand UO_2384 (O_2384,N_24318,N_24736);
nor UO_2385 (O_2385,N_23324,N_23951);
nand UO_2386 (O_2386,N_24359,N_23349);
xnor UO_2387 (O_2387,N_24088,N_23431);
nor UO_2388 (O_2388,N_22783,N_23436);
and UO_2389 (O_2389,N_23622,N_24106);
xor UO_2390 (O_2390,N_23821,N_23211);
xor UO_2391 (O_2391,N_22671,N_24291);
and UO_2392 (O_2392,N_24519,N_23164);
nor UO_2393 (O_2393,N_23073,N_23295);
nand UO_2394 (O_2394,N_22714,N_23321);
nor UO_2395 (O_2395,N_23662,N_24201);
nor UO_2396 (O_2396,N_23901,N_22807);
nand UO_2397 (O_2397,N_24666,N_23699);
nand UO_2398 (O_2398,N_23626,N_24107);
nand UO_2399 (O_2399,N_23577,N_24893);
xor UO_2400 (O_2400,N_24143,N_23283);
nand UO_2401 (O_2401,N_24106,N_24612);
xor UO_2402 (O_2402,N_24679,N_22978);
xnor UO_2403 (O_2403,N_24507,N_22932);
and UO_2404 (O_2404,N_22940,N_24612);
nor UO_2405 (O_2405,N_24453,N_24619);
and UO_2406 (O_2406,N_22503,N_24893);
xor UO_2407 (O_2407,N_24924,N_22855);
or UO_2408 (O_2408,N_23710,N_22669);
or UO_2409 (O_2409,N_22583,N_24662);
xnor UO_2410 (O_2410,N_23680,N_22589);
or UO_2411 (O_2411,N_23937,N_22585);
nor UO_2412 (O_2412,N_23619,N_24787);
nand UO_2413 (O_2413,N_24632,N_24398);
or UO_2414 (O_2414,N_23785,N_24559);
xnor UO_2415 (O_2415,N_24184,N_22519);
nor UO_2416 (O_2416,N_23504,N_22981);
or UO_2417 (O_2417,N_24574,N_24449);
or UO_2418 (O_2418,N_23742,N_23263);
or UO_2419 (O_2419,N_23696,N_22831);
nand UO_2420 (O_2420,N_24135,N_22930);
nand UO_2421 (O_2421,N_23557,N_24071);
or UO_2422 (O_2422,N_22976,N_24951);
or UO_2423 (O_2423,N_24372,N_23018);
or UO_2424 (O_2424,N_24655,N_22742);
or UO_2425 (O_2425,N_24054,N_24079);
or UO_2426 (O_2426,N_24301,N_22619);
and UO_2427 (O_2427,N_24766,N_24778);
nor UO_2428 (O_2428,N_24008,N_24805);
and UO_2429 (O_2429,N_23161,N_22894);
nand UO_2430 (O_2430,N_23896,N_22747);
xnor UO_2431 (O_2431,N_22629,N_23116);
or UO_2432 (O_2432,N_23482,N_23477);
xor UO_2433 (O_2433,N_24213,N_23939);
or UO_2434 (O_2434,N_23994,N_23078);
xor UO_2435 (O_2435,N_24005,N_24163);
or UO_2436 (O_2436,N_23713,N_24052);
nor UO_2437 (O_2437,N_22663,N_22783);
xor UO_2438 (O_2438,N_24090,N_23381);
or UO_2439 (O_2439,N_23462,N_24385);
nand UO_2440 (O_2440,N_24349,N_24671);
and UO_2441 (O_2441,N_23187,N_22666);
and UO_2442 (O_2442,N_24365,N_23405);
or UO_2443 (O_2443,N_23911,N_24940);
nand UO_2444 (O_2444,N_23441,N_23714);
or UO_2445 (O_2445,N_24360,N_23955);
nor UO_2446 (O_2446,N_22982,N_22932);
nand UO_2447 (O_2447,N_24450,N_22895);
xnor UO_2448 (O_2448,N_23887,N_24461);
nor UO_2449 (O_2449,N_23985,N_24595);
or UO_2450 (O_2450,N_23782,N_23641);
or UO_2451 (O_2451,N_23874,N_23935);
and UO_2452 (O_2452,N_23610,N_22665);
or UO_2453 (O_2453,N_23442,N_22979);
nor UO_2454 (O_2454,N_24148,N_23894);
xor UO_2455 (O_2455,N_24974,N_23422);
and UO_2456 (O_2456,N_23509,N_24931);
and UO_2457 (O_2457,N_23904,N_23145);
nand UO_2458 (O_2458,N_24326,N_24292);
xnor UO_2459 (O_2459,N_23568,N_23108);
and UO_2460 (O_2460,N_23038,N_23331);
xnor UO_2461 (O_2461,N_24195,N_23034);
or UO_2462 (O_2462,N_23177,N_23539);
and UO_2463 (O_2463,N_24315,N_23073);
xnor UO_2464 (O_2464,N_24161,N_23452);
xnor UO_2465 (O_2465,N_23305,N_22503);
or UO_2466 (O_2466,N_24916,N_24343);
and UO_2467 (O_2467,N_24305,N_24674);
nor UO_2468 (O_2468,N_24797,N_24510);
nand UO_2469 (O_2469,N_23454,N_24122);
and UO_2470 (O_2470,N_24091,N_23934);
xor UO_2471 (O_2471,N_23425,N_24798);
nand UO_2472 (O_2472,N_24823,N_24102);
and UO_2473 (O_2473,N_24232,N_24100);
or UO_2474 (O_2474,N_22979,N_22641);
nor UO_2475 (O_2475,N_22837,N_24578);
xor UO_2476 (O_2476,N_23154,N_22938);
nor UO_2477 (O_2477,N_23306,N_22621);
and UO_2478 (O_2478,N_24213,N_24209);
or UO_2479 (O_2479,N_24075,N_23250);
xor UO_2480 (O_2480,N_23012,N_23294);
and UO_2481 (O_2481,N_23450,N_23808);
and UO_2482 (O_2482,N_24726,N_24577);
xnor UO_2483 (O_2483,N_23666,N_22562);
or UO_2484 (O_2484,N_24663,N_24462);
and UO_2485 (O_2485,N_23541,N_23235);
and UO_2486 (O_2486,N_22745,N_24826);
nor UO_2487 (O_2487,N_24242,N_24218);
xnor UO_2488 (O_2488,N_24141,N_23867);
and UO_2489 (O_2489,N_24291,N_23811);
or UO_2490 (O_2490,N_24975,N_22503);
nand UO_2491 (O_2491,N_24234,N_23826);
and UO_2492 (O_2492,N_24023,N_24411);
nand UO_2493 (O_2493,N_22635,N_23252);
xor UO_2494 (O_2494,N_22661,N_23178);
nor UO_2495 (O_2495,N_23404,N_23398);
xor UO_2496 (O_2496,N_23310,N_24536);
nand UO_2497 (O_2497,N_23226,N_24444);
and UO_2498 (O_2498,N_24894,N_24487);
nand UO_2499 (O_2499,N_24873,N_24115);
nand UO_2500 (O_2500,N_23683,N_23524);
nor UO_2501 (O_2501,N_23528,N_24391);
or UO_2502 (O_2502,N_23734,N_24875);
or UO_2503 (O_2503,N_24437,N_24122);
or UO_2504 (O_2504,N_24439,N_24240);
xnor UO_2505 (O_2505,N_24799,N_23933);
and UO_2506 (O_2506,N_22560,N_24364);
nor UO_2507 (O_2507,N_23994,N_22640);
nor UO_2508 (O_2508,N_22691,N_23545);
nor UO_2509 (O_2509,N_23811,N_23676);
nand UO_2510 (O_2510,N_24370,N_24139);
xor UO_2511 (O_2511,N_22992,N_22609);
nor UO_2512 (O_2512,N_23579,N_23448);
nor UO_2513 (O_2513,N_24618,N_24648);
xor UO_2514 (O_2514,N_24393,N_22654);
and UO_2515 (O_2515,N_23510,N_23429);
or UO_2516 (O_2516,N_24059,N_22542);
xor UO_2517 (O_2517,N_23009,N_24895);
nor UO_2518 (O_2518,N_23861,N_22605);
nand UO_2519 (O_2519,N_23055,N_22705);
nand UO_2520 (O_2520,N_24041,N_23350);
and UO_2521 (O_2521,N_24012,N_23259);
xnor UO_2522 (O_2522,N_23489,N_24698);
nor UO_2523 (O_2523,N_22944,N_23322);
or UO_2524 (O_2524,N_24669,N_23211);
and UO_2525 (O_2525,N_23580,N_23025);
or UO_2526 (O_2526,N_24583,N_24123);
nor UO_2527 (O_2527,N_22998,N_22654);
nand UO_2528 (O_2528,N_23750,N_23335);
nand UO_2529 (O_2529,N_23855,N_23165);
nor UO_2530 (O_2530,N_24323,N_24234);
nor UO_2531 (O_2531,N_24271,N_23888);
and UO_2532 (O_2532,N_23502,N_24517);
xor UO_2533 (O_2533,N_23804,N_22823);
or UO_2534 (O_2534,N_22867,N_22600);
nor UO_2535 (O_2535,N_23929,N_22802);
or UO_2536 (O_2536,N_24380,N_24101);
nand UO_2537 (O_2537,N_24347,N_24258);
or UO_2538 (O_2538,N_24162,N_23381);
xnor UO_2539 (O_2539,N_24079,N_23167);
and UO_2540 (O_2540,N_24742,N_23130);
xor UO_2541 (O_2541,N_24581,N_23407);
xnor UO_2542 (O_2542,N_24003,N_22522);
nor UO_2543 (O_2543,N_24364,N_23366);
nor UO_2544 (O_2544,N_23395,N_24052);
nand UO_2545 (O_2545,N_24739,N_22826);
xor UO_2546 (O_2546,N_24549,N_23483);
nor UO_2547 (O_2547,N_24529,N_23902);
nand UO_2548 (O_2548,N_23298,N_23658);
xnor UO_2549 (O_2549,N_23499,N_23790);
or UO_2550 (O_2550,N_22711,N_24819);
nand UO_2551 (O_2551,N_23121,N_24583);
or UO_2552 (O_2552,N_24599,N_24906);
xor UO_2553 (O_2553,N_22698,N_23760);
and UO_2554 (O_2554,N_24922,N_24759);
xnor UO_2555 (O_2555,N_23625,N_23020);
nand UO_2556 (O_2556,N_23185,N_24733);
xor UO_2557 (O_2557,N_24050,N_24066);
nor UO_2558 (O_2558,N_23652,N_23233);
nor UO_2559 (O_2559,N_24102,N_22946);
nor UO_2560 (O_2560,N_24606,N_22789);
nand UO_2561 (O_2561,N_23706,N_23795);
nand UO_2562 (O_2562,N_24160,N_24359);
and UO_2563 (O_2563,N_23500,N_23354);
or UO_2564 (O_2564,N_24852,N_24893);
nor UO_2565 (O_2565,N_22694,N_23023);
or UO_2566 (O_2566,N_24043,N_23095);
nor UO_2567 (O_2567,N_24858,N_24339);
nand UO_2568 (O_2568,N_22680,N_22861);
nor UO_2569 (O_2569,N_23407,N_22845);
xor UO_2570 (O_2570,N_23248,N_24461);
and UO_2571 (O_2571,N_24455,N_24199);
and UO_2572 (O_2572,N_23534,N_24351);
xnor UO_2573 (O_2573,N_23246,N_22887);
xnor UO_2574 (O_2574,N_24399,N_22892);
nor UO_2575 (O_2575,N_24282,N_23070);
or UO_2576 (O_2576,N_24116,N_24486);
or UO_2577 (O_2577,N_24397,N_23080);
and UO_2578 (O_2578,N_23415,N_22972);
nor UO_2579 (O_2579,N_22757,N_23358);
nand UO_2580 (O_2580,N_24310,N_24387);
nand UO_2581 (O_2581,N_23676,N_23485);
nand UO_2582 (O_2582,N_24526,N_23137);
and UO_2583 (O_2583,N_22577,N_24070);
or UO_2584 (O_2584,N_24748,N_24869);
nand UO_2585 (O_2585,N_23636,N_24298);
xor UO_2586 (O_2586,N_23484,N_23259);
nor UO_2587 (O_2587,N_23233,N_22924);
xnor UO_2588 (O_2588,N_23629,N_23676);
and UO_2589 (O_2589,N_24025,N_24101);
or UO_2590 (O_2590,N_22640,N_24843);
and UO_2591 (O_2591,N_24055,N_23612);
nor UO_2592 (O_2592,N_22874,N_23304);
nand UO_2593 (O_2593,N_23956,N_22749);
and UO_2594 (O_2594,N_23225,N_23943);
xor UO_2595 (O_2595,N_23013,N_24685);
or UO_2596 (O_2596,N_24107,N_24383);
and UO_2597 (O_2597,N_24837,N_24058);
nand UO_2598 (O_2598,N_24258,N_23768);
nand UO_2599 (O_2599,N_23015,N_24190);
or UO_2600 (O_2600,N_23738,N_23648);
xnor UO_2601 (O_2601,N_23421,N_23175);
nor UO_2602 (O_2602,N_24857,N_24572);
nand UO_2603 (O_2603,N_22959,N_24179);
and UO_2604 (O_2604,N_24845,N_24608);
nand UO_2605 (O_2605,N_24390,N_22701);
nand UO_2606 (O_2606,N_24752,N_23501);
or UO_2607 (O_2607,N_24457,N_22929);
nand UO_2608 (O_2608,N_23800,N_24917);
or UO_2609 (O_2609,N_24145,N_23656);
and UO_2610 (O_2610,N_23903,N_24696);
or UO_2611 (O_2611,N_22774,N_22811);
nor UO_2612 (O_2612,N_24990,N_23992);
and UO_2613 (O_2613,N_22663,N_23987);
or UO_2614 (O_2614,N_22946,N_24674);
and UO_2615 (O_2615,N_22902,N_23212);
xnor UO_2616 (O_2616,N_24411,N_23539);
nand UO_2617 (O_2617,N_22750,N_23893);
nand UO_2618 (O_2618,N_23622,N_22523);
or UO_2619 (O_2619,N_24850,N_24903);
or UO_2620 (O_2620,N_22572,N_23237);
nand UO_2621 (O_2621,N_22932,N_24074);
or UO_2622 (O_2622,N_24463,N_23921);
or UO_2623 (O_2623,N_23536,N_24636);
nor UO_2624 (O_2624,N_24706,N_23888);
nor UO_2625 (O_2625,N_22818,N_22744);
nand UO_2626 (O_2626,N_23708,N_24363);
and UO_2627 (O_2627,N_23522,N_23073);
and UO_2628 (O_2628,N_23701,N_22965);
nand UO_2629 (O_2629,N_23670,N_24430);
and UO_2630 (O_2630,N_23952,N_23381);
and UO_2631 (O_2631,N_24988,N_24385);
and UO_2632 (O_2632,N_23318,N_23470);
xnor UO_2633 (O_2633,N_24156,N_22596);
or UO_2634 (O_2634,N_23080,N_24719);
and UO_2635 (O_2635,N_23907,N_24573);
and UO_2636 (O_2636,N_22553,N_24152);
and UO_2637 (O_2637,N_23579,N_22505);
or UO_2638 (O_2638,N_24722,N_24555);
xor UO_2639 (O_2639,N_23472,N_23985);
nand UO_2640 (O_2640,N_22814,N_23603);
or UO_2641 (O_2641,N_24355,N_23218);
and UO_2642 (O_2642,N_24685,N_24709);
nor UO_2643 (O_2643,N_22954,N_22866);
xnor UO_2644 (O_2644,N_24580,N_24666);
xnor UO_2645 (O_2645,N_23892,N_24912);
nand UO_2646 (O_2646,N_23735,N_23027);
nor UO_2647 (O_2647,N_23556,N_22788);
nand UO_2648 (O_2648,N_24564,N_22867);
and UO_2649 (O_2649,N_24501,N_22558);
nor UO_2650 (O_2650,N_23097,N_23138);
nand UO_2651 (O_2651,N_24370,N_24543);
and UO_2652 (O_2652,N_24411,N_23317);
or UO_2653 (O_2653,N_24572,N_24160);
nor UO_2654 (O_2654,N_24796,N_23851);
and UO_2655 (O_2655,N_23034,N_24156);
and UO_2656 (O_2656,N_23308,N_24054);
and UO_2657 (O_2657,N_23045,N_23875);
nor UO_2658 (O_2658,N_24288,N_24683);
or UO_2659 (O_2659,N_22535,N_24497);
nor UO_2660 (O_2660,N_24594,N_23264);
and UO_2661 (O_2661,N_23053,N_23295);
xnor UO_2662 (O_2662,N_24257,N_23726);
nor UO_2663 (O_2663,N_23855,N_23475);
nand UO_2664 (O_2664,N_22974,N_24440);
xor UO_2665 (O_2665,N_24313,N_24629);
nand UO_2666 (O_2666,N_23159,N_24622);
nand UO_2667 (O_2667,N_23784,N_23774);
xnor UO_2668 (O_2668,N_24941,N_23809);
xor UO_2669 (O_2669,N_23857,N_23333);
xor UO_2670 (O_2670,N_24950,N_23081);
or UO_2671 (O_2671,N_23688,N_23924);
xnor UO_2672 (O_2672,N_23890,N_24279);
nand UO_2673 (O_2673,N_23895,N_23519);
and UO_2674 (O_2674,N_24196,N_22913);
xnor UO_2675 (O_2675,N_24802,N_22560);
xor UO_2676 (O_2676,N_23205,N_23023);
nor UO_2677 (O_2677,N_24935,N_22903);
or UO_2678 (O_2678,N_24641,N_24256);
nand UO_2679 (O_2679,N_22763,N_24748);
and UO_2680 (O_2680,N_24243,N_23445);
or UO_2681 (O_2681,N_22992,N_24106);
xnor UO_2682 (O_2682,N_23151,N_22730);
or UO_2683 (O_2683,N_22516,N_23775);
and UO_2684 (O_2684,N_23843,N_23918);
or UO_2685 (O_2685,N_23732,N_22980);
and UO_2686 (O_2686,N_22802,N_24733);
nand UO_2687 (O_2687,N_24013,N_24002);
or UO_2688 (O_2688,N_23951,N_24592);
and UO_2689 (O_2689,N_22816,N_23607);
xnor UO_2690 (O_2690,N_22943,N_22807);
nand UO_2691 (O_2691,N_24652,N_24270);
nor UO_2692 (O_2692,N_24865,N_23436);
nand UO_2693 (O_2693,N_23325,N_24776);
nand UO_2694 (O_2694,N_22975,N_23126);
xor UO_2695 (O_2695,N_22653,N_23352);
nand UO_2696 (O_2696,N_23223,N_22808);
or UO_2697 (O_2697,N_24714,N_24731);
nand UO_2698 (O_2698,N_23374,N_23742);
nand UO_2699 (O_2699,N_24618,N_23504);
nor UO_2700 (O_2700,N_22742,N_24250);
xor UO_2701 (O_2701,N_23386,N_24705);
xnor UO_2702 (O_2702,N_23551,N_23685);
and UO_2703 (O_2703,N_23200,N_22620);
and UO_2704 (O_2704,N_24977,N_22595);
and UO_2705 (O_2705,N_24769,N_23167);
nand UO_2706 (O_2706,N_24556,N_23137);
or UO_2707 (O_2707,N_24417,N_24641);
nor UO_2708 (O_2708,N_24092,N_23205);
nor UO_2709 (O_2709,N_24986,N_23238);
or UO_2710 (O_2710,N_24829,N_23089);
nand UO_2711 (O_2711,N_23934,N_24510);
xnor UO_2712 (O_2712,N_24705,N_22927);
nor UO_2713 (O_2713,N_23163,N_22969);
nor UO_2714 (O_2714,N_23973,N_23208);
and UO_2715 (O_2715,N_22851,N_24380);
nand UO_2716 (O_2716,N_23655,N_24668);
and UO_2717 (O_2717,N_23914,N_24560);
nand UO_2718 (O_2718,N_23394,N_24511);
or UO_2719 (O_2719,N_23186,N_22883);
xnor UO_2720 (O_2720,N_23060,N_24411);
and UO_2721 (O_2721,N_23569,N_24853);
nand UO_2722 (O_2722,N_23261,N_22974);
and UO_2723 (O_2723,N_23697,N_23549);
xor UO_2724 (O_2724,N_23520,N_24624);
or UO_2725 (O_2725,N_23114,N_23121);
or UO_2726 (O_2726,N_22506,N_24672);
xnor UO_2727 (O_2727,N_23403,N_23929);
nor UO_2728 (O_2728,N_23075,N_22800);
and UO_2729 (O_2729,N_23817,N_23414);
xnor UO_2730 (O_2730,N_23473,N_24148);
xnor UO_2731 (O_2731,N_22817,N_24802);
nor UO_2732 (O_2732,N_24556,N_23699);
nor UO_2733 (O_2733,N_23604,N_23965);
or UO_2734 (O_2734,N_24232,N_23470);
and UO_2735 (O_2735,N_23231,N_22664);
nor UO_2736 (O_2736,N_24205,N_22870);
nand UO_2737 (O_2737,N_23021,N_24097);
xor UO_2738 (O_2738,N_24491,N_23099);
or UO_2739 (O_2739,N_24724,N_24532);
nand UO_2740 (O_2740,N_24870,N_23466);
nor UO_2741 (O_2741,N_23536,N_24263);
or UO_2742 (O_2742,N_22688,N_22630);
and UO_2743 (O_2743,N_23056,N_23695);
xor UO_2744 (O_2744,N_24566,N_23813);
or UO_2745 (O_2745,N_23158,N_24996);
nor UO_2746 (O_2746,N_23231,N_24121);
and UO_2747 (O_2747,N_24604,N_23669);
and UO_2748 (O_2748,N_22667,N_23718);
or UO_2749 (O_2749,N_24125,N_23338);
nand UO_2750 (O_2750,N_23692,N_22634);
nand UO_2751 (O_2751,N_24922,N_23112);
nor UO_2752 (O_2752,N_24296,N_22839);
nor UO_2753 (O_2753,N_23200,N_23063);
xnor UO_2754 (O_2754,N_23788,N_24161);
or UO_2755 (O_2755,N_24842,N_24050);
xnor UO_2756 (O_2756,N_23757,N_24440);
nor UO_2757 (O_2757,N_24444,N_23092);
xor UO_2758 (O_2758,N_24496,N_23324);
nor UO_2759 (O_2759,N_23049,N_23335);
nor UO_2760 (O_2760,N_23267,N_23891);
xnor UO_2761 (O_2761,N_23833,N_24583);
or UO_2762 (O_2762,N_23980,N_22733);
nor UO_2763 (O_2763,N_23088,N_22570);
or UO_2764 (O_2764,N_24535,N_24524);
nor UO_2765 (O_2765,N_24652,N_22661);
or UO_2766 (O_2766,N_24913,N_24605);
and UO_2767 (O_2767,N_24941,N_23149);
or UO_2768 (O_2768,N_23197,N_23842);
nand UO_2769 (O_2769,N_24071,N_24271);
and UO_2770 (O_2770,N_23632,N_22601);
or UO_2771 (O_2771,N_24453,N_24079);
xnor UO_2772 (O_2772,N_24938,N_22708);
xnor UO_2773 (O_2773,N_24956,N_23433);
xor UO_2774 (O_2774,N_23926,N_22752);
nor UO_2775 (O_2775,N_22866,N_23245);
nor UO_2776 (O_2776,N_22766,N_22924);
nor UO_2777 (O_2777,N_23320,N_24200);
or UO_2778 (O_2778,N_22751,N_22876);
nor UO_2779 (O_2779,N_22762,N_24875);
and UO_2780 (O_2780,N_24330,N_23803);
and UO_2781 (O_2781,N_23851,N_24434);
xnor UO_2782 (O_2782,N_24699,N_24994);
nand UO_2783 (O_2783,N_23942,N_23974);
nor UO_2784 (O_2784,N_23611,N_24589);
or UO_2785 (O_2785,N_24831,N_24453);
xor UO_2786 (O_2786,N_24508,N_24950);
xor UO_2787 (O_2787,N_23512,N_22844);
or UO_2788 (O_2788,N_23480,N_23229);
nand UO_2789 (O_2789,N_24225,N_24002);
nor UO_2790 (O_2790,N_23953,N_24049);
nand UO_2791 (O_2791,N_22660,N_24629);
nand UO_2792 (O_2792,N_23826,N_24589);
nor UO_2793 (O_2793,N_24853,N_23341);
nor UO_2794 (O_2794,N_24137,N_24202);
or UO_2795 (O_2795,N_23864,N_23180);
xnor UO_2796 (O_2796,N_23884,N_22712);
nand UO_2797 (O_2797,N_23913,N_22576);
nand UO_2798 (O_2798,N_24776,N_23026);
nand UO_2799 (O_2799,N_23304,N_23638);
or UO_2800 (O_2800,N_24501,N_24428);
nor UO_2801 (O_2801,N_22990,N_24061);
nand UO_2802 (O_2802,N_24485,N_24780);
nand UO_2803 (O_2803,N_22539,N_23002);
and UO_2804 (O_2804,N_24360,N_23638);
nor UO_2805 (O_2805,N_23933,N_24166);
or UO_2806 (O_2806,N_24716,N_24884);
and UO_2807 (O_2807,N_22962,N_22605);
xor UO_2808 (O_2808,N_24520,N_24218);
nor UO_2809 (O_2809,N_23604,N_23823);
xnor UO_2810 (O_2810,N_23830,N_24639);
xnor UO_2811 (O_2811,N_23344,N_23915);
nand UO_2812 (O_2812,N_22532,N_23102);
and UO_2813 (O_2813,N_23947,N_23687);
nor UO_2814 (O_2814,N_23433,N_23519);
and UO_2815 (O_2815,N_23536,N_22839);
nor UO_2816 (O_2816,N_23061,N_22743);
and UO_2817 (O_2817,N_22939,N_24570);
nand UO_2818 (O_2818,N_22941,N_22751);
xor UO_2819 (O_2819,N_22820,N_24190);
nor UO_2820 (O_2820,N_22772,N_22832);
and UO_2821 (O_2821,N_23816,N_23416);
nor UO_2822 (O_2822,N_22836,N_23940);
or UO_2823 (O_2823,N_23175,N_22862);
xor UO_2824 (O_2824,N_24028,N_22736);
xor UO_2825 (O_2825,N_23101,N_23143);
nand UO_2826 (O_2826,N_23282,N_23609);
or UO_2827 (O_2827,N_24262,N_23609);
or UO_2828 (O_2828,N_23921,N_24597);
and UO_2829 (O_2829,N_23110,N_23780);
xor UO_2830 (O_2830,N_23101,N_23624);
or UO_2831 (O_2831,N_23218,N_23842);
and UO_2832 (O_2832,N_24321,N_24718);
nand UO_2833 (O_2833,N_24448,N_24105);
nand UO_2834 (O_2834,N_24998,N_23504);
nand UO_2835 (O_2835,N_24898,N_22558);
nand UO_2836 (O_2836,N_23580,N_24519);
nand UO_2837 (O_2837,N_24908,N_23352);
nor UO_2838 (O_2838,N_24208,N_22727);
and UO_2839 (O_2839,N_23771,N_22617);
nand UO_2840 (O_2840,N_22722,N_24845);
and UO_2841 (O_2841,N_24304,N_23607);
or UO_2842 (O_2842,N_24606,N_23850);
nor UO_2843 (O_2843,N_24894,N_23431);
and UO_2844 (O_2844,N_24004,N_24605);
nor UO_2845 (O_2845,N_23298,N_24277);
nor UO_2846 (O_2846,N_24342,N_24359);
nand UO_2847 (O_2847,N_23052,N_23168);
nand UO_2848 (O_2848,N_23122,N_23378);
nor UO_2849 (O_2849,N_24206,N_23036);
xor UO_2850 (O_2850,N_22871,N_22841);
and UO_2851 (O_2851,N_23575,N_22707);
xor UO_2852 (O_2852,N_23361,N_24336);
and UO_2853 (O_2853,N_24679,N_23150);
nand UO_2854 (O_2854,N_23351,N_24503);
and UO_2855 (O_2855,N_24349,N_24448);
xnor UO_2856 (O_2856,N_24431,N_24425);
or UO_2857 (O_2857,N_24823,N_24213);
xor UO_2858 (O_2858,N_23976,N_22641);
xnor UO_2859 (O_2859,N_23406,N_24088);
or UO_2860 (O_2860,N_24957,N_22975);
xor UO_2861 (O_2861,N_22934,N_23738);
nand UO_2862 (O_2862,N_24820,N_24810);
nor UO_2863 (O_2863,N_24287,N_22745);
and UO_2864 (O_2864,N_23907,N_23759);
nor UO_2865 (O_2865,N_24665,N_24191);
xnor UO_2866 (O_2866,N_24670,N_24252);
and UO_2867 (O_2867,N_24209,N_23601);
or UO_2868 (O_2868,N_22881,N_24017);
nor UO_2869 (O_2869,N_24650,N_22718);
or UO_2870 (O_2870,N_23531,N_24715);
nor UO_2871 (O_2871,N_23095,N_22699);
nand UO_2872 (O_2872,N_24969,N_24932);
nor UO_2873 (O_2873,N_23073,N_23728);
and UO_2874 (O_2874,N_22618,N_23983);
or UO_2875 (O_2875,N_24453,N_24122);
or UO_2876 (O_2876,N_24347,N_24977);
or UO_2877 (O_2877,N_24284,N_24434);
nor UO_2878 (O_2878,N_24259,N_23208);
or UO_2879 (O_2879,N_23951,N_23430);
and UO_2880 (O_2880,N_24459,N_23892);
and UO_2881 (O_2881,N_24841,N_23176);
or UO_2882 (O_2882,N_23588,N_24666);
or UO_2883 (O_2883,N_24948,N_24857);
nor UO_2884 (O_2884,N_24395,N_23765);
nand UO_2885 (O_2885,N_23365,N_22996);
nand UO_2886 (O_2886,N_24343,N_23427);
xnor UO_2887 (O_2887,N_24875,N_24532);
and UO_2888 (O_2888,N_23521,N_23502);
nor UO_2889 (O_2889,N_24462,N_23675);
and UO_2890 (O_2890,N_23800,N_24990);
nand UO_2891 (O_2891,N_22556,N_22574);
and UO_2892 (O_2892,N_23599,N_24190);
or UO_2893 (O_2893,N_24254,N_23708);
and UO_2894 (O_2894,N_23691,N_23122);
nor UO_2895 (O_2895,N_23690,N_24993);
and UO_2896 (O_2896,N_23932,N_23940);
and UO_2897 (O_2897,N_22810,N_24347);
nand UO_2898 (O_2898,N_22896,N_23644);
or UO_2899 (O_2899,N_24370,N_24885);
nand UO_2900 (O_2900,N_23558,N_22647);
nand UO_2901 (O_2901,N_23158,N_24641);
or UO_2902 (O_2902,N_22662,N_24156);
and UO_2903 (O_2903,N_22924,N_22864);
or UO_2904 (O_2904,N_23087,N_24860);
xor UO_2905 (O_2905,N_23902,N_24060);
nor UO_2906 (O_2906,N_24174,N_23248);
or UO_2907 (O_2907,N_22660,N_22946);
and UO_2908 (O_2908,N_24352,N_24323);
xor UO_2909 (O_2909,N_24827,N_24520);
xnor UO_2910 (O_2910,N_23498,N_24369);
nor UO_2911 (O_2911,N_22576,N_24657);
and UO_2912 (O_2912,N_24992,N_24383);
or UO_2913 (O_2913,N_23059,N_24890);
xnor UO_2914 (O_2914,N_23691,N_22642);
nor UO_2915 (O_2915,N_24611,N_24574);
or UO_2916 (O_2916,N_22788,N_23586);
and UO_2917 (O_2917,N_24891,N_22928);
nor UO_2918 (O_2918,N_22866,N_22651);
and UO_2919 (O_2919,N_24224,N_22820);
and UO_2920 (O_2920,N_22997,N_22995);
and UO_2921 (O_2921,N_24784,N_24562);
and UO_2922 (O_2922,N_24123,N_23609);
nand UO_2923 (O_2923,N_23276,N_23547);
nand UO_2924 (O_2924,N_23332,N_24797);
or UO_2925 (O_2925,N_24664,N_24963);
or UO_2926 (O_2926,N_23285,N_22956);
xor UO_2927 (O_2927,N_23126,N_23677);
nor UO_2928 (O_2928,N_24322,N_22603);
and UO_2929 (O_2929,N_23982,N_23570);
nor UO_2930 (O_2930,N_22533,N_22895);
and UO_2931 (O_2931,N_24798,N_24820);
nand UO_2932 (O_2932,N_23479,N_23607);
nor UO_2933 (O_2933,N_23928,N_22969);
nor UO_2934 (O_2934,N_23426,N_23934);
xnor UO_2935 (O_2935,N_23745,N_23507);
xnor UO_2936 (O_2936,N_24202,N_24004);
nand UO_2937 (O_2937,N_24658,N_24899);
and UO_2938 (O_2938,N_24125,N_24172);
or UO_2939 (O_2939,N_24133,N_23880);
nor UO_2940 (O_2940,N_23294,N_24094);
xnor UO_2941 (O_2941,N_23500,N_24163);
nor UO_2942 (O_2942,N_22666,N_24667);
and UO_2943 (O_2943,N_24594,N_22854);
or UO_2944 (O_2944,N_22914,N_24413);
and UO_2945 (O_2945,N_22649,N_24297);
nor UO_2946 (O_2946,N_23571,N_24826);
or UO_2947 (O_2947,N_24765,N_23767);
xor UO_2948 (O_2948,N_23229,N_24599);
or UO_2949 (O_2949,N_23951,N_23841);
xnor UO_2950 (O_2950,N_23362,N_24333);
and UO_2951 (O_2951,N_22595,N_23024);
nand UO_2952 (O_2952,N_23896,N_22808);
nand UO_2953 (O_2953,N_22857,N_23530);
nor UO_2954 (O_2954,N_23738,N_22999);
or UO_2955 (O_2955,N_23131,N_23414);
or UO_2956 (O_2956,N_22749,N_24018);
or UO_2957 (O_2957,N_24667,N_22722);
nor UO_2958 (O_2958,N_22886,N_23823);
or UO_2959 (O_2959,N_23535,N_24655);
nor UO_2960 (O_2960,N_23073,N_22844);
and UO_2961 (O_2961,N_24992,N_24532);
xnor UO_2962 (O_2962,N_22578,N_24537);
or UO_2963 (O_2963,N_22694,N_23462);
and UO_2964 (O_2964,N_23210,N_23892);
or UO_2965 (O_2965,N_23942,N_24939);
and UO_2966 (O_2966,N_22785,N_23760);
nand UO_2967 (O_2967,N_22558,N_23310);
nand UO_2968 (O_2968,N_22663,N_24590);
nand UO_2969 (O_2969,N_22985,N_23523);
or UO_2970 (O_2970,N_22651,N_24611);
nand UO_2971 (O_2971,N_22656,N_24891);
nor UO_2972 (O_2972,N_23759,N_23520);
and UO_2973 (O_2973,N_24191,N_24141);
xor UO_2974 (O_2974,N_24272,N_24402);
or UO_2975 (O_2975,N_24716,N_22906);
nand UO_2976 (O_2976,N_23647,N_24047);
nand UO_2977 (O_2977,N_24817,N_23442);
nor UO_2978 (O_2978,N_24864,N_24812);
or UO_2979 (O_2979,N_22608,N_23524);
and UO_2980 (O_2980,N_24527,N_22600);
xnor UO_2981 (O_2981,N_23125,N_22832);
nor UO_2982 (O_2982,N_24063,N_24250);
nor UO_2983 (O_2983,N_24844,N_24436);
and UO_2984 (O_2984,N_22722,N_23310);
xnor UO_2985 (O_2985,N_24814,N_23219);
nand UO_2986 (O_2986,N_24150,N_24211);
xor UO_2987 (O_2987,N_22553,N_22875);
nor UO_2988 (O_2988,N_23947,N_24806);
or UO_2989 (O_2989,N_24367,N_22680);
and UO_2990 (O_2990,N_22855,N_22836);
nor UO_2991 (O_2991,N_23310,N_24030);
nand UO_2992 (O_2992,N_23409,N_22670);
nor UO_2993 (O_2993,N_22998,N_23190);
or UO_2994 (O_2994,N_23589,N_24088);
nand UO_2995 (O_2995,N_23615,N_24561);
and UO_2996 (O_2996,N_22678,N_24363);
xor UO_2997 (O_2997,N_23001,N_23575);
nor UO_2998 (O_2998,N_22870,N_23196);
nor UO_2999 (O_2999,N_23747,N_24229);
endmodule