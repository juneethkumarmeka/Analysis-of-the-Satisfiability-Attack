module basic_3000_30000_3500_50_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_1353,In_404);
or U1 (N_1,In_172,In_1031);
or U2 (N_2,In_219,In_2981);
nand U3 (N_3,In_323,In_2656);
nor U4 (N_4,In_2887,In_1938);
or U5 (N_5,In_448,In_2795);
nor U6 (N_6,In_2180,In_2149);
nand U7 (N_7,In_594,In_1725);
xnor U8 (N_8,In_773,In_805);
nand U9 (N_9,In_1127,In_2097);
or U10 (N_10,In_1825,In_442);
nand U11 (N_11,In_359,In_2895);
or U12 (N_12,In_2218,In_80);
and U13 (N_13,In_100,In_622);
and U14 (N_14,In_1060,In_971);
xor U15 (N_15,In_1873,In_322);
nor U16 (N_16,In_2142,In_2379);
xnor U17 (N_17,In_2181,In_2444);
xnor U18 (N_18,In_24,In_2605);
xnor U19 (N_19,In_874,In_904);
nor U20 (N_20,In_538,In_454);
xnor U21 (N_21,In_2223,In_2320);
xnor U22 (N_22,In_736,In_1231);
and U23 (N_23,In_1993,In_38);
xor U24 (N_24,In_2517,In_1775);
nand U25 (N_25,In_2297,In_2588);
nand U26 (N_26,In_869,In_483);
and U27 (N_27,In_124,In_2041);
or U28 (N_28,In_1126,In_276);
nand U29 (N_29,In_2075,In_1878);
xor U30 (N_30,In_1483,In_2693);
and U31 (N_31,In_539,In_777);
or U32 (N_32,In_400,In_1448);
or U33 (N_33,In_2827,In_149);
nor U34 (N_34,In_1558,In_102);
xnor U35 (N_35,In_1970,In_2234);
and U36 (N_36,In_2987,In_785);
or U37 (N_37,In_1250,In_192);
nand U38 (N_38,In_2138,In_1947);
nand U39 (N_39,In_1169,In_2799);
nand U40 (N_40,In_356,In_593);
and U41 (N_41,In_2586,In_2720);
or U42 (N_42,In_30,In_909);
nor U43 (N_43,In_851,In_2617);
or U44 (N_44,In_1113,In_677);
xnor U45 (N_45,In_1147,In_2269);
or U46 (N_46,In_1685,In_486);
and U47 (N_47,In_1515,In_1210);
nor U48 (N_48,In_2897,In_667);
or U49 (N_49,In_1859,In_2811);
nand U50 (N_50,In_2859,In_1764);
and U51 (N_51,In_2106,In_74);
nand U52 (N_52,In_2336,In_2900);
or U53 (N_53,In_1111,In_673);
xor U54 (N_54,In_2791,In_1084);
nand U55 (N_55,In_843,In_1156);
nand U56 (N_56,In_1344,In_1914);
or U57 (N_57,In_2738,In_2330);
or U58 (N_58,In_2716,In_2454);
and U59 (N_59,In_2189,In_1062);
or U60 (N_60,In_902,In_547);
or U61 (N_61,In_202,In_2660);
and U62 (N_62,In_576,In_1753);
or U63 (N_63,In_792,In_1415);
xnor U64 (N_64,In_2115,In_227);
and U65 (N_65,In_760,In_1423);
and U66 (N_66,In_580,In_2564);
nand U67 (N_67,In_1861,In_1308);
and U68 (N_68,In_599,In_1939);
nand U69 (N_69,In_1659,In_1220);
nor U70 (N_70,In_2099,In_469);
or U71 (N_71,In_1891,In_1583);
xor U72 (N_72,In_974,In_372);
nand U73 (N_73,In_1851,In_1459);
nand U74 (N_74,In_1841,In_2945);
xnor U75 (N_75,In_1066,In_2748);
nand U76 (N_76,In_1472,In_885);
nor U77 (N_77,In_2882,In_1000);
nand U78 (N_78,In_746,In_1789);
and U79 (N_79,In_2028,In_21);
xnor U80 (N_80,In_2346,In_724);
nand U81 (N_81,In_1979,In_595);
and U82 (N_82,In_2674,In_2764);
nor U83 (N_83,In_1586,In_2035);
or U84 (N_84,In_685,In_1886);
xnor U85 (N_85,In_684,In_98);
and U86 (N_86,In_2808,In_551);
and U87 (N_87,In_2440,In_549);
nor U88 (N_88,In_1040,In_765);
nand U89 (N_89,In_2348,In_1893);
xor U90 (N_90,In_883,In_2102);
and U91 (N_91,In_528,In_387);
nor U92 (N_92,In_875,In_888);
and U93 (N_93,In_2151,In_2428);
nand U94 (N_94,In_1114,In_7);
nand U95 (N_95,In_1826,In_1957);
xor U96 (N_96,In_68,In_317);
nor U97 (N_97,In_1416,In_1296);
nor U98 (N_98,In_589,In_1517);
xor U99 (N_99,In_2015,In_2876);
xnor U100 (N_100,In_312,In_1740);
nor U101 (N_101,In_775,In_476);
nor U102 (N_102,In_876,In_2094);
or U103 (N_103,In_2146,In_2689);
nand U104 (N_104,In_1604,In_334);
and U105 (N_105,In_2017,In_1014);
or U106 (N_106,In_250,In_2541);
nor U107 (N_107,In_2825,In_1866);
nor U108 (N_108,In_1161,In_54);
xnor U109 (N_109,In_852,In_2435);
nand U110 (N_110,In_121,In_893);
nand U111 (N_111,In_348,In_1976);
nor U112 (N_112,In_982,In_1363);
xnor U113 (N_113,In_2512,In_2641);
nor U114 (N_114,In_1240,In_1817);
xnor U115 (N_115,In_627,In_847);
nand U116 (N_116,In_2554,In_2830);
nand U117 (N_117,In_2123,In_1034);
or U118 (N_118,In_737,In_744);
or U119 (N_119,In_2177,In_1253);
nand U120 (N_120,In_1802,In_510);
nor U121 (N_121,In_1499,In_2083);
xnor U122 (N_122,In_373,In_2531);
and U123 (N_123,In_1830,In_2804);
nor U124 (N_124,In_1036,In_862);
and U125 (N_125,In_1911,In_641);
nor U126 (N_126,In_505,In_2315);
nor U127 (N_127,In_1862,In_22);
or U128 (N_128,In_2031,In_2621);
xnor U129 (N_129,In_329,In_2359);
nand U130 (N_130,In_2418,In_1904);
or U131 (N_131,In_2152,In_650);
xnor U132 (N_132,In_2194,In_2487);
or U133 (N_133,In_567,In_1853);
nand U134 (N_134,In_1567,In_2137);
nor U135 (N_135,In_1394,In_1838);
xor U136 (N_136,In_1987,In_1063);
nor U137 (N_137,In_2979,In_1058);
or U138 (N_138,In_2204,In_1310);
or U139 (N_139,In_1117,In_2148);
xor U140 (N_140,In_1566,In_808);
xnor U141 (N_141,In_1053,In_2150);
nor U142 (N_142,In_50,In_2597);
xor U143 (N_143,In_273,In_2378);
and U144 (N_144,In_42,In_71);
nand U145 (N_145,In_919,In_190);
nand U146 (N_146,In_2861,In_1379);
nor U147 (N_147,In_2666,In_1529);
and U148 (N_148,In_2547,In_2778);
xor U149 (N_149,In_1283,In_1008);
or U150 (N_150,In_1724,In_1457);
nor U151 (N_151,In_1626,In_2991);
and U152 (N_152,In_705,In_1004);
and U153 (N_153,In_704,In_1446);
xor U154 (N_154,In_393,In_363);
and U155 (N_155,In_2686,In_940);
nor U156 (N_156,In_2479,In_88);
nor U157 (N_157,In_2345,In_1143);
nor U158 (N_158,In_1346,In_258);
nor U159 (N_159,In_2854,In_1164);
nor U160 (N_160,In_2712,In_2626);
nor U161 (N_161,In_2236,In_1577);
and U162 (N_162,In_79,In_503);
and U163 (N_163,In_1440,In_2971);
nand U164 (N_164,In_1167,In_2461);
nor U165 (N_165,In_544,In_1769);
and U166 (N_166,In_1624,In_35);
and U167 (N_167,In_1872,In_1612);
nand U168 (N_168,In_206,In_1432);
nor U169 (N_169,In_1497,In_1528);
or U170 (N_170,In_520,In_2601);
nand U171 (N_171,In_645,In_2697);
or U172 (N_172,In_1622,In_1295);
xnor U173 (N_173,In_2376,In_892);
xor U174 (N_174,In_2749,In_166);
xnor U175 (N_175,In_1700,In_630);
nand U176 (N_176,In_129,In_2121);
xnor U177 (N_177,In_1565,In_1162);
and U178 (N_178,In_2019,In_1067);
xnor U179 (N_179,In_434,In_864);
nor U180 (N_180,In_1888,In_1803);
nor U181 (N_181,In_2871,In_176);
and U182 (N_182,In_164,In_2216);
nand U183 (N_183,In_76,In_2091);
nor U184 (N_184,In_2253,In_2924);
or U185 (N_185,In_577,In_2679);
and U186 (N_186,In_299,In_887);
nor U187 (N_187,In_212,In_1356);
nor U188 (N_188,In_144,In_119);
or U189 (N_189,In_588,In_162);
and U190 (N_190,In_1367,In_288);
nand U191 (N_191,In_1901,In_307);
nand U192 (N_192,In_686,In_1555);
nor U193 (N_193,In_2340,In_456);
and U194 (N_194,In_522,In_2286);
nor U195 (N_195,In_2200,In_265);
nor U196 (N_196,In_2630,In_2309);
nor U197 (N_197,In_1476,In_1083);
and U198 (N_198,In_2168,In_2821);
nand U199 (N_199,In_492,In_1050);
xnor U200 (N_200,In_2439,In_1504);
xor U201 (N_201,In_656,In_1300);
nand U202 (N_202,In_40,In_2129);
or U203 (N_203,In_327,In_1696);
and U204 (N_204,In_2657,In_1784);
xor U205 (N_205,In_2460,In_2777);
or U206 (N_206,In_2172,In_1549);
or U207 (N_207,In_839,In_1465);
and U208 (N_208,In_1159,In_374);
nor U209 (N_209,In_1695,In_1179);
or U210 (N_210,In_871,In_936);
xnor U211 (N_211,In_568,In_699);
nor U212 (N_212,In_301,In_2619);
or U213 (N_213,In_2604,In_1928);
and U214 (N_214,In_421,In_2308);
nor U215 (N_215,In_1548,In_617);
nor U216 (N_216,In_1967,In_2362);
xnor U217 (N_217,In_2134,In_1191);
or U218 (N_218,In_2759,In_1322);
nand U219 (N_219,In_2555,In_2769);
or U220 (N_220,In_2721,In_972);
and U221 (N_221,In_1994,In_504);
or U222 (N_222,In_826,In_2751);
and U223 (N_223,In_975,In_1675);
nor U224 (N_224,In_2493,In_2767);
or U225 (N_225,In_2516,In_908);
xor U226 (N_226,In_2976,In_1896);
nand U227 (N_227,In_2544,In_412);
nand U228 (N_228,In_2277,In_722);
nor U229 (N_229,In_93,In_799);
xor U230 (N_230,In_1209,In_2029);
nand U231 (N_231,In_23,In_1899);
xor U232 (N_232,In_1048,In_2207);
and U233 (N_233,In_1936,In_2704);
or U234 (N_234,In_1706,In_2488);
or U235 (N_235,In_712,In_377);
xor U236 (N_236,In_2325,In_2353);
nor U237 (N_237,In_1213,In_794);
nand U238 (N_238,In_753,In_2703);
xnor U239 (N_239,In_2539,In_2628);
or U240 (N_240,In_1368,In_281);
nor U241 (N_241,In_1238,In_786);
xnor U242 (N_242,In_94,In_1389);
nand U243 (N_243,In_795,In_2483);
nand U244 (N_244,In_1252,In_1441);
or U245 (N_245,In_822,In_2245);
xor U246 (N_246,In_2990,In_613);
nor U247 (N_247,In_1520,In_1846);
or U248 (N_248,In_1332,In_845);
or U249 (N_249,In_330,In_2062);
nor U250 (N_250,In_1687,In_1350);
and U251 (N_251,In_644,In_2725);
and U252 (N_252,In_2765,In_560);
or U253 (N_253,In_734,In_2685);
and U254 (N_254,In_311,In_1436);
nor U255 (N_255,In_1949,In_2288);
xor U256 (N_256,In_1510,In_1788);
or U257 (N_257,In_1076,In_2451);
and U258 (N_258,In_2910,In_44);
nand U259 (N_259,In_222,In_452);
nor U260 (N_260,In_2989,In_1154);
nor U261 (N_261,In_1297,In_2219);
xor U262 (N_262,In_1087,In_17);
nor U263 (N_263,In_2230,In_1171);
nand U264 (N_264,In_2073,In_468);
nor U265 (N_265,In_815,In_376);
nor U266 (N_266,In_2665,In_221);
nor U267 (N_267,In_1197,In_1487);
nor U268 (N_268,In_137,In_466);
nand U269 (N_269,In_918,In_1991);
nor U270 (N_270,In_475,In_810);
nor U271 (N_271,In_1038,In_2124);
xor U272 (N_272,In_184,In_106);
nand U273 (N_273,In_2065,In_1969);
and U274 (N_274,In_2728,In_171);
xor U275 (N_275,In_2143,In_1015);
or U276 (N_276,In_178,In_1698);
xor U277 (N_277,In_1425,In_1829);
nor U278 (N_278,In_639,In_579);
and U279 (N_279,In_267,In_1224);
xnor U280 (N_280,In_981,In_565);
nor U281 (N_281,In_1261,In_229);
xnor U282 (N_282,In_1324,In_2321);
or U283 (N_283,In_2045,In_2495);
xor U284 (N_284,In_881,In_2783);
nor U285 (N_285,In_592,In_2009);
or U286 (N_286,In_241,In_2633);
nor U287 (N_287,In_1214,In_2581);
and U288 (N_288,In_514,In_635);
and U289 (N_289,In_1274,In_1597);
xor U290 (N_290,In_1581,In_2875);
or U291 (N_291,In_2888,In_2217);
nand U292 (N_292,In_2179,In_185);
or U293 (N_293,In_2242,In_1544);
and U294 (N_294,In_1285,In_1494);
nand U295 (N_295,In_2585,In_1180);
or U296 (N_296,In_420,In_2477);
and U297 (N_297,In_1046,In_2937);
or U298 (N_298,In_2879,In_2314);
or U299 (N_299,In_2915,In_1184);
and U300 (N_300,In_1516,In_1124);
nor U301 (N_301,In_2747,In_1902);
and U302 (N_302,In_1682,In_2188);
or U303 (N_303,In_1730,In_177);
and U304 (N_304,In_1455,In_1424);
or U305 (N_305,In_260,In_2154);
nand U306 (N_306,In_850,In_1560);
xnor U307 (N_307,In_437,In_2835);
and U308 (N_308,In_727,In_1837);
nor U309 (N_309,In_621,In_415);
and U310 (N_310,In_1467,In_1381);
and U311 (N_311,In_1676,In_1621);
and U312 (N_312,In_2774,In_659);
or U313 (N_313,In_2886,In_1550);
nor U314 (N_314,In_1139,In_274);
or U315 (N_315,In_2710,In_2868);
nor U316 (N_316,In_803,In_1017);
nand U317 (N_317,In_796,In_2452);
nor U318 (N_318,In_153,In_2350);
xor U319 (N_319,In_1506,In_2468);
nand U320 (N_320,In_2145,In_2923);
nand U321 (N_321,In_1832,In_2476);
or U322 (N_322,In_2675,In_944);
nor U323 (N_323,In_1168,In_2011);
nor U324 (N_324,In_264,In_2515);
and U325 (N_325,In_2251,In_1318);
xnor U326 (N_326,In_2926,In_1992);
or U327 (N_327,In_1140,In_2190);
nor U328 (N_328,In_662,In_2948);
nor U329 (N_329,In_2241,In_941);
or U330 (N_330,In_2607,In_2104);
nand U331 (N_331,In_812,In_761);
nor U332 (N_332,In_1648,In_1236);
or U333 (N_333,In_1406,In_1307);
or U334 (N_334,In_825,In_679);
and U335 (N_335,In_2670,In_2212);
nor U336 (N_336,In_1972,In_1664);
and U337 (N_337,In_1847,In_1690);
and U338 (N_338,In_298,In_1473);
and U339 (N_339,In_333,In_590);
or U340 (N_340,In_1092,In_2920);
and U341 (N_341,In_2566,In_1807);
nor U342 (N_342,In_2687,In_1962);
nand U343 (N_343,In_1320,In_2756);
nand U344 (N_344,In_427,In_2438);
nand U345 (N_345,In_601,In_2732);
nor U346 (N_346,In_411,In_2785);
and U347 (N_347,In_2611,In_1141);
and U348 (N_348,In_1396,In_745);
or U349 (N_349,In_1632,In_905);
and U350 (N_350,In_1105,In_1875);
and U351 (N_351,In_695,In_251);
nor U352 (N_352,In_2006,In_2231);
xor U353 (N_353,In_2205,In_1605);
xor U354 (N_354,In_2147,In_757);
nor U355 (N_355,In_134,In_2946);
or U356 (N_356,In_457,In_2263);
nand U357 (N_357,In_2482,In_1718);
or U358 (N_358,In_2908,In_604);
or U359 (N_359,In_968,In_1848);
and U360 (N_360,In_1865,In_2239);
or U361 (N_361,In_1010,In_1172);
nand U362 (N_362,In_467,In_2387);
or U363 (N_363,In_654,In_2889);
nand U364 (N_364,In_535,In_436);
and U365 (N_365,In_2537,In_226);
xnor U366 (N_366,In_1811,In_1923);
nor U367 (N_367,In_1248,In_945);
nor U368 (N_368,In_1311,In_65);
nor U369 (N_369,In_1611,In_543);
and U370 (N_370,In_2443,In_1630);
nand U371 (N_371,In_548,In_83);
or U372 (N_372,In_75,In_2402);
nand U373 (N_373,In_1086,In_256);
xnor U374 (N_374,In_506,In_1655);
and U375 (N_375,In_47,In_25);
or U376 (N_376,In_2414,In_383);
xnor U377 (N_377,In_1391,In_986);
nand U378 (N_378,In_2007,In_1265);
and U379 (N_379,In_2316,In_1226);
nand U380 (N_380,In_976,In_523);
nand U381 (N_381,In_189,In_2629);
nor U382 (N_382,In_2691,In_2650);
nand U383 (N_383,In_880,In_2553);
nor U384 (N_384,In_1735,In_2141);
or U385 (N_385,In_1175,In_903);
nor U386 (N_386,In_2044,In_2227);
xor U387 (N_387,In_2762,In_1026);
xor U388 (N_388,In_2036,In_1070);
nor U389 (N_389,In_315,In_2433);
nor U390 (N_390,In_2425,In_950);
nand U391 (N_391,In_2499,In_2939);
nor U392 (N_392,In_2296,In_2614);
nand U393 (N_393,In_1178,In_438);
nand U394 (N_394,In_2930,In_2892);
nor U395 (N_395,In_337,In_1654);
or U396 (N_396,In_354,In_2415);
nor U397 (N_397,In_357,In_390);
and U398 (N_398,In_1591,In_818);
xor U399 (N_399,In_2742,In_953);
nand U400 (N_400,In_1688,In_2815);
xnor U401 (N_401,In_2240,In_1816);
xnor U402 (N_402,In_756,In_1892);
nand U403 (N_403,In_101,In_2549);
nand U404 (N_404,In_1618,In_648);
and U405 (N_405,In_2467,In_2118);
and U406 (N_406,In_1575,In_2513);
nor U407 (N_407,In_1326,In_447);
nor U408 (N_408,In_1374,In_403);
or U409 (N_409,In_2463,In_2661);
xnor U410 (N_410,In_1671,In_2828);
and U411 (N_411,In_2349,In_1025);
nor U412 (N_412,In_1943,In_1944);
nor U413 (N_413,In_1500,In_2802);
xnor U414 (N_414,In_748,In_1961);
xnor U415 (N_415,In_2978,In_1203);
or U416 (N_416,In_2833,In_114);
xor U417 (N_417,In_1699,In_1431);
or U418 (N_418,In_2426,In_2088);
or U419 (N_419,In_1995,In_70);
or U420 (N_420,In_1745,In_1708);
and U421 (N_421,In_1068,In_2519);
nor U422 (N_422,In_424,In_1247);
and U423 (N_423,In_1585,In_2453);
nor U424 (N_424,In_1475,In_2388);
or U425 (N_425,In_1433,In_423);
nand U426 (N_426,In_66,In_672);
xor U427 (N_427,In_1372,In_2022);
nand U428 (N_428,In_2956,In_702);
nand U429 (N_429,In_159,In_1762);
or U430 (N_430,In_2410,In_798);
or U431 (N_431,In_1439,In_1375);
nand U432 (N_432,In_602,In_2819);
and U433 (N_433,In_2883,In_130);
and U434 (N_434,In_2954,In_1578);
xnor U435 (N_435,In_1937,In_208);
nand U436 (N_436,In_1819,In_2702);
nand U437 (N_437,In_1794,In_1376);
nor U438 (N_438,In_1409,In_1312);
nor U439 (N_439,In_1098,In_2925);
xor U440 (N_440,In_1704,In_2140);
nand U441 (N_441,In_245,In_15);
xnor U442 (N_442,In_2786,In_788);
and U443 (N_443,In_2891,In_1080);
xnor U444 (N_444,In_2341,In_2540);
and U445 (N_445,In_2470,In_1119);
and U446 (N_446,In_470,In_120);
or U447 (N_447,In_1109,In_2175);
or U448 (N_448,In_1369,In_2668);
nand U449 (N_449,In_623,In_2911);
nand U450 (N_450,In_2906,In_2663);
and U451 (N_451,In_1402,In_170);
nand U452 (N_452,In_2333,In_325);
or U453 (N_453,In_61,In_674);
and U454 (N_454,In_1047,In_1857);
or U455 (N_455,In_1713,In_1397);
xnor U456 (N_456,In_1634,In_2589);
nor U457 (N_457,In_1952,In_1395);
and U458 (N_458,In_2773,In_413);
nor U459 (N_459,In_2775,In_1966);
xnor U460 (N_460,In_145,In_1259);
or U461 (N_461,In_2355,In_2061);
nor U462 (N_462,In_28,In_2842);
and U463 (N_463,In_1731,In_2964);
nor U464 (N_464,In_872,In_2127);
nor U465 (N_465,In_1044,In_683);
nand U466 (N_466,In_2448,In_1201);
nand U467 (N_467,In_148,In_2529);
and U468 (N_468,In_873,In_2730);
nor U469 (N_469,In_2135,In_462);
nor U470 (N_470,In_1001,In_1712);
xnor U471 (N_471,In_2580,In_2021);
nand U472 (N_472,In_988,In_205);
or U473 (N_473,In_1849,In_2546);
xor U474 (N_474,In_1741,In_1470);
xnor U475 (N_475,In_1027,In_2182);
or U476 (N_476,In_2165,In_1759);
xnor U477 (N_477,In_651,In_277);
or U478 (N_478,In_328,In_2536);
xor U479 (N_479,In_688,In_1960);
or U480 (N_480,In_801,In_782);
or U481 (N_481,In_789,In_2932);
xnor U482 (N_482,In_1069,In_709);
xnor U483 (N_483,In_2059,In_1204);
and U484 (N_484,In_152,In_2642);
xor U485 (N_485,In_2763,In_2708);
nand U486 (N_486,In_1288,In_1625);
xor U487 (N_487,In_2105,In_1920);
xnor U488 (N_488,In_557,In_1427);
or U489 (N_489,In_966,In_2327);
nor U490 (N_490,In_1103,In_675);
nand U491 (N_491,In_2858,In_633);
or U492 (N_492,In_2865,In_1884);
xor U493 (N_493,In_542,In_2281);
nor U494 (N_494,In_819,In_179);
xnor U495 (N_495,In_2046,In_1777);
xor U496 (N_496,In_2736,In_77);
xnor U497 (N_497,In_2707,In_1480);
nand U498 (N_498,In_750,In_581);
xor U499 (N_499,In_1852,In_1466);
nand U500 (N_500,In_1129,In_2119);
and U501 (N_501,In_853,In_1384);
nand U502 (N_502,In_2037,In_859);
nand U503 (N_503,In_2429,In_45);
nor U504 (N_504,In_1254,In_2744);
or U505 (N_505,In_2896,In_1812);
xnor U506 (N_506,In_1187,In_1533);
or U507 (N_507,In_2995,In_2796);
nand U508 (N_508,In_2199,In_1953);
or U509 (N_509,In_477,In_2399);
or U510 (N_510,In_1138,In_511);
or U511 (N_511,In_496,In_930);
xor U512 (N_512,In_571,In_2636);
xnor U513 (N_513,In_1948,In_2583);
nor U514 (N_514,In_2056,In_787);
xor U515 (N_515,In_1106,In_2820);
or U516 (N_516,In_2643,In_2780);
xnor U517 (N_517,In_1192,In_598);
nor U518 (N_518,In_341,In_2064);
or U519 (N_519,In_2416,In_1919);
and U520 (N_520,In_2922,In_2983);
xor U521 (N_521,In_916,In_2855);
or U522 (N_522,In_1279,In_2186);
nand U523 (N_523,In_181,In_2282);
and U524 (N_524,In_2381,In_1828);
and U525 (N_525,In_2620,In_287);
and U526 (N_526,In_1758,In_895);
nor U527 (N_527,In_2645,In_2191);
or U528 (N_528,In_1883,In_586);
nor U529 (N_529,In_1215,In_203);
xnor U530 (N_530,In_2054,In_1243);
and U531 (N_531,In_1323,In_1592);
nor U532 (N_532,In_1365,In_2974);
or U533 (N_533,In_2653,In_1107);
or U534 (N_534,In_2401,In_620);
and U535 (N_535,In_2184,In_116);
nand U536 (N_536,In_591,In_2012);
and U537 (N_537,In_827,In_1881);
or U538 (N_538,In_835,In_2466);
xor U539 (N_539,In_2718,In_96);
and U540 (N_540,In_283,In_303);
nor U541 (N_541,In_1909,In_1195);
nand U542 (N_542,In_143,In_781);
nand U543 (N_543,In_914,In_2085);
xor U544 (N_544,In_1940,In_1508);
or U545 (N_545,In_1325,In_554);
or U546 (N_546,In_1756,In_2265);
nand U547 (N_547,In_2694,In_938);
nand U548 (N_548,In_1145,In_358);
nand U549 (N_549,In_2696,In_248);
nand U550 (N_550,In_2268,In_2214);
nor U551 (N_551,In_898,In_175);
and U552 (N_552,In_573,In_210);
or U553 (N_553,In_1562,In_946);
xor U554 (N_554,In_830,In_2542);
nand U555 (N_555,In_1462,In_1669);
xor U556 (N_556,In_855,In_29);
xnor U557 (N_557,In_1744,In_2558);
or U558 (N_558,In_371,In_1352);
nor U559 (N_559,In_1527,In_2113);
nor U560 (N_560,In_1118,In_561);
and U561 (N_561,In_402,In_951);
xor U562 (N_562,In_209,In_2001);
nor U563 (N_563,In_1752,In_811);
xnor U564 (N_564,In_2985,In_1347);
nor U565 (N_565,In_122,In_2446);
xnor U566 (N_566,In_2916,In_2016);
nor U567 (N_567,In_2382,In_1925);
or U568 (N_568,In_1458,In_1786);
nand U569 (N_569,In_2005,In_278);
xor U570 (N_570,In_2408,In_2706);
or U571 (N_571,In_1678,In_2806);
nand U572 (N_572,In_2631,In_1442);
and U573 (N_573,In_1964,In_142);
or U574 (N_574,In_1132,In_628);
or U575 (N_575,In_1620,In_729);
xor U576 (N_576,In_1211,In_2404);
and U577 (N_577,In_2867,In_485);
xor U578 (N_578,In_763,In_2684);
and U579 (N_579,In_814,In_562);
and U580 (N_580,In_2612,In_2723);
xnor U581 (N_581,In_1673,In_1278);
nand U582 (N_582,In_1403,In_196);
nand U583 (N_583,In_1999,In_2364);
nand U584 (N_584,In_365,In_894);
nand U585 (N_585,In_1407,In_2396);
nand U586 (N_586,In_2445,In_1496);
and U587 (N_587,In_2050,In_2369);
nand U588 (N_588,In_2436,In_1094);
xor U589 (N_589,In_1763,In_1077);
and U590 (N_590,In_133,In_2081);
nand U591 (N_591,In_2422,In_1182);
or U592 (N_592,In_2174,In_1383);
xnor U593 (N_593,In_193,In_1387);
and U594 (N_594,In_558,In_886);
xor U595 (N_595,In_1413,In_611);
nand U596 (N_596,In_2794,In_1163);
and U597 (N_597,In_2904,In_754);
nor U598 (N_598,In_280,In_2862);
and U599 (N_599,In_2018,In_2421);
and U600 (N_600,N_20,In_1233);
and U601 (N_601,N_411,N_433);
nor U602 (N_602,In_671,In_2587);
nor U603 (N_603,N_291,In_316);
nand U604 (N_604,In_2158,In_2750);
and U605 (N_605,In_1543,N_596);
xnor U606 (N_606,N_322,In_2111);
or U607 (N_607,In_2255,In_1398);
nand U608 (N_608,N_110,N_266);
or U609 (N_609,N_262,In_347);
nand U610 (N_610,In_1055,In_837);
nor U611 (N_611,In_1879,In_2596);
nand U612 (N_612,In_681,N_577);
or U613 (N_613,In_1418,N_540);
or U614 (N_614,In_1286,N_76);
and U615 (N_615,In_1573,In_1411);
nand U616 (N_616,In_2776,In_2274);
and U617 (N_617,N_422,N_89);
nor U618 (N_618,In_1073,In_2500);
or U619 (N_619,In_246,In_1490);
or U620 (N_620,In_2561,In_2905);
nor U621 (N_621,In_2449,In_2260);
nor U622 (N_622,In_2571,In_999);
nand U623 (N_623,In_2846,In_1299);
and U624 (N_624,In_844,In_254);
xnor U625 (N_625,In_417,N_559);
and U626 (N_626,In_2818,In_2502);
or U627 (N_627,In_2677,In_2033);
or U628 (N_628,N_133,N_210);
xnor U629 (N_629,In_739,N_228);
and U630 (N_630,In_198,N_315);
nor U631 (N_631,In_1056,N_551);
and U632 (N_632,In_2623,N_357);
nand U633 (N_633,In_2729,In_1007);
nand U634 (N_634,In_1485,In_1085);
nor U635 (N_635,In_95,In_1366);
nor U636 (N_636,N_269,In_132);
xor U637 (N_637,In_546,N_408);
nor U638 (N_638,In_2089,N_55);
xnor U639 (N_639,In_1033,N_242);
xnor U640 (N_640,In_2455,In_2823);
and U641 (N_641,In_296,In_2481);
xor U642 (N_642,In_2919,In_537);
xor U643 (N_643,In_429,N_509);
and U644 (N_644,In_1190,In_2984);
nor U645 (N_645,N_84,In_497);
nand U646 (N_646,In_1821,N_80);
nand U647 (N_647,N_531,In_1343);
nand U648 (N_648,In_2552,In_1900);
xnor U649 (N_649,In_2312,N_169);
xor U650 (N_650,In_2573,In_2366);
nand U651 (N_651,N_403,In_2616);
nand U652 (N_652,In_927,In_2724);
and U653 (N_653,In_1390,N_384);
nor U654 (N_654,In_2510,In_2683);
nand U655 (N_655,N_191,N_152);
xnor U656 (N_656,N_97,In_678);
and U657 (N_657,In_1232,In_1743);
nand U658 (N_658,N_120,In_2167);
or U659 (N_659,In_806,In_1804);
nor U660 (N_660,In_1061,In_1222);
xor U661 (N_661,N_387,In_1249);
nand U662 (N_662,In_2944,In_2244);
nand U663 (N_663,In_67,In_2100);
nand U664 (N_664,In_715,N_42);
or U665 (N_665,In_706,In_933);
or U666 (N_666,N_455,In_407);
xor U667 (N_667,N_353,In_1329);
xor U668 (N_668,In_382,In_821);
nor U669 (N_669,In_1747,In_2909);
nor U670 (N_670,In_995,In_2535);
or U671 (N_671,In_957,In_489);
xnor U672 (N_672,In_603,In_446);
and U673 (N_673,In_540,In_2584);
and U674 (N_674,In_2013,In_987);
and U675 (N_675,In_2824,In_2365);
nor U676 (N_676,N_63,In_1963);
xnor U677 (N_677,N_424,In_2010);
xor U678 (N_678,In_2681,N_440);
xor U679 (N_679,In_2568,In_780);
nand U680 (N_680,In_1557,N_447);
xor U681 (N_681,In_1041,N_416);
xnor U682 (N_682,In_285,In_2508);
xnor U683 (N_683,In_1929,In_1521);
or U684 (N_684,N_25,In_131);
xor U685 (N_685,N_473,N_91);
nor U686 (N_686,In_244,In_2163);
nand U687 (N_687,In_896,N_108);
nor U688 (N_688,In_735,In_1737);
and U689 (N_689,N_218,In_2144);
xor U690 (N_690,In_861,In_770);
and U691 (N_691,In_1155,N_464);
nand U692 (N_692,In_1607,In_2960);
or U693 (N_693,In_1373,N_556);
nor U694 (N_694,In_2430,In_1166);
nand U695 (N_695,N_501,In_1910);
and U696 (N_696,In_740,In_2248);
nor U697 (N_697,In_2068,In_1647);
nor U698 (N_698,In_2624,N_591);
nand U699 (N_699,In_2270,In_2090);
xor U700 (N_700,In_1684,In_570);
or U701 (N_701,In_2550,In_127);
nand U702 (N_702,In_1013,N_241);
and U703 (N_703,In_2069,N_156);
xor U704 (N_704,In_1043,N_140);
or U705 (N_705,N_128,In_2084);
nand U706 (N_706,N_581,In_2726);
xor U707 (N_707,In_959,In_218);
nand U708 (N_708,In_1072,N_153);
or U709 (N_709,In_2688,In_1855);
xor U710 (N_710,In_2328,In_431);
or U711 (N_711,In_508,N_407);
nor U712 (N_712,N_74,N_230);
xor U713 (N_713,N_359,In_778);
or U714 (N_714,In_2790,N_261);
nand U715 (N_715,In_1791,In_2881);
nand U716 (N_716,In_1890,N_507);
xor U717 (N_717,In_1785,In_2999);
nor U718 (N_718,In_1280,In_33);
xnor U719 (N_719,N_255,In_1498);
nor U720 (N_720,In_1680,In_1951);
or U721 (N_721,N_530,In_2599);
nor U722 (N_722,N_151,In_751);
nor U723 (N_723,N_503,In_1932);
nor U724 (N_724,N_206,In_878);
nand U725 (N_725,In_2695,In_2202);
or U726 (N_726,N_563,N_176);
nand U727 (N_727,N_160,In_2740);
or U728 (N_728,In_2947,In_1217);
nor U729 (N_729,In_2988,In_2548);
nor U730 (N_730,In_955,In_2052);
xor U731 (N_731,In_993,In_1774);
or U732 (N_732,In_1016,In_1600);
nor U733 (N_733,In_2257,In_2262);
and U734 (N_734,In_2109,In_2651);
nand U735 (N_735,In_2112,In_682);
and U736 (N_736,N_355,In_2996);
and U737 (N_737,N_101,In_297);
nand U738 (N_738,In_2485,N_94);
nand U739 (N_739,In_1404,In_634);
nor U740 (N_740,N_227,In_1188);
nand U741 (N_741,In_1723,In_690);
or U742 (N_742,In_758,N_282);
xor U743 (N_743,In_1633,In_2514);
and U744 (N_744,In_1594,In_2162);
and U745 (N_745,In_2,N_61);
or U746 (N_746,In_1551,N_198);
or U747 (N_747,In_998,N_532);
nor U748 (N_748,In_1136,In_2249);
and U749 (N_749,In_1151,In_1580);
xnor U750 (N_750,In_2159,In_13);
nand U751 (N_751,In_1935,In_1609);
and U752 (N_752,In_289,In_2417);
nor U753 (N_753,In_922,In_2278);
and U754 (N_754,In_2375,In_1091);
nand U755 (N_755,In_2898,In_1831);
nand U756 (N_756,N_47,In_6);
xor U757 (N_757,N_232,N_253);
or U758 (N_758,In_1702,N_572);
and U759 (N_759,In_670,In_2225);
and U760 (N_760,In_1328,N_550);
and U761 (N_761,In_2816,In_2673);
nand U762 (N_762,In_2283,In_1385);
xnor U763 (N_763,In_2579,N_78);
nand U764 (N_764,In_657,In_1637);
xnor U765 (N_765,In_2928,In_2298);
and U766 (N_766,In_841,N_90);
xor U767 (N_767,In_1727,N_522);
xnor U768 (N_768,In_1524,N_158);
and U769 (N_769,In_86,In_609);
or U770 (N_770,N_111,In_385);
nand U771 (N_771,N_413,In_156);
nor U772 (N_772,In_478,In_1787);
and U773 (N_773,In_494,In_1885);
nor U774 (N_774,N_248,N_425);
and U775 (N_775,In_1531,N_516);
or U776 (N_776,N_14,N_44);
or U777 (N_777,N_366,In_1709);
xnor U778 (N_778,In_2080,In_361);
nand U779 (N_779,In_2678,In_1656);
nor U780 (N_780,In_891,In_191);
and U781 (N_781,In_2096,N_363);
nand U782 (N_782,In_631,In_2938);
nand U783 (N_783,In_2313,In_2504);
nor U784 (N_784,In_732,N_568);
nor U785 (N_785,In_1257,In_533);
nor U786 (N_786,In_1836,N_290);
xnor U787 (N_787,In_1477,In_324);
or U788 (N_788,N_356,N_490);
and U789 (N_789,In_2761,In_151);
xor U790 (N_790,N_130,In_5);
nor U791 (N_791,In_692,In_527);
or U792 (N_792,N_460,In_515);
xor U793 (N_793,In_2380,In_157);
nand U794 (N_794,In_349,In_791);
or U795 (N_795,In_1160,In_2852);
and U796 (N_796,In_2955,N_166);
or U797 (N_797,N_341,In_2047);
and U798 (N_798,In_1464,N_50);
nand U799 (N_799,In_2048,N_595);
and U800 (N_800,In_2176,In_31);
xnor U801 (N_801,In_85,In_1054);
or U802 (N_802,In_2635,In_2731);
nor U803 (N_803,N_121,N_43);
nand U804 (N_804,In_332,In_141);
nand U805 (N_805,In_1509,In_391);
or U806 (N_806,In_2847,In_2639);
nand U807 (N_807,In_2518,In_2338);
nor U808 (N_808,In_2306,In_168);
xor U809 (N_809,In_2638,In_1984);
and U810 (N_810,In_473,In_1364);
and U811 (N_811,In_243,In_1023);
and U812 (N_812,In_2373,In_2437);
or U813 (N_813,In_1239,N_35);
or U814 (N_814,In_664,In_948);
or U815 (N_815,In_1463,N_267);
nand U816 (N_816,N_268,In_2848);
and U817 (N_817,In_752,In_1608);
nand U818 (N_818,In_963,In_701);
or U819 (N_819,N_336,In_1200);
nand U820 (N_820,N_428,In_1443);
or U821 (N_821,In_235,In_2735);
nor U822 (N_822,In_1643,In_2335);
nor U823 (N_823,N_102,N_542);
nand U824 (N_824,In_768,In_994);
nand U825 (N_825,In_2822,In_985);
xnor U826 (N_826,N_498,In_2781);
nand U827 (N_827,In_925,In_755);
and U828 (N_828,In_1750,In_284);
and U829 (N_829,In_1493,In_899);
xor U830 (N_830,N_337,N_217);
nand U831 (N_831,In_1130,In_1658);
and U832 (N_832,In_529,In_1212);
or U833 (N_833,In_2860,In_2784);
xor U834 (N_834,In_1714,In_1351);
nor U835 (N_835,N_395,In_614);
nor U836 (N_836,In_58,N_429);
and U837 (N_837,In_1754,In_879);
xnor U838 (N_838,In_924,In_465);
and U839 (N_839,In_1334,In_2511);
nor U840 (N_840,In_1749,N_339);
nor U841 (N_841,In_1778,N_34);
and U842 (N_842,In_292,In_2658);
nor U843 (N_843,In_2950,In_1734);
nand U844 (N_844,In_2371,N_442);
nand U845 (N_845,In_112,In_12);
and U846 (N_846,In_1313,In_1456);
xnor U847 (N_847,In_870,In_1864);
or U848 (N_848,In_487,In_366);
nor U849 (N_849,In_1627,In_2959);
nand U850 (N_850,In_2498,In_1020);
nor U851 (N_851,In_279,In_1152);
or U852 (N_852,In_1903,In_1946);
and U853 (N_853,In_625,N_11);
nand U854 (N_854,In_62,In_2053);
or U855 (N_855,In_1386,In_1613);
or U856 (N_856,In_1123,N_476);
or U857 (N_857,In_1309,In_2169);
nor U858 (N_858,In_1768,In_379);
or U859 (N_859,N_427,In_668);
and U860 (N_860,In_583,In_110);
and U861 (N_861,In_1294,In_1660);
and U862 (N_862,In_2567,In_2574);
or U863 (N_863,N_53,In_2506);
and U864 (N_864,In_2475,In_458);
xnor U865 (N_865,In_1773,In_2259);
and U866 (N_866,In_605,In_1761);
nor U867 (N_867,In_713,In_2845);
xor U868 (N_868,In_2841,In_967);
and U869 (N_869,In_1088,In_2357);
and U870 (N_870,In_1635,N_325);
and U871 (N_871,N_419,In_1926);
or U872 (N_872,In_1793,N_124);
xnor U873 (N_873,In_2800,In_1641);
and U874 (N_874,In_2305,In_1636);
xnor U875 (N_875,In_1339,N_149);
and U876 (N_876,In_636,N_148);
nor U877 (N_877,In_217,N_298);
xor U878 (N_878,In_2318,N_238);
xnor U879 (N_879,In_2077,N_420);
nand U880 (N_880,In_55,N_434);
or U881 (N_881,In_680,N_86);
nand U882 (N_882,In_2992,In_840);
nand U883 (N_883,In_1335,N_441);
nand U884 (N_884,N_229,In_890);
or U885 (N_885,In_2193,In_51);
and U886 (N_886,In_619,N_483);
and U887 (N_887,In_772,In_1733);
and U888 (N_888,In_2980,N_181);
nor U889 (N_889,In_237,In_2869);
and U890 (N_890,N_358,In_2532);
or U891 (N_891,In_1277,In_921);
nand U892 (N_892,In_1382,In_1867);
xnor U893 (N_893,In_1380,N_141);
and U894 (N_894,In_2672,In_2299);
or U895 (N_895,In_2690,N_36);
nor U896 (N_896,N_304,In_1271);
and U897 (N_897,In_2782,N_18);
nor U898 (N_898,In_2195,In_2238);
or U899 (N_899,N_9,In_1301);
and U900 (N_900,In_232,N_334);
nor U901 (N_901,N_244,In_1051);
nor U902 (N_902,In_1338,N_95);
nand U903 (N_903,In_2368,N_66);
nor U904 (N_904,In_553,N_443);
nor U905 (N_905,In_2003,In_730);
or U906 (N_906,N_349,In_1757);
nor U907 (N_907,In_741,In_1579);
and U908 (N_908,In_1795,In_1445);
nor U909 (N_909,In_2002,In_1593);
nor U910 (N_910,In_2505,N_475);
or U911 (N_911,N_396,In_111);
and U912 (N_912,In_247,In_2462);
or U913 (N_913,N_514,In_1985);
or U914 (N_914,In_1833,In_2247);
nand U915 (N_915,In_384,In_1572);
and U916 (N_916,In_1125,In_2344);
nor U917 (N_917,N_564,In_216);
nand U918 (N_918,In_138,N_466);
or U919 (N_919,In_2563,In_1345);
or U920 (N_920,In_807,In_1629);
or U921 (N_921,In_1679,In_1924);
and U922 (N_922,N_159,In_2809);
nor U923 (N_923,In_375,In_2839);
nor U924 (N_924,In_2640,N_96);
and U925 (N_925,In_1541,In_2793);
nand U926 (N_926,In_10,In_1717);
xnor U927 (N_927,In_1894,N_144);
xnor U928 (N_928,In_1719,In_1681);
or U929 (N_929,N_309,In_136);
and U930 (N_930,In_63,In_2400);
and U931 (N_931,In_2326,In_46);
and U932 (N_932,In_2880,In_2864);
nand U933 (N_933,In_1358,In_2431);
or U934 (N_934,In_261,In_1071);
nand U935 (N_935,In_2256,In_1460);
and U936 (N_936,In_1823,N_161);
nand U937 (N_937,In_2560,N_444);
nand U938 (N_938,In_717,In_552);
and U939 (N_939,N_257,In_2831);
or U940 (N_940,In_716,In_2131);
nand U941 (N_941,N_239,In_1505);
and U942 (N_942,N_528,In_20);
nor U943 (N_943,In_1799,In_200);
nand U944 (N_944,In_1616,In_1649);
xor U945 (N_945,In_728,In_2067);
and U946 (N_946,In_1858,In_1223);
or U947 (N_947,N_252,In_793);
nand U948 (N_948,N_71,In_64);
and U949 (N_949,In_2078,In_774);
or U950 (N_950,In_449,In_2722);
and U951 (N_951,In_809,In_2086);
nor U952 (N_952,In_1554,N_87);
nor U953 (N_953,In_2060,In_2473);
nor U954 (N_954,N_287,N_406);
or U955 (N_955,In_225,In_1536);
or U956 (N_956,In_1601,N_352);
xor U957 (N_957,In_126,N_372);
nor U958 (N_958,In_1539,N_389);
xor U959 (N_959,N_318,N_404);
and U960 (N_960,In_135,N_126);
nand U961 (N_961,In_2412,In_1530);
nand U962 (N_962,In_802,N_397);
nand U963 (N_963,In_2741,N_10);
nor U964 (N_964,N_211,In_2472);
or U965 (N_965,In_512,In_1198);
or U966 (N_966,In_1589,In_882);
or U967 (N_967,In_643,In_911);
xnor U968 (N_968,N_297,N_197);
xnor U969 (N_969,In_2442,In_2715);
or U970 (N_970,In_743,N_462);
nand U971 (N_971,In_1042,In_271);
and U972 (N_972,In_1582,In_2680);
nor U973 (N_973,N_414,In_877);
nor U974 (N_974,In_1662,N_571);
nand U975 (N_975,N_583,In_2038);
nor U976 (N_976,In_1024,In_2289);
or U977 (N_977,N_569,In_2226);
nand U978 (N_978,In_1081,In_2004);
and U979 (N_979,N_163,In_2646);
xnor U980 (N_980,N_209,In_220);
nor U981 (N_981,In_1868,In_2074);
or U982 (N_982,N_171,In_1905);
and U983 (N_983,In_1186,In_990);
xor U984 (N_984,In_109,N_558);
or U985 (N_985,In_72,In_69);
xor U986 (N_986,In_2287,N_202);
and U987 (N_987,In_1546,In_1619);
nor U988 (N_988,In_2569,In_2471);
xor U989 (N_989,N_69,In_2456);
xor U990 (N_990,In_519,In_723);
nor U991 (N_991,In_1451,In_1438);
xor U992 (N_992,N_520,N_329);
nand U993 (N_993,In_1291,In_37);
or U994 (N_994,In_2840,In_48);
nor U995 (N_995,In_1552,In_1854);
nand U996 (N_996,N_3,In_1912);
and U997 (N_997,In_2323,In_2931);
xor U998 (N_998,N_31,In_860);
nor U999 (N_999,In_0,In_1563);
nand U1000 (N_1000,In_2874,In_2853);
xor U1001 (N_1001,N_346,In_2295);
xor U1002 (N_1002,In_836,N_578);
nand U1003 (N_1003,In_2863,In_900);
xnor U1004 (N_1004,In_2057,In_550);
or U1005 (N_1005,N_28,In_2739);
nand U1006 (N_1006,N_579,In_201);
nand U1007 (N_1007,In_1644,In_616);
nand U1008 (N_1008,In_719,In_2424);
nor U1009 (N_1009,In_700,N_243);
xor U1010 (N_1010,N_49,N_454);
xor U1011 (N_1011,In_842,In_2595);
and U1012 (N_1012,In_1783,In_2358);
nand U1013 (N_1013,In_2807,In_749);
nor U1014 (N_1014,In_401,N_180);
or U1015 (N_1015,In_517,N_430);
and U1016 (N_1016,In_1898,In_1908);
or U1017 (N_1017,In_2484,In_541);
and U1018 (N_1018,In_733,N_342);
xnor U1019 (N_1019,N_597,In_1736);
nor U1020 (N_1020,In_163,In_2766);
or U1021 (N_1021,In_1599,In_566);
nand U1022 (N_1022,N_565,In_2884);
or U1023 (N_1023,In_1983,In_1694);
nand U1024 (N_1024,In_2304,In_410);
and U1025 (N_1025,In_574,N_538);
nor U1026 (N_1026,In_1045,In_1059);
nand U1027 (N_1027,In_1906,In_1289);
xnor U1028 (N_1028,In_2975,In_1856);
and U1029 (N_1029,In_1792,In_2049);
nand U1030 (N_1030,In_1942,N_251);
and U1031 (N_1031,In_2625,In_2040);
or U1032 (N_1032,N_54,N_281);
xor U1033 (N_1033,In_1990,In_1272);
xor U1034 (N_1034,In_2901,In_2125);
nor U1035 (N_1035,N_512,N_360);
or U1036 (N_1036,N_59,In_1537);
nor U1037 (N_1037,In_2538,In_2943);
nand U1038 (N_1038,In_817,In_624);
xnor U1039 (N_1039,N_453,N_375);
nand U1040 (N_1040,In_1617,In_300);
or U1041 (N_1041,In_125,N_477);
and U1042 (N_1042,In_2753,In_2071);
xnor U1043 (N_1043,N_392,In_2043);
nor U1044 (N_1044,In_534,In_1739);
nand U1045 (N_1045,In_2832,In_2164);
xnor U1046 (N_1046,In_1181,N_409);
and U1047 (N_1047,N_548,N_212);
and U1048 (N_1048,In_49,In_965);
or U1049 (N_1049,In_866,In_1766);
or U1050 (N_1050,In_2136,In_19);
and U1051 (N_1051,In_1269,In_1065);
nor U1052 (N_1052,In_2520,In_2116);
xor U1053 (N_1053,N_70,In_694);
nor U1054 (N_1054,In_2669,In_865);
nand U1055 (N_1055,In_2221,In_502);
or U1056 (N_1056,In_1474,In_1645);
nor U1057 (N_1057,In_253,In_1079);
or U1058 (N_1058,In_2565,N_82);
and U1059 (N_1059,In_2185,In_199);
xnor U1060 (N_1060,In_430,In_1765);
or U1061 (N_1061,In_9,N_2);
or U1062 (N_1062,N_23,In_2079);
and U1063 (N_1063,In_459,In_1437);
nor U1064 (N_1064,In_2171,In_14);
or U1065 (N_1065,N_226,In_1298);
nand U1066 (N_1066,In_2405,In_2570);
nor U1067 (N_1067,In_2676,In_2409);
xnor U1068 (N_1068,In_291,In_2372);
xor U1069 (N_1069,N_274,In_1760);
nor U1070 (N_1070,In_2447,In_1362);
xor U1071 (N_1071,In_1447,In_2324);
nand U1072 (N_1072,N_472,In_2501);
or U1073 (N_1073,In_917,N_165);
nand U1074 (N_1074,In_1378,In_1755);
and U1075 (N_1075,In_2907,In_1193);
nor U1076 (N_1076,In_392,In_2386);
xor U1077 (N_1077,In_397,In_2878);
nor U1078 (N_1078,In_398,N_585);
and U1079 (N_1079,In_1806,In_2294);
xnor U1080 (N_1080,In_500,In_2590);
xnor U1081 (N_1081,In_1400,In_1064);
or U1082 (N_1082,In_884,N_13);
nor U1083 (N_1083,N_310,In_295);
and U1084 (N_1084,In_714,In_2622);
xnor U1085 (N_1085,In_1561,In_2664);
nor U1086 (N_1086,In_3,In_1315);
or U1087 (N_1087,In_1275,In_2393);
nor U1088 (N_1088,In_1144,N_458);
and U1089 (N_1089,In_1697,In_1954);
nor U1090 (N_1090,In_1246,In_493);
and U1091 (N_1091,In_405,In_2792);
nor U1092 (N_1092,N_112,In_1421);
or U1093 (N_1093,In_2507,N_340);
and U1094 (N_1094,In_1907,N_173);
xor U1095 (N_1095,In_1603,In_2395);
xnor U1096 (N_1096,In_2114,In_2877);
xnor U1097 (N_1097,In_2492,In_1);
xor U1098 (N_1098,In_1844,In_1229);
or U1099 (N_1099,N_533,N_527);
xnor U1100 (N_1100,N_319,In_1392);
xor U1101 (N_1101,N_179,In_2652);
nand U1102 (N_1102,In_160,In_784);
xor U1103 (N_1103,In_996,In_428);
and U1104 (N_1104,N_247,In_646);
nor U1105 (N_1105,In_2994,In_2894);
xor U1106 (N_1106,In_1330,In_1715);
and U1107 (N_1107,In_1518,N_549);
nand U1108 (N_1108,In_2027,In_2302);
xnor U1109 (N_1109,N_505,In_2322);
nand U1110 (N_1110,In_1978,In_2183);
nor U1111 (N_1111,In_2465,N_65);
and U1112 (N_1112,In_2949,In_2496);
nor U1113 (N_1113,In_1522,In_2603);
nor U1114 (N_1114,N_109,In_60);
nand U1115 (N_1115,N_320,N_330);
xnor U1116 (N_1116,In_2235,In_513);
or U1117 (N_1117,In_368,N_52);
and U1118 (N_1118,In_1827,In_1417);
nor U1119 (N_1119,In_1174,In_1030);
nor U1120 (N_1120,In_932,In_16);
and U1121 (N_1121,In_422,N_215);
nand U1122 (N_1122,In_2480,In_2733);
or U1123 (N_1123,In_204,In_1495);
or U1124 (N_1124,In_691,In_1638);
nand U1125 (N_1125,In_450,In_2812);
nand U1126 (N_1126,N_1,N_525);
nor U1127 (N_1127,In_1800,N_24);
or U1128 (N_1128,In_174,In_395);
nor U1129 (N_1129,In_282,N_4);
nor U1130 (N_1130,In_1921,In_169);
nor U1131 (N_1131,N_106,In_81);
nand U1132 (N_1132,In_721,In_73);
and U1133 (N_1133,In_769,N_415);
and U1134 (N_1134,In_1194,N_348);
or U1135 (N_1135,N_271,In_1242);
and U1136 (N_1136,In_207,In_2902);
xor U1137 (N_1137,In_2598,In_2745);
xnor U1138 (N_1138,In_2843,N_450);
nor U1139 (N_1139,In_1078,In_2743);
nand U1140 (N_1140,N_324,In_1453);
or U1141 (N_1141,In_2403,In_2801);
or U1142 (N_1142,N_276,In_1221);
and U1143 (N_1143,N_326,In_1918);
or U1144 (N_1144,N_374,N_284);
nor U1145 (N_1145,N_394,In_443);
xnor U1146 (N_1146,In_1877,In_2837);
nand U1147 (N_1147,N_21,In_97);
nand U1148 (N_1148,In_1547,In_2899);
xor U1149 (N_1149,In_2076,In_84);
and U1150 (N_1150,In_1241,N_33);
nor U1151 (N_1151,N_546,In_2173);
or U1152 (N_1152,In_1691,In_1631);
and U1153 (N_1153,N_260,N_136);
nand U1154 (N_1154,In_742,In_663);
nor U1155 (N_1155,In_103,In_983);
nand U1156 (N_1156,N_380,N_321);
nor U1157 (N_1157,In_2367,In_1701);
or U1158 (N_1158,In_2441,In_707);
nand U1159 (N_1159,In_834,In_2940);
xor U1160 (N_1160,In_1052,In_173);
or U1161 (N_1161,In_2758,In_1874);
or U1162 (N_1162,In_2961,In_2098);
and U1163 (N_1163,In_501,In_564);
or U1164 (N_1164,In_1478,In_649);
nand U1165 (N_1165,N_484,In_1360);
xnor U1166 (N_1166,N_172,In_640);
nor U1167 (N_1167,In_257,In_2222);
and U1168 (N_1168,In_367,In_1149);
nor U1169 (N_1169,N_137,In_150);
xor U1170 (N_1170,In_321,N_224);
nor U1171 (N_1171,N_237,In_2213);
nor U1172 (N_1172,In_1202,In_2873);
xor U1173 (N_1173,In_2521,In_2233);
nand U1174 (N_1174,In_1405,In_11);
nor U1175 (N_1175,In_2836,In_2128);
xnor U1176 (N_1176,In_790,N_311);
xnor U1177 (N_1177,In_451,In_647);
nor U1178 (N_1178,In_1813,In_381);
or U1179 (N_1179,N_272,In_1606);
nor U1180 (N_1180,In_2337,In_99);
nor U1181 (N_1181,In_302,In_600);
and U1182 (N_1182,In_396,In_531);
or U1183 (N_1183,In_1615,In_89);
and U1184 (N_1184,N_275,In_346);
or U1185 (N_1185,N_288,In_2458);
nor U1186 (N_1186,N_154,N_383);
and U1187 (N_1187,In_824,N_201);
nand U1188 (N_1188,In_530,In_1461);
nand U1189 (N_1189,In_1484,In_1165);
or U1190 (N_1190,N_361,In_1158);
xnor U1191 (N_1191,N_222,In_1721);
nor U1192 (N_1192,In_828,In_2391);
nor U1193 (N_1193,In_652,In_36);
nand U1194 (N_1194,In_2533,In_2527);
and U1195 (N_1195,In_992,N_145);
or U1196 (N_1196,N_51,In_1227);
nor U1197 (N_1197,In_2593,N_296);
and U1198 (N_1198,In_849,In_215);
or U1199 (N_1199,In_2392,In_2711);
or U1200 (N_1200,In_1568,In_2107);
or U1201 (N_1201,N_1146,N_1002);
nor U1202 (N_1202,N_178,In_2095);
and U1203 (N_1203,In_1880,In_2293);
nand U1204 (N_1204,In_2755,In_2303);
nor U1205 (N_1205,N_887,In_2273);
or U1206 (N_1206,N_977,In_676);
and U1207 (N_1207,In_2427,In_2024);
nand U1208 (N_1208,In_2319,In_1120);
and U1209 (N_1209,N_937,In_2374);
nand U1210 (N_1210,In_2885,N_386);
and U1211 (N_1211,In_344,In_820);
nand U1212 (N_1212,N_586,N_1145);
and U1213 (N_1213,In_1377,N_371);
nor U1214 (N_1214,N_1074,In_2556);
and U1215 (N_1215,N_557,N_1123);
or U1216 (N_1216,N_435,N_589);
nand U1217 (N_1217,N_1163,In_378);
xnor U1218 (N_1218,N_702,N_587);
xnor U1219 (N_1219,N_760,N_46);
and U1220 (N_1220,N_713,N_1135);
nand U1221 (N_1221,N_142,In_509);
nand U1222 (N_1222,N_647,N_676);
and U1223 (N_1223,In_587,N_608);
nor U1224 (N_1224,N_1154,N_367);
and U1225 (N_1225,N_799,N_1101);
xor U1226 (N_1226,In_471,N_784);
nor U1227 (N_1227,In_2014,In_2671);
xor U1228 (N_1228,N_867,In_1115);
nand U1229 (N_1229,In_1479,In_1122);
nand U1230 (N_1230,N_1041,N_1055);
nand U1231 (N_1231,In_1183,N_706);
or U1232 (N_1232,N_1025,N_491);
and U1233 (N_1233,In_1284,N_645);
nor U1234 (N_1234,N_365,N_646);
nor U1235 (N_1235,N_911,N_689);
or U1236 (N_1236,N_916,N_780);
and U1237 (N_1237,In_1640,N_1042);
nor U1238 (N_1238,N_904,N_767);
nand U1239 (N_1239,N_785,In_2093);
nor U1240 (N_1240,N_1037,In_1121);
nand U1241 (N_1241,N_666,N_1095);
or U1242 (N_1242,In_762,N_1152);
nor U1243 (N_1243,N_553,In_1933);
nand U1244 (N_1244,N_417,In_2872);
or U1245 (N_1245,N_1059,N_1138);
nand U1246 (N_1246,In_1208,In_2525);
and U1247 (N_1247,N_1071,N_961);
nor U1248 (N_1248,In_726,In_612);
nor U1249 (N_1249,N_439,N_696);
or U1250 (N_1250,In_1728,In_2958);
or U1251 (N_1251,In_660,N_727);
xnor U1252 (N_1252,N_293,In_1770);
nand U1253 (N_1253,In_1150,N_625);
or U1254 (N_1254,In_78,In_1588);
nor U1255 (N_1255,N_1147,N_1064);
nand U1256 (N_1256,In_2838,In_2963);
nor U1257 (N_1257,In_432,N_1133);
or U1258 (N_1258,In_1981,N_1081);
or U1259 (N_1259,N_614,In_238);
or U1260 (N_1260,N_1089,In_214);
nor U1261 (N_1261,N_620,N_738);
nand U1262 (N_1262,N_1118,N_987);
nor U1263 (N_1263,N_979,In_2192);
nand U1264 (N_1264,N_364,N_279);
nor U1265 (N_1265,N_1184,N_740);
or U1266 (N_1266,N_81,In_2788);
nor U1267 (N_1267,N_914,In_2384);
and U1268 (N_1268,In_1146,In_186);
or U1269 (N_1269,N_519,N_100);
nor U1270 (N_1270,In_1268,In_2803);
xnor U1271 (N_1271,N_1020,N_193);
nand U1272 (N_1272,N_912,In_1576);
or U1273 (N_1273,In_1748,N_203);
nand U1274 (N_1274,In_1790,N_1040);
nor U1275 (N_1275,N_539,In_848);
or U1276 (N_1276,In_167,In_1090);
nand U1277 (N_1277,N_661,In_1449);
nor U1278 (N_1278,In_499,N_690);
or U1279 (N_1279,In_2275,In_165);
nand U1280 (N_1280,In_2576,N_1039);
nor U1281 (N_1281,In_943,N_350);
and U1282 (N_1282,In_2575,In_2737);
nor U1283 (N_1283,N_452,N_612);
nor U1284 (N_1284,In_813,In_56);
or U1285 (N_1285,In_569,N_584);
or U1286 (N_1286,N_657,N_915);
or U1287 (N_1287,In_1354,In_545);
xor U1288 (N_1288,N_438,In_1435);
nand U1289 (N_1289,N_976,In_2101);
nor U1290 (N_1290,In_1584,In_954);
and U1291 (N_1291,In_263,N_231);
and U1292 (N_1292,In_414,N_731);
xnor U1293 (N_1293,N_400,N_536);
nand U1294 (N_1294,N_995,In_2394);
or U1295 (N_1295,N_1157,N_1088);
or U1296 (N_1296,In_351,In_290);
nand U1297 (N_1297,In_1282,N_611);
nor U1298 (N_1298,N_186,N_83);
nor U1299 (N_1299,N_245,N_967);
nand U1300 (N_1300,In_1915,In_2692);
nor U1301 (N_1301,In_1556,In_2258);
and U1302 (N_1302,In_408,N_680);
and U1303 (N_1303,In_889,In_224);
xor U1304 (N_1304,N_27,In_1839);
xnor U1305 (N_1305,In_863,In_1218);
or U1306 (N_1306,N_468,N_632);
and U1307 (N_1307,N_840,In_829);
and U1308 (N_1308,In_2360,In_2228);
or U1309 (N_1309,In_1523,N_0);
or U1310 (N_1310,In_912,N_908);
xnor U1311 (N_1311,N_988,N_199);
or U1312 (N_1312,N_923,In_2130);
xnor U1313 (N_1313,In_1860,N_993);
nand U1314 (N_1314,N_877,In_2072);
and U1315 (N_1315,In_1359,N_779);
and U1316 (N_1316,In_1082,N_432);
or U1317 (N_1317,In_2494,In_57);
and U1318 (N_1318,In_910,In_1642);
xnor U1319 (N_1319,In_1798,N_1060);
and U1320 (N_1320,In_262,In_2967);
nor U1321 (N_1321,N_959,In_1692);
nand U1322 (N_1322,N_560,In_696);
xor U1323 (N_1323,In_1153,In_1393);
nor U1324 (N_1324,In_139,N_306);
nand U1325 (N_1325,In_26,N_878);
and U1326 (N_1326,In_2459,In_1780);
and U1327 (N_1327,In_2229,N_1048);
and U1328 (N_1328,N_872,N_129);
and U1329 (N_1329,N_629,In_2246);
or U1330 (N_1330,In_455,N_1137);
and U1331 (N_1331,In_1255,In_1032);
nor U1332 (N_1332,N_1141,In_563);
nand U1333 (N_1333,In_1005,N_942);
nor U1334 (N_1334,In_731,N_889);
nor U1335 (N_1335,In_2139,In_2082);
nor U1336 (N_1336,In_831,In_406);
and U1337 (N_1337,N_1080,N_1029);
or U1338 (N_1338,In_1371,N_1117);
nor U1339 (N_1339,In_507,N_746);
xnor U1340 (N_1340,N_943,In_2215);
and U1341 (N_1341,N_749,In_2627);
and U1342 (N_1342,N_622,In_867);
nand U1343 (N_1343,In_1596,In_2122);
nand U1344 (N_1344,N_881,N_1109);
nor U1345 (N_1345,In_1650,N_1032);
and U1346 (N_1346,In_1037,N_922);
or U1347 (N_1347,In_1355,In_2432);
nand U1348 (N_1348,In_2198,N_547);
or U1349 (N_1349,In_2942,N_873);
or U1350 (N_1350,N_1180,N_263);
nand U1351 (N_1351,N_240,N_816);
xor U1352 (N_1352,In_2935,N_861);
and U1353 (N_1353,In_1767,In_1361);
and U1354 (N_1354,N_1077,In_2701);
nor U1355 (N_1355,N_98,In_1931);
or U1356 (N_1356,In_1469,In_2654);
and U1357 (N_1357,N_651,N_1104);
or U1358 (N_1358,N_280,N_105);
xor U1359 (N_1359,In_2317,In_1287);
and U1360 (N_1360,In_490,N_143);
and U1361 (N_1361,N_1153,In_418);
nor U1362 (N_1362,In_1244,In_1317);
or U1363 (N_1363,In_270,In_188);
nand U1364 (N_1364,In_1093,N_728);
nor U1365 (N_1365,N_1127,In_2667);
or U1366 (N_1366,N_890,In_1316);
nor U1367 (N_1367,In_2903,N_642);
and U1368 (N_1368,N_235,In_582);
xnor U1369 (N_1369,In_147,In_239);
or U1370 (N_1370,In_82,In_2030);
xor U1371 (N_1371,N_1150,N_775);
xnor U1372 (N_1372,In_1670,In_816);
and U1373 (N_1373,In_606,In_269);
xor U1374 (N_1374,In_104,In_2760);
and U1375 (N_1375,In_2406,In_857);
and U1376 (N_1376,N_833,In_2300);
nor U1377 (N_1377,In_1982,N_469);
and U1378 (N_1378,N_58,In_572);
nand U1379 (N_1379,N_1144,N_619);
nand U1380 (N_1380,N_463,In_1148);
and U1381 (N_1381,N_511,N_828);
and U1382 (N_1382,In_1157,In_1131);
or U1383 (N_1383,In_2243,N_628);
nor U1384 (N_1384,In_2264,N_37);
and U1385 (N_1385,N_333,N_535);
nand U1386 (N_1386,N_1047,In_1965);
or U1387 (N_1387,In_2951,N_495);
nand U1388 (N_1388,In_1021,N_504);
xnor U1389 (N_1389,In_140,N_673);
and U1390 (N_1390,In_2787,N_721);
nand U1391 (N_1391,In_1100,In_2058);
and U1392 (N_1392,N_418,In_1534);
nor U1393 (N_1393,N_704,In_2423);
nor U1394 (N_1394,In_2953,N_1112);
and U1395 (N_1395,In_708,In_2377);
and U1396 (N_1396,N_846,In_53);
xor U1397 (N_1397,In_687,N_896);
or U1398 (N_1398,In_2609,In_1022);
nor U1399 (N_1399,In_2020,In_1110);
nand U1400 (N_1400,N_855,In_1651);
nor U1401 (N_1401,N_116,N_377);
xnor U1402 (N_1402,N_1036,In_2343);
and U1403 (N_1403,In_440,In_1519);
nor U1404 (N_1404,N_286,N_29);
nand U1405 (N_1405,In_41,In_2224);
nand U1406 (N_1406,N_362,N_1015);
nor U1407 (N_1407,In_1251,In_1998);
and U1408 (N_1408,In_1842,In_1801);
and U1409 (N_1409,N_950,In_2413);
and U1410 (N_1410,N_825,In_1834);
nor U1411 (N_1411,N_939,N_544);
nor U1412 (N_1412,In_1571,N_182);
xor U1413 (N_1413,N_800,In_1820);
nor U1414 (N_1414,In_1977,N_1010);
nor U1415 (N_1415,In_2232,N_502);
and U1416 (N_1416,N_849,In_1414);
xor U1417 (N_1417,In_907,N_853);
nand U1418 (N_1418,In_2757,N_644);
nor U1419 (N_1419,In_2153,N_947);
xor U1420 (N_1420,In_1491,N_928);
xor U1421 (N_1421,In_698,N_277);
xnor U1422 (N_1422,In_926,N_552);
nor U1423 (N_1423,In_2591,In_1327);
nor U1424 (N_1424,N_593,N_88);
nand U1425 (N_1425,In_59,N_1197);
nand U1426 (N_1426,N_308,N_842);
and U1427 (N_1427,In_2000,N_38);
nor U1428 (N_1428,N_667,In_2397);
nand U1429 (N_1429,N_841,N_845);
xnor U1430 (N_1430,N_933,In_961);
nor U1431 (N_1431,In_2849,In_607);
and U1432 (N_1432,In_1331,In_2254);
nor U1433 (N_1433,N_999,N_641);
or U1434 (N_1434,In_1545,N_1134);
nand U1435 (N_1435,In_1818,N_264);
nor U1436 (N_1436,N_697,In_1540);
nor U1437 (N_1437,N_521,In_1419);
xnor U1438 (N_1438,N_513,N_789);
or U1439 (N_1439,In_2912,In_1930);
and U1440 (N_1440,In_1018,N_823);
xor U1441 (N_1441,N_660,In_2363);
nand U1442 (N_1442,In_2727,N_683);
nor U1443 (N_1443,In_18,N_104);
xor U1444 (N_1444,In_1108,N_941);
or U1445 (N_1445,In_353,N_1191);
nor U1446 (N_1446,In_1781,N_64);
nor U1447 (N_1447,In_1959,N_748);
and U1448 (N_1448,N_772,In_308);
xor U1449 (N_1449,N_886,In_858);
nor U1450 (N_1450,N_698,N_763);
xor U1451 (N_1451,N_795,N_678);
nor U1452 (N_1452,In_1370,In_1559);
xor U1453 (N_1453,In_213,In_1006);
xnor U1454 (N_1454,In_340,In_1646);
nor U1455 (N_1455,In_1796,In_1101);
nor U1456 (N_1456,In_158,In_1610);
xnor U1457 (N_1457,In_2042,In_1011);
and U1458 (N_1458,N_1051,In_107);
nand U1459 (N_1459,N_194,In_1677);
or U1460 (N_1460,N_876,In_868);
nand U1461 (N_1461,In_2551,In_360);
nor U1462 (N_1462,In_294,N_770);
xnor U1463 (N_1463,N_603,N_307);
or U1464 (N_1464,In_1683,In_2709);
xor U1465 (N_1465,In_2659,In_463);
xnor U1466 (N_1466,In_444,N_493);
nor U1467 (N_1467,N_1181,N_488);
nand U1468 (N_1468,In_305,N_481);
or U1469 (N_1469,In_2419,N_606);
nor U1470 (N_1470,N_654,N_294);
nand U1471 (N_1471,In_484,In_275);
xnor U1472 (N_1472,N_200,N_794);
nand U1473 (N_1473,In_1989,N_26);
nand U1474 (N_1474,N_436,N_966);
xor U1475 (N_1475,N_157,N_638);
nor U1476 (N_1476,In_637,N_837);
nor U1477 (N_1477,In_1574,N_688);
and U1478 (N_1478,N_712,N_630);
and U1479 (N_1479,N_1106,In_973);
and U1480 (N_1480,In_389,In_409);
or U1481 (N_1481,N_1185,N_978);
nand U1482 (N_1482,In_969,N_847);
nor U1483 (N_1483,In_2952,In_1262);
nor U1484 (N_1484,In_1412,N_1189);
nor U1485 (N_1485,N_1188,In_1602);
and U1486 (N_1486,In_1840,In_1028);
or U1487 (N_1487,N_776,N_1170);
or U1488 (N_1488,In_2170,In_2126);
and U1489 (N_1489,N_931,In_923);
or U1490 (N_1490,N_1093,In_2389);
and U1491 (N_1491,In_1810,In_425);
xor U1492 (N_1492,In_2307,N_827);
and U1493 (N_1493,In_2933,In_2934);
and U1494 (N_1494,N_1034,In_1974);
nand U1495 (N_1495,N_32,N_1079);
nor U1496 (N_1496,In_804,In_655);
nor U1497 (N_1497,In_2209,In_2354);
or U1498 (N_1498,In_27,In_464);
or U1499 (N_1499,N_250,N_285);
nor U1500 (N_1500,In_2110,N_997);
xor U1501 (N_1501,N_72,N_624);
xor U1502 (N_1502,N_664,N_829);
xor U1503 (N_1503,In_934,N_580);
nand U1504 (N_1504,In_1468,N_401);
and U1505 (N_1505,N_45,N_984);
or U1506 (N_1506,In_342,N_190);
and U1507 (N_1507,N_843,N_750);
nand U1508 (N_1508,In_658,In_610);
nand U1509 (N_1509,In_1705,In_2301);
xnor U1510 (N_1510,In_1542,In_380);
and U1511 (N_1511,N_146,N_85);
xnor U1512 (N_1512,In_2699,In_1009);
nor U1513 (N_1513,N_1173,N_574);
nand U1514 (N_1514,In_2632,In_90);
nand U1515 (N_1515,N_119,N_1014);
nor U1516 (N_1516,N_343,In_2370);
nor U1517 (N_1517,In_1276,In_1674);
nor U1518 (N_1518,In_661,N_650);
or U1519 (N_1519,In_1206,In_2973);
xor U1520 (N_1520,In_1452,N_771);
or U1521 (N_1521,In_1895,In_2850);
and U1522 (N_1522,In_2734,In_653);
nand U1523 (N_1523,N_457,In_2434);
nor U1524 (N_1524,N_6,N_1066);
and U1525 (N_1525,In_1290,In_1003);
and U1526 (N_1526,N_982,In_1850);
xor U1527 (N_1527,In_1281,N_700);
and U1528 (N_1528,In_2491,N_860);
and U1529 (N_1529,In_2649,In_2292);
xor U1530 (N_1530,N_499,N_663);
nand U1531 (N_1531,N_1140,In_249);
nor U1532 (N_1532,In_2714,In_1388);
or U1533 (N_1533,N_924,In_39);
nand U1534 (N_1534,N_1151,In_228);
and U1535 (N_1535,N_900,N_1130);
and U1536 (N_1536,N_314,In_1955);
and U1537 (N_1537,In_2577,N_48);
or U1538 (N_1538,In_1661,In_2746);
xor U1539 (N_1539,N_1190,In_1941);
nand U1540 (N_1540,N_737,N_561);
nand U1541 (N_1541,N_1126,In_2310);
xnor U1542 (N_1542,N_289,In_1207);
and U1543 (N_1543,N_117,N_636);
xor U1544 (N_1544,N_627,N_302);
or U1545 (N_1545,N_1178,N_1160);
or U1546 (N_1546,N_617,In_2361);
and U1547 (N_1547,N_446,In_1302);
and U1548 (N_1548,In_1039,N_1161);
nor U1549 (N_1549,In_1225,In_2166);
and U1550 (N_1550,N_719,N_175);
and U1551 (N_1551,In_958,In_776);
nand U1552 (N_1552,N_1090,N_1022);
or U1553 (N_1553,N_769,N_1061);
xor U1554 (N_1554,In_445,In_1897);
nand U1555 (N_1555,N_1046,N_1091);
nor U1556 (N_1556,In_1587,In_767);
or U1557 (N_1557,In_272,In_632);
nand U1558 (N_1558,N_162,N_761);
xor U1559 (N_1559,In_710,In_252);
nor U1560 (N_1560,N_1023,In_2092);
or U1561 (N_1561,In_2557,In_2267);
or U1562 (N_1562,In_1196,N_185);
or U1563 (N_1563,In_2965,N_968);
nor U1564 (N_1564,N_723,In_1809);
and U1565 (N_1565,In_2592,N_368);
nand U1566 (N_1566,In_1945,N_265);
nand U1567 (N_1567,N_859,In_1751);
and U1568 (N_1568,In_195,N_312);
or U1569 (N_1569,N_534,N_936);
and U1570 (N_1570,N_945,N_835);
nor U1571 (N_1571,In_1410,In_942);
nor U1572 (N_1572,N_373,In_521);
or U1573 (N_1573,In_416,In_1104);
xnor U1574 (N_1574,In_1996,In_1450);
and U1575 (N_1575,N_1053,N_485);
nand U1576 (N_1576,In_1482,N_891);
or U1577 (N_1577,N_806,N_195);
nor U1578 (N_1578,In_1012,N_710);
nand U1579 (N_1579,In_146,N_1085);
and U1580 (N_1580,N_410,N_1131);
nor U1581 (N_1581,N_449,N_150);
nand U1582 (N_1582,N_956,N_103);
and U1583 (N_1583,N_753,In_1137);
nor U1584 (N_1584,N_1003,N_57);
xnor U1585 (N_1585,N_691,N_465);
nor U1586 (N_1586,In_2276,N_1124);
or U1587 (N_1587,In_2509,N_986);
or U1588 (N_1588,In_2120,N_382);
or U1589 (N_1589,In_725,N_631);
and U1590 (N_1590,N_1070,In_1507);
and U1591 (N_1591,N_1063,N_1008);
or U1592 (N_1592,In_230,N_940);
nand U1593 (N_1593,N_451,In_1988);
nand U1594 (N_1594,N_715,N_1084);
or U1595 (N_1595,In_1408,In_2970);
nor U1596 (N_1596,In_345,In_1337);
or U1597 (N_1597,In_1958,In_913);
nand U1598 (N_1598,N_545,In_2351);
or U1599 (N_1599,In_559,In_970);
or U1600 (N_1600,In_2698,N_1072);
or U1601 (N_1601,N_898,N_927);
nor U1602 (N_1602,N_273,N_598);
nand U1603 (N_1603,In_2717,In_2927);
nand U1604 (N_1604,N_677,N_221);
or U1605 (N_1605,In_2600,N_990);
nor U1606 (N_1606,N_701,In_2602);
and U1607 (N_1607,N_566,N_883);
nor U1608 (N_1608,N_134,N_635);
or U1609 (N_1609,In_355,N_616);
or U1610 (N_1610,N_1083,In_779);
nor U1611 (N_1611,N_75,In_479);
nand U1612 (N_1612,In_2797,N_17);
and U1613 (N_1613,N_735,N_1012);
xnor U1614 (N_1614,N_1094,In_1771);
or U1615 (N_1615,In_1822,In_915);
nand U1616 (N_1616,N_113,In_618);
nor U1617 (N_1617,N_796,N_695);
and U1618 (N_1618,N_653,N_497);
or U1619 (N_1619,In_352,In_689);
or U1620 (N_1620,N_164,In_1420);
nand U1621 (N_1621,In_2606,In_304);
nor U1622 (N_1622,N_270,N_487);
or U1623 (N_1623,N_998,In_2197);
nor U1624 (N_1624,In_197,N_777);
or U1625 (N_1625,N_756,N_991);
and U1626 (N_1626,N_405,In_2280);
and U1627 (N_1627,N_381,In_1135);
xor U1628 (N_1628,In_441,N_1024);
nand U1629 (N_1629,In_2608,N_345);
nor U1630 (N_1630,In_1340,N_467);
xnor U1631 (N_1631,In_532,N_219);
or U1632 (N_1632,N_658,N_951);
nand U1633 (N_1633,N_1052,In_1263);
or U1634 (N_1634,In_720,N_742);
xnor U1635 (N_1635,N_1027,N_1132);
nand U1636 (N_1636,In_223,N_214);
and U1637 (N_1637,N_246,N_1057);
nor U1638 (N_1638,In_8,N_717);
or U1639 (N_1639,N_139,N_813);
and U1640 (N_1640,In_669,N_332);
xor U1641 (N_1641,In_314,In_1173);
xor U1642 (N_1642,N_850,N_851);
nor U1643 (N_1643,In_491,In_2772);
nand U1644 (N_1644,In_2250,In_1089);
and U1645 (N_1645,In_1199,N_724);
nand U1646 (N_1646,In_1710,N_30);
or U1647 (N_1647,N_838,N_917);
nor U1648 (N_1648,In_2523,In_2490);
or U1649 (N_1649,In_615,N_177);
xor U1650 (N_1650,In_693,In_4);
and U1651 (N_1651,N_1049,N_518);
nand U1652 (N_1652,N_774,N_949);
and U1653 (N_1653,N_1098,N_1167);
and U1654 (N_1654,In_1237,N_819);
xnor U1655 (N_1655,N_744,N_1062);
or U1656 (N_1656,N_15,N_745);
xnor U1657 (N_1657,N_768,N_1045);
nor U1658 (N_1658,In_1401,N_299);
nand U1659 (N_1659,N_894,In_2522);
nand U1660 (N_1660,N_901,In_1916);
or U1661 (N_1661,In_2817,In_1422);
or U1662 (N_1662,In_211,N_1001);
xor U1663 (N_1663,In_1703,In_1776);
nor U1664 (N_1664,N_5,In_2644);
nor U1665 (N_1665,In_2103,In_233);
or U1666 (N_1666,In_2342,In_2977);
nand U1667 (N_1667,N_1009,N_1076);
nand U1668 (N_1668,In_231,N_809);
and U1669 (N_1669,In_1968,In_1720);
nand U1670 (N_1670,N_623,N_613);
or U1671 (N_1671,In_1973,In_2705);
and U1672 (N_1672,In_2032,In_1797);
nand U1673 (N_1673,N_541,In_718);
or U1674 (N_1674,In_526,N_996);
or U1675 (N_1675,In_1782,N_170);
and U1676 (N_1676,In_800,In_2331);
nor U1677 (N_1677,In_1489,In_1726);
or U1678 (N_1678,In_2578,N_810);
or U1679 (N_1679,N_1005,N_787);
nor U1680 (N_1680,In_2334,N_925);
nand U1681 (N_1681,In_2398,In_453);
nand U1682 (N_1682,N_910,N_369);
xor U1683 (N_1683,N_969,N_786);
or U1684 (N_1684,In_1824,In_1913);
and U1685 (N_1685,In_833,In_1511);
xor U1686 (N_1686,In_2339,In_2856);
nand U1687 (N_1687,In_2618,In_2087);
nand U1688 (N_1688,N_1196,N_788);
xnor U1689 (N_1689,N_857,In_1526);
nor U1690 (N_1690,N_965,In_1742);
xnor U1691 (N_1691,In_1956,N_524);
xnor U1692 (N_1692,In_665,In_2768);
nand U1693 (N_1693,In_1917,N_972);
nand U1694 (N_1694,N_1114,N_757);
xnor U1695 (N_1695,In_846,N_921);
and U1696 (N_1696,In_1835,In_1950);
xnor U1697 (N_1697,N_378,N_954);
nor U1698 (N_1698,N_981,N_456);
nand U1699 (N_1699,In_460,N_863);
or U1700 (N_1700,In_2572,In_518);
nand U1701 (N_1701,N_1013,N_138);
and U1702 (N_1702,N_734,N_718);
nand U1703 (N_1703,N_694,N_431);
or U1704 (N_1704,In_2279,In_832);
or U1705 (N_1705,N_681,N_316);
or U1706 (N_1706,N_839,N_803);
nand U1707 (N_1707,In_2918,N_555);
or U1708 (N_1708,In_2713,N_637);
xnor U1709 (N_1709,N_755,In_480);
nand U1710 (N_1710,N_765,In_350);
nor U1711 (N_1711,In_2157,In_313);
and U1712 (N_1712,N_953,In_2615);
and U1713 (N_1713,In_1303,In_2285);
xnor U1714 (N_1714,N_751,N_1087);
or U1715 (N_1715,In_2798,In_2070);
and U1716 (N_1716,In_2770,N_811);
nand U1717 (N_1717,N_605,In_1870);
nor U1718 (N_1718,In_2291,N_1019);
nor U1719 (N_1719,N_283,N_1026);
xor U1720 (N_1720,In_394,In_266);
or U1721 (N_1721,N_1169,In_1711);
nand U1722 (N_1722,In_854,N_670);
or U1723 (N_1723,N_743,In_331);
xor U1724 (N_1724,N_711,N_1166);
and U1725 (N_1725,In_771,N_1175);
nor U1726 (N_1726,In_310,N_836);
and U1727 (N_1727,N_672,N_155);
or U1728 (N_1728,N_884,In_2203);
or U1729 (N_1729,In_2826,In_182);
nand U1730 (N_1730,N_354,N_402);
or U1731 (N_1731,N_707,N_754);
nand U1732 (N_1732,In_1657,N_892);
nand U1733 (N_1733,N_412,N_935);
nand U1734 (N_1734,N_92,In_1553);
nor U1735 (N_1735,In_388,N_610);
nand U1736 (N_1736,In_920,In_2051);
nand U1737 (N_1737,In_2528,N_870);
nor U1738 (N_1738,N_682,N_906);
nand U1739 (N_1739,In_1333,In_91);
nor U1740 (N_1740,In_2450,In_2779);
nor U1741 (N_1741,N_187,In_2161);
nand U1742 (N_1742,N_722,In_1341);
xor U1743 (N_1743,In_2420,In_1057);
xnor U1744 (N_1744,In_1319,N_1165);
nor U1745 (N_1745,N_1171,In_2390);
nor U1746 (N_1746,In_666,N_1174);
or U1747 (N_1747,In_1170,In_1738);
xnor U1748 (N_1748,In_1454,N_331);
nor U1749 (N_1749,N_994,N_223);
xnor U1750 (N_1750,In_1488,In_2993);
xnor U1751 (N_1751,N_189,N_426);
nand U1752 (N_1752,In_2866,N_1069);
or U1753 (N_1753,In_2771,N_1121);
and U1754 (N_1754,N_687,N_975);
xnor U1755 (N_1755,N_897,In_1707);
nor U1756 (N_1756,In_991,N_871);
nand U1757 (N_1757,In_1035,In_956);
xor U1758 (N_1758,In_1871,N_669);
nor U1759 (N_1759,In_1348,In_2754);
or U1760 (N_1760,In_978,N_1176);
and U1761 (N_1761,N_665,In_1434);
or U1762 (N_1762,N_639,N_56);
xnor U1763 (N_1763,In_1429,In_2613);
and U1764 (N_1764,In_2634,N_679);
nor U1765 (N_1765,N_804,In_1779);
or U1766 (N_1766,In_1665,N_609);
xnor U1767 (N_1767,N_720,N_588);
or U1768 (N_1768,N_844,N_254);
nor U1769 (N_1769,In_309,N_699);
and U1770 (N_1770,In_1177,N_486);
or U1771 (N_1771,In_2206,N_1100);
nand U1772 (N_1772,N_726,N_1172);
nor U1773 (N_1773,In_1481,N_1018);
xor U1774 (N_1774,N_708,In_2997);
or U1775 (N_1775,N_895,In_115);
nor U1776 (N_1776,N_808,N_899);
nor U1777 (N_1777,In_939,N_882);
and U1778 (N_1778,In_259,N_93);
nor U1779 (N_1779,N_492,In_2352);
and U1780 (N_1780,N_907,In_1889);
or U1781 (N_1781,N_854,N_338);
or U1782 (N_1782,N_798,N_868);
or U1783 (N_1783,In_2196,N_758);
or U1784 (N_1784,In_2272,N_973);
xnor U1785 (N_1785,N_60,In_2156);
nand U1786 (N_1786,In_797,In_370);
nor U1787 (N_1787,In_1444,In_711);
xnor U1788 (N_1788,N_576,In_2789);
xor U1789 (N_1789,N_590,In_1569);
nor U1790 (N_1790,N_1016,N_344);
and U1791 (N_1791,N_573,In_1869);
xor U1792 (N_1792,N_1183,In_2385);
or U1793 (N_1793,N_1125,N_1102);
nor U1794 (N_1794,In_426,In_1668);
and U1795 (N_1795,In_92,In_2023);
nand U1796 (N_1796,In_536,N_543);
nor U1797 (N_1797,In_1845,N_764);
xnor U1798 (N_1798,N_125,In_2025);
xor U1799 (N_1799,N_762,N_393);
nand U1800 (N_1800,In_2829,N_1143);
nand U1801 (N_1801,N_1735,N_1754);
and U1802 (N_1802,N_79,In_2026);
xnor U1803 (N_1803,N_1477,N_1658);
and U1804 (N_1804,N_1213,N_1260);
and U1805 (N_1805,N_1685,N_1695);
nand U1806 (N_1806,N_506,N_1356);
and U1807 (N_1807,N_1442,N_1757);
xor U1808 (N_1808,N_295,N_741);
nand U1809 (N_1809,N_1352,N_1669);
and U1810 (N_1810,In_1260,N_1119);
or U1811 (N_1811,N_1044,N_1323);
or U1812 (N_1812,In_155,N_1788);
or U1813 (N_1813,In_1270,N_1110);
or U1814 (N_1814,In_629,In_1808);
nor U1815 (N_1815,N_1222,N_1456);
and U1816 (N_1816,N_1766,N_470);
nand U1817 (N_1817,N_388,N_123);
nor U1818 (N_1818,N_1200,In_1628);
and U1819 (N_1819,N_626,N_77);
and U1820 (N_1820,N_1238,N_1711);
nand U1821 (N_1821,N_1455,N_1475);
and U1822 (N_1822,In_362,N_1299);
and U1823 (N_1823,In_1570,N_1116);
or U1824 (N_1824,N_1795,N_1743);
xor U1825 (N_1825,N_1715,N_1778);
nand U1826 (N_1826,N_1496,N_131);
xor U1827 (N_1827,N_1564,N_1306);
nor U1828 (N_1828,In_1514,In_2489);
or U1829 (N_1829,N_1347,N_1082);
or U1830 (N_1830,N_1258,N_1759);
xnor U1831 (N_1831,In_642,N_1350);
and U1832 (N_1832,In_2543,N_1211);
or U1833 (N_1833,N_1679,N_1334);
xor U1834 (N_1834,N_1791,N_1248);
nor U1835 (N_1835,N_1775,N_562);
or U1836 (N_1836,N_1724,In_823);
or U1837 (N_1837,In_474,N_1179);
or U1838 (N_1838,N_920,N_1629);
nor U1839 (N_1839,N_1731,N_1096);
and U1840 (N_1840,N_1291,N_183);
or U1841 (N_1841,N_1635,In_2805);
nand U1842 (N_1842,In_838,N_1302);
nor U1843 (N_1843,N_1610,N_930);
or U1844 (N_1844,N_1276,N_1528);
nand U1845 (N_1845,N_1214,N_39);
nand U1846 (N_1846,N_714,N_184);
nand U1847 (N_1847,In_1342,N_1758);
or U1848 (N_1848,In_2610,N_1220);
and U1849 (N_1849,In_180,In_364);
nor U1850 (N_1850,N_1377,In_949);
and U1851 (N_1851,N_1259,N_1557);
nor U1852 (N_1852,N_1343,N_1483);
nor U1853 (N_1853,N_213,N_621);
nor U1854 (N_1854,N_323,N_1329);
or U1855 (N_1855,N_1623,In_1019);
nor U1856 (N_1856,In_386,N_1753);
nor U1857 (N_1857,N_1453,N_1490);
nor U1858 (N_1858,N_952,N_1750);
and U1859 (N_1859,N_1644,N_1253);
nor U1860 (N_1860,N_1634,N_1529);
or U1861 (N_1861,N_1492,N_196);
or U1862 (N_1862,N_703,In_1430);
nor U1863 (N_1863,N_1544,N_1747);
or U1864 (N_1864,In_52,N_652);
or U1865 (N_1865,In_2857,In_2407);
nand U1866 (N_1866,N_1000,N_478);
nand U1867 (N_1867,In_2682,N_1767);
nand U1868 (N_1868,In_108,N_1493);
or U1869 (N_1869,N_1129,N_929);
nor U1870 (N_1870,N_1043,In_2411);
nor U1871 (N_1871,In_369,N_1355);
xnor U1872 (N_1872,N_205,In_1049);
nand U1873 (N_1873,In_1116,N_1700);
nor U1874 (N_1874,N_1581,N_634);
and U1875 (N_1875,N_1627,In_488);
or U1876 (N_1876,N_1781,N_1502);
nor U1877 (N_1877,In_1219,In_1492);
nor U1878 (N_1878,In_1815,N_1626);
nand U1879 (N_1879,N_1317,N_1463);
xor U1880 (N_1880,N_1338,In_1653);
or U1881 (N_1881,N_370,N_1421);
xnor U1882 (N_1882,In_525,N_1537);
xor U1883 (N_1883,N_736,N_615);
or U1884 (N_1884,N_1381,In_516);
xor U1885 (N_1885,N_1498,N_1384);
nor U1886 (N_1886,N_1727,N_234);
xnor U1887 (N_1887,In_1503,In_234);
nand U1888 (N_1888,N_1774,N_1702);
or U1889 (N_1889,In_1134,In_764);
nor U1890 (N_1890,N_1663,N_1408);
and U1891 (N_1891,N_1748,N_1360);
nand U1892 (N_1892,N_1282,N_1568);
or U1893 (N_1893,In_1293,N_1289);
xor U1894 (N_1894,N_494,N_1136);
nor U1895 (N_1895,N_204,N_1641);
and U1896 (N_1896,N_814,N_1676);
nor U1897 (N_1897,N_1785,In_989);
or U1898 (N_1898,N_1357,In_1666);
nand U1899 (N_1899,N_1570,N_1389);
xor U1900 (N_1900,In_2962,N_1086);
nand U1901 (N_1901,N_1538,N_1501);
nor U1902 (N_1902,In_1205,N_1591);
nand U1903 (N_1903,N_1675,N_875);
xor U1904 (N_1904,N_671,N_1742);
xor U1905 (N_1905,N_1558,N_570);
xnor U1906 (N_1906,In_1614,N_1420);
nand U1907 (N_1907,N_1684,In_419);
nand U1908 (N_1908,N_1726,In_1336);
or U1909 (N_1909,N_313,In_268);
and U1910 (N_1910,N_643,N_1304);
nor U1911 (N_1911,N_1633,N_107);
xnor U1912 (N_1912,In_1639,N_1478);
nand U1913 (N_1913,N_1680,N_1651);
xnor U1914 (N_1914,N_1031,N_1017);
nand U1915 (N_1915,N_1749,N_1733);
nand U1916 (N_1916,In_187,N_99);
and U1917 (N_1917,N_934,N_1278);
or U1918 (N_1918,In_962,N_1670);
nor U1919 (N_1919,In_123,In_1266);
or U1920 (N_1920,N_1553,N_1409);
or U1921 (N_1921,In_1971,N_258);
xor U1922 (N_1922,In_2752,N_1551);
and U1923 (N_1923,N_1321,N_1033);
nand U1924 (N_1924,N_1364,N_1387);
or U1925 (N_1925,N_1092,In_2814);
or U1926 (N_1926,N_1790,N_1257);
nand U1927 (N_1927,N_16,N_1107);
or U1928 (N_1928,N_1438,N_303);
or U1929 (N_1929,In_2719,In_1099);
nand U1930 (N_1930,N_1782,In_1975);
nand U1931 (N_1931,N_1745,N_1552);
nor U1932 (N_1932,N_1432,N_391);
nor U1933 (N_1933,N_1628,In_2066);
xnor U1934 (N_1934,N_604,N_1313);
xor U1935 (N_1935,N_1264,N_1556);
nor U1936 (N_1936,N_1280,N_974);
nor U1937 (N_1937,N_1296,N_1729);
or U1938 (N_1938,N_1097,N_1307);
nand U1939 (N_1939,In_2266,N_1507);
and U1940 (N_1940,N_1513,N_1476);
and U1941 (N_1941,N_1208,In_1772);
nand U1942 (N_1942,N_1430,In_1258);
and U1943 (N_1943,N_1450,N_1740);
nor U1944 (N_1944,N_1607,N_662);
xor U1945 (N_1945,N_685,In_1729);
nor U1946 (N_1946,N_1228,N_1525);
or U1947 (N_1947,N_1373,N_1416);
nand U1948 (N_1948,N_684,N_1674);
xor U1949 (N_1949,N_1325,In_2311);
or U1950 (N_1950,N_1227,N_317);
nor U1951 (N_1951,N_716,N_1439);
nand U1952 (N_1952,N_1598,N_1688);
or U1953 (N_1953,In_1512,N_582);
and U1954 (N_1954,In_1663,In_2383);
nor U1955 (N_1955,N_858,In_2893);
or U1956 (N_1956,N_1630,N_1314);
xor U1957 (N_1957,N_67,N_1667);
and U1958 (N_1958,N_1472,N_1288);
nor U1959 (N_1959,N_1761,N_1569);
nand U1960 (N_1960,N_791,N_1590);
xor U1961 (N_1961,N_376,N_1148);
and U1962 (N_1962,N_602,N_905);
nor U1963 (N_1963,In_236,N_192);
nor U1964 (N_1964,In_897,N_592);
nand U1965 (N_1965,In_2545,N_508);
nand U1966 (N_1966,N_1687,N_1233);
and U1967 (N_1967,N_1369,N_1186);
nand U1968 (N_1968,N_1799,N_1494);
xor U1969 (N_1969,N_805,N_1275);
and U1970 (N_1970,N_1612,N_618);
or U1971 (N_1971,N_902,N_1699);
nor U1972 (N_1972,N_385,N_1194);
nand U1973 (N_1973,N_832,N_1252);
and U1974 (N_1974,N_1520,In_2957);
xnor U1975 (N_1975,In_2834,N_732);
nand U1976 (N_1976,N_1298,N_114);
nand U1977 (N_1977,N_278,N_1366);
or U1978 (N_1978,N_421,N_500);
nand U1979 (N_1979,N_1458,N_964);
nor U1980 (N_1980,In_2063,In_2034);
nand U1981 (N_1981,In_1513,N_379);
or U1982 (N_1982,N_1358,N_797);
xor U1983 (N_1983,N_659,N_1508);
xor U1984 (N_1984,N_1536,N_1187);
and U1985 (N_1985,N_1719,N_1593);
xor U1986 (N_1986,N_1444,N_824);
nor U1987 (N_1987,In_1228,N_1225);
xnor U1988 (N_1988,N_970,N_1504);
nor U1989 (N_1989,N_1054,In_937);
nor U1990 (N_1990,N_1479,N_1301);
and U1991 (N_1991,N_305,In_399);
xnor U1992 (N_1992,N_1489,N_1353);
xnor U1993 (N_1993,N_1466,In_2559);
xnor U1994 (N_1994,N_1696,N_649);
xnor U1995 (N_1995,In_1185,N_1368);
nand U1996 (N_1996,N_1115,In_2662);
or U1997 (N_1997,N_1659,N_729);
xor U1998 (N_1998,N_526,In_286);
and U1999 (N_1999,N_1682,N_1279);
or U2000 (N_2000,In_1722,In_336);
or U2001 (N_2001,N_8,N_1424);
nor U2002 (N_2002,N_1058,In_597);
or U2003 (N_2003,In_977,N_1604);
nor U2004 (N_2004,N_1370,N_1499);
xor U2005 (N_2005,N_1309,N_1293);
nand U2006 (N_2006,N_1707,In_161);
nor U2007 (N_2007,In_997,N_1263);
xor U2008 (N_2008,N_1266,In_578);
nand U2009 (N_2009,N_1269,N_1796);
xnor U2010 (N_2010,N_1155,N_705);
xor U2011 (N_2011,N_1565,N_1485);
and U2012 (N_2012,In_2594,N_1511);
and U2013 (N_2013,N_1336,N_1531);
xor U2014 (N_2014,N_537,In_2201);
xnor U2015 (N_2015,N_1392,N_1500);
xnor U2016 (N_2016,N_1433,N_1237);
or U2017 (N_2017,N_880,N_1789);
or U2018 (N_2018,N_960,In_306);
nor U2019 (N_2019,N_1534,N_1065);
and U2020 (N_2020,N_1595,N_445);
or U2021 (N_2021,N_1464,N_554);
nand U2022 (N_2022,In_118,N_1639);
and U2023 (N_2023,In_984,N_68);
nand U2024 (N_2024,In_1686,N_1717);
nor U2025 (N_2025,N_1240,In_343);
nand U2026 (N_2026,N_1596,In_1716);
nor U2027 (N_2027,N_1561,N_1666);
xnor U2028 (N_2028,N_1397,N_1541);
nand U2029 (N_2029,N_1539,In_439);
or U2030 (N_2030,N_1524,N_1262);
or U2031 (N_2031,N_783,N_1202);
nor U2032 (N_2032,In_1882,N_1371);
nor U2033 (N_2033,N_208,N_983);
and U2034 (N_2034,N_1467,N_1547);
nand U2035 (N_2035,N_1247,N_1621);
xnor U2036 (N_2036,In_2972,N_1349);
xnor U2037 (N_2037,N_1787,N_1158);
xnor U2038 (N_2038,N_471,N_1756);
or U2039 (N_2039,N_1120,N_1677);
or U2040 (N_2040,In_1525,N_792);
nor U2041 (N_2041,N_1792,N_1075);
nor U2042 (N_2042,N_122,N_1793);
nand U2043 (N_2043,N_1449,N_1650);
or U2044 (N_2044,N_1103,N_1218);
or U2045 (N_2045,N_888,N_1393);
nor U2046 (N_2046,N_1241,N_1391);
and U2047 (N_2047,N_174,N_607);
or U2048 (N_2048,N_1625,In_1096);
or U2049 (N_2049,N_1254,N_1067);
xor U2050 (N_2050,In_2210,In_524);
and U2051 (N_2051,N_1156,In_2284);
or U2052 (N_2052,In_2700,N_1471);
xnor U2053 (N_2053,N_856,N_1705);
nand U2054 (N_2054,N_1798,In_2913);
nand U2055 (N_2055,N_301,N_135);
nor U2056 (N_2056,N_1693,N_1689);
nor U2057 (N_2057,N_1533,N_1770);
nand U2058 (N_2058,N_980,N_1506);
or U2059 (N_2059,In_2844,In_596);
or U2060 (N_2060,N_1580,N_1412);
nand U2061 (N_2061,In_338,In_2982);
and U2062 (N_2062,N_1571,N_1737);
xor U2063 (N_2063,N_1436,N_1209);
and U2064 (N_2064,N_1779,In_1234);
or U2065 (N_2065,In_2117,N_233);
or U2066 (N_2066,N_1021,In_1029);
xnor U2067 (N_2067,N_1710,N_1643);
nor U2068 (N_2068,N_1235,N_496);
and U2069 (N_2069,N_1177,In_1652);
and U2070 (N_2070,N_1562,N_1305);
nor U2071 (N_2071,N_1512,In_1863);
nor U2072 (N_2072,N_390,N_1327);
nor U2073 (N_2073,N_766,In_194);
nor U2074 (N_2074,N_1243,In_1304);
or U2075 (N_2075,N_1422,N_1786);
nor U2076 (N_2076,In_2211,N_1128);
nand U2077 (N_2077,In_2457,N_1540);
nand U2078 (N_2078,In_1876,N_1330);
or U2079 (N_2079,In_1934,In_2008);
and U2080 (N_2080,N_328,In_1095);
nor U2081 (N_2081,N_1193,In_1598);
nor U2082 (N_2082,In_2208,In_2464);
or U2083 (N_2083,In_43,N_674);
and U2084 (N_2084,N_1509,N_292);
nor U2085 (N_2085,N_147,N_1548);
nand U2086 (N_2086,N_1668,N_1256);
nand U2087 (N_2087,N_1671,N_1073);
and U2088 (N_2088,N_1440,In_697);
nor U2089 (N_2089,N_1618,N_73);
and U2090 (N_2090,N_1470,N_1611);
nand U2091 (N_2091,N_1532,N_1741);
nand U2092 (N_2092,N_1772,In_1805);
nand U2093 (N_2093,N_437,In_931);
or U2094 (N_2094,In_1176,N_19);
and U2095 (N_2095,In_575,N_1390);
and U2096 (N_2096,N_1744,In_1321);
xnor U2097 (N_2097,N_1346,In_1235);
nor U2098 (N_2098,N_459,In_2914);
nor U2099 (N_2099,N_1105,N_971);
or U2100 (N_2100,N_1405,In_2936);
xnor U2101 (N_2101,In_1667,N_903);
xor U2102 (N_2102,In_1997,N_725);
xor U2103 (N_2103,In_2237,N_1708);
nor U2104 (N_2104,N_1426,In_154);
nand U2105 (N_2105,In_2478,N_1099);
nand U2106 (N_2106,N_1261,N_1242);
and U2107 (N_2107,N_575,N_1681);
and U2108 (N_2108,N_821,N_1411);
xnor U2109 (N_2109,N_802,N_1441);
nand U2110 (N_2110,N_1543,N_1311);
nor U2111 (N_2111,In_183,In_2261);
or U2112 (N_2112,In_964,N_1376);
or U2113 (N_2113,In_585,N_127);
nor U2114 (N_2114,N_1605,N_479);
nor U2115 (N_2115,N_1510,N_1703);
or U2116 (N_2116,N_1586,N_1122);
and U2117 (N_2117,N_236,N_1763);
xor U2118 (N_2118,N_1443,N_801);
or U2119 (N_2119,N_1584,N_1139);
xnor U2120 (N_2120,N_1686,N_1312);
nor U2121 (N_2121,In_1980,N_1712);
nand U2122 (N_2122,In_2469,N_633);
or U2123 (N_2123,In_113,In_1230);
or U2124 (N_2124,N_1078,N_1035);
nor U2125 (N_2125,In_928,N_820);
nor U2126 (N_2126,N_1704,N_1339);
or U2127 (N_2127,In_1471,N_1481);
and U2128 (N_2128,In_240,In_1814);
nand U2129 (N_2129,In_766,In_856);
xor U2130 (N_2130,N_1515,N_1505);
and U2131 (N_2131,N_7,N_1578);
or U2132 (N_2132,In_2220,N_686);
nand U2133 (N_2133,N_790,N_831);
nor U2134 (N_2134,N_1652,N_529);
nor U2135 (N_2135,N_655,In_255);
nand U2136 (N_2136,N_709,In_2039);
nor U2137 (N_2137,N_1473,In_2851);
xor U2138 (N_2138,N_1324,N_188);
nand U2139 (N_2139,In_1693,N_1713);
nand U2140 (N_2140,N_600,N_1028);
xor U2141 (N_2141,In_556,In_495);
nand U2142 (N_2142,N_1410,N_773);
and U2143 (N_2143,N_1582,In_2356);
or U2144 (N_2144,In_320,In_2647);
xor U2145 (N_2145,N_1162,N_1574);
nor U2146 (N_2146,N_1613,In_2969);
and U2147 (N_2147,N_1270,N_1287);
and U2148 (N_2148,In_1306,N_1435);
nor U2149 (N_2149,N_1230,N_1245);
and U2150 (N_2150,N_1624,N_1217);
nor U2151 (N_2151,In_2813,N_1657);
nor U2152 (N_2152,In_935,N_865);
or U2153 (N_2153,In_608,N_1206);
nand U2154 (N_2154,N_1739,N_1638);
or U2155 (N_2155,N_1589,N_480);
xor U2156 (N_2156,N_1318,N_1056);
nor U2157 (N_2157,In_1349,In_2966);
nand U2158 (N_2158,N_1283,N_1503);
nand U2159 (N_2159,N_225,N_1399);
and U2160 (N_2160,N_1606,In_2160);
xnor U2161 (N_2161,In_1927,N_778);
or U2162 (N_2162,N_781,N_1068);
nor U2163 (N_2163,In_1314,N_848);
or U2164 (N_2164,N_1457,In_2941);
and U2165 (N_2165,In_1672,N_1546);
nor U2166 (N_2166,N_1375,N_1587);
xor U2167 (N_2167,N_1362,N_1723);
nor U2168 (N_2168,In_1074,N_1521);
xor U2169 (N_2169,In_1887,N_300);
and U2170 (N_2170,N_1428,In_979);
xnor U2171 (N_2171,N_1030,N_1760);
xnor U2172 (N_2172,N_938,N_1231);
and U2173 (N_2173,N_1622,N_826);
nor U2174 (N_2174,In_1590,N_1469);
nand U2175 (N_2175,N_913,N_1431);
xnor U2176 (N_2176,N_1404,N_1672);
or U2177 (N_2177,N_1567,In_1746);
and U2178 (N_2178,In_1142,In_1292);
or U2179 (N_2179,In_1399,N_1199);
nor U2180 (N_2180,N_1446,N_216);
nand U2181 (N_2181,N_1284,N_1365);
nand U2182 (N_2182,N_1006,N_1342);
nor U2183 (N_2183,N_926,N_1322);
nand U2184 (N_2184,N_1482,N_1550);
nand U2185 (N_2185,N_1563,In_2271);
and U2186 (N_2186,N_1007,N_62);
xor U2187 (N_2187,N_1461,N_1487);
nor U2188 (N_2188,N_1694,N_1661);
or U2189 (N_2189,N_1542,N_1204);
or U2190 (N_2190,N_1219,N_1691);
nand U2191 (N_2191,N_1718,In_1532);
or U2192 (N_2192,In_2133,N_1285);
or U2193 (N_2193,N_1447,In_2108);
nor U2194 (N_2194,N_733,N_1486);
xnor U2195 (N_2195,In_1623,N_510);
or U2196 (N_2196,In_117,In_1922);
and U2197 (N_2197,N_1223,N_1654);
xnor U2198 (N_2198,N_1730,In_1075);
nand U2199 (N_2199,N_1380,In_1732);
nor U2200 (N_2200,In_1538,In_1245);
and U2201 (N_2201,N_1491,N_168);
or U2202 (N_2202,N_1277,N_1769);
and U2203 (N_2203,N_1452,N_693);
nor U2204 (N_2204,N_1328,N_1374);
and U2205 (N_2205,In_2526,N_866);
and U2206 (N_2206,N_1771,N_1768);
nand U2207 (N_2207,N_1720,N_1549);
nor U2208 (N_2208,N_1011,N_1236);
nor U2209 (N_2209,In_87,N_692);
or U2210 (N_2210,N_1514,N_1545);
and U2211 (N_2211,N_1738,N_1265);
and U2212 (N_2212,N_1221,In_1133);
nand U2213 (N_2213,N_1215,In_2290);
nor U2214 (N_2214,N_523,N_1602);
nand U2215 (N_2215,N_118,In_2252);
or U2216 (N_2216,N_879,N_818);
or U2217 (N_2217,N_1272,N_1149);
nor U2218 (N_2218,In_1426,N_1205);
and U2219 (N_2219,N_1560,N_1414);
xnor U2220 (N_2220,N_1319,N_1646);
nor U2221 (N_2221,N_259,N_423);
nor U2222 (N_2222,N_1394,In_2810);
nor U2223 (N_2223,N_668,N_1600);
nand U2224 (N_2224,N_822,N_1454);
nor U2225 (N_2225,N_1614,N_793);
and U2226 (N_2226,N_1752,In_2524);
or U2227 (N_2227,N_1673,In_584);
nand U2228 (N_2228,N_1348,N_599);
nor U2229 (N_2229,N_1794,N_398);
nand U2230 (N_2230,N_752,N_1320);
nor U2231 (N_2231,N_1212,N_1649);
and U2232 (N_2232,In_1689,N_1488);
xnor U2233 (N_2233,N_1619,N_1755);
nor U2234 (N_2234,In_433,N_963);
nor U2235 (N_2235,N_1732,N_1367);
or U2236 (N_2236,N_567,N_1579);
and U2237 (N_2237,N_1239,In_339);
or U2238 (N_2238,N_1555,N_1573);
or U2239 (N_2239,N_1725,N_1337);
nand U2240 (N_2240,N_448,N_1372);
nor U2241 (N_2241,N_1168,N_1300);
nand U2242 (N_2242,N_474,N_1403);
xor U2243 (N_2243,N_1425,N_1519);
and U2244 (N_2244,N_852,N_1396);
nor U2245 (N_2245,N_1697,N_1297);
and U2246 (N_2246,N_167,In_960);
nand U2247 (N_2247,N_1530,N_1734);
xor U2248 (N_2248,N_220,N_1692);
and U2249 (N_2249,N_1645,In_128);
and U2250 (N_2250,N_1229,In_929);
nand U2251 (N_2251,In_2132,In_2968);
or U2252 (N_2252,N_1004,N_1664);
xor U2253 (N_2253,N_958,N_1255);
or U2254 (N_2254,N_249,In_318);
or U2255 (N_2255,N_909,In_1128);
and U2256 (N_2256,N_1575,N_1698);
nand U2257 (N_2257,In_34,N_932);
and U2258 (N_2258,N_918,N_1361);
xnor U2259 (N_2259,N_812,N_1597);
and U2260 (N_2260,N_1388,In_2187);
nand U2261 (N_2261,N_1113,N_461);
or U2262 (N_2262,In_2648,In_482);
and U2263 (N_2263,N_1251,N_1216);
xnor U2264 (N_2264,N_1341,N_1751);
or U2265 (N_2265,N_1273,N_1721);
and U2266 (N_2266,N_955,In_2870);
nor U2267 (N_2267,N_1417,In_2530);
or U2268 (N_2268,N_759,N_1419);
nand U2269 (N_2269,N_256,N_1292);
and U2270 (N_2270,N_957,N_1678);
xor U2271 (N_2271,N_1407,N_1268);
xor U2272 (N_2272,N_1653,N_1303);
or U2273 (N_2273,N_1728,N_1647);
nand U2274 (N_2274,In_1256,In_2474);
nor U2275 (N_2275,In_1595,In_2986);
xnor U2276 (N_2276,In_1097,N_1592);
and U2277 (N_2277,N_1660,N_1648);
nand U2278 (N_2278,In_293,N_1784);
and U2279 (N_2279,N_1326,In_2998);
nand U2280 (N_2280,N_919,N_1655);
xnor U2281 (N_2281,N_946,N_40);
nand U2282 (N_2282,N_1182,In_1216);
nand U2283 (N_2283,In_32,N_517);
nand U2284 (N_2284,N_1451,N_1401);
or U2285 (N_2285,N_1773,N_1386);
nand U2286 (N_2286,N_1345,In_1305);
and U2287 (N_2287,N_1797,N_1516);
xor U2288 (N_2288,N_1354,N_1701);
or U2289 (N_2289,N_985,N_1585);
nor U2290 (N_2290,N_1378,In_2582);
nor U2291 (N_2291,N_944,N_874);
nor U2292 (N_2292,N_1406,N_1429);
xnor U2293 (N_2293,N_482,N_1246);
nor U2294 (N_2294,N_1497,In_319);
or U2295 (N_2295,N_1535,N_1437);
or U2296 (N_2296,N_1783,N_817);
nor U2297 (N_2297,In_980,N_648);
nand U2298 (N_2298,In_472,In_2503);
nor U2299 (N_2299,N_1459,N_1716);
xnor U2300 (N_2300,N_893,N_1722);
and U2301 (N_2301,N_115,N_1640);
xnor U2302 (N_2302,In_1112,In_555);
xnor U2303 (N_2303,N_1777,N_1460);
or U2304 (N_2304,N_1210,N_1316);
and U2305 (N_2305,In_906,N_1274);
xnor U2306 (N_2306,N_1526,N_41);
or U2307 (N_2307,N_1359,N_1468);
xnor U2308 (N_2308,N_1332,N_1495);
nand U2309 (N_2309,N_1038,In_738);
or U2310 (N_2310,N_675,In_1986);
nor U2311 (N_2311,N_1207,N_1637);
xor U2312 (N_2312,N_1527,N_489);
and U2313 (N_2313,N_1142,N_1617);
nand U2314 (N_2314,N_1402,In_1486);
nor U2315 (N_2315,In_2055,In_2329);
xor U2316 (N_2316,N_1413,N_1195);
or U2317 (N_2317,N_1108,N_1434);
xnor U2318 (N_2318,N_640,N_1267);
and U2319 (N_2319,N_1599,N_1331);
nand U2320 (N_2320,N_1423,N_1566);
xor U2321 (N_2321,N_12,In_2332);
or U2322 (N_2322,N_885,N_1295);
or U2323 (N_2323,In_1535,N_1780);
or U2324 (N_2324,N_1465,In_1501);
nand U2325 (N_2325,N_1445,N_1249);
and U2326 (N_2326,In_2534,N_1714);
nand U2327 (N_2327,In_747,In_2497);
nor U2328 (N_2328,N_1290,N_1333);
and U2329 (N_2329,N_1764,N_399);
nor U2330 (N_2330,N_1554,N_347);
nor U2331 (N_2331,In_2917,N_1111);
and U2332 (N_2332,N_1400,N_1615);
xnor U2333 (N_2333,N_1636,In_1002);
xnor U2334 (N_2334,N_992,N_1363);
or U2335 (N_2335,In_105,In_1273);
or U2336 (N_2336,N_1308,In_335);
and U2337 (N_2337,N_1344,N_864);
nand U2338 (N_2338,N_830,In_2486);
xor U2339 (N_2339,N_1577,In_626);
nand U2340 (N_2340,N_834,In_703);
xor U2341 (N_2341,N_1050,N_1765);
xnor U2342 (N_2342,N_1395,In_2347);
or U2343 (N_2343,N_327,In_498);
nand U2344 (N_2344,N_1642,N_1522);
and U2345 (N_2345,N_1631,N_1706);
nand U2346 (N_2346,N_1683,N_1559);
nor U2347 (N_2347,In_1189,N_1418);
xor U2348 (N_2348,N_1517,N_132);
nor U2349 (N_2349,N_515,N_1480);
nor U2350 (N_2350,N_1690,N_1294);
nand U2351 (N_2351,In_242,N_1462);
xnor U2352 (N_2352,N_1762,In_759);
or U2353 (N_2353,N_1340,N_1379);
nor U2354 (N_2354,N_1576,N_656);
nor U2355 (N_2355,In_481,N_1198);
nand U2356 (N_2356,N_1608,N_1594);
xor U2357 (N_2357,N_22,N_335);
nand U2358 (N_2358,N_1609,N_1385);
and U2359 (N_2359,N_1620,N_1656);
nor U2360 (N_2360,N_1234,In_2178);
and U2361 (N_2361,N_1351,N_1665);
or U2362 (N_2362,N_782,N_1281);
or U2363 (N_2363,N_1286,N_594);
nor U2364 (N_2364,N_1448,In_947);
xor U2365 (N_2365,N_1271,N_1583);
and U2366 (N_2366,In_901,In_2655);
nor U2367 (N_2367,N_1383,In_326);
xor U2368 (N_2368,N_1232,In_1357);
and U2369 (N_2369,N_747,N_1226);
or U2370 (N_2370,N_1588,N_601);
nand U2371 (N_2371,N_807,In_952);
nand U2372 (N_2372,N_207,N_1164);
nor U2373 (N_2373,In_638,N_989);
nand U2374 (N_2374,In_461,N_948);
and U2375 (N_2375,N_1632,N_1523);
or U2376 (N_2376,N_1474,In_2155);
xor U2377 (N_2377,N_1601,N_1662);
nor U2378 (N_2378,N_1603,N_1315);
nand U2379 (N_2379,In_2890,N_1736);
xor U2380 (N_2380,N_1224,N_1484);
or U2381 (N_2381,In_1843,N_1203);
nor U2382 (N_2382,N_962,In_1564);
nand U2383 (N_2383,N_1335,N_1572);
nand U2384 (N_2384,N_1518,N_1250);
and U2385 (N_2385,N_1192,In_2929);
xnor U2386 (N_2386,N_1398,N_862);
or U2387 (N_2387,N_1310,N_1709);
and U2388 (N_2388,N_730,In_1102);
xnor U2389 (N_2389,N_1746,N_1776);
and U2390 (N_2390,N_1244,N_739);
xnor U2391 (N_2391,N_815,N_1415);
nor U2392 (N_2392,In_1428,N_1201);
nand U2393 (N_2393,N_1616,N_351);
or U2394 (N_2394,N_1427,N_1382);
nor U2395 (N_2395,In_783,N_1159);
xnor U2396 (N_2396,In_1264,In_1267);
xnor U2397 (N_2397,In_2921,In_2637);
and U2398 (N_2398,N_869,In_2562);
or U2399 (N_2399,In_1502,In_435);
and U2400 (N_2400,N_2289,N_1972);
xnor U2401 (N_2401,N_1808,N_2333);
or U2402 (N_2402,N_1907,N_2164);
nand U2403 (N_2403,N_1878,N_2154);
nor U2404 (N_2404,N_2203,N_2005);
xor U2405 (N_2405,N_2373,N_2184);
nand U2406 (N_2406,N_2023,N_1847);
or U2407 (N_2407,N_2063,N_2363);
nand U2408 (N_2408,N_1855,N_2351);
or U2409 (N_2409,N_2198,N_2220);
xnor U2410 (N_2410,N_2369,N_1897);
nor U2411 (N_2411,N_2194,N_2051);
and U2412 (N_2412,N_2045,N_2152);
nand U2413 (N_2413,N_2179,N_2095);
nand U2414 (N_2414,N_2276,N_2293);
nand U2415 (N_2415,N_2034,N_2271);
nand U2416 (N_2416,N_2167,N_2129);
and U2417 (N_2417,N_2102,N_2116);
nor U2418 (N_2418,N_2245,N_1813);
and U2419 (N_2419,N_1862,N_2089);
and U2420 (N_2420,N_2191,N_1900);
xnor U2421 (N_2421,N_1964,N_1817);
nor U2422 (N_2422,N_2066,N_1837);
xnor U2423 (N_2423,N_2026,N_2357);
xnor U2424 (N_2424,N_2285,N_2278);
or U2425 (N_2425,N_2071,N_1903);
nand U2426 (N_2426,N_2320,N_2170);
or U2427 (N_2427,N_2042,N_2379);
xnor U2428 (N_2428,N_2321,N_1984);
nand U2429 (N_2429,N_2099,N_2027);
and U2430 (N_2430,N_2368,N_1927);
or U2431 (N_2431,N_2165,N_2061);
nand U2432 (N_2432,N_2062,N_2308);
nand U2433 (N_2433,N_2094,N_2145);
or U2434 (N_2434,N_2262,N_1871);
and U2435 (N_2435,N_2228,N_2181);
nor U2436 (N_2436,N_1938,N_2134);
nand U2437 (N_2437,N_2012,N_2307);
xor U2438 (N_2438,N_2113,N_2097);
xor U2439 (N_2439,N_1835,N_2013);
xnor U2440 (N_2440,N_1844,N_2079);
and U2441 (N_2441,N_1962,N_2038);
nand U2442 (N_2442,N_1956,N_2234);
and U2443 (N_2443,N_1807,N_1821);
nor U2444 (N_2444,N_2310,N_2052);
and U2445 (N_2445,N_2033,N_2081);
nor U2446 (N_2446,N_2330,N_2139);
and U2447 (N_2447,N_2096,N_2201);
nor U2448 (N_2448,N_1815,N_2117);
xnor U2449 (N_2449,N_1993,N_1830);
nor U2450 (N_2450,N_2315,N_2016);
xnor U2451 (N_2451,N_2252,N_2190);
and U2452 (N_2452,N_1831,N_2270);
and U2453 (N_2453,N_1905,N_1967);
or U2454 (N_2454,N_1850,N_2173);
and U2455 (N_2455,N_2107,N_2251);
or U2456 (N_2456,N_2003,N_2207);
nor U2457 (N_2457,N_1805,N_2199);
nor U2458 (N_2458,N_1978,N_1969);
nor U2459 (N_2459,N_2290,N_1932);
or U2460 (N_2460,N_2312,N_2223);
nor U2461 (N_2461,N_2339,N_2215);
and U2462 (N_2462,N_1886,N_1985);
xnor U2463 (N_2463,N_1957,N_2280);
or U2464 (N_2464,N_2247,N_2160);
xor U2465 (N_2465,N_2316,N_2216);
nor U2466 (N_2466,N_2058,N_1914);
xor U2467 (N_2467,N_2273,N_1874);
nand U2468 (N_2468,N_2287,N_2159);
or U2469 (N_2469,N_1823,N_2263);
or U2470 (N_2470,N_2070,N_1864);
nand U2471 (N_2471,N_2233,N_1918);
nand U2472 (N_2472,N_2187,N_2153);
and U2473 (N_2473,N_1877,N_2031);
nand U2474 (N_2474,N_2217,N_1977);
or U2475 (N_2475,N_2317,N_2246);
nand U2476 (N_2476,N_1802,N_1951);
nand U2477 (N_2477,N_1992,N_2382);
or U2478 (N_2478,N_2327,N_2050);
xnor U2479 (N_2479,N_1856,N_2225);
and U2480 (N_2480,N_2200,N_2142);
and U2481 (N_2481,N_1942,N_2298);
xnor U2482 (N_2482,N_1888,N_2296);
nor U2483 (N_2483,N_1820,N_2218);
and U2484 (N_2484,N_1987,N_2349);
or U2485 (N_2485,N_2390,N_2162);
xnor U2486 (N_2486,N_2137,N_2323);
nor U2487 (N_2487,N_1828,N_2021);
xnor U2488 (N_2488,N_2185,N_2178);
nor U2489 (N_2489,N_1958,N_2138);
or U2490 (N_2490,N_1960,N_2224);
xor U2491 (N_2491,N_2146,N_2014);
xnor U2492 (N_2492,N_1902,N_2073);
xor U2493 (N_2493,N_1885,N_2020);
and U2494 (N_2494,N_1946,N_2255);
and U2495 (N_2495,N_2193,N_2337);
nor U2496 (N_2496,N_1843,N_2334);
or U2497 (N_2497,N_2221,N_2157);
nand U2498 (N_2498,N_2105,N_1804);
and U2499 (N_2499,N_1838,N_1944);
nor U2500 (N_2500,N_2158,N_1822);
or U2501 (N_2501,N_2206,N_2074);
nor U2502 (N_2502,N_2143,N_1814);
xnor U2503 (N_2503,N_2387,N_2300);
and U2504 (N_2504,N_2378,N_2318);
and U2505 (N_2505,N_1827,N_1923);
or U2506 (N_2506,N_2226,N_2366);
xor U2507 (N_2507,N_1916,N_2098);
nor U2508 (N_2508,N_2001,N_1806);
nor U2509 (N_2509,N_1921,N_2056);
and U2510 (N_2510,N_1858,N_1935);
or U2511 (N_2511,N_2172,N_2186);
or U2512 (N_2512,N_1895,N_2305);
xnor U2513 (N_2513,N_2077,N_2384);
nand U2514 (N_2514,N_2135,N_1928);
and U2515 (N_2515,N_1976,N_2344);
nand U2516 (N_2516,N_1904,N_1950);
nor U2517 (N_2517,N_1968,N_1981);
or U2518 (N_2518,N_2332,N_1997);
nor U2519 (N_2519,N_2261,N_2372);
nand U2520 (N_2520,N_2037,N_2303);
or U2521 (N_2521,N_1911,N_2364);
or U2522 (N_2522,N_2044,N_2377);
or U2523 (N_2523,N_2248,N_1970);
nand U2524 (N_2524,N_2313,N_2018);
xor U2525 (N_2525,N_2359,N_2348);
xnor U2526 (N_2526,N_2314,N_1999);
or U2527 (N_2527,N_1873,N_1833);
or U2528 (N_2528,N_1990,N_2189);
xor U2529 (N_2529,N_2171,N_1824);
nor U2530 (N_2530,N_2028,N_2163);
nand U2531 (N_2531,N_1979,N_2148);
nand U2532 (N_2532,N_2385,N_2370);
nor U2533 (N_2533,N_2072,N_2383);
xnor U2534 (N_2534,N_1819,N_2115);
xor U2535 (N_2535,N_1860,N_1901);
xnor U2536 (N_2536,N_2149,N_2010);
nand U2537 (N_2537,N_1925,N_1961);
xor U2538 (N_2538,N_1915,N_2168);
and U2539 (N_2539,N_1971,N_2029);
nor U2540 (N_2540,N_1879,N_2268);
nand U2541 (N_2541,N_2264,N_1883);
xnor U2542 (N_2542,N_2078,N_2202);
and U2543 (N_2543,N_1834,N_2030);
and U2544 (N_2544,N_2311,N_2043);
nand U2545 (N_2545,N_2294,N_2389);
and U2546 (N_2546,N_2241,N_2249);
xnor U2547 (N_2547,N_2182,N_2120);
xor U2548 (N_2548,N_1913,N_2108);
xor U2549 (N_2549,N_2101,N_1924);
nand U2550 (N_2550,N_2065,N_2125);
xor U2551 (N_2551,N_1800,N_2331);
and U2552 (N_2552,N_2046,N_2068);
or U2553 (N_2553,N_2324,N_2150);
or U2554 (N_2554,N_2002,N_2380);
and U2555 (N_2555,N_2269,N_2151);
or U2556 (N_2556,N_1842,N_1892);
or U2557 (N_2557,N_2000,N_1832);
xnor U2558 (N_2558,N_2092,N_1893);
nor U2559 (N_2559,N_2192,N_1943);
nand U2560 (N_2560,N_2292,N_2393);
nor U2561 (N_2561,N_2176,N_2397);
nor U2562 (N_2562,N_2136,N_2110);
and U2563 (N_2563,N_2040,N_1930);
xnor U2564 (N_2564,N_1933,N_1965);
nor U2565 (N_2565,N_2375,N_1884);
nor U2566 (N_2566,N_2242,N_2039);
nor U2567 (N_2567,N_1934,N_1909);
and U2568 (N_2568,N_2286,N_1840);
and U2569 (N_2569,N_2265,N_2231);
nand U2570 (N_2570,N_2212,N_2222);
or U2571 (N_2571,N_2282,N_2067);
xor U2572 (N_2572,N_2362,N_1896);
or U2573 (N_2573,N_1857,N_2253);
and U2574 (N_2574,N_2205,N_2347);
nand U2575 (N_2575,N_2259,N_1975);
nor U2576 (N_2576,N_2007,N_2343);
xnor U2577 (N_2577,N_1917,N_1811);
xnor U2578 (N_2578,N_2376,N_1929);
or U2579 (N_2579,N_2237,N_2360);
and U2580 (N_2580,N_2087,N_2340);
or U2581 (N_2581,N_1863,N_2111);
nand U2582 (N_2582,N_2175,N_2197);
and U2583 (N_2583,N_2085,N_2213);
nor U2584 (N_2584,N_2036,N_2180);
and U2585 (N_2585,N_2121,N_1899);
nand U2586 (N_2586,N_2141,N_1980);
nand U2587 (N_2587,N_1866,N_2283);
or U2588 (N_2588,N_2080,N_2304);
nor U2589 (N_2589,N_2391,N_2358);
nor U2590 (N_2590,N_2024,N_1836);
nor U2591 (N_2591,N_1989,N_1998);
nand U2592 (N_2592,N_2356,N_2353);
nor U2593 (N_2593,N_2183,N_2338);
or U2594 (N_2594,N_1949,N_2196);
xnor U2595 (N_2595,N_1829,N_2302);
nand U2596 (N_2596,N_2124,N_2133);
nand U2597 (N_2597,N_2100,N_1880);
or U2598 (N_2598,N_1891,N_2301);
nor U2599 (N_2599,N_2188,N_2035);
nor U2600 (N_2600,N_1996,N_2395);
nor U2601 (N_2601,N_2250,N_2214);
xor U2602 (N_2602,N_1941,N_2341);
xnor U2603 (N_2603,N_1955,N_2367);
and U2604 (N_2604,N_2104,N_1849);
nand U2605 (N_2605,N_2309,N_1887);
or U2606 (N_2606,N_1825,N_2054);
and U2607 (N_2607,N_2156,N_2335);
and U2608 (N_2608,N_2266,N_2239);
nand U2609 (N_2609,N_1991,N_2230);
nor U2610 (N_2610,N_2392,N_1846);
and U2611 (N_2611,N_1926,N_2049);
nor U2612 (N_2612,N_1851,N_1910);
xnor U2613 (N_2613,N_1974,N_1859);
xnor U2614 (N_2614,N_2281,N_2275);
or U2615 (N_2615,N_2048,N_2090);
and U2616 (N_2616,N_2254,N_2106);
xor U2617 (N_2617,N_1810,N_1845);
nand U2618 (N_2618,N_2279,N_1939);
and U2619 (N_2619,N_1853,N_1931);
nor U2620 (N_2620,N_1912,N_2082);
and U2621 (N_2621,N_2060,N_1936);
xnor U2622 (N_2622,N_2386,N_1945);
xnor U2623 (N_2623,N_1890,N_2299);
and U2624 (N_2624,N_1865,N_1963);
xnor U2625 (N_2625,N_1983,N_2346);
xor U2626 (N_2626,N_2277,N_2064);
nor U2627 (N_2627,N_2004,N_1852);
nand U2628 (N_2628,N_2329,N_2238);
nand U2629 (N_2629,N_2122,N_2053);
nand U2630 (N_2630,N_2227,N_1812);
xnor U2631 (N_2631,N_2174,N_1986);
nand U2632 (N_2632,N_2126,N_2144);
xnor U2633 (N_2633,N_2019,N_2394);
nor U2634 (N_2634,N_1994,N_1867);
nand U2635 (N_2635,N_1882,N_2345);
or U2636 (N_2636,N_2244,N_1816);
nor U2637 (N_2637,N_2272,N_2009);
or U2638 (N_2638,N_2008,N_1919);
nor U2639 (N_2639,N_2209,N_2088);
nor U2640 (N_2640,N_1875,N_2059);
and U2641 (N_2641,N_2119,N_1937);
xnor U2642 (N_2642,N_1841,N_2161);
xor U2643 (N_2643,N_2295,N_2219);
nor U2644 (N_2644,N_1872,N_2123);
xor U2645 (N_2645,N_2155,N_2083);
xnor U2646 (N_2646,N_1898,N_1868);
nor U2647 (N_2647,N_1948,N_1848);
nor U2648 (N_2648,N_1947,N_2328);
and U2649 (N_2649,N_2118,N_2130);
nor U2650 (N_2650,N_1826,N_2006);
nand U2651 (N_2651,N_2075,N_2256);
xnor U2652 (N_2652,N_2204,N_2232);
or U2653 (N_2653,N_2131,N_2210);
and U2654 (N_2654,N_1809,N_2211);
or U2655 (N_2655,N_1988,N_1995);
or U2656 (N_2656,N_2326,N_2169);
or U2657 (N_2657,N_1894,N_2235);
and U2658 (N_2658,N_1906,N_1940);
xnor U2659 (N_2659,N_2274,N_2022);
xnor U2660 (N_2660,N_2288,N_2147);
xor U2661 (N_2661,N_2091,N_2381);
xnor U2662 (N_2662,N_2396,N_2195);
xnor U2663 (N_2663,N_2355,N_2055);
or U2664 (N_2664,N_1966,N_2127);
xor U2665 (N_2665,N_2297,N_1870);
or U2666 (N_2666,N_2374,N_1953);
xor U2667 (N_2667,N_2365,N_1881);
nor U2668 (N_2668,N_2140,N_2011);
nor U2669 (N_2669,N_2257,N_2258);
or U2670 (N_2670,N_2015,N_2086);
and U2671 (N_2671,N_2032,N_1869);
nand U2672 (N_2672,N_2291,N_2319);
and U2673 (N_2673,N_1908,N_1803);
nand U2674 (N_2674,N_1959,N_2371);
nor U2675 (N_2675,N_2076,N_2166);
or U2676 (N_2676,N_2025,N_1973);
nand U2677 (N_2677,N_2354,N_2399);
nor U2678 (N_2678,N_1920,N_2114);
or U2679 (N_2679,N_2112,N_2236);
xnor U2680 (N_2680,N_2267,N_2084);
and U2681 (N_2681,N_2240,N_2306);
and U2682 (N_2682,N_1861,N_1952);
nand U2683 (N_2683,N_1801,N_2229);
xnor U2684 (N_2684,N_2350,N_2069);
and U2685 (N_2685,N_2128,N_2284);
nor U2686 (N_2686,N_2017,N_2132);
nor U2687 (N_2687,N_2398,N_1982);
nor U2688 (N_2688,N_1922,N_2361);
nor U2689 (N_2689,N_2342,N_2336);
nand U2690 (N_2690,N_2057,N_1954);
or U2691 (N_2691,N_2208,N_2322);
and U2692 (N_2692,N_1854,N_1839);
and U2693 (N_2693,N_1889,N_2388);
nand U2694 (N_2694,N_2041,N_2260);
and U2695 (N_2695,N_2243,N_1818);
nor U2696 (N_2696,N_2352,N_2093);
xnor U2697 (N_2697,N_2177,N_2103);
nand U2698 (N_2698,N_2109,N_2325);
or U2699 (N_2699,N_2047,N_1876);
nor U2700 (N_2700,N_1984,N_1983);
or U2701 (N_2701,N_1910,N_2010);
nand U2702 (N_2702,N_2309,N_2278);
xor U2703 (N_2703,N_2260,N_1960);
xnor U2704 (N_2704,N_1878,N_2380);
and U2705 (N_2705,N_2235,N_2175);
nand U2706 (N_2706,N_1903,N_2305);
xnor U2707 (N_2707,N_2035,N_1833);
and U2708 (N_2708,N_2045,N_2231);
nand U2709 (N_2709,N_2250,N_2103);
or U2710 (N_2710,N_2340,N_1977);
and U2711 (N_2711,N_1832,N_2025);
and U2712 (N_2712,N_1963,N_2331);
and U2713 (N_2713,N_2305,N_1933);
or U2714 (N_2714,N_2214,N_1880);
nor U2715 (N_2715,N_2357,N_2358);
nand U2716 (N_2716,N_2168,N_2163);
or U2717 (N_2717,N_1854,N_2023);
nand U2718 (N_2718,N_1833,N_2334);
xnor U2719 (N_2719,N_1840,N_2241);
or U2720 (N_2720,N_2046,N_2027);
nand U2721 (N_2721,N_1881,N_2330);
nand U2722 (N_2722,N_2304,N_1965);
xor U2723 (N_2723,N_2325,N_1861);
and U2724 (N_2724,N_2097,N_2041);
nand U2725 (N_2725,N_2076,N_2365);
nor U2726 (N_2726,N_1963,N_2095);
or U2727 (N_2727,N_1994,N_2348);
nor U2728 (N_2728,N_2027,N_1973);
nand U2729 (N_2729,N_2314,N_1891);
or U2730 (N_2730,N_1959,N_1802);
nand U2731 (N_2731,N_1887,N_2272);
or U2732 (N_2732,N_2200,N_2031);
or U2733 (N_2733,N_2369,N_2165);
and U2734 (N_2734,N_2332,N_2126);
and U2735 (N_2735,N_2324,N_2173);
or U2736 (N_2736,N_2126,N_1929);
or U2737 (N_2737,N_2077,N_2390);
nor U2738 (N_2738,N_1946,N_2284);
nor U2739 (N_2739,N_2217,N_1973);
and U2740 (N_2740,N_2328,N_1939);
or U2741 (N_2741,N_2348,N_1881);
nor U2742 (N_2742,N_2085,N_2353);
nor U2743 (N_2743,N_2245,N_2142);
and U2744 (N_2744,N_1858,N_1902);
xnor U2745 (N_2745,N_2256,N_1973);
and U2746 (N_2746,N_1810,N_2090);
nor U2747 (N_2747,N_2160,N_2171);
nand U2748 (N_2748,N_2322,N_2168);
nor U2749 (N_2749,N_2099,N_2341);
nand U2750 (N_2750,N_1974,N_1936);
nand U2751 (N_2751,N_2224,N_2169);
nor U2752 (N_2752,N_2389,N_2218);
or U2753 (N_2753,N_2183,N_2299);
nor U2754 (N_2754,N_2256,N_2107);
nor U2755 (N_2755,N_1851,N_2222);
nor U2756 (N_2756,N_2093,N_2161);
xnor U2757 (N_2757,N_2054,N_2231);
and U2758 (N_2758,N_2301,N_1879);
xnor U2759 (N_2759,N_1805,N_1917);
or U2760 (N_2760,N_2288,N_2113);
and U2761 (N_2761,N_2089,N_2062);
xnor U2762 (N_2762,N_1942,N_2358);
or U2763 (N_2763,N_2392,N_1812);
and U2764 (N_2764,N_2208,N_2329);
or U2765 (N_2765,N_2178,N_2396);
and U2766 (N_2766,N_2329,N_2397);
and U2767 (N_2767,N_2239,N_2137);
nor U2768 (N_2768,N_2061,N_2030);
xnor U2769 (N_2769,N_2158,N_2183);
xnor U2770 (N_2770,N_2011,N_2251);
and U2771 (N_2771,N_1978,N_2045);
nand U2772 (N_2772,N_2104,N_2002);
nand U2773 (N_2773,N_1839,N_1838);
or U2774 (N_2774,N_1901,N_2390);
nor U2775 (N_2775,N_1845,N_2028);
nand U2776 (N_2776,N_1855,N_1801);
nor U2777 (N_2777,N_1975,N_2383);
xnor U2778 (N_2778,N_2121,N_2107);
nor U2779 (N_2779,N_2173,N_2012);
or U2780 (N_2780,N_1831,N_2192);
xor U2781 (N_2781,N_1874,N_2196);
and U2782 (N_2782,N_2178,N_1971);
xnor U2783 (N_2783,N_2247,N_2131);
and U2784 (N_2784,N_2028,N_1990);
and U2785 (N_2785,N_2208,N_1927);
or U2786 (N_2786,N_2052,N_2255);
and U2787 (N_2787,N_1866,N_2379);
and U2788 (N_2788,N_1992,N_2379);
and U2789 (N_2789,N_1923,N_2121);
or U2790 (N_2790,N_2112,N_2008);
nand U2791 (N_2791,N_1971,N_1932);
or U2792 (N_2792,N_1842,N_1831);
or U2793 (N_2793,N_1916,N_1925);
nand U2794 (N_2794,N_2114,N_2090);
nor U2795 (N_2795,N_2229,N_1956);
nor U2796 (N_2796,N_2050,N_2133);
or U2797 (N_2797,N_2248,N_1897);
or U2798 (N_2798,N_2067,N_2360);
xnor U2799 (N_2799,N_2235,N_1880);
and U2800 (N_2800,N_2021,N_2161);
nor U2801 (N_2801,N_2292,N_2357);
xnor U2802 (N_2802,N_2234,N_1845);
nor U2803 (N_2803,N_1903,N_1965);
and U2804 (N_2804,N_2153,N_1893);
nand U2805 (N_2805,N_1869,N_1868);
or U2806 (N_2806,N_2060,N_2251);
and U2807 (N_2807,N_2197,N_2155);
nor U2808 (N_2808,N_2074,N_2224);
nand U2809 (N_2809,N_2057,N_1869);
xor U2810 (N_2810,N_2053,N_2252);
and U2811 (N_2811,N_2346,N_1932);
nor U2812 (N_2812,N_1834,N_1953);
nand U2813 (N_2813,N_1859,N_2041);
or U2814 (N_2814,N_1888,N_1947);
nand U2815 (N_2815,N_2352,N_2356);
and U2816 (N_2816,N_1994,N_1992);
or U2817 (N_2817,N_2324,N_1945);
or U2818 (N_2818,N_2040,N_2047);
or U2819 (N_2819,N_2316,N_2205);
and U2820 (N_2820,N_1875,N_1963);
and U2821 (N_2821,N_1844,N_2247);
nor U2822 (N_2822,N_1832,N_1856);
nor U2823 (N_2823,N_2320,N_2363);
xnor U2824 (N_2824,N_2210,N_1953);
or U2825 (N_2825,N_2329,N_2361);
and U2826 (N_2826,N_2059,N_2297);
xor U2827 (N_2827,N_2080,N_2039);
or U2828 (N_2828,N_2087,N_1859);
nor U2829 (N_2829,N_1807,N_2399);
or U2830 (N_2830,N_2330,N_2208);
or U2831 (N_2831,N_1930,N_2167);
nor U2832 (N_2832,N_1895,N_2111);
nor U2833 (N_2833,N_2203,N_1881);
nand U2834 (N_2834,N_1974,N_2217);
nor U2835 (N_2835,N_2228,N_2337);
nand U2836 (N_2836,N_2318,N_1989);
nor U2837 (N_2837,N_2217,N_2322);
xor U2838 (N_2838,N_2235,N_1951);
nand U2839 (N_2839,N_2366,N_1955);
and U2840 (N_2840,N_2268,N_2369);
nand U2841 (N_2841,N_2261,N_2060);
or U2842 (N_2842,N_2124,N_2102);
xor U2843 (N_2843,N_2238,N_2363);
or U2844 (N_2844,N_1956,N_2335);
and U2845 (N_2845,N_1892,N_1818);
or U2846 (N_2846,N_2126,N_2308);
or U2847 (N_2847,N_2140,N_2326);
and U2848 (N_2848,N_1822,N_2012);
nand U2849 (N_2849,N_2237,N_2076);
or U2850 (N_2850,N_1891,N_1832);
and U2851 (N_2851,N_2222,N_2237);
nand U2852 (N_2852,N_2288,N_2262);
xor U2853 (N_2853,N_1838,N_2250);
nor U2854 (N_2854,N_2048,N_1992);
xnor U2855 (N_2855,N_2192,N_2232);
nand U2856 (N_2856,N_2044,N_2234);
nand U2857 (N_2857,N_2051,N_2036);
nor U2858 (N_2858,N_2058,N_2084);
and U2859 (N_2859,N_2277,N_2099);
or U2860 (N_2860,N_1925,N_2176);
xor U2861 (N_2861,N_1890,N_2149);
or U2862 (N_2862,N_2209,N_2213);
xnor U2863 (N_2863,N_1991,N_1828);
or U2864 (N_2864,N_2316,N_1800);
or U2865 (N_2865,N_2182,N_2298);
or U2866 (N_2866,N_1806,N_2129);
and U2867 (N_2867,N_2399,N_1996);
xor U2868 (N_2868,N_2075,N_1905);
or U2869 (N_2869,N_2283,N_2030);
nor U2870 (N_2870,N_1977,N_2171);
and U2871 (N_2871,N_2108,N_1905);
nor U2872 (N_2872,N_2280,N_1855);
or U2873 (N_2873,N_1858,N_2115);
and U2874 (N_2874,N_2118,N_1898);
and U2875 (N_2875,N_2279,N_2333);
or U2876 (N_2876,N_2345,N_2106);
xnor U2877 (N_2877,N_2379,N_1841);
xor U2878 (N_2878,N_1985,N_2184);
nor U2879 (N_2879,N_1866,N_1908);
and U2880 (N_2880,N_2099,N_2367);
nor U2881 (N_2881,N_2371,N_1873);
nand U2882 (N_2882,N_2151,N_1979);
xor U2883 (N_2883,N_2248,N_2014);
nor U2884 (N_2884,N_2340,N_1878);
and U2885 (N_2885,N_1975,N_1935);
xor U2886 (N_2886,N_1857,N_1919);
nand U2887 (N_2887,N_2277,N_1841);
and U2888 (N_2888,N_1899,N_2136);
and U2889 (N_2889,N_2186,N_1890);
xnor U2890 (N_2890,N_2082,N_2266);
or U2891 (N_2891,N_2319,N_2233);
or U2892 (N_2892,N_2023,N_2263);
and U2893 (N_2893,N_2128,N_2240);
or U2894 (N_2894,N_2296,N_2342);
and U2895 (N_2895,N_2325,N_2343);
xor U2896 (N_2896,N_2090,N_2343);
or U2897 (N_2897,N_2210,N_2348);
or U2898 (N_2898,N_1862,N_2224);
nor U2899 (N_2899,N_2337,N_2241);
nor U2900 (N_2900,N_2084,N_2306);
xor U2901 (N_2901,N_1868,N_1845);
nand U2902 (N_2902,N_1985,N_2075);
nor U2903 (N_2903,N_1907,N_1929);
nand U2904 (N_2904,N_2266,N_1972);
nor U2905 (N_2905,N_2236,N_1889);
nand U2906 (N_2906,N_2375,N_2061);
or U2907 (N_2907,N_1929,N_2112);
xor U2908 (N_2908,N_1803,N_1857);
xnor U2909 (N_2909,N_2148,N_1965);
xor U2910 (N_2910,N_1909,N_1835);
or U2911 (N_2911,N_2386,N_2355);
or U2912 (N_2912,N_1984,N_1838);
nand U2913 (N_2913,N_1989,N_1804);
xnor U2914 (N_2914,N_2271,N_2128);
xor U2915 (N_2915,N_2159,N_2151);
or U2916 (N_2916,N_1873,N_2206);
nand U2917 (N_2917,N_1846,N_2090);
xor U2918 (N_2918,N_2174,N_2130);
xnor U2919 (N_2919,N_2080,N_2302);
and U2920 (N_2920,N_2022,N_1904);
nand U2921 (N_2921,N_2101,N_2363);
or U2922 (N_2922,N_2387,N_2389);
nor U2923 (N_2923,N_2150,N_2247);
xor U2924 (N_2924,N_2252,N_2316);
nor U2925 (N_2925,N_1902,N_2168);
xnor U2926 (N_2926,N_2061,N_2351);
and U2927 (N_2927,N_2030,N_1849);
nand U2928 (N_2928,N_1921,N_2315);
or U2929 (N_2929,N_1995,N_2134);
nand U2930 (N_2930,N_1841,N_1911);
nand U2931 (N_2931,N_2326,N_1978);
xnor U2932 (N_2932,N_1838,N_2297);
nor U2933 (N_2933,N_1804,N_2346);
or U2934 (N_2934,N_2065,N_2100);
xor U2935 (N_2935,N_2138,N_1849);
and U2936 (N_2936,N_2056,N_2220);
nand U2937 (N_2937,N_2047,N_2059);
nand U2938 (N_2938,N_2142,N_2154);
or U2939 (N_2939,N_1823,N_2369);
xnor U2940 (N_2940,N_2366,N_1945);
and U2941 (N_2941,N_2035,N_1990);
and U2942 (N_2942,N_2081,N_2063);
nand U2943 (N_2943,N_1836,N_2041);
and U2944 (N_2944,N_2219,N_2130);
nor U2945 (N_2945,N_1848,N_1976);
or U2946 (N_2946,N_1891,N_2308);
nand U2947 (N_2947,N_2362,N_2352);
or U2948 (N_2948,N_1818,N_2209);
and U2949 (N_2949,N_2163,N_2206);
and U2950 (N_2950,N_2318,N_2184);
xnor U2951 (N_2951,N_2378,N_2255);
or U2952 (N_2952,N_2261,N_1914);
xnor U2953 (N_2953,N_2269,N_2099);
xnor U2954 (N_2954,N_2000,N_1999);
and U2955 (N_2955,N_1939,N_2271);
xnor U2956 (N_2956,N_2221,N_1935);
nand U2957 (N_2957,N_1830,N_2258);
nor U2958 (N_2958,N_2225,N_2344);
nor U2959 (N_2959,N_1889,N_2310);
xor U2960 (N_2960,N_1852,N_2071);
or U2961 (N_2961,N_2016,N_2280);
nor U2962 (N_2962,N_2048,N_2178);
and U2963 (N_2963,N_2320,N_1914);
and U2964 (N_2964,N_2070,N_2178);
nor U2965 (N_2965,N_2179,N_2397);
xor U2966 (N_2966,N_2399,N_1971);
and U2967 (N_2967,N_2350,N_1969);
nand U2968 (N_2968,N_2166,N_2164);
nor U2969 (N_2969,N_2025,N_1841);
or U2970 (N_2970,N_2187,N_2110);
xor U2971 (N_2971,N_2290,N_2242);
and U2972 (N_2972,N_2154,N_2268);
nand U2973 (N_2973,N_1854,N_1964);
nand U2974 (N_2974,N_2317,N_1801);
xnor U2975 (N_2975,N_1844,N_2043);
nor U2976 (N_2976,N_2202,N_1823);
xnor U2977 (N_2977,N_2223,N_1859);
and U2978 (N_2978,N_1975,N_1852);
or U2979 (N_2979,N_2077,N_1998);
nor U2980 (N_2980,N_2094,N_2081);
and U2981 (N_2981,N_2201,N_1852);
xor U2982 (N_2982,N_2146,N_2229);
or U2983 (N_2983,N_2365,N_2332);
or U2984 (N_2984,N_2359,N_2355);
or U2985 (N_2985,N_2019,N_1990);
nand U2986 (N_2986,N_1967,N_2126);
nor U2987 (N_2987,N_2322,N_2132);
nand U2988 (N_2988,N_2332,N_2239);
and U2989 (N_2989,N_2234,N_2249);
nor U2990 (N_2990,N_2398,N_1833);
and U2991 (N_2991,N_2267,N_1869);
and U2992 (N_2992,N_2025,N_2119);
nor U2993 (N_2993,N_1912,N_2213);
nand U2994 (N_2994,N_2291,N_2210);
nand U2995 (N_2995,N_2054,N_2083);
or U2996 (N_2996,N_1833,N_1889);
or U2997 (N_2997,N_2166,N_2336);
and U2998 (N_2998,N_1942,N_2108);
or U2999 (N_2999,N_2300,N_2277);
or U3000 (N_3000,N_2432,N_2916);
nand U3001 (N_3001,N_2798,N_2549);
nand U3002 (N_3002,N_2438,N_2466);
xnor U3003 (N_3003,N_2627,N_2846);
nand U3004 (N_3004,N_2858,N_2845);
xor U3005 (N_3005,N_2642,N_2987);
xnor U3006 (N_3006,N_2459,N_2476);
nand U3007 (N_3007,N_2494,N_2553);
nand U3008 (N_3008,N_2910,N_2779);
nor U3009 (N_3009,N_2555,N_2656);
and U3010 (N_3010,N_2850,N_2436);
nor U3011 (N_3011,N_2412,N_2733);
or U3012 (N_3012,N_2566,N_2613);
or U3013 (N_3013,N_2948,N_2870);
nand U3014 (N_3014,N_2588,N_2983);
xor U3015 (N_3015,N_2737,N_2478);
nand U3016 (N_3016,N_2554,N_2672);
nor U3017 (N_3017,N_2712,N_2471);
or U3018 (N_3018,N_2986,N_2865);
nor U3019 (N_3019,N_2723,N_2594);
xnor U3020 (N_3020,N_2702,N_2938);
and U3021 (N_3021,N_2450,N_2664);
nand U3022 (N_3022,N_2603,N_2626);
nand U3023 (N_3023,N_2568,N_2463);
and U3024 (N_3024,N_2659,N_2449);
xnor U3025 (N_3025,N_2468,N_2631);
nand U3026 (N_3026,N_2762,N_2913);
or U3027 (N_3027,N_2602,N_2473);
or U3028 (N_3028,N_2457,N_2467);
nor U3029 (N_3029,N_2743,N_2915);
nand U3030 (N_3030,N_2978,N_2559);
or U3031 (N_3031,N_2958,N_2666);
or U3032 (N_3032,N_2851,N_2734);
and U3033 (N_3033,N_2618,N_2639);
and U3034 (N_3034,N_2847,N_2498);
nand U3035 (N_3035,N_2722,N_2608);
xnor U3036 (N_3036,N_2887,N_2867);
and U3037 (N_3037,N_2590,N_2953);
nor U3038 (N_3038,N_2932,N_2726);
nand U3039 (N_3039,N_2576,N_2655);
xor U3040 (N_3040,N_2804,N_2748);
and U3041 (N_3041,N_2877,N_2944);
xnor U3042 (N_3042,N_2721,N_2534);
or U3043 (N_3043,N_2786,N_2869);
nor U3044 (N_3044,N_2751,N_2413);
nor U3045 (N_3045,N_2415,N_2660);
xor U3046 (N_3046,N_2556,N_2647);
and U3047 (N_3047,N_2897,N_2483);
nand U3048 (N_3048,N_2581,N_2907);
or U3049 (N_3049,N_2765,N_2605);
and U3050 (N_3050,N_2946,N_2426);
or U3051 (N_3051,N_2538,N_2580);
nor U3052 (N_3052,N_2492,N_2678);
nor U3053 (N_3053,N_2652,N_2550);
xor U3054 (N_3054,N_2451,N_2452);
nor U3055 (N_3055,N_2911,N_2552);
xnor U3056 (N_3056,N_2782,N_2753);
xor U3057 (N_3057,N_2788,N_2919);
xnor U3058 (N_3058,N_2690,N_2925);
xnor U3059 (N_3059,N_2914,N_2419);
xor U3060 (N_3060,N_2515,N_2713);
xnor U3061 (N_3061,N_2674,N_2711);
and U3062 (N_3062,N_2527,N_2885);
nand U3063 (N_3063,N_2661,N_2805);
or U3064 (N_3064,N_2417,N_2866);
xnor U3065 (N_3065,N_2774,N_2439);
or U3066 (N_3066,N_2745,N_2884);
xor U3067 (N_3067,N_2518,N_2902);
nand U3068 (N_3068,N_2536,N_2638);
nor U3069 (N_3069,N_2771,N_2571);
nand U3070 (N_3070,N_2640,N_2669);
xor U3071 (N_3071,N_2604,N_2500);
or U3072 (N_3072,N_2755,N_2826);
nand U3073 (N_3073,N_2773,N_2569);
nor U3074 (N_3074,N_2828,N_2908);
or U3075 (N_3075,N_2617,N_2942);
or U3076 (N_3076,N_2474,N_2906);
nand U3077 (N_3077,N_2587,N_2738);
and U3078 (N_3078,N_2584,N_2757);
nand U3079 (N_3079,N_2514,N_2684);
nand U3080 (N_3080,N_2614,N_2863);
xor U3081 (N_3081,N_2752,N_2448);
nor U3082 (N_3082,N_2917,N_2420);
and U3083 (N_3083,N_2951,N_2957);
nand U3084 (N_3084,N_2790,N_2504);
nand U3085 (N_3085,N_2470,N_2645);
nor U3086 (N_3086,N_2636,N_2969);
nor U3087 (N_3087,N_2543,N_2905);
and U3088 (N_3088,N_2434,N_2896);
nor U3089 (N_3089,N_2704,N_2489);
nand U3090 (N_3090,N_2505,N_2533);
nor U3091 (N_3091,N_2763,N_2521);
nand U3092 (N_3092,N_2873,N_2565);
and U3093 (N_3093,N_2881,N_2698);
nand U3094 (N_3094,N_2528,N_2993);
and U3095 (N_3095,N_2675,N_2551);
xor U3096 (N_3096,N_2747,N_2522);
and U3097 (N_3097,N_2813,N_2864);
or U3098 (N_3098,N_2807,N_2435);
or U3099 (N_3099,N_2563,N_2720);
nand U3100 (N_3100,N_2988,N_2834);
xor U3101 (N_3101,N_2431,N_2546);
or U3102 (N_3102,N_2796,N_2530);
xnor U3103 (N_3103,N_2802,N_2837);
or U3104 (N_3104,N_2517,N_2954);
and U3105 (N_3105,N_2888,N_2776);
nand U3106 (N_3106,N_2511,N_2760);
and U3107 (N_3107,N_2572,N_2985);
or U3108 (N_3108,N_2519,N_2484);
and U3109 (N_3109,N_2730,N_2840);
or U3110 (N_3110,N_2650,N_2818);
xor U3111 (N_3111,N_2831,N_2524);
xnor U3112 (N_3112,N_2815,N_2510);
nand U3113 (N_3113,N_2692,N_2593);
or U3114 (N_3114,N_2405,N_2899);
and U3115 (N_3115,N_2477,N_2653);
or U3116 (N_3116,N_2564,N_2795);
nand U3117 (N_3117,N_2497,N_2822);
nand U3118 (N_3118,N_2507,N_2461);
xnor U3119 (N_3119,N_2544,N_2673);
xor U3120 (N_3120,N_2783,N_2615);
xor U3121 (N_3121,N_2689,N_2874);
nor U3122 (N_3122,N_2794,N_2844);
nor U3123 (N_3123,N_2716,N_2641);
and U3124 (N_3124,N_2838,N_2956);
nor U3125 (N_3125,N_2663,N_2693);
nand U3126 (N_3126,N_2761,N_2715);
or U3127 (N_3127,N_2637,N_2422);
nand U3128 (N_3128,N_2982,N_2814);
nand U3129 (N_3129,N_2547,N_2445);
nor U3130 (N_3130,N_2425,N_2890);
nand U3131 (N_3131,N_2630,N_2941);
nor U3132 (N_3132,N_2930,N_2525);
xnor U3133 (N_3133,N_2597,N_2537);
and U3134 (N_3134,N_2410,N_2975);
and U3135 (N_3135,N_2931,N_2924);
and U3136 (N_3136,N_2749,N_2853);
or U3137 (N_3137,N_2622,N_2973);
nor U3138 (N_3138,N_2950,N_2769);
and U3139 (N_3139,N_2456,N_2400);
or U3140 (N_3140,N_2531,N_2574);
and U3141 (N_3141,N_2812,N_2895);
or U3142 (N_3142,N_2454,N_2775);
xor U3143 (N_3143,N_2406,N_2465);
nand U3144 (N_3144,N_2872,N_2800);
nor U3145 (N_3145,N_2539,N_2703);
xor U3146 (N_3146,N_2854,N_2441);
or U3147 (N_3147,N_2778,N_2770);
and U3148 (N_3148,N_2827,N_2408);
or U3149 (N_3149,N_2810,N_2922);
nor U3150 (N_3150,N_2596,N_2947);
xnor U3151 (N_3151,N_2859,N_2933);
nand U3152 (N_3152,N_2725,N_2570);
and U3153 (N_3153,N_2823,N_2981);
nor U3154 (N_3154,N_2861,N_2876);
and U3155 (N_3155,N_2404,N_2485);
nor U3156 (N_3156,N_2526,N_2789);
nor U3157 (N_3157,N_2430,N_2599);
nor U3158 (N_3158,N_2535,N_2621);
xor U3159 (N_3159,N_2513,N_2735);
xor U3160 (N_3160,N_2740,N_2829);
nor U3161 (N_3161,N_2964,N_2423);
and U3162 (N_3162,N_2416,N_2680);
or U3163 (N_3163,N_2729,N_2756);
nor U3164 (N_3164,N_2857,N_2889);
nor U3165 (N_3165,N_2633,N_2839);
and U3166 (N_3166,N_2414,N_2793);
nand U3167 (N_3167,N_2480,N_2764);
nand U3168 (N_3168,N_2442,N_2443);
and U3169 (N_3169,N_2634,N_2998);
and U3170 (N_3170,N_2479,N_2825);
and U3171 (N_3171,N_2741,N_2742);
nand U3172 (N_3172,N_2971,N_2582);
xor U3173 (N_3173,N_2512,N_2992);
or U3174 (N_3174,N_2830,N_2462);
xor U3175 (N_3175,N_2671,N_2900);
and U3176 (N_3176,N_2646,N_2523);
or U3177 (N_3177,N_2424,N_2696);
or U3178 (N_3178,N_2785,N_2488);
or U3179 (N_3179,N_2901,N_2609);
xor U3180 (N_3180,N_2836,N_2959);
nor U3181 (N_3181,N_2894,N_2968);
nor U3182 (N_3182,N_2643,N_2583);
and U3183 (N_3183,N_2799,N_2868);
and U3184 (N_3184,N_2990,N_2632);
nor U3185 (N_3185,N_2573,N_2682);
or U3186 (N_3186,N_2841,N_2991);
or U3187 (N_3187,N_2677,N_2589);
or U3188 (N_3188,N_2548,N_2952);
xnor U3189 (N_3189,N_2852,N_2440);
nor U3190 (N_3190,N_2880,N_2475);
nand U3191 (N_3191,N_2903,N_2598);
nand U3192 (N_3192,N_2979,N_2921);
nand U3193 (N_3193,N_2999,N_2705);
xnor U3194 (N_3194,N_2706,N_2487);
xnor U3195 (N_3195,N_2965,N_2411);
nand U3196 (N_3196,N_2777,N_2739);
and U3197 (N_3197,N_2665,N_2961);
and U3198 (N_3198,N_2912,N_2649);
xor U3199 (N_3199,N_2648,N_2995);
xnor U3200 (N_3200,N_2699,N_2508);
nand U3201 (N_3201,N_2586,N_2695);
or U3202 (N_3202,N_2821,N_2429);
and U3203 (N_3203,N_2700,N_2444);
xnor U3204 (N_3204,N_2835,N_2433);
and U3205 (N_3205,N_2491,N_2898);
nor U3206 (N_3206,N_2437,N_2849);
xor U3207 (N_3207,N_2681,N_2620);
xnor U3208 (N_3208,N_2601,N_2832);
nand U3209 (N_3209,N_2808,N_2472);
and U3210 (N_3210,N_2501,N_2878);
or U3211 (N_3211,N_2532,N_2927);
or U3212 (N_3212,N_2670,N_2893);
nor U3213 (N_3213,N_2974,N_2623);
xnor U3214 (N_3214,N_2676,N_2509);
nand U3215 (N_3215,N_2616,N_2862);
nor U3216 (N_3216,N_2685,N_2455);
and U3217 (N_3217,N_2600,N_2579);
nor U3218 (N_3218,N_2486,N_2803);
nand U3219 (N_3219,N_2791,N_2994);
nor U3220 (N_3220,N_2750,N_2575);
nor U3221 (N_3221,N_2736,N_2819);
xor U3222 (N_3222,N_2909,N_2401);
or U3223 (N_3223,N_2833,N_2628);
nor U3224 (N_3224,N_2679,N_2686);
and U3225 (N_3225,N_2506,N_2654);
nand U3226 (N_3226,N_2662,N_2939);
xor U3227 (N_3227,N_2935,N_2883);
or U3228 (N_3228,N_2731,N_2781);
nand U3229 (N_3229,N_2976,N_2447);
nor U3230 (N_3230,N_2784,N_2611);
nor U3231 (N_3231,N_2855,N_2403);
nor U3232 (N_3232,N_2806,N_2972);
nor U3233 (N_3233,N_2694,N_2824);
nand U3234 (N_3234,N_2945,N_2561);
xnor U3235 (N_3235,N_2493,N_2949);
nand U3236 (N_3236,N_2934,N_2520);
nand U3237 (N_3237,N_2962,N_2820);
nor U3238 (N_3238,N_2892,N_2427);
and U3239 (N_3239,N_2635,N_2502);
or U3240 (N_3240,N_2918,N_2929);
or U3241 (N_3241,N_2651,N_2926);
nor U3242 (N_3242,N_2464,N_2529);
xnor U3243 (N_3243,N_2904,N_2708);
or U3244 (N_3244,N_2607,N_2567);
nand U3245 (N_3245,N_2503,N_2469);
or U3246 (N_3246,N_2481,N_2746);
nor U3247 (N_3247,N_2707,N_2591);
and U3248 (N_3248,N_2516,N_2545);
or U3249 (N_3249,N_2817,N_2458);
nor U3250 (N_3250,N_2595,N_2714);
or U3251 (N_3251,N_2923,N_2848);
and U3252 (N_3252,N_2658,N_2710);
nor U3253 (N_3253,N_2732,N_2882);
and U3254 (N_3254,N_2936,N_2767);
nand U3255 (N_3255,N_2792,N_2963);
nand U3256 (N_3256,N_2816,N_2970);
xnor U3257 (N_3257,N_2667,N_2871);
or U3258 (N_3258,N_2728,N_2560);
nand U3259 (N_3259,N_2562,N_2809);
and U3260 (N_3260,N_2407,N_2754);
and U3261 (N_3261,N_2612,N_2446);
nand U3262 (N_3262,N_2719,N_2801);
nor U3263 (N_3263,N_2490,N_2625);
or U3264 (N_3264,N_2557,N_2709);
and U3265 (N_3265,N_2940,N_2418);
nand U3266 (N_3266,N_2683,N_2717);
or U3267 (N_3267,N_2768,N_2943);
xnor U3268 (N_3268,N_2928,N_2668);
xor U3269 (N_3269,N_2453,N_2758);
nor U3270 (N_3270,N_2701,N_2920);
nor U3271 (N_3271,N_2421,N_2787);
or U3272 (N_3272,N_2697,N_2409);
xor U3273 (N_3273,N_2860,N_2955);
or U3274 (N_3274,N_2402,N_2937);
nor U3275 (N_3275,N_2657,N_2691);
nor U3276 (N_3276,N_2496,N_2879);
nor U3277 (N_3277,N_2499,N_2724);
nor U3278 (N_3278,N_2606,N_2843);
nor U3279 (N_3279,N_2960,N_2577);
or U3280 (N_3280,N_2585,N_2856);
and U3281 (N_3281,N_2629,N_2610);
nor U3282 (N_3282,N_2541,N_2482);
and U3283 (N_3283,N_2984,N_2578);
xor U3284 (N_3284,N_2989,N_2891);
nand U3285 (N_3285,N_2688,N_2966);
nor U3286 (N_3286,N_2540,N_2811);
nand U3287 (N_3287,N_2780,N_2980);
nor U3288 (N_3288,N_2624,N_2428);
and U3289 (N_3289,N_2558,N_2766);
and U3290 (N_3290,N_2842,N_2727);
nand U3291 (N_3291,N_2772,N_2644);
nor U3292 (N_3292,N_2718,N_2967);
nand U3293 (N_3293,N_2687,N_2759);
or U3294 (N_3294,N_2619,N_2592);
nand U3295 (N_3295,N_2542,N_2797);
nor U3296 (N_3296,N_2460,N_2875);
xor U3297 (N_3297,N_2996,N_2977);
nor U3298 (N_3298,N_2744,N_2997);
nor U3299 (N_3299,N_2495,N_2886);
or U3300 (N_3300,N_2963,N_2459);
xor U3301 (N_3301,N_2549,N_2472);
and U3302 (N_3302,N_2840,N_2744);
or U3303 (N_3303,N_2734,N_2676);
nand U3304 (N_3304,N_2903,N_2871);
and U3305 (N_3305,N_2400,N_2993);
and U3306 (N_3306,N_2734,N_2808);
nor U3307 (N_3307,N_2815,N_2871);
xnor U3308 (N_3308,N_2793,N_2564);
and U3309 (N_3309,N_2683,N_2672);
nand U3310 (N_3310,N_2991,N_2585);
nor U3311 (N_3311,N_2424,N_2490);
and U3312 (N_3312,N_2491,N_2654);
xor U3313 (N_3313,N_2870,N_2556);
or U3314 (N_3314,N_2925,N_2704);
or U3315 (N_3315,N_2659,N_2952);
nor U3316 (N_3316,N_2541,N_2811);
and U3317 (N_3317,N_2874,N_2934);
nand U3318 (N_3318,N_2831,N_2958);
and U3319 (N_3319,N_2958,N_2717);
or U3320 (N_3320,N_2805,N_2745);
nor U3321 (N_3321,N_2860,N_2529);
and U3322 (N_3322,N_2650,N_2754);
nand U3323 (N_3323,N_2613,N_2598);
xor U3324 (N_3324,N_2648,N_2694);
nor U3325 (N_3325,N_2549,N_2565);
xor U3326 (N_3326,N_2461,N_2545);
xor U3327 (N_3327,N_2845,N_2409);
xnor U3328 (N_3328,N_2984,N_2588);
or U3329 (N_3329,N_2622,N_2907);
nand U3330 (N_3330,N_2493,N_2675);
and U3331 (N_3331,N_2466,N_2410);
and U3332 (N_3332,N_2522,N_2563);
xnor U3333 (N_3333,N_2579,N_2946);
or U3334 (N_3334,N_2608,N_2733);
or U3335 (N_3335,N_2658,N_2630);
nand U3336 (N_3336,N_2777,N_2571);
nand U3337 (N_3337,N_2820,N_2402);
or U3338 (N_3338,N_2895,N_2574);
xnor U3339 (N_3339,N_2962,N_2831);
nor U3340 (N_3340,N_2740,N_2701);
or U3341 (N_3341,N_2563,N_2462);
or U3342 (N_3342,N_2410,N_2477);
nand U3343 (N_3343,N_2632,N_2941);
or U3344 (N_3344,N_2800,N_2974);
nand U3345 (N_3345,N_2924,N_2456);
xnor U3346 (N_3346,N_2742,N_2758);
xor U3347 (N_3347,N_2446,N_2543);
or U3348 (N_3348,N_2513,N_2516);
or U3349 (N_3349,N_2867,N_2691);
xor U3350 (N_3350,N_2573,N_2690);
nor U3351 (N_3351,N_2750,N_2452);
nand U3352 (N_3352,N_2902,N_2668);
nor U3353 (N_3353,N_2438,N_2602);
nand U3354 (N_3354,N_2765,N_2939);
xnor U3355 (N_3355,N_2783,N_2909);
xnor U3356 (N_3356,N_2982,N_2634);
nor U3357 (N_3357,N_2913,N_2685);
or U3358 (N_3358,N_2837,N_2751);
nand U3359 (N_3359,N_2608,N_2926);
or U3360 (N_3360,N_2741,N_2563);
and U3361 (N_3361,N_2818,N_2580);
xor U3362 (N_3362,N_2589,N_2656);
xnor U3363 (N_3363,N_2512,N_2466);
nor U3364 (N_3364,N_2883,N_2684);
nor U3365 (N_3365,N_2609,N_2948);
or U3366 (N_3366,N_2913,N_2601);
xor U3367 (N_3367,N_2833,N_2437);
or U3368 (N_3368,N_2702,N_2591);
nand U3369 (N_3369,N_2419,N_2754);
nor U3370 (N_3370,N_2932,N_2593);
nor U3371 (N_3371,N_2650,N_2812);
nor U3372 (N_3372,N_2985,N_2750);
nor U3373 (N_3373,N_2477,N_2458);
xnor U3374 (N_3374,N_2421,N_2805);
xor U3375 (N_3375,N_2675,N_2527);
or U3376 (N_3376,N_2932,N_2807);
xor U3377 (N_3377,N_2515,N_2771);
nor U3378 (N_3378,N_2768,N_2853);
or U3379 (N_3379,N_2655,N_2888);
nor U3380 (N_3380,N_2692,N_2823);
or U3381 (N_3381,N_2475,N_2989);
xnor U3382 (N_3382,N_2815,N_2773);
and U3383 (N_3383,N_2876,N_2447);
nand U3384 (N_3384,N_2977,N_2411);
or U3385 (N_3385,N_2530,N_2895);
nor U3386 (N_3386,N_2515,N_2588);
nand U3387 (N_3387,N_2608,N_2888);
nand U3388 (N_3388,N_2746,N_2508);
and U3389 (N_3389,N_2762,N_2944);
or U3390 (N_3390,N_2494,N_2834);
nand U3391 (N_3391,N_2615,N_2855);
xnor U3392 (N_3392,N_2925,N_2628);
nor U3393 (N_3393,N_2951,N_2779);
nand U3394 (N_3394,N_2963,N_2414);
or U3395 (N_3395,N_2896,N_2920);
or U3396 (N_3396,N_2441,N_2402);
nand U3397 (N_3397,N_2881,N_2888);
nand U3398 (N_3398,N_2589,N_2609);
or U3399 (N_3399,N_2910,N_2613);
or U3400 (N_3400,N_2833,N_2533);
or U3401 (N_3401,N_2764,N_2407);
xnor U3402 (N_3402,N_2440,N_2522);
nand U3403 (N_3403,N_2927,N_2517);
and U3404 (N_3404,N_2944,N_2783);
nand U3405 (N_3405,N_2457,N_2971);
and U3406 (N_3406,N_2747,N_2816);
nand U3407 (N_3407,N_2560,N_2998);
nor U3408 (N_3408,N_2682,N_2413);
or U3409 (N_3409,N_2718,N_2860);
or U3410 (N_3410,N_2973,N_2509);
or U3411 (N_3411,N_2911,N_2987);
nand U3412 (N_3412,N_2979,N_2720);
or U3413 (N_3413,N_2679,N_2631);
nand U3414 (N_3414,N_2970,N_2857);
xor U3415 (N_3415,N_2727,N_2530);
nand U3416 (N_3416,N_2982,N_2666);
nand U3417 (N_3417,N_2789,N_2567);
or U3418 (N_3418,N_2671,N_2514);
or U3419 (N_3419,N_2613,N_2753);
xnor U3420 (N_3420,N_2748,N_2810);
or U3421 (N_3421,N_2403,N_2814);
nand U3422 (N_3422,N_2531,N_2957);
nor U3423 (N_3423,N_2629,N_2488);
or U3424 (N_3424,N_2543,N_2609);
xor U3425 (N_3425,N_2465,N_2557);
and U3426 (N_3426,N_2777,N_2674);
nand U3427 (N_3427,N_2840,N_2435);
nand U3428 (N_3428,N_2709,N_2809);
nand U3429 (N_3429,N_2712,N_2978);
nand U3430 (N_3430,N_2499,N_2897);
xor U3431 (N_3431,N_2998,N_2997);
nand U3432 (N_3432,N_2924,N_2842);
and U3433 (N_3433,N_2879,N_2753);
nor U3434 (N_3434,N_2677,N_2769);
xnor U3435 (N_3435,N_2436,N_2514);
or U3436 (N_3436,N_2571,N_2514);
nor U3437 (N_3437,N_2426,N_2707);
nand U3438 (N_3438,N_2702,N_2712);
xor U3439 (N_3439,N_2841,N_2873);
or U3440 (N_3440,N_2526,N_2694);
and U3441 (N_3441,N_2669,N_2650);
nor U3442 (N_3442,N_2499,N_2578);
xnor U3443 (N_3443,N_2446,N_2532);
or U3444 (N_3444,N_2500,N_2643);
xnor U3445 (N_3445,N_2766,N_2618);
nor U3446 (N_3446,N_2800,N_2447);
or U3447 (N_3447,N_2547,N_2776);
nor U3448 (N_3448,N_2914,N_2736);
and U3449 (N_3449,N_2800,N_2675);
or U3450 (N_3450,N_2809,N_2457);
xor U3451 (N_3451,N_2871,N_2983);
or U3452 (N_3452,N_2657,N_2491);
xor U3453 (N_3453,N_2625,N_2874);
xnor U3454 (N_3454,N_2845,N_2562);
or U3455 (N_3455,N_2874,N_2603);
and U3456 (N_3456,N_2654,N_2504);
or U3457 (N_3457,N_2598,N_2531);
nand U3458 (N_3458,N_2800,N_2695);
nor U3459 (N_3459,N_2444,N_2542);
nor U3460 (N_3460,N_2679,N_2585);
xor U3461 (N_3461,N_2869,N_2880);
nand U3462 (N_3462,N_2829,N_2907);
nor U3463 (N_3463,N_2439,N_2530);
and U3464 (N_3464,N_2472,N_2485);
nand U3465 (N_3465,N_2591,N_2935);
xor U3466 (N_3466,N_2628,N_2913);
or U3467 (N_3467,N_2779,N_2471);
and U3468 (N_3468,N_2642,N_2426);
and U3469 (N_3469,N_2824,N_2791);
or U3470 (N_3470,N_2757,N_2599);
nand U3471 (N_3471,N_2577,N_2537);
xor U3472 (N_3472,N_2495,N_2674);
and U3473 (N_3473,N_2588,N_2972);
and U3474 (N_3474,N_2553,N_2548);
nor U3475 (N_3475,N_2773,N_2456);
or U3476 (N_3476,N_2461,N_2547);
nand U3477 (N_3477,N_2680,N_2987);
nor U3478 (N_3478,N_2585,N_2528);
xnor U3479 (N_3479,N_2859,N_2523);
and U3480 (N_3480,N_2577,N_2918);
xnor U3481 (N_3481,N_2431,N_2628);
nor U3482 (N_3482,N_2971,N_2799);
nand U3483 (N_3483,N_2999,N_2792);
or U3484 (N_3484,N_2953,N_2487);
or U3485 (N_3485,N_2609,N_2498);
nor U3486 (N_3486,N_2656,N_2786);
nand U3487 (N_3487,N_2521,N_2680);
and U3488 (N_3488,N_2838,N_2793);
nand U3489 (N_3489,N_2445,N_2820);
or U3490 (N_3490,N_2741,N_2623);
and U3491 (N_3491,N_2969,N_2725);
nor U3492 (N_3492,N_2850,N_2468);
and U3493 (N_3493,N_2700,N_2990);
xor U3494 (N_3494,N_2985,N_2711);
xor U3495 (N_3495,N_2565,N_2983);
xnor U3496 (N_3496,N_2476,N_2818);
and U3497 (N_3497,N_2482,N_2927);
xnor U3498 (N_3498,N_2585,N_2511);
nand U3499 (N_3499,N_2983,N_2591);
and U3500 (N_3500,N_2706,N_2743);
and U3501 (N_3501,N_2964,N_2880);
nand U3502 (N_3502,N_2684,N_2656);
nand U3503 (N_3503,N_2452,N_2778);
nand U3504 (N_3504,N_2626,N_2452);
nor U3505 (N_3505,N_2512,N_2495);
nand U3506 (N_3506,N_2926,N_2579);
xnor U3507 (N_3507,N_2510,N_2470);
or U3508 (N_3508,N_2984,N_2453);
or U3509 (N_3509,N_2423,N_2667);
and U3510 (N_3510,N_2411,N_2819);
or U3511 (N_3511,N_2579,N_2605);
and U3512 (N_3512,N_2566,N_2838);
and U3513 (N_3513,N_2592,N_2741);
xnor U3514 (N_3514,N_2774,N_2702);
or U3515 (N_3515,N_2575,N_2712);
or U3516 (N_3516,N_2553,N_2511);
or U3517 (N_3517,N_2976,N_2410);
and U3518 (N_3518,N_2591,N_2592);
xor U3519 (N_3519,N_2703,N_2726);
xor U3520 (N_3520,N_2435,N_2781);
or U3521 (N_3521,N_2961,N_2765);
nand U3522 (N_3522,N_2635,N_2584);
and U3523 (N_3523,N_2673,N_2518);
nand U3524 (N_3524,N_2601,N_2565);
nor U3525 (N_3525,N_2949,N_2756);
or U3526 (N_3526,N_2758,N_2978);
or U3527 (N_3527,N_2461,N_2864);
xnor U3528 (N_3528,N_2455,N_2906);
or U3529 (N_3529,N_2702,N_2949);
nor U3530 (N_3530,N_2728,N_2806);
nand U3531 (N_3531,N_2554,N_2713);
and U3532 (N_3532,N_2602,N_2973);
xor U3533 (N_3533,N_2765,N_2659);
or U3534 (N_3534,N_2722,N_2832);
nor U3535 (N_3535,N_2437,N_2507);
and U3536 (N_3536,N_2414,N_2573);
nand U3537 (N_3537,N_2756,N_2609);
xnor U3538 (N_3538,N_2803,N_2540);
nor U3539 (N_3539,N_2524,N_2983);
xnor U3540 (N_3540,N_2731,N_2821);
xnor U3541 (N_3541,N_2924,N_2784);
nand U3542 (N_3542,N_2494,N_2536);
or U3543 (N_3543,N_2624,N_2670);
or U3544 (N_3544,N_2713,N_2719);
xnor U3545 (N_3545,N_2440,N_2513);
or U3546 (N_3546,N_2942,N_2445);
or U3547 (N_3547,N_2517,N_2863);
and U3548 (N_3548,N_2454,N_2805);
nand U3549 (N_3549,N_2618,N_2977);
xor U3550 (N_3550,N_2973,N_2460);
nor U3551 (N_3551,N_2668,N_2995);
nor U3552 (N_3552,N_2557,N_2676);
nand U3553 (N_3553,N_2960,N_2965);
or U3554 (N_3554,N_2604,N_2487);
nand U3555 (N_3555,N_2979,N_2744);
or U3556 (N_3556,N_2656,N_2707);
or U3557 (N_3557,N_2587,N_2835);
xor U3558 (N_3558,N_2813,N_2655);
or U3559 (N_3559,N_2416,N_2887);
xor U3560 (N_3560,N_2694,N_2937);
and U3561 (N_3561,N_2506,N_2513);
nor U3562 (N_3562,N_2549,N_2506);
xnor U3563 (N_3563,N_2732,N_2822);
xnor U3564 (N_3564,N_2839,N_2612);
and U3565 (N_3565,N_2660,N_2653);
and U3566 (N_3566,N_2818,N_2736);
nand U3567 (N_3567,N_2908,N_2867);
and U3568 (N_3568,N_2961,N_2414);
nor U3569 (N_3569,N_2614,N_2540);
nor U3570 (N_3570,N_2420,N_2790);
and U3571 (N_3571,N_2564,N_2610);
nor U3572 (N_3572,N_2960,N_2672);
and U3573 (N_3573,N_2998,N_2928);
nand U3574 (N_3574,N_2765,N_2555);
nor U3575 (N_3575,N_2586,N_2909);
or U3576 (N_3576,N_2966,N_2992);
and U3577 (N_3577,N_2584,N_2626);
nand U3578 (N_3578,N_2957,N_2544);
nor U3579 (N_3579,N_2752,N_2540);
nand U3580 (N_3580,N_2581,N_2488);
xnor U3581 (N_3581,N_2844,N_2834);
and U3582 (N_3582,N_2988,N_2999);
or U3583 (N_3583,N_2539,N_2756);
nor U3584 (N_3584,N_2527,N_2571);
xor U3585 (N_3585,N_2888,N_2507);
or U3586 (N_3586,N_2747,N_2914);
and U3587 (N_3587,N_2565,N_2839);
nand U3588 (N_3588,N_2527,N_2725);
and U3589 (N_3589,N_2568,N_2999);
xor U3590 (N_3590,N_2897,N_2458);
and U3591 (N_3591,N_2974,N_2811);
xor U3592 (N_3592,N_2500,N_2735);
nand U3593 (N_3593,N_2603,N_2512);
nor U3594 (N_3594,N_2852,N_2996);
nor U3595 (N_3595,N_2507,N_2643);
and U3596 (N_3596,N_2761,N_2736);
nor U3597 (N_3597,N_2872,N_2789);
xor U3598 (N_3598,N_2874,N_2794);
nand U3599 (N_3599,N_2662,N_2460);
nor U3600 (N_3600,N_3141,N_3383);
nand U3601 (N_3601,N_3581,N_3245);
or U3602 (N_3602,N_3167,N_3177);
nor U3603 (N_3603,N_3487,N_3423);
or U3604 (N_3604,N_3284,N_3330);
nor U3605 (N_3605,N_3565,N_3143);
and U3606 (N_3606,N_3094,N_3080);
and U3607 (N_3607,N_3260,N_3077);
and U3608 (N_3608,N_3180,N_3058);
and U3609 (N_3609,N_3113,N_3116);
xor U3610 (N_3610,N_3578,N_3041);
xor U3611 (N_3611,N_3365,N_3569);
nor U3612 (N_3612,N_3033,N_3158);
xor U3613 (N_3613,N_3082,N_3222);
nand U3614 (N_3614,N_3079,N_3530);
nand U3615 (N_3615,N_3430,N_3376);
xor U3616 (N_3616,N_3134,N_3480);
nor U3617 (N_3617,N_3050,N_3303);
or U3618 (N_3618,N_3521,N_3479);
nor U3619 (N_3619,N_3542,N_3321);
nand U3620 (N_3620,N_3380,N_3357);
nor U3621 (N_3621,N_3200,N_3329);
nor U3622 (N_3622,N_3121,N_3154);
xor U3623 (N_3623,N_3316,N_3492);
nand U3624 (N_3624,N_3532,N_3211);
xnor U3625 (N_3625,N_3131,N_3318);
nor U3626 (N_3626,N_3510,N_3571);
nand U3627 (N_3627,N_3101,N_3025);
xnor U3628 (N_3628,N_3468,N_3074);
xnor U3629 (N_3629,N_3105,N_3499);
nand U3630 (N_3630,N_3460,N_3442);
nand U3631 (N_3631,N_3297,N_3439);
nand U3632 (N_3632,N_3241,N_3411);
nor U3633 (N_3633,N_3298,N_3497);
nand U3634 (N_3634,N_3202,N_3014);
nor U3635 (N_3635,N_3336,N_3166);
nor U3636 (N_3636,N_3465,N_3300);
nand U3637 (N_3637,N_3562,N_3308);
and U3638 (N_3638,N_3396,N_3013);
or U3639 (N_3639,N_3547,N_3496);
or U3640 (N_3640,N_3512,N_3185);
nor U3641 (N_3641,N_3556,N_3037);
or U3642 (N_3642,N_3389,N_3020);
and U3643 (N_3643,N_3086,N_3559);
nand U3644 (N_3644,N_3433,N_3520);
nand U3645 (N_3645,N_3119,N_3215);
xnor U3646 (N_3646,N_3428,N_3341);
nand U3647 (N_3647,N_3395,N_3440);
xnor U3648 (N_3648,N_3238,N_3507);
and U3649 (N_3649,N_3282,N_3247);
xnor U3650 (N_3650,N_3490,N_3504);
or U3651 (N_3651,N_3089,N_3124);
nor U3652 (N_3652,N_3372,N_3159);
nor U3653 (N_3653,N_3043,N_3534);
nand U3654 (N_3654,N_3466,N_3432);
nand U3655 (N_3655,N_3481,N_3107);
nand U3656 (N_3656,N_3386,N_3059);
nand U3657 (N_3657,N_3262,N_3566);
and U3658 (N_3658,N_3355,N_3498);
and U3659 (N_3659,N_3312,N_3589);
nor U3660 (N_3660,N_3172,N_3168);
or U3661 (N_3661,N_3213,N_3067);
and U3662 (N_3662,N_3276,N_3135);
nor U3663 (N_3663,N_3580,N_3413);
nor U3664 (N_3664,N_3563,N_3391);
nand U3665 (N_3665,N_3403,N_3036);
and U3666 (N_3666,N_3017,N_3169);
nand U3667 (N_3667,N_3431,N_3579);
nor U3668 (N_3668,N_3174,N_3047);
nor U3669 (N_3669,N_3127,N_3418);
nor U3670 (N_3670,N_3148,N_3553);
nand U3671 (N_3671,N_3065,N_3505);
nand U3672 (N_3672,N_3449,N_3333);
or U3673 (N_3673,N_3390,N_3593);
and U3674 (N_3674,N_3406,N_3339);
xor U3675 (N_3675,N_3452,N_3206);
xnor U3676 (N_3676,N_3026,N_3191);
xnor U3677 (N_3677,N_3083,N_3334);
or U3678 (N_3678,N_3155,N_3299);
xnor U3679 (N_3679,N_3209,N_3558);
xnor U3680 (N_3680,N_3275,N_3181);
nor U3681 (N_3681,N_3427,N_3595);
or U3682 (N_3682,N_3332,N_3438);
and U3683 (N_3683,N_3235,N_3228);
or U3684 (N_3684,N_3108,N_3529);
nand U3685 (N_3685,N_3269,N_3021);
xnor U3686 (N_3686,N_3404,N_3560);
nor U3687 (N_3687,N_3443,N_3236);
or U3688 (N_3688,N_3220,N_3258);
nor U3689 (N_3689,N_3522,N_3313);
and U3690 (N_3690,N_3016,N_3103);
nand U3691 (N_3691,N_3271,N_3212);
nand U3692 (N_3692,N_3374,N_3267);
nand U3693 (N_3693,N_3062,N_3118);
or U3694 (N_3694,N_3204,N_3295);
or U3695 (N_3695,N_3445,N_3296);
or U3696 (N_3696,N_3182,N_3464);
and U3697 (N_3697,N_3458,N_3585);
nand U3698 (N_3698,N_3599,N_3249);
nor U3699 (N_3699,N_3109,N_3388);
nor U3700 (N_3700,N_3156,N_3576);
nand U3701 (N_3701,N_3231,N_3369);
nor U3702 (N_3702,N_3291,N_3123);
xnor U3703 (N_3703,N_3410,N_3470);
xnor U3704 (N_3704,N_3268,N_3347);
nand U3705 (N_3705,N_3409,N_3052);
nand U3706 (N_3706,N_3527,N_3243);
nor U3707 (N_3707,N_3461,N_3183);
nand U3708 (N_3708,N_3574,N_3517);
nor U3709 (N_3709,N_3533,N_3005);
xnor U3710 (N_3710,N_3320,N_3032);
or U3711 (N_3711,N_3264,N_3484);
nor U3712 (N_3712,N_3494,N_3371);
nor U3713 (N_3713,N_3352,N_3583);
nand U3714 (N_3714,N_3392,N_3144);
nand U3715 (N_3715,N_3188,N_3309);
or U3716 (N_3716,N_3394,N_3099);
nor U3717 (N_3717,N_3035,N_3225);
or U3718 (N_3718,N_3071,N_3535);
nand U3719 (N_3719,N_3425,N_3214);
xor U3720 (N_3720,N_3591,N_3474);
or U3721 (N_3721,N_3278,N_3230);
nor U3722 (N_3722,N_3338,N_3179);
nand U3723 (N_3723,N_3457,N_3205);
or U3724 (N_3724,N_3543,N_3250);
nor U3725 (N_3725,N_3328,N_3597);
xor U3726 (N_3726,N_3375,N_3592);
nand U3727 (N_3727,N_3596,N_3463);
nand U3728 (N_3728,N_3501,N_3381);
and U3729 (N_3729,N_3049,N_3417);
nand U3730 (N_3730,N_3459,N_3126);
and U3731 (N_3731,N_3160,N_3051);
nor U3732 (N_3732,N_3359,N_3146);
and U3733 (N_3733,N_3324,N_3584);
or U3734 (N_3734,N_3446,N_3045);
and U3735 (N_3735,N_3069,N_3340);
or U3736 (N_3736,N_3518,N_3493);
and U3737 (N_3737,N_3286,N_3454);
nand U3738 (N_3738,N_3248,N_3531);
nand U3739 (N_3739,N_3254,N_3010);
nor U3740 (N_3740,N_3450,N_3219);
nor U3741 (N_3741,N_3007,N_3216);
xnor U3742 (N_3742,N_3437,N_3472);
and U3743 (N_3743,N_3024,N_3218);
nand U3744 (N_3744,N_3102,N_3057);
and U3745 (N_3745,N_3110,N_3598);
and U3746 (N_3746,N_3223,N_3112);
nor U3747 (N_3747,N_3537,N_3421);
nand U3748 (N_3748,N_3053,N_3467);
nand U3749 (N_3749,N_3162,N_3055);
xor U3750 (N_3750,N_3149,N_3195);
or U3751 (N_3751,N_3471,N_3373);
nor U3752 (N_3752,N_3420,N_3070);
nand U3753 (N_3753,N_3039,N_3265);
or U3754 (N_3754,N_3003,N_3226);
xor U3755 (N_3755,N_3367,N_3536);
nand U3756 (N_3756,N_3190,N_3462);
or U3757 (N_3757,N_3257,N_3561);
and U3758 (N_3758,N_3034,N_3317);
nand U3759 (N_3759,N_3551,N_3064);
xnor U3760 (N_3760,N_3201,N_3519);
and U3761 (N_3761,N_3489,N_3364);
or U3762 (N_3762,N_3028,N_3273);
nor U3763 (N_3763,N_3042,N_3436);
nor U3764 (N_3764,N_3000,N_3416);
or U3765 (N_3765,N_3186,N_3502);
and U3766 (N_3766,N_3076,N_3319);
nor U3767 (N_3767,N_3526,N_3277);
or U3768 (N_3768,N_3397,N_3019);
nor U3769 (N_3769,N_3165,N_3544);
xor U3770 (N_3770,N_3322,N_3500);
or U3771 (N_3771,N_3572,N_3353);
or U3772 (N_3772,N_3444,N_3046);
or U3773 (N_3773,N_3424,N_3068);
xor U3774 (N_3774,N_3337,N_3304);
or U3775 (N_3775,N_3491,N_3414);
nor U3776 (N_3776,N_3582,N_3060);
and U3777 (N_3777,N_3075,N_3577);
nor U3778 (N_3778,N_3161,N_3163);
or U3779 (N_3779,N_3385,N_3040);
xor U3780 (N_3780,N_3187,N_3157);
xor U3781 (N_3781,N_3233,N_3279);
xor U3782 (N_3782,N_3259,N_3125);
xor U3783 (N_3783,N_3266,N_3311);
and U3784 (N_3784,N_3176,N_3590);
xnor U3785 (N_3785,N_3557,N_3356);
and U3786 (N_3786,N_3448,N_3227);
or U3787 (N_3787,N_3221,N_3066);
xor U3788 (N_3788,N_3244,N_3054);
nand U3789 (N_3789,N_3012,N_3088);
and U3790 (N_3790,N_3111,N_3350);
nand U3791 (N_3791,N_3198,N_3027);
nand U3792 (N_3792,N_3085,N_3384);
nor U3793 (N_3793,N_3242,N_3594);
or U3794 (N_3794,N_3587,N_3325);
xor U3795 (N_3795,N_3239,N_3008);
nor U3796 (N_3796,N_3173,N_3415);
and U3797 (N_3797,N_3129,N_3253);
nor U3798 (N_3798,N_3570,N_3096);
nand U3799 (N_3799,N_3031,N_3004);
or U3800 (N_3800,N_3128,N_3150);
or U3801 (N_3801,N_3117,N_3514);
xor U3802 (N_3802,N_3084,N_3555);
and U3803 (N_3803,N_3274,N_3140);
or U3804 (N_3804,N_3270,N_3545);
xnor U3805 (N_3805,N_3192,N_3335);
nor U3806 (N_3806,N_3314,N_3554);
nand U3807 (N_3807,N_3175,N_3546);
and U3808 (N_3808,N_3525,N_3237);
nor U3809 (N_3809,N_3002,N_3151);
and U3810 (N_3810,N_3009,N_3379);
nand U3811 (N_3811,N_3208,N_3511);
nand U3812 (N_3812,N_3048,N_3358);
nand U3813 (N_3813,N_3001,N_3306);
and U3814 (N_3814,N_3038,N_3132);
nor U3815 (N_3815,N_3366,N_3399);
nand U3816 (N_3816,N_3368,N_3104);
nor U3817 (N_3817,N_3293,N_3139);
nor U3818 (N_3818,N_3184,N_3261);
nor U3819 (N_3819,N_3018,N_3283);
xor U3820 (N_3820,N_3568,N_3344);
or U3821 (N_3821,N_3255,N_3029);
nand U3822 (N_3822,N_3073,N_3170);
nor U3823 (N_3823,N_3097,N_3130);
xnor U3824 (N_3824,N_3441,N_3199);
or U3825 (N_3825,N_3289,N_3246);
or U3826 (N_3826,N_3091,N_3538);
xor U3827 (N_3827,N_3092,N_3370);
and U3828 (N_3828,N_3217,N_3363);
and U3829 (N_3829,N_3072,N_3061);
or U3830 (N_3830,N_3400,N_3539);
or U3831 (N_3831,N_3426,N_3345);
or U3832 (N_3832,N_3056,N_3145);
nand U3833 (N_3833,N_3194,N_3469);
and U3834 (N_3834,N_3288,N_3022);
xnor U3835 (N_3835,N_3203,N_3164);
xor U3836 (N_3836,N_3509,N_3152);
nand U3837 (N_3837,N_3407,N_3564);
nand U3838 (N_3838,N_3354,N_3290);
xnor U3839 (N_3839,N_3343,N_3234);
nor U3840 (N_3840,N_3434,N_3224);
nand U3841 (N_3841,N_3095,N_3310);
or U3842 (N_3842,N_3435,N_3292);
xor U3843 (N_3843,N_3252,N_3412);
nor U3844 (N_3844,N_3323,N_3307);
nor U3845 (N_3845,N_3477,N_3361);
nor U3846 (N_3846,N_3302,N_3567);
nand U3847 (N_3847,N_3342,N_3408);
nand U3848 (N_3848,N_3515,N_3106);
nor U3849 (N_3849,N_3136,N_3456);
nor U3850 (N_3850,N_3137,N_3011);
and U3851 (N_3851,N_3475,N_3488);
or U3852 (N_3852,N_3473,N_3478);
nor U3853 (N_3853,N_3524,N_3147);
or U3854 (N_3854,N_3287,N_3513);
nor U3855 (N_3855,N_3210,N_3232);
nor U3856 (N_3856,N_3405,N_3528);
and U3857 (N_3857,N_3015,N_3482);
nor U3858 (N_3858,N_3122,N_3301);
nor U3859 (N_3859,N_3360,N_3081);
nor U3860 (N_3860,N_3193,N_3090);
xnor U3861 (N_3861,N_3171,N_3196);
xnor U3862 (N_3862,N_3093,N_3348);
and U3863 (N_3863,N_3401,N_3387);
nand U3864 (N_3864,N_3429,N_3280);
nand U3865 (N_3865,N_3455,N_3550);
and U3866 (N_3866,N_3447,N_3326);
and U3867 (N_3867,N_3063,N_3588);
nand U3868 (N_3868,N_3315,N_3351);
xnor U3869 (N_3869,N_3281,N_3207);
xor U3870 (N_3870,N_3115,N_3023);
xor U3871 (N_3871,N_3100,N_3251);
or U3872 (N_3872,N_3495,N_3503);
and U3873 (N_3873,N_3138,N_3044);
nor U3874 (N_3874,N_3142,N_3006);
nand U3875 (N_3875,N_3516,N_3541);
nor U3876 (N_3876,N_3398,N_3272);
nor U3877 (N_3877,N_3549,N_3382);
xor U3878 (N_3878,N_3575,N_3153);
or U3879 (N_3879,N_3586,N_3256);
xnor U3880 (N_3880,N_3240,N_3331);
nand U3881 (N_3881,N_3178,N_3285);
nand U3882 (N_3882,N_3393,N_3552);
nand U3883 (N_3883,N_3419,N_3114);
nor U3884 (N_3884,N_3305,N_3346);
and U3885 (N_3885,N_3189,N_3483);
and U3886 (N_3886,N_3540,N_3548);
or U3887 (N_3887,N_3485,N_3197);
and U3888 (N_3888,N_3263,N_3087);
and U3889 (N_3889,N_3229,N_3030);
and U3890 (N_3890,N_3506,N_3508);
xnor U3891 (N_3891,N_3573,N_3402);
xnor U3892 (N_3892,N_3098,N_3327);
xor U3893 (N_3893,N_3378,N_3133);
xnor U3894 (N_3894,N_3078,N_3377);
or U3895 (N_3895,N_3453,N_3422);
nor U3896 (N_3896,N_3476,N_3362);
and U3897 (N_3897,N_3349,N_3294);
xnor U3898 (N_3898,N_3486,N_3120);
and U3899 (N_3899,N_3451,N_3523);
and U3900 (N_3900,N_3098,N_3397);
nor U3901 (N_3901,N_3488,N_3191);
and U3902 (N_3902,N_3422,N_3172);
nor U3903 (N_3903,N_3022,N_3584);
nand U3904 (N_3904,N_3081,N_3547);
xor U3905 (N_3905,N_3295,N_3128);
and U3906 (N_3906,N_3358,N_3089);
and U3907 (N_3907,N_3455,N_3214);
nand U3908 (N_3908,N_3115,N_3344);
nor U3909 (N_3909,N_3303,N_3562);
or U3910 (N_3910,N_3382,N_3513);
xnor U3911 (N_3911,N_3553,N_3049);
nor U3912 (N_3912,N_3460,N_3409);
or U3913 (N_3913,N_3311,N_3107);
nand U3914 (N_3914,N_3356,N_3348);
nor U3915 (N_3915,N_3146,N_3096);
nand U3916 (N_3916,N_3106,N_3360);
and U3917 (N_3917,N_3097,N_3117);
nand U3918 (N_3918,N_3012,N_3582);
nor U3919 (N_3919,N_3168,N_3202);
xor U3920 (N_3920,N_3599,N_3038);
nor U3921 (N_3921,N_3072,N_3082);
and U3922 (N_3922,N_3460,N_3555);
xnor U3923 (N_3923,N_3592,N_3586);
and U3924 (N_3924,N_3382,N_3597);
or U3925 (N_3925,N_3040,N_3523);
nand U3926 (N_3926,N_3167,N_3592);
nand U3927 (N_3927,N_3411,N_3033);
and U3928 (N_3928,N_3141,N_3475);
or U3929 (N_3929,N_3527,N_3177);
nor U3930 (N_3930,N_3183,N_3174);
nand U3931 (N_3931,N_3001,N_3385);
xnor U3932 (N_3932,N_3111,N_3201);
nor U3933 (N_3933,N_3260,N_3185);
nor U3934 (N_3934,N_3142,N_3479);
nor U3935 (N_3935,N_3196,N_3270);
nor U3936 (N_3936,N_3382,N_3586);
nand U3937 (N_3937,N_3308,N_3028);
and U3938 (N_3938,N_3275,N_3228);
nand U3939 (N_3939,N_3458,N_3421);
or U3940 (N_3940,N_3316,N_3272);
or U3941 (N_3941,N_3238,N_3543);
or U3942 (N_3942,N_3375,N_3192);
xor U3943 (N_3943,N_3477,N_3137);
or U3944 (N_3944,N_3218,N_3537);
or U3945 (N_3945,N_3319,N_3479);
xor U3946 (N_3946,N_3489,N_3349);
nor U3947 (N_3947,N_3316,N_3389);
nor U3948 (N_3948,N_3314,N_3219);
xor U3949 (N_3949,N_3304,N_3538);
nand U3950 (N_3950,N_3139,N_3318);
xor U3951 (N_3951,N_3518,N_3051);
xnor U3952 (N_3952,N_3158,N_3560);
nor U3953 (N_3953,N_3496,N_3318);
or U3954 (N_3954,N_3578,N_3554);
nor U3955 (N_3955,N_3296,N_3591);
nor U3956 (N_3956,N_3557,N_3445);
xor U3957 (N_3957,N_3096,N_3536);
xor U3958 (N_3958,N_3114,N_3167);
xnor U3959 (N_3959,N_3417,N_3175);
nor U3960 (N_3960,N_3385,N_3553);
or U3961 (N_3961,N_3565,N_3433);
nor U3962 (N_3962,N_3265,N_3289);
xnor U3963 (N_3963,N_3109,N_3545);
and U3964 (N_3964,N_3032,N_3532);
nand U3965 (N_3965,N_3516,N_3360);
nor U3966 (N_3966,N_3594,N_3237);
xnor U3967 (N_3967,N_3140,N_3514);
or U3968 (N_3968,N_3259,N_3227);
xnor U3969 (N_3969,N_3411,N_3051);
and U3970 (N_3970,N_3426,N_3209);
and U3971 (N_3971,N_3102,N_3170);
or U3972 (N_3972,N_3310,N_3534);
nand U3973 (N_3973,N_3073,N_3171);
xor U3974 (N_3974,N_3548,N_3169);
and U3975 (N_3975,N_3408,N_3070);
or U3976 (N_3976,N_3391,N_3392);
or U3977 (N_3977,N_3310,N_3013);
nor U3978 (N_3978,N_3000,N_3067);
nor U3979 (N_3979,N_3348,N_3554);
and U3980 (N_3980,N_3497,N_3164);
xor U3981 (N_3981,N_3596,N_3273);
or U3982 (N_3982,N_3308,N_3451);
nand U3983 (N_3983,N_3229,N_3078);
or U3984 (N_3984,N_3003,N_3048);
and U3985 (N_3985,N_3321,N_3049);
nand U3986 (N_3986,N_3588,N_3573);
and U3987 (N_3987,N_3093,N_3390);
nor U3988 (N_3988,N_3591,N_3471);
xnor U3989 (N_3989,N_3323,N_3325);
or U3990 (N_3990,N_3317,N_3584);
nand U3991 (N_3991,N_3551,N_3311);
and U3992 (N_3992,N_3144,N_3377);
or U3993 (N_3993,N_3390,N_3546);
nor U3994 (N_3994,N_3357,N_3304);
nor U3995 (N_3995,N_3104,N_3164);
or U3996 (N_3996,N_3589,N_3314);
xnor U3997 (N_3997,N_3139,N_3410);
nor U3998 (N_3998,N_3338,N_3298);
xnor U3999 (N_3999,N_3456,N_3581);
or U4000 (N_4000,N_3489,N_3101);
or U4001 (N_4001,N_3391,N_3403);
and U4002 (N_4002,N_3177,N_3343);
nor U4003 (N_4003,N_3192,N_3227);
and U4004 (N_4004,N_3226,N_3597);
nor U4005 (N_4005,N_3109,N_3506);
nor U4006 (N_4006,N_3537,N_3318);
nor U4007 (N_4007,N_3326,N_3413);
and U4008 (N_4008,N_3379,N_3166);
xor U4009 (N_4009,N_3560,N_3286);
xnor U4010 (N_4010,N_3355,N_3491);
and U4011 (N_4011,N_3541,N_3468);
xnor U4012 (N_4012,N_3474,N_3347);
and U4013 (N_4013,N_3283,N_3324);
nor U4014 (N_4014,N_3334,N_3252);
nor U4015 (N_4015,N_3126,N_3106);
or U4016 (N_4016,N_3165,N_3281);
xor U4017 (N_4017,N_3549,N_3011);
nor U4018 (N_4018,N_3049,N_3146);
or U4019 (N_4019,N_3292,N_3448);
nand U4020 (N_4020,N_3404,N_3486);
xor U4021 (N_4021,N_3076,N_3180);
nor U4022 (N_4022,N_3312,N_3262);
and U4023 (N_4023,N_3162,N_3362);
xnor U4024 (N_4024,N_3297,N_3598);
nand U4025 (N_4025,N_3245,N_3055);
nor U4026 (N_4026,N_3201,N_3506);
and U4027 (N_4027,N_3347,N_3269);
xnor U4028 (N_4028,N_3404,N_3193);
or U4029 (N_4029,N_3379,N_3266);
nand U4030 (N_4030,N_3335,N_3534);
nand U4031 (N_4031,N_3083,N_3091);
xnor U4032 (N_4032,N_3457,N_3350);
nand U4033 (N_4033,N_3486,N_3356);
nand U4034 (N_4034,N_3269,N_3259);
and U4035 (N_4035,N_3133,N_3429);
or U4036 (N_4036,N_3573,N_3232);
or U4037 (N_4037,N_3063,N_3220);
and U4038 (N_4038,N_3425,N_3131);
nor U4039 (N_4039,N_3527,N_3484);
or U4040 (N_4040,N_3468,N_3308);
and U4041 (N_4041,N_3318,N_3075);
and U4042 (N_4042,N_3114,N_3299);
nand U4043 (N_4043,N_3267,N_3142);
nor U4044 (N_4044,N_3294,N_3173);
nor U4045 (N_4045,N_3551,N_3416);
nand U4046 (N_4046,N_3174,N_3296);
and U4047 (N_4047,N_3089,N_3409);
and U4048 (N_4048,N_3371,N_3403);
or U4049 (N_4049,N_3351,N_3324);
and U4050 (N_4050,N_3507,N_3034);
and U4051 (N_4051,N_3223,N_3585);
and U4052 (N_4052,N_3555,N_3372);
xnor U4053 (N_4053,N_3135,N_3464);
nor U4054 (N_4054,N_3565,N_3357);
nor U4055 (N_4055,N_3102,N_3079);
and U4056 (N_4056,N_3541,N_3146);
or U4057 (N_4057,N_3099,N_3461);
xor U4058 (N_4058,N_3565,N_3364);
and U4059 (N_4059,N_3378,N_3171);
xor U4060 (N_4060,N_3543,N_3205);
nor U4061 (N_4061,N_3272,N_3147);
nand U4062 (N_4062,N_3508,N_3575);
and U4063 (N_4063,N_3430,N_3369);
or U4064 (N_4064,N_3552,N_3452);
xor U4065 (N_4065,N_3068,N_3130);
nand U4066 (N_4066,N_3475,N_3162);
or U4067 (N_4067,N_3177,N_3389);
nor U4068 (N_4068,N_3028,N_3016);
nor U4069 (N_4069,N_3136,N_3294);
or U4070 (N_4070,N_3343,N_3166);
xnor U4071 (N_4071,N_3476,N_3029);
xnor U4072 (N_4072,N_3185,N_3013);
and U4073 (N_4073,N_3093,N_3535);
nand U4074 (N_4074,N_3413,N_3377);
and U4075 (N_4075,N_3413,N_3335);
and U4076 (N_4076,N_3364,N_3285);
nand U4077 (N_4077,N_3371,N_3130);
nand U4078 (N_4078,N_3436,N_3448);
xnor U4079 (N_4079,N_3447,N_3383);
xor U4080 (N_4080,N_3326,N_3320);
xnor U4081 (N_4081,N_3109,N_3174);
nand U4082 (N_4082,N_3460,N_3590);
xor U4083 (N_4083,N_3076,N_3285);
and U4084 (N_4084,N_3230,N_3154);
nor U4085 (N_4085,N_3071,N_3502);
or U4086 (N_4086,N_3598,N_3188);
and U4087 (N_4087,N_3090,N_3157);
and U4088 (N_4088,N_3478,N_3348);
xor U4089 (N_4089,N_3517,N_3570);
nor U4090 (N_4090,N_3022,N_3403);
and U4091 (N_4091,N_3037,N_3433);
nor U4092 (N_4092,N_3562,N_3547);
or U4093 (N_4093,N_3152,N_3149);
xnor U4094 (N_4094,N_3119,N_3293);
nand U4095 (N_4095,N_3061,N_3599);
or U4096 (N_4096,N_3513,N_3174);
nor U4097 (N_4097,N_3241,N_3177);
xor U4098 (N_4098,N_3099,N_3170);
and U4099 (N_4099,N_3063,N_3296);
nand U4100 (N_4100,N_3412,N_3532);
nor U4101 (N_4101,N_3435,N_3082);
nor U4102 (N_4102,N_3018,N_3010);
xor U4103 (N_4103,N_3012,N_3527);
nor U4104 (N_4104,N_3135,N_3333);
and U4105 (N_4105,N_3499,N_3204);
and U4106 (N_4106,N_3246,N_3348);
or U4107 (N_4107,N_3336,N_3527);
xnor U4108 (N_4108,N_3059,N_3459);
xor U4109 (N_4109,N_3196,N_3277);
or U4110 (N_4110,N_3493,N_3142);
nor U4111 (N_4111,N_3590,N_3376);
or U4112 (N_4112,N_3441,N_3014);
nor U4113 (N_4113,N_3578,N_3424);
or U4114 (N_4114,N_3414,N_3533);
or U4115 (N_4115,N_3530,N_3097);
and U4116 (N_4116,N_3358,N_3577);
nor U4117 (N_4117,N_3123,N_3075);
nand U4118 (N_4118,N_3160,N_3100);
or U4119 (N_4119,N_3176,N_3536);
and U4120 (N_4120,N_3002,N_3334);
nor U4121 (N_4121,N_3593,N_3074);
nor U4122 (N_4122,N_3419,N_3597);
nor U4123 (N_4123,N_3454,N_3186);
and U4124 (N_4124,N_3403,N_3439);
nand U4125 (N_4125,N_3265,N_3426);
nor U4126 (N_4126,N_3384,N_3454);
and U4127 (N_4127,N_3335,N_3319);
nand U4128 (N_4128,N_3522,N_3415);
or U4129 (N_4129,N_3510,N_3186);
nor U4130 (N_4130,N_3541,N_3593);
and U4131 (N_4131,N_3386,N_3258);
or U4132 (N_4132,N_3125,N_3116);
nand U4133 (N_4133,N_3177,N_3087);
and U4134 (N_4134,N_3422,N_3436);
xor U4135 (N_4135,N_3235,N_3510);
nor U4136 (N_4136,N_3593,N_3447);
and U4137 (N_4137,N_3537,N_3004);
xor U4138 (N_4138,N_3416,N_3152);
and U4139 (N_4139,N_3209,N_3300);
xnor U4140 (N_4140,N_3575,N_3143);
nand U4141 (N_4141,N_3128,N_3550);
nand U4142 (N_4142,N_3443,N_3382);
xor U4143 (N_4143,N_3173,N_3074);
and U4144 (N_4144,N_3206,N_3371);
or U4145 (N_4145,N_3369,N_3479);
nand U4146 (N_4146,N_3489,N_3351);
or U4147 (N_4147,N_3408,N_3109);
and U4148 (N_4148,N_3553,N_3220);
nand U4149 (N_4149,N_3544,N_3415);
and U4150 (N_4150,N_3276,N_3465);
and U4151 (N_4151,N_3004,N_3391);
or U4152 (N_4152,N_3241,N_3013);
nand U4153 (N_4153,N_3373,N_3595);
xnor U4154 (N_4154,N_3164,N_3076);
xor U4155 (N_4155,N_3294,N_3582);
nor U4156 (N_4156,N_3334,N_3358);
xor U4157 (N_4157,N_3440,N_3014);
nor U4158 (N_4158,N_3146,N_3456);
nor U4159 (N_4159,N_3271,N_3470);
and U4160 (N_4160,N_3068,N_3134);
or U4161 (N_4161,N_3417,N_3302);
and U4162 (N_4162,N_3173,N_3254);
and U4163 (N_4163,N_3282,N_3331);
nand U4164 (N_4164,N_3517,N_3181);
or U4165 (N_4165,N_3067,N_3239);
or U4166 (N_4166,N_3317,N_3122);
or U4167 (N_4167,N_3243,N_3363);
and U4168 (N_4168,N_3567,N_3358);
xnor U4169 (N_4169,N_3336,N_3050);
and U4170 (N_4170,N_3587,N_3458);
xnor U4171 (N_4171,N_3046,N_3105);
xnor U4172 (N_4172,N_3246,N_3411);
xnor U4173 (N_4173,N_3564,N_3567);
nor U4174 (N_4174,N_3428,N_3382);
or U4175 (N_4175,N_3552,N_3326);
xnor U4176 (N_4176,N_3154,N_3299);
nand U4177 (N_4177,N_3167,N_3357);
or U4178 (N_4178,N_3144,N_3451);
nor U4179 (N_4179,N_3052,N_3433);
and U4180 (N_4180,N_3153,N_3309);
or U4181 (N_4181,N_3140,N_3225);
or U4182 (N_4182,N_3469,N_3238);
nand U4183 (N_4183,N_3456,N_3331);
xnor U4184 (N_4184,N_3464,N_3060);
or U4185 (N_4185,N_3159,N_3597);
and U4186 (N_4186,N_3560,N_3247);
and U4187 (N_4187,N_3107,N_3100);
nor U4188 (N_4188,N_3408,N_3493);
nand U4189 (N_4189,N_3114,N_3427);
nor U4190 (N_4190,N_3296,N_3126);
nor U4191 (N_4191,N_3501,N_3303);
nand U4192 (N_4192,N_3558,N_3212);
xnor U4193 (N_4193,N_3321,N_3368);
xnor U4194 (N_4194,N_3312,N_3465);
nand U4195 (N_4195,N_3473,N_3056);
nand U4196 (N_4196,N_3587,N_3334);
nand U4197 (N_4197,N_3257,N_3322);
nor U4198 (N_4198,N_3471,N_3068);
and U4199 (N_4199,N_3159,N_3205);
and U4200 (N_4200,N_3717,N_4035);
xnor U4201 (N_4201,N_4185,N_3987);
and U4202 (N_4202,N_3664,N_4013);
and U4203 (N_4203,N_3866,N_3846);
nand U4204 (N_4204,N_3756,N_3891);
and U4205 (N_4205,N_3665,N_4106);
or U4206 (N_4206,N_4045,N_4002);
xnor U4207 (N_4207,N_4149,N_3610);
nor U4208 (N_4208,N_3948,N_4082);
and U4209 (N_4209,N_3822,N_3649);
xor U4210 (N_4210,N_3735,N_4078);
xnor U4211 (N_4211,N_3788,N_3787);
or U4212 (N_4212,N_3913,N_3967);
xnor U4213 (N_4213,N_3950,N_4086);
xnor U4214 (N_4214,N_4003,N_3922);
nand U4215 (N_4215,N_4054,N_4069);
or U4216 (N_4216,N_3994,N_3900);
or U4217 (N_4217,N_4197,N_3702);
nand U4218 (N_4218,N_3766,N_4148);
and U4219 (N_4219,N_4083,N_3616);
xor U4220 (N_4220,N_3736,N_4088);
nand U4221 (N_4221,N_4066,N_3984);
nand U4222 (N_4222,N_3689,N_3957);
or U4223 (N_4223,N_3751,N_3976);
and U4224 (N_4224,N_3731,N_3612);
and U4225 (N_4225,N_4025,N_3601);
nor U4226 (N_4226,N_3892,N_4181);
and U4227 (N_4227,N_3924,N_3627);
nor U4228 (N_4228,N_3739,N_3770);
and U4229 (N_4229,N_3973,N_4028);
and U4230 (N_4230,N_3843,N_3602);
or U4231 (N_4231,N_3930,N_3647);
nand U4232 (N_4232,N_3865,N_3870);
or U4233 (N_4233,N_3943,N_3896);
xor U4234 (N_4234,N_3841,N_4107);
or U4235 (N_4235,N_3845,N_3884);
or U4236 (N_4236,N_4017,N_3722);
xor U4237 (N_4237,N_4116,N_3942);
and U4238 (N_4238,N_3615,N_3693);
or U4239 (N_4239,N_3810,N_4122);
xor U4240 (N_4240,N_3772,N_3874);
and U4241 (N_4241,N_3868,N_4170);
nand U4242 (N_4242,N_4022,N_4060);
or U4243 (N_4243,N_4141,N_4196);
or U4244 (N_4244,N_4135,N_3740);
and U4245 (N_4245,N_3911,N_4043);
xor U4246 (N_4246,N_3919,N_3645);
nand U4247 (N_4247,N_4194,N_4114);
nand U4248 (N_4248,N_3652,N_3655);
and U4249 (N_4249,N_3659,N_4038);
and U4250 (N_4250,N_3904,N_4010);
nand U4251 (N_4251,N_4031,N_3691);
nand U4252 (N_4252,N_3660,N_4128);
and U4253 (N_4253,N_4095,N_3672);
xor U4254 (N_4254,N_4130,N_4187);
nand U4255 (N_4255,N_3642,N_3630);
nand U4256 (N_4256,N_3864,N_3949);
or U4257 (N_4257,N_3638,N_3928);
nand U4258 (N_4258,N_4015,N_4112);
nor U4259 (N_4259,N_3695,N_3869);
or U4260 (N_4260,N_4072,N_4090);
nand U4261 (N_4261,N_4065,N_3859);
or U4262 (N_4262,N_3901,N_3873);
xnor U4263 (N_4263,N_4137,N_3975);
xnor U4264 (N_4264,N_4008,N_4174);
xor U4265 (N_4265,N_3726,N_3754);
or U4266 (N_4266,N_3785,N_3643);
or U4267 (N_4267,N_3879,N_4146);
xor U4268 (N_4268,N_3636,N_3742);
nor U4269 (N_4269,N_3666,N_4100);
or U4270 (N_4270,N_4094,N_4076);
xor U4271 (N_4271,N_3600,N_4092);
nor U4272 (N_4272,N_3966,N_4063);
xnor U4273 (N_4273,N_4004,N_4189);
nor U4274 (N_4274,N_3906,N_3982);
nand U4275 (N_4275,N_4079,N_4037);
nand U4276 (N_4276,N_3737,N_4198);
xnor U4277 (N_4277,N_4191,N_3799);
and U4278 (N_4278,N_3923,N_4144);
nand U4279 (N_4279,N_3881,N_3708);
xnor U4280 (N_4280,N_4177,N_3793);
or U4281 (N_4281,N_4160,N_3686);
and U4282 (N_4282,N_4000,N_3993);
nand U4283 (N_4283,N_3831,N_4140);
nor U4284 (N_4284,N_3953,N_4009);
nor U4285 (N_4285,N_4077,N_3646);
and U4286 (N_4286,N_3741,N_4166);
nor U4287 (N_4287,N_3607,N_3935);
or U4288 (N_4288,N_3821,N_4154);
xor U4289 (N_4289,N_4131,N_3794);
nor U4290 (N_4290,N_3764,N_3803);
xor U4291 (N_4291,N_3941,N_4171);
xor U4292 (N_4292,N_4162,N_3974);
xnor U4293 (N_4293,N_3947,N_3637);
and U4294 (N_4294,N_3675,N_4121);
xor U4295 (N_4295,N_3639,N_4005);
xnor U4296 (N_4296,N_3763,N_3914);
or U4297 (N_4297,N_4142,N_4178);
nor U4298 (N_4298,N_4110,N_4026);
or U4299 (N_4299,N_3789,N_3872);
or U4300 (N_4300,N_3700,N_3828);
nor U4301 (N_4301,N_3867,N_3680);
and U4302 (N_4302,N_3929,N_3832);
or U4303 (N_4303,N_4019,N_3743);
xor U4304 (N_4304,N_4195,N_4097);
nand U4305 (N_4305,N_4176,N_4012);
nand U4306 (N_4306,N_3813,N_4071);
nand U4307 (N_4307,N_4027,N_3997);
nor U4308 (N_4308,N_3818,N_3698);
nand U4309 (N_4309,N_3651,N_3815);
nand U4310 (N_4310,N_3856,N_3768);
nand U4311 (N_4311,N_3678,N_3852);
and U4312 (N_4312,N_3885,N_4042);
nor U4313 (N_4313,N_3747,N_4024);
nor U4314 (N_4314,N_4052,N_3724);
xnor U4315 (N_4315,N_3980,N_3677);
nor U4316 (N_4316,N_4123,N_3902);
xnor U4317 (N_4317,N_3862,N_3886);
xor U4318 (N_4318,N_3844,N_3688);
or U4319 (N_4319,N_3728,N_4074);
or U4320 (N_4320,N_3623,N_3851);
nand U4321 (N_4321,N_4014,N_4108);
nand U4322 (N_4322,N_4081,N_3632);
xor U4323 (N_4323,N_4132,N_3959);
nor U4324 (N_4324,N_3985,N_3738);
nand U4325 (N_4325,N_3807,N_3916);
xnor U4326 (N_4326,N_3762,N_3991);
and U4327 (N_4327,N_3781,N_4030);
and U4328 (N_4328,N_4041,N_4039);
and U4329 (N_4329,N_4125,N_3628);
nand U4330 (N_4330,N_3779,N_4073);
nand U4331 (N_4331,N_4186,N_3617);
nor U4332 (N_4332,N_3667,N_3979);
xnor U4333 (N_4333,N_3988,N_3631);
and U4334 (N_4334,N_4057,N_3806);
xor U4335 (N_4335,N_4127,N_3661);
nand U4336 (N_4336,N_4151,N_4175);
and U4337 (N_4337,N_4085,N_3909);
nand U4338 (N_4338,N_4104,N_3671);
nor U4339 (N_4339,N_4118,N_3709);
nand U4340 (N_4340,N_3774,N_3907);
and U4341 (N_4341,N_3790,N_3719);
nor U4342 (N_4342,N_3965,N_3771);
xnor U4343 (N_4343,N_3658,N_4034);
and U4344 (N_4344,N_3773,N_3725);
xnor U4345 (N_4345,N_3877,N_3895);
or U4346 (N_4346,N_3836,N_3707);
and U4347 (N_4347,N_4109,N_3710);
nand U4348 (N_4348,N_3972,N_3621);
and U4349 (N_4349,N_3669,N_4029);
or U4350 (N_4350,N_3618,N_3931);
nor U4351 (N_4351,N_3795,N_3955);
nor U4352 (N_4352,N_3687,N_3606);
or U4353 (N_4353,N_3977,N_4099);
or U4354 (N_4354,N_3921,N_4150);
and U4355 (N_4355,N_3752,N_3854);
and U4356 (N_4356,N_3641,N_3937);
nand U4357 (N_4357,N_4093,N_3760);
xnor U4358 (N_4358,N_4064,N_3603);
and U4359 (N_4359,N_3918,N_4105);
xor U4360 (N_4360,N_3634,N_3926);
nand U4361 (N_4361,N_3826,N_3614);
nor U4362 (N_4362,N_3681,N_3734);
xor U4363 (N_4363,N_3920,N_3968);
nand U4364 (N_4364,N_3940,N_3712);
xor U4365 (N_4365,N_4129,N_4138);
nand U4366 (N_4366,N_4193,N_4070);
and U4367 (N_4367,N_3780,N_3871);
xor U4368 (N_4368,N_4169,N_3858);
nand U4369 (N_4369,N_3855,N_3750);
or U4370 (N_4370,N_4059,N_4120);
xnor U4371 (N_4371,N_4001,N_3847);
xor U4372 (N_4372,N_3932,N_3744);
and U4373 (N_4373,N_3808,N_3765);
or U4374 (N_4374,N_3767,N_3829);
nand U4375 (N_4375,N_3668,N_3888);
nand U4376 (N_4376,N_3823,N_4040);
xnor U4377 (N_4377,N_3848,N_3833);
and U4378 (N_4378,N_3696,N_3777);
xor U4379 (N_4379,N_3811,N_4192);
and U4380 (N_4380,N_4155,N_4020);
nand U4381 (N_4381,N_3620,N_3798);
nor U4382 (N_4382,N_3969,N_4096);
or U4383 (N_4383,N_4068,N_4152);
and U4384 (N_4384,N_3624,N_3662);
nand U4385 (N_4385,N_3746,N_3878);
or U4386 (N_4386,N_3897,N_4180);
nor U4387 (N_4387,N_3999,N_3748);
or U4388 (N_4388,N_3648,N_3983);
xnor U4389 (N_4389,N_4033,N_3749);
xor U4390 (N_4390,N_4133,N_4048);
nand U4391 (N_4391,N_3755,N_3730);
or U4392 (N_4392,N_3653,N_3608);
or U4393 (N_4393,N_4143,N_3758);
and U4394 (N_4394,N_4053,N_3805);
nor U4395 (N_4395,N_4156,N_3650);
nor U4396 (N_4396,N_3804,N_3611);
and U4397 (N_4397,N_4134,N_3761);
nand U4398 (N_4398,N_3654,N_3729);
or U4399 (N_4399,N_3899,N_3694);
xnor U4400 (N_4400,N_4190,N_3908);
nor U4401 (N_4401,N_3640,N_3989);
or U4402 (N_4402,N_4006,N_3990);
and U4403 (N_4403,N_3697,N_3715);
or U4404 (N_4404,N_4016,N_3626);
and U4405 (N_4405,N_3850,N_4145);
and U4406 (N_4406,N_3721,N_3622);
nor U4407 (N_4407,N_3759,N_3882);
or U4408 (N_4408,N_4113,N_4050);
or U4409 (N_4409,N_3946,N_3625);
or U4410 (N_4410,N_3819,N_3915);
or U4411 (N_4411,N_3889,N_3961);
or U4412 (N_4412,N_3863,N_4182);
or U4413 (N_4413,N_4139,N_3676);
or U4414 (N_4414,N_3732,N_3861);
nand U4415 (N_4415,N_3786,N_4055);
or U4416 (N_4416,N_4044,N_4172);
nand U4417 (N_4417,N_3692,N_3934);
and U4418 (N_4418,N_4167,N_3938);
nand U4419 (N_4419,N_3784,N_4089);
nor U4420 (N_4420,N_3883,N_4087);
and U4421 (N_4421,N_3998,N_3830);
nor U4422 (N_4422,N_3842,N_4183);
nand U4423 (N_4423,N_4056,N_4188);
xor U4424 (N_4424,N_3825,N_3939);
nor U4425 (N_4425,N_4179,N_3605);
and U4426 (N_4426,N_3894,N_3701);
nand U4427 (N_4427,N_3933,N_4051);
xnor U4428 (N_4428,N_3682,N_3778);
and U4429 (N_4429,N_4098,N_3705);
and U4430 (N_4430,N_3797,N_3776);
xor U4431 (N_4431,N_3753,N_3876);
and U4432 (N_4432,N_3782,N_3917);
or U4433 (N_4433,N_3820,N_4018);
or U4434 (N_4434,N_4061,N_4119);
or U4435 (N_4435,N_3952,N_4126);
xnor U4436 (N_4436,N_3995,N_4136);
xnor U4437 (N_4437,N_3714,N_3898);
or U4438 (N_4438,N_3853,N_3690);
nor U4439 (N_4439,N_3887,N_3809);
and U4440 (N_4440,N_4023,N_3962);
and U4441 (N_4441,N_3733,N_3633);
xor U4442 (N_4442,N_3880,N_4199);
nor U4443 (N_4443,N_3910,N_4147);
xnor U4444 (N_4444,N_3604,N_4117);
xor U4445 (N_4445,N_3912,N_3699);
xor U4446 (N_4446,N_3890,N_3860);
xnor U4447 (N_4447,N_3963,N_3849);
nand U4448 (N_4448,N_3775,N_3663);
or U4449 (N_4449,N_3679,N_3857);
xor U4450 (N_4450,N_3657,N_3656);
or U4451 (N_4451,N_4058,N_3817);
nor U4452 (N_4452,N_3703,N_3893);
or U4453 (N_4453,N_4159,N_4047);
and U4454 (N_4454,N_3816,N_3981);
and U4455 (N_4455,N_4080,N_3796);
nand U4456 (N_4456,N_4184,N_3619);
nand U4457 (N_4457,N_4157,N_4032);
nand U4458 (N_4458,N_3684,N_3840);
nand U4459 (N_4459,N_3951,N_4062);
xnor U4460 (N_4460,N_3683,N_3903);
xnor U4461 (N_4461,N_3720,N_3769);
nor U4462 (N_4462,N_4046,N_4124);
xnor U4463 (N_4463,N_3716,N_4158);
and U4464 (N_4464,N_4067,N_3670);
nor U4465 (N_4465,N_4161,N_3644);
nand U4466 (N_4466,N_3970,N_3783);
nor U4467 (N_4467,N_4075,N_4168);
and U4468 (N_4468,N_3727,N_3945);
or U4469 (N_4469,N_3814,N_3838);
or U4470 (N_4470,N_3875,N_3824);
nand U4471 (N_4471,N_4102,N_4036);
nand U4472 (N_4472,N_4103,N_3685);
nor U4473 (N_4473,N_4091,N_3837);
and U4474 (N_4474,N_4115,N_3812);
xnor U4475 (N_4475,N_4011,N_3834);
xnor U4476 (N_4476,N_3954,N_3927);
or U4477 (N_4477,N_3706,N_3723);
and U4478 (N_4478,N_3792,N_3801);
or U4479 (N_4479,N_4049,N_4173);
xor U4480 (N_4480,N_3613,N_3704);
and U4481 (N_4481,N_3673,N_3986);
nor U4482 (N_4482,N_3791,N_3971);
nand U4483 (N_4483,N_3996,N_3800);
nor U4484 (N_4484,N_3958,N_3674);
xnor U4485 (N_4485,N_3960,N_4084);
or U4486 (N_4486,N_3964,N_3711);
nand U4487 (N_4487,N_4021,N_3718);
or U4488 (N_4488,N_3936,N_3713);
and U4489 (N_4489,N_3802,N_3745);
or U4490 (N_4490,N_3925,N_4163);
xnor U4491 (N_4491,N_3992,N_3835);
nor U4492 (N_4492,N_3978,N_3944);
nor U4493 (N_4493,N_3827,N_4101);
xnor U4494 (N_4494,N_3905,N_3629);
nand U4495 (N_4495,N_3635,N_4165);
nand U4496 (N_4496,N_3757,N_4164);
xnor U4497 (N_4497,N_3956,N_4153);
and U4498 (N_4498,N_4111,N_3609);
nor U4499 (N_4499,N_3839,N_4007);
nor U4500 (N_4500,N_3944,N_4166);
nand U4501 (N_4501,N_3691,N_3606);
xnor U4502 (N_4502,N_4036,N_3859);
nor U4503 (N_4503,N_3637,N_3937);
or U4504 (N_4504,N_4159,N_3755);
nor U4505 (N_4505,N_3703,N_3921);
nand U4506 (N_4506,N_4018,N_3772);
and U4507 (N_4507,N_3959,N_4022);
nand U4508 (N_4508,N_4097,N_3989);
xnor U4509 (N_4509,N_3825,N_4106);
nor U4510 (N_4510,N_4129,N_4024);
and U4511 (N_4511,N_3922,N_3974);
and U4512 (N_4512,N_3968,N_3795);
xnor U4513 (N_4513,N_3683,N_3805);
or U4514 (N_4514,N_4052,N_4121);
nor U4515 (N_4515,N_3631,N_4024);
nor U4516 (N_4516,N_3672,N_4076);
or U4517 (N_4517,N_3846,N_3835);
and U4518 (N_4518,N_3634,N_3784);
nand U4519 (N_4519,N_4027,N_4039);
nand U4520 (N_4520,N_3994,N_4027);
and U4521 (N_4521,N_3980,N_4130);
nor U4522 (N_4522,N_4135,N_3943);
nor U4523 (N_4523,N_3744,N_3844);
nor U4524 (N_4524,N_3927,N_4057);
nand U4525 (N_4525,N_3865,N_3906);
xnor U4526 (N_4526,N_3794,N_4024);
nand U4527 (N_4527,N_4165,N_3890);
xor U4528 (N_4528,N_4050,N_4143);
xnor U4529 (N_4529,N_3649,N_3700);
and U4530 (N_4530,N_4151,N_3611);
xor U4531 (N_4531,N_3905,N_4102);
nor U4532 (N_4532,N_4113,N_4019);
nand U4533 (N_4533,N_3946,N_3774);
and U4534 (N_4534,N_4015,N_3973);
nand U4535 (N_4535,N_4132,N_3683);
xnor U4536 (N_4536,N_3783,N_3774);
nor U4537 (N_4537,N_4060,N_4002);
and U4538 (N_4538,N_4153,N_3729);
xnor U4539 (N_4539,N_3839,N_3834);
or U4540 (N_4540,N_3804,N_3963);
nor U4541 (N_4541,N_4083,N_4054);
and U4542 (N_4542,N_3914,N_3747);
or U4543 (N_4543,N_4050,N_3686);
or U4544 (N_4544,N_4007,N_3707);
xor U4545 (N_4545,N_3634,N_4113);
or U4546 (N_4546,N_3722,N_4015);
nor U4547 (N_4547,N_3663,N_4090);
xnor U4548 (N_4548,N_4062,N_3903);
xor U4549 (N_4549,N_4162,N_4064);
nor U4550 (N_4550,N_4003,N_3783);
xor U4551 (N_4551,N_3995,N_4009);
nor U4552 (N_4552,N_3887,N_3838);
and U4553 (N_4553,N_3800,N_4016);
and U4554 (N_4554,N_4192,N_3790);
nor U4555 (N_4555,N_3738,N_4096);
nand U4556 (N_4556,N_3685,N_3643);
xnor U4557 (N_4557,N_3890,N_4171);
nand U4558 (N_4558,N_3751,N_4158);
and U4559 (N_4559,N_3671,N_4092);
and U4560 (N_4560,N_3859,N_3664);
nand U4561 (N_4561,N_4101,N_4174);
xnor U4562 (N_4562,N_3958,N_4150);
xnor U4563 (N_4563,N_3667,N_3649);
or U4564 (N_4564,N_3851,N_4069);
xor U4565 (N_4565,N_4143,N_3719);
xor U4566 (N_4566,N_4180,N_3878);
or U4567 (N_4567,N_3987,N_3992);
and U4568 (N_4568,N_3958,N_3826);
xor U4569 (N_4569,N_3842,N_4012);
xor U4570 (N_4570,N_3748,N_3636);
nor U4571 (N_4571,N_4061,N_3830);
xor U4572 (N_4572,N_3617,N_3974);
nor U4573 (N_4573,N_3733,N_3895);
nor U4574 (N_4574,N_3900,N_3714);
nand U4575 (N_4575,N_3736,N_3627);
and U4576 (N_4576,N_4176,N_3679);
and U4577 (N_4577,N_3975,N_4182);
and U4578 (N_4578,N_4153,N_3928);
and U4579 (N_4579,N_4114,N_4003);
nand U4580 (N_4580,N_4036,N_3692);
xnor U4581 (N_4581,N_3802,N_3985);
nand U4582 (N_4582,N_3935,N_4038);
xnor U4583 (N_4583,N_4082,N_3850);
xor U4584 (N_4584,N_3941,N_3783);
xor U4585 (N_4585,N_4086,N_3966);
nand U4586 (N_4586,N_3819,N_3880);
and U4587 (N_4587,N_3681,N_4124);
and U4588 (N_4588,N_3930,N_3798);
and U4589 (N_4589,N_4111,N_3928);
and U4590 (N_4590,N_4162,N_3746);
or U4591 (N_4591,N_3905,N_3723);
nand U4592 (N_4592,N_4192,N_3995);
nor U4593 (N_4593,N_3803,N_3704);
xor U4594 (N_4594,N_4014,N_3710);
nand U4595 (N_4595,N_3781,N_3971);
nor U4596 (N_4596,N_3699,N_4172);
xor U4597 (N_4597,N_4003,N_3770);
nor U4598 (N_4598,N_4077,N_3909);
nor U4599 (N_4599,N_3848,N_3973);
nand U4600 (N_4600,N_3772,N_3815);
nor U4601 (N_4601,N_3871,N_4050);
nand U4602 (N_4602,N_3804,N_3750);
nor U4603 (N_4603,N_4017,N_3791);
xor U4604 (N_4604,N_3915,N_3922);
and U4605 (N_4605,N_4091,N_4026);
or U4606 (N_4606,N_3670,N_3958);
nand U4607 (N_4607,N_3910,N_3922);
or U4608 (N_4608,N_4161,N_3950);
and U4609 (N_4609,N_4167,N_3651);
and U4610 (N_4610,N_4129,N_3755);
nand U4611 (N_4611,N_4123,N_4090);
nor U4612 (N_4612,N_3855,N_3905);
nor U4613 (N_4613,N_3712,N_3612);
nand U4614 (N_4614,N_4066,N_3657);
nor U4615 (N_4615,N_3822,N_3674);
nand U4616 (N_4616,N_3729,N_4084);
nor U4617 (N_4617,N_3817,N_3921);
xor U4618 (N_4618,N_3675,N_3836);
nand U4619 (N_4619,N_4189,N_3819);
and U4620 (N_4620,N_3757,N_3708);
nand U4621 (N_4621,N_3912,N_4198);
or U4622 (N_4622,N_3932,N_3875);
and U4623 (N_4623,N_3940,N_3779);
and U4624 (N_4624,N_3746,N_4068);
nor U4625 (N_4625,N_3827,N_3916);
nand U4626 (N_4626,N_4061,N_4107);
nand U4627 (N_4627,N_3849,N_3681);
xnor U4628 (N_4628,N_4058,N_4017);
and U4629 (N_4629,N_3872,N_3699);
nand U4630 (N_4630,N_4122,N_3925);
nor U4631 (N_4631,N_4003,N_3643);
nor U4632 (N_4632,N_3864,N_4171);
and U4633 (N_4633,N_3714,N_3747);
nor U4634 (N_4634,N_4141,N_3860);
or U4635 (N_4635,N_3926,N_4018);
or U4636 (N_4636,N_4024,N_3935);
nand U4637 (N_4637,N_3825,N_4045);
or U4638 (N_4638,N_4069,N_3755);
nor U4639 (N_4639,N_3845,N_4147);
or U4640 (N_4640,N_3681,N_3656);
nor U4641 (N_4641,N_3718,N_4041);
nor U4642 (N_4642,N_4055,N_3670);
xor U4643 (N_4643,N_3980,N_3972);
xnor U4644 (N_4644,N_3675,N_3986);
xnor U4645 (N_4645,N_3646,N_4140);
or U4646 (N_4646,N_4156,N_3741);
xnor U4647 (N_4647,N_3710,N_4191);
nor U4648 (N_4648,N_3927,N_4020);
xor U4649 (N_4649,N_3883,N_4172);
nor U4650 (N_4650,N_3971,N_3919);
and U4651 (N_4651,N_4082,N_3805);
or U4652 (N_4652,N_3840,N_4118);
xor U4653 (N_4653,N_3878,N_3763);
xor U4654 (N_4654,N_3663,N_4061);
nand U4655 (N_4655,N_3886,N_3939);
and U4656 (N_4656,N_3636,N_3738);
and U4657 (N_4657,N_4156,N_4158);
nand U4658 (N_4658,N_4174,N_3629);
nand U4659 (N_4659,N_3651,N_3691);
xor U4660 (N_4660,N_3699,N_3893);
nand U4661 (N_4661,N_3824,N_4051);
or U4662 (N_4662,N_3772,N_4014);
or U4663 (N_4663,N_4149,N_4157);
nand U4664 (N_4664,N_4065,N_4186);
nor U4665 (N_4665,N_3792,N_3667);
nor U4666 (N_4666,N_3899,N_4053);
or U4667 (N_4667,N_4057,N_3732);
or U4668 (N_4668,N_3988,N_3857);
nor U4669 (N_4669,N_3817,N_3823);
nor U4670 (N_4670,N_3903,N_3771);
xnor U4671 (N_4671,N_3932,N_3974);
nor U4672 (N_4672,N_3837,N_4019);
and U4673 (N_4673,N_3906,N_3782);
and U4674 (N_4674,N_3911,N_4065);
xnor U4675 (N_4675,N_4052,N_4110);
nor U4676 (N_4676,N_4033,N_3901);
or U4677 (N_4677,N_3949,N_3832);
or U4678 (N_4678,N_4150,N_4181);
or U4679 (N_4679,N_4157,N_3805);
nand U4680 (N_4680,N_3953,N_3618);
xor U4681 (N_4681,N_4035,N_4106);
nor U4682 (N_4682,N_4138,N_4105);
nand U4683 (N_4683,N_3920,N_3825);
xnor U4684 (N_4684,N_4013,N_3814);
or U4685 (N_4685,N_4102,N_4198);
xor U4686 (N_4686,N_3958,N_3875);
or U4687 (N_4687,N_4134,N_3698);
nor U4688 (N_4688,N_4061,N_3605);
and U4689 (N_4689,N_4097,N_4076);
xor U4690 (N_4690,N_3904,N_4170);
xor U4691 (N_4691,N_3640,N_4153);
nand U4692 (N_4692,N_3736,N_3852);
and U4693 (N_4693,N_3920,N_3646);
xnor U4694 (N_4694,N_3876,N_4013);
xnor U4695 (N_4695,N_4198,N_4010);
nand U4696 (N_4696,N_4058,N_4162);
xnor U4697 (N_4697,N_3825,N_3866);
xor U4698 (N_4698,N_4069,N_3893);
or U4699 (N_4699,N_3677,N_3715);
and U4700 (N_4700,N_4013,N_4190);
nor U4701 (N_4701,N_3627,N_4170);
nor U4702 (N_4702,N_3896,N_3706);
nand U4703 (N_4703,N_3780,N_3704);
nand U4704 (N_4704,N_3726,N_3894);
or U4705 (N_4705,N_3814,N_4069);
or U4706 (N_4706,N_3721,N_4087);
or U4707 (N_4707,N_3861,N_4123);
nand U4708 (N_4708,N_3743,N_3811);
xor U4709 (N_4709,N_4086,N_3601);
or U4710 (N_4710,N_3916,N_3837);
nand U4711 (N_4711,N_4199,N_3608);
nor U4712 (N_4712,N_3620,N_3857);
nand U4713 (N_4713,N_4078,N_3779);
nand U4714 (N_4714,N_3888,N_4149);
xnor U4715 (N_4715,N_3661,N_4184);
xnor U4716 (N_4716,N_4059,N_3868);
nand U4717 (N_4717,N_3844,N_3900);
or U4718 (N_4718,N_3873,N_4061);
or U4719 (N_4719,N_4097,N_3743);
xor U4720 (N_4720,N_3850,N_4059);
nor U4721 (N_4721,N_3963,N_3643);
and U4722 (N_4722,N_4187,N_3926);
nor U4723 (N_4723,N_3936,N_3682);
nand U4724 (N_4724,N_4006,N_3792);
nor U4725 (N_4725,N_3667,N_4009);
and U4726 (N_4726,N_3844,N_3782);
nand U4727 (N_4727,N_3838,N_3670);
nand U4728 (N_4728,N_3995,N_3886);
xor U4729 (N_4729,N_3787,N_3651);
and U4730 (N_4730,N_3613,N_4149);
and U4731 (N_4731,N_4129,N_4187);
and U4732 (N_4732,N_3892,N_3696);
nand U4733 (N_4733,N_3654,N_4145);
nand U4734 (N_4734,N_3784,N_4016);
nand U4735 (N_4735,N_3813,N_3723);
xnor U4736 (N_4736,N_3828,N_4174);
xnor U4737 (N_4737,N_3758,N_4178);
or U4738 (N_4738,N_3865,N_3619);
xnor U4739 (N_4739,N_3881,N_3843);
and U4740 (N_4740,N_3997,N_4154);
or U4741 (N_4741,N_3988,N_4083);
nand U4742 (N_4742,N_4003,N_3904);
or U4743 (N_4743,N_3746,N_4131);
nand U4744 (N_4744,N_3701,N_4002);
or U4745 (N_4745,N_3600,N_3766);
or U4746 (N_4746,N_3750,N_3623);
nand U4747 (N_4747,N_4121,N_3941);
and U4748 (N_4748,N_3691,N_3960);
xor U4749 (N_4749,N_3746,N_3818);
nand U4750 (N_4750,N_3939,N_4048);
nand U4751 (N_4751,N_3844,N_4150);
and U4752 (N_4752,N_3730,N_4191);
or U4753 (N_4753,N_3995,N_4180);
xnor U4754 (N_4754,N_4003,N_3624);
nand U4755 (N_4755,N_4162,N_3662);
or U4756 (N_4756,N_3994,N_3930);
or U4757 (N_4757,N_4161,N_3666);
nand U4758 (N_4758,N_4129,N_3743);
xor U4759 (N_4759,N_3760,N_3704);
or U4760 (N_4760,N_4115,N_3641);
nor U4761 (N_4761,N_4167,N_3801);
xor U4762 (N_4762,N_4064,N_3914);
nand U4763 (N_4763,N_4154,N_3765);
or U4764 (N_4764,N_3888,N_3925);
or U4765 (N_4765,N_4026,N_3693);
nor U4766 (N_4766,N_3753,N_3605);
and U4767 (N_4767,N_3665,N_4120);
xor U4768 (N_4768,N_4016,N_4050);
xor U4769 (N_4769,N_3721,N_3609);
xnor U4770 (N_4770,N_3894,N_3781);
or U4771 (N_4771,N_4112,N_3951);
and U4772 (N_4772,N_3951,N_4078);
nor U4773 (N_4773,N_4112,N_3631);
nor U4774 (N_4774,N_4032,N_3703);
and U4775 (N_4775,N_3959,N_3984);
nor U4776 (N_4776,N_3788,N_4152);
xor U4777 (N_4777,N_3842,N_4051);
and U4778 (N_4778,N_3948,N_3798);
and U4779 (N_4779,N_4102,N_3937);
or U4780 (N_4780,N_3826,N_4164);
nand U4781 (N_4781,N_3972,N_4157);
nand U4782 (N_4782,N_3810,N_3780);
nand U4783 (N_4783,N_3975,N_3816);
nor U4784 (N_4784,N_3916,N_3647);
or U4785 (N_4785,N_3707,N_4054);
or U4786 (N_4786,N_4184,N_3703);
and U4787 (N_4787,N_3600,N_3747);
or U4788 (N_4788,N_3600,N_4044);
or U4789 (N_4789,N_4036,N_3776);
xor U4790 (N_4790,N_3894,N_3999);
nor U4791 (N_4791,N_4115,N_3633);
xor U4792 (N_4792,N_3964,N_4062);
or U4793 (N_4793,N_3837,N_3784);
or U4794 (N_4794,N_3714,N_3706);
or U4795 (N_4795,N_4137,N_4115);
nor U4796 (N_4796,N_3637,N_3945);
and U4797 (N_4797,N_3851,N_3684);
xor U4798 (N_4798,N_3788,N_4146);
or U4799 (N_4799,N_3601,N_4162);
xnor U4800 (N_4800,N_4334,N_4488);
nor U4801 (N_4801,N_4264,N_4744);
nand U4802 (N_4802,N_4711,N_4709);
xor U4803 (N_4803,N_4246,N_4462);
or U4804 (N_4804,N_4511,N_4553);
and U4805 (N_4805,N_4693,N_4594);
and U4806 (N_4806,N_4662,N_4733);
xor U4807 (N_4807,N_4249,N_4208);
or U4808 (N_4808,N_4243,N_4395);
nor U4809 (N_4809,N_4292,N_4466);
nand U4810 (N_4810,N_4342,N_4298);
xnor U4811 (N_4811,N_4477,N_4384);
or U4812 (N_4812,N_4233,N_4541);
xor U4813 (N_4813,N_4286,N_4781);
nor U4814 (N_4814,N_4452,N_4371);
nor U4815 (N_4815,N_4281,N_4280);
and U4816 (N_4816,N_4418,N_4390);
xnor U4817 (N_4817,N_4603,N_4235);
nor U4818 (N_4818,N_4760,N_4643);
nand U4819 (N_4819,N_4649,N_4204);
nor U4820 (N_4820,N_4627,N_4473);
or U4821 (N_4821,N_4729,N_4338);
or U4822 (N_4822,N_4593,N_4561);
or U4823 (N_4823,N_4546,N_4383);
xor U4824 (N_4824,N_4721,N_4279);
xnor U4825 (N_4825,N_4312,N_4258);
or U4826 (N_4826,N_4524,N_4660);
nor U4827 (N_4827,N_4534,N_4588);
and U4828 (N_4828,N_4745,N_4317);
nor U4829 (N_4829,N_4429,N_4426);
nand U4830 (N_4830,N_4407,N_4444);
or U4831 (N_4831,N_4360,N_4658);
and U4832 (N_4832,N_4367,N_4387);
nand U4833 (N_4833,N_4295,N_4589);
nand U4834 (N_4834,N_4366,N_4691);
and U4835 (N_4835,N_4369,N_4346);
nor U4836 (N_4836,N_4726,N_4609);
nand U4837 (N_4837,N_4764,N_4372);
nor U4838 (N_4838,N_4758,N_4552);
nor U4839 (N_4839,N_4720,N_4459);
xor U4840 (N_4840,N_4463,N_4308);
xnor U4841 (N_4841,N_4499,N_4618);
or U4842 (N_4842,N_4613,N_4453);
xor U4843 (N_4843,N_4650,N_4778);
nand U4844 (N_4844,N_4261,N_4450);
and U4845 (N_4845,N_4419,N_4651);
nor U4846 (N_4846,N_4333,N_4748);
nor U4847 (N_4847,N_4297,N_4211);
or U4848 (N_4848,N_4277,N_4590);
nand U4849 (N_4849,N_4388,N_4700);
and U4850 (N_4850,N_4492,N_4275);
nor U4851 (N_4851,N_4447,N_4486);
xor U4852 (N_4852,N_4610,N_4697);
nor U4853 (N_4853,N_4451,N_4667);
nand U4854 (N_4854,N_4528,N_4596);
nand U4855 (N_4855,N_4519,N_4647);
nor U4856 (N_4856,N_4494,N_4508);
xnor U4857 (N_4857,N_4737,N_4248);
xnor U4858 (N_4858,N_4547,N_4227);
or U4859 (N_4859,N_4558,N_4740);
or U4860 (N_4860,N_4685,N_4717);
or U4861 (N_4861,N_4747,N_4457);
and U4862 (N_4862,N_4762,N_4584);
xor U4863 (N_4863,N_4202,N_4291);
or U4864 (N_4864,N_4708,N_4676);
nor U4865 (N_4865,N_4704,N_4795);
and U4866 (N_4866,N_4785,N_4771);
and U4867 (N_4867,N_4699,N_4485);
nor U4868 (N_4868,N_4670,N_4322);
xor U4869 (N_4869,N_4751,N_4430);
and U4870 (N_4870,N_4607,N_4644);
nand U4871 (N_4871,N_4784,N_4560);
nor U4872 (N_4872,N_4757,N_4501);
nor U4873 (N_4873,N_4329,N_4365);
nand U4874 (N_4874,N_4688,N_4648);
nand U4875 (N_4875,N_4780,N_4272);
nand U4876 (N_4876,N_4743,N_4398);
nand U4877 (N_4877,N_4544,N_4624);
xor U4878 (N_4878,N_4428,N_4496);
xor U4879 (N_4879,N_4305,N_4680);
nor U4880 (N_4880,N_4702,N_4682);
and U4881 (N_4881,N_4422,N_4380);
and U4882 (N_4882,N_4223,N_4537);
nor U4883 (N_4883,N_4514,N_4799);
and U4884 (N_4884,N_4331,N_4659);
and U4885 (N_4885,N_4504,N_4483);
xnor U4886 (N_4886,N_4516,N_4475);
nand U4887 (N_4887,N_4738,N_4563);
nand U4888 (N_4888,N_4414,N_4727);
and U4889 (N_4889,N_4472,N_4489);
nor U4890 (N_4890,N_4728,N_4340);
and U4891 (N_4891,N_4311,N_4424);
nand U4892 (N_4892,N_4569,N_4797);
or U4893 (N_4893,N_4361,N_4580);
nor U4894 (N_4894,N_4539,N_4262);
nand U4895 (N_4895,N_4595,N_4782);
nand U4896 (N_4896,N_4548,N_4374);
nor U4897 (N_4897,N_4621,N_4776);
or U4898 (N_4898,N_4756,N_4266);
and U4899 (N_4899,N_4313,N_4214);
and U4900 (N_4900,N_4455,N_4218);
and U4901 (N_4901,N_4671,N_4578);
xnor U4902 (N_4902,N_4723,N_4517);
xor U4903 (N_4903,N_4283,N_4399);
nor U4904 (N_4904,N_4349,N_4336);
nand U4905 (N_4905,N_4217,N_4495);
and U4906 (N_4906,N_4716,N_4210);
or U4907 (N_4907,N_4714,N_4343);
or U4908 (N_4908,N_4385,N_4386);
or U4909 (N_4909,N_4611,N_4479);
nand U4910 (N_4910,N_4456,N_4432);
nand U4911 (N_4911,N_4228,N_4646);
nor U4912 (N_4912,N_4521,N_4482);
and U4913 (N_4913,N_4545,N_4206);
nand U4914 (N_4914,N_4557,N_4410);
nand U4915 (N_4915,N_4656,N_4209);
or U4916 (N_4916,N_4412,N_4309);
nor U4917 (N_4917,N_4695,N_4765);
nand U4918 (N_4918,N_4420,N_4260);
or U4919 (N_4919,N_4710,N_4592);
nor U4920 (N_4920,N_4774,N_4348);
or U4921 (N_4921,N_4755,N_4379);
xnor U4922 (N_4922,N_4350,N_4319);
xnor U4923 (N_4923,N_4265,N_4318);
nand U4924 (N_4924,N_4294,N_4600);
nand U4925 (N_4925,N_4375,N_4427);
or U4926 (N_4926,N_4400,N_4612);
nor U4927 (N_4927,N_4796,N_4268);
nor U4928 (N_4928,N_4798,N_4619);
and U4929 (N_4929,N_4397,N_4257);
nor U4930 (N_4930,N_4622,N_4777);
and U4931 (N_4931,N_4351,N_4523);
xnor U4932 (N_4932,N_4289,N_4377);
nand U4933 (N_4933,N_4373,N_4672);
or U4934 (N_4934,N_4299,N_4635);
xnor U4935 (N_4935,N_4357,N_4454);
and U4936 (N_4936,N_4417,N_4431);
and U4937 (N_4937,N_4703,N_4527);
nor U4938 (N_4938,N_4789,N_4315);
xnor U4939 (N_4939,N_4719,N_4438);
or U4940 (N_4940,N_4555,N_4220);
and U4941 (N_4941,N_4241,N_4582);
xnor U4942 (N_4942,N_4389,N_4628);
xnor U4943 (N_4943,N_4677,N_4476);
nor U4944 (N_4944,N_4290,N_4363);
nand U4945 (N_4945,N_4436,N_4240);
or U4946 (N_4946,N_4421,N_4435);
and U4947 (N_4947,N_4219,N_4341);
nor U4948 (N_4948,N_4378,N_4730);
and U4949 (N_4949,N_4347,N_4411);
nor U4950 (N_4950,N_4376,N_4718);
and U4951 (N_4951,N_4330,N_4259);
xnor U4952 (N_4952,N_4274,N_4530);
nand U4953 (N_4953,N_4467,N_4254);
xnor U4954 (N_4954,N_4559,N_4657);
xnor U4955 (N_4955,N_4696,N_4679);
xor U4956 (N_4956,N_4278,N_4749);
nor U4957 (N_4957,N_4474,N_4250);
and U4958 (N_4958,N_4532,N_4484);
xor U4959 (N_4959,N_4538,N_4352);
nor U4960 (N_4960,N_4581,N_4323);
xor U4961 (N_4961,N_4692,N_4353);
and U4962 (N_4962,N_4630,N_4626);
xor U4963 (N_4963,N_4509,N_4724);
nand U4964 (N_4964,N_4437,N_4549);
nand U4965 (N_4965,N_4675,N_4324);
nor U4966 (N_4966,N_4345,N_4326);
xnor U4967 (N_4967,N_4481,N_4402);
or U4968 (N_4968,N_4480,N_4470);
or U4969 (N_4969,N_4713,N_4792);
nor U4970 (N_4970,N_4478,N_4736);
nand U4971 (N_4971,N_4786,N_4238);
or U4972 (N_4972,N_4753,N_4271);
nor U4973 (N_4973,N_4464,N_4614);
and U4974 (N_4974,N_4567,N_4715);
or U4975 (N_4975,N_4734,N_4779);
nor U4976 (N_4976,N_4296,N_4449);
nor U4977 (N_4977,N_4328,N_4631);
xor U4978 (N_4978,N_4602,N_4406);
and U4979 (N_4979,N_4766,N_4510);
nand U4980 (N_4980,N_4641,N_4344);
nand U4981 (N_4981,N_4768,N_4556);
and U4982 (N_4982,N_4629,N_4393);
xor U4983 (N_4983,N_4225,N_4304);
or U4984 (N_4984,N_4321,N_4314);
nand U4985 (N_4985,N_4458,N_4415);
or U4986 (N_4986,N_4433,N_4722);
nor U4987 (N_4987,N_4498,N_4741);
and U4988 (N_4988,N_4645,N_4276);
and U4989 (N_4989,N_4597,N_4526);
and U4990 (N_4990,N_4502,N_4306);
nor U4991 (N_4991,N_4623,N_4448);
and U4992 (N_4992,N_4769,N_4663);
or U4993 (N_4993,N_4423,N_4687);
nor U4994 (N_4994,N_4655,N_4543);
xor U4995 (N_4995,N_4636,N_4587);
xor U4996 (N_4996,N_4790,N_4242);
xnor U4997 (N_4997,N_4392,N_4673);
nand U4998 (N_4998,N_4794,N_4568);
nand U4999 (N_4999,N_4533,N_4752);
xor U5000 (N_5000,N_4226,N_4763);
nor U5001 (N_5001,N_4540,N_4368);
or U5002 (N_5002,N_4301,N_4471);
and U5003 (N_5003,N_4245,N_4574);
and U5004 (N_5004,N_4791,N_4640);
nand U5005 (N_5005,N_4576,N_4601);
nand U5006 (N_5006,N_4773,N_4591);
nand U5007 (N_5007,N_4579,N_4221);
nand U5008 (N_5008,N_4571,N_4566);
nand U5009 (N_5009,N_4633,N_4637);
nor U5010 (N_5010,N_4490,N_4302);
nor U5011 (N_5011,N_4772,N_4707);
and U5012 (N_5012,N_4525,N_4403);
xor U5013 (N_5013,N_4487,N_4513);
nor U5014 (N_5014,N_4531,N_4535);
and U5015 (N_5015,N_4354,N_4701);
nor U5016 (N_5016,N_4251,N_4269);
nor U5017 (N_5017,N_4750,N_4287);
nor U5018 (N_5018,N_4775,N_4493);
xor U5019 (N_5019,N_4500,N_4689);
nand U5020 (N_5020,N_4668,N_4263);
xor U5021 (N_5021,N_4237,N_4732);
or U5022 (N_5022,N_4585,N_4536);
nand U5023 (N_5023,N_4408,N_4382);
and U5024 (N_5024,N_4683,N_4270);
or U5025 (N_5025,N_4577,N_4739);
xnor U5026 (N_5026,N_4506,N_4586);
nand U5027 (N_5027,N_4507,N_4664);
nand U5028 (N_5028,N_4231,N_4273);
nor U5029 (N_5029,N_4761,N_4573);
and U5030 (N_5030,N_4698,N_4222);
xor U5031 (N_5031,N_4327,N_4207);
xnor U5032 (N_5032,N_4599,N_4212);
or U5033 (N_5033,N_4616,N_4783);
and U5034 (N_5034,N_4445,N_4416);
nor U5035 (N_5035,N_4200,N_4370);
nand U5036 (N_5036,N_4460,N_4332);
nor U5037 (N_5037,N_4520,N_4468);
and U5038 (N_5038,N_4632,N_4608);
and U5039 (N_5039,N_4572,N_4554);
nand U5040 (N_5040,N_4665,N_4356);
or U5041 (N_5041,N_4583,N_4355);
xnor U5042 (N_5042,N_4767,N_4731);
or U5043 (N_5043,N_4497,N_4446);
xor U5044 (N_5044,N_4620,N_4793);
nand U5045 (N_5045,N_4282,N_4300);
or U5046 (N_5046,N_4391,N_4247);
xor U5047 (N_5047,N_4604,N_4439);
and U5048 (N_5048,N_4401,N_4503);
nand U5049 (N_5049,N_4230,N_4316);
nor U5050 (N_5050,N_4425,N_4652);
and U5051 (N_5051,N_4255,N_4605);
and U5052 (N_5052,N_4381,N_4201);
and U5053 (N_5053,N_4310,N_4686);
or U5054 (N_5054,N_4303,N_4642);
nand U5055 (N_5055,N_4267,N_4404);
nor U5056 (N_5056,N_4770,N_4551);
nor U5057 (N_5057,N_4213,N_4615);
and U5058 (N_5058,N_4788,N_4690);
or U5059 (N_5059,N_4565,N_4654);
nor U5060 (N_5060,N_4694,N_4606);
or U5061 (N_5061,N_4746,N_4505);
nand U5062 (N_5062,N_4742,N_4522);
nand U5063 (N_5063,N_4542,N_4203);
nor U5064 (N_5064,N_4413,N_4678);
xor U5065 (N_5065,N_4252,N_4442);
or U5066 (N_5066,N_4216,N_4285);
xnor U5067 (N_5067,N_4653,N_4441);
nand U5068 (N_5068,N_4759,N_4224);
and U5069 (N_5069,N_4512,N_4725);
xnor U5070 (N_5070,N_4735,N_4706);
or U5071 (N_5071,N_4253,N_4625);
or U5072 (N_5072,N_4409,N_4617);
nor U5073 (N_5073,N_4434,N_4681);
xor U5074 (N_5074,N_4661,N_4754);
nor U5075 (N_5075,N_4575,N_4491);
or U5076 (N_5076,N_4320,N_4712);
and U5077 (N_5077,N_4244,N_4205);
nor U5078 (N_5078,N_4669,N_4564);
and U5079 (N_5079,N_4284,N_4364);
nand U5080 (N_5080,N_4518,N_4234);
or U5081 (N_5081,N_4443,N_4666);
nor U5082 (N_5082,N_4339,N_4337);
or U5083 (N_5083,N_4288,N_4529);
and U5084 (N_5084,N_4236,N_4405);
xnor U5085 (N_5085,N_4335,N_4515);
xor U5086 (N_5086,N_4570,N_4239);
and U5087 (N_5087,N_4598,N_4232);
or U5088 (N_5088,N_4440,N_4394);
nand U5089 (N_5089,N_4550,N_4256);
or U5090 (N_5090,N_4293,N_4562);
and U5091 (N_5091,N_4787,N_4229);
nand U5092 (N_5092,N_4396,N_4461);
nand U5093 (N_5093,N_4325,N_4359);
nand U5094 (N_5094,N_4638,N_4639);
nand U5095 (N_5095,N_4358,N_4684);
or U5096 (N_5096,N_4307,N_4469);
or U5097 (N_5097,N_4215,N_4674);
nand U5098 (N_5098,N_4362,N_4705);
or U5099 (N_5099,N_4465,N_4634);
xor U5100 (N_5100,N_4306,N_4472);
xnor U5101 (N_5101,N_4404,N_4695);
nor U5102 (N_5102,N_4334,N_4769);
or U5103 (N_5103,N_4620,N_4647);
nor U5104 (N_5104,N_4529,N_4741);
and U5105 (N_5105,N_4524,N_4529);
xnor U5106 (N_5106,N_4616,N_4437);
nor U5107 (N_5107,N_4751,N_4322);
nand U5108 (N_5108,N_4727,N_4498);
nand U5109 (N_5109,N_4341,N_4731);
nand U5110 (N_5110,N_4684,N_4554);
nand U5111 (N_5111,N_4410,N_4781);
nor U5112 (N_5112,N_4538,N_4422);
nand U5113 (N_5113,N_4671,N_4763);
nand U5114 (N_5114,N_4230,N_4381);
nand U5115 (N_5115,N_4741,N_4467);
and U5116 (N_5116,N_4420,N_4641);
nor U5117 (N_5117,N_4510,N_4463);
xnor U5118 (N_5118,N_4684,N_4406);
or U5119 (N_5119,N_4355,N_4423);
nor U5120 (N_5120,N_4277,N_4464);
nand U5121 (N_5121,N_4262,N_4524);
xnor U5122 (N_5122,N_4642,N_4492);
xnor U5123 (N_5123,N_4243,N_4350);
and U5124 (N_5124,N_4473,N_4430);
nor U5125 (N_5125,N_4599,N_4355);
and U5126 (N_5126,N_4216,N_4502);
and U5127 (N_5127,N_4626,N_4690);
xor U5128 (N_5128,N_4533,N_4370);
nor U5129 (N_5129,N_4388,N_4233);
nand U5130 (N_5130,N_4298,N_4799);
xnor U5131 (N_5131,N_4319,N_4690);
nor U5132 (N_5132,N_4683,N_4722);
xnor U5133 (N_5133,N_4239,N_4261);
nand U5134 (N_5134,N_4326,N_4558);
xnor U5135 (N_5135,N_4712,N_4799);
or U5136 (N_5136,N_4751,N_4259);
nand U5137 (N_5137,N_4473,N_4484);
nor U5138 (N_5138,N_4478,N_4689);
and U5139 (N_5139,N_4203,N_4550);
nor U5140 (N_5140,N_4359,N_4604);
nor U5141 (N_5141,N_4617,N_4230);
and U5142 (N_5142,N_4461,N_4272);
xor U5143 (N_5143,N_4624,N_4635);
xnor U5144 (N_5144,N_4477,N_4483);
nand U5145 (N_5145,N_4648,N_4352);
and U5146 (N_5146,N_4679,N_4706);
and U5147 (N_5147,N_4258,N_4313);
nand U5148 (N_5148,N_4494,N_4488);
nand U5149 (N_5149,N_4589,N_4283);
and U5150 (N_5150,N_4582,N_4320);
or U5151 (N_5151,N_4513,N_4574);
nor U5152 (N_5152,N_4721,N_4362);
nor U5153 (N_5153,N_4519,N_4494);
or U5154 (N_5154,N_4726,N_4708);
and U5155 (N_5155,N_4355,N_4731);
nor U5156 (N_5156,N_4703,N_4327);
or U5157 (N_5157,N_4479,N_4296);
nor U5158 (N_5158,N_4392,N_4422);
nor U5159 (N_5159,N_4521,N_4214);
or U5160 (N_5160,N_4339,N_4222);
xnor U5161 (N_5161,N_4398,N_4301);
xnor U5162 (N_5162,N_4236,N_4205);
nand U5163 (N_5163,N_4710,N_4569);
nor U5164 (N_5164,N_4274,N_4762);
nor U5165 (N_5165,N_4447,N_4455);
or U5166 (N_5166,N_4320,N_4554);
nor U5167 (N_5167,N_4410,N_4690);
nand U5168 (N_5168,N_4576,N_4677);
nand U5169 (N_5169,N_4263,N_4701);
nor U5170 (N_5170,N_4304,N_4291);
xor U5171 (N_5171,N_4329,N_4239);
xor U5172 (N_5172,N_4525,N_4663);
nor U5173 (N_5173,N_4231,N_4788);
and U5174 (N_5174,N_4504,N_4595);
nor U5175 (N_5175,N_4489,N_4243);
and U5176 (N_5176,N_4659,N_4454);
or U5177 (N_5177,N_4466,N_4759);
nand U5178 (N_5178,N_4691,N_4462);
and U5179 (N_5179,N_4760,N_4592);
and U5180 (N_5180,N_4592,N_4614);
xnor U5181 (N_5181,N_4507,N_4583);
nand U5182 (N_5182,N_4727,N_4422);
xor U5183 (N_5183,N_4781,N_4338);
and U5184 (N_5184,N_4635,N_4707);
and U5185 (N_5185,N_4317,N_4273);
nand U5186 (N_5186,N_4203,N_4236);
or U5187 (N_5187,N_4538,N_4349);
and U5188 (N_5188,N_4606,N_4211);
nand U5189 (N_5189,N_4211,N_4355);
xnor U5190 (N_5190,N_4345,N_4481);
nor U5191 (N_5191,N_4205,N_4576);
xnor U5192 (N_5192,N_4662,N_4353);
nand U5193 (N_5193,N_4311,N_4487);
nor U5194 (N_5194,N_4271,N_4583);
nand U5195 (N_5195,N_4681,N_4377);
xor U5196 (N_5196,N_4641,N_4676);
or U5197 (N_5197,N_4314,N_4270);
nor U5198 (N_5198,N_4231,N_4699);
and U5199 (N_5199,N_4364,N_4505);
nor U5200 (N_5200,N_4370,N_4534);
and U5201 (N_5201,N_4679,N_4667);
xor U5202 (N_5202,N_4631,N_4661);
nor U5203 (N_5203,N_4723,N_4703);
nor U5204 (N_5204,N_4498,N_4385);
or U5205 (N_5205,N_4225,N_4238);
nor U5206 (N_5206,N_4763,N_4355);
nand U5207 (N_5207,N_4488,N_4430);
nand U5208 (N_5208,N_4728,N_4622);
xnor U5209 (N_5209,N_4522,N_4345);
nor U5210 (N_5210,N_4741,N_4625);
and U5211 (N_5211,N_4591,N_4742);
nor U5212 (N_5212,N_4519,N_4347);
xnor U5213 (N_5213,N_4461,N_4260);
xor U5214 (N_5214,N_4426,N_4600);
and U5215 (N_5215,N_4481,N_4252);
xor U5216 (N_5216,N_4268,N_4326);
nand U5217 (N_5217,N_4630,N_4572);
nor U5218 (N_5218,N_4243,N_4483);
nand U5219 (N_5219,N_4242,N_4424);
and U5220 (N_5220,N_4368,N_4571);
xnor U5221 (N_5221,N_4501,N_4752);
and U5222 (N_5222,N_4553,N_4388);
nand U5223 (N_5223,N_4321,N_4787);
xor U5224 (N_5224,N_4362,N_4219);
and U5225 (N_5225,N_4742,N_4581);
nor U5226 (N_5226,N_4687,N_4258);
xnor U5227 (N_5227,N_4775,N_4436);
xor U5228 (N_5228,N_4643,N_4272);
or U5229 (N_5229,N_4274,N_4287);
nor U5230 (N_5230,N_4658,N_4299);
xor U5231 (N_5231,N_4787,N_4389);
and U5232 (N_5232,N_4468,N_4542);
or U5233 (N_5233,N_4249,N_4509);
nor U5234 (N_5234,N_4277,N_4700);
or U5235 (N_5235,N_4598,N_4441);
xnor U5236 (N_5236,N_4703,N_4793);
nand U5237 (N_5237,N_4713,N_4320);
or U5238 (N_5238,N_4552,N_4223);
and U5239 (N_5239,N_4272,N_4331);
or U5240 (N_5240,N_4699,N_4267);
and U5241 (N_5241,N_4225,N_4221);
or U5242 (N_5242,N_4264,N_4397);
nor U5243 (N_5243,N_4478,N_4539);
xor U5244 (N_5244,N_4694,N_4529);
nor U5245 (N_5245,N_4577,N_4319);
nor U5246 (N_5246,N_4427,N_4354);
and U5247 (N_5247,N_4525,N_4352);
nand U5248 (N_5248,N_4675,N_4711);
or U5249 (N_5249,N_4523,N_4310);
nor U5250 (N_5250,N_4567,N_4764);
or U5251 (N_5251,N_4233,N_4356);
and U5252 (N_5252,N_4315,N_4667);
or U5253 (N_5253,N_4731,N_4556);
nor U5254 (N_5254,N_4478,N_4290);
and U5255 (N_5255,N_4347,N_4491);
or U5256 (N_5256,N_4444,N_4389);
or U5257 (N_5257,N_4473,N_4477);
or U5258 (N_5258,N_4785,N_4641);
or U5259 (N_5259,N_4393,N_4607);
or U5260 (N_5260,N_4781,N_4473);
nor U5261 (N_5261,N_4225,N_4678);
nor U5262 (N_5262,N_4292,N_4405);
nor U5263 (N_5263,N_4797,N_4416);
nor U5264 (N_5264,N_4553,N_4728);
xor U5265 (N_5265,N_4446,N_4382);
nor U5266 (N_5266,N_4776,N_4346);
or U5267 (N_5267,N_4388,N_4748);
nand U5268 (N_5268,N_4250,N_4791);
nand U5269 (N_5269,N_4418,N_4506);
and U5270 (N_5270,N_4505,N_4652);
or U5271 (N_5271,N_4590,N_4304);
nor U5272 (N_5272,N_4482,N_4477);
xnor U5273 (N_5273,N_4275,N_4248);
or U5274 (N_5274,N_4775,N_4718);
nor U5275 (N_5275,N_4353,N_4425);
nand U5276 (N_5276,N_4321,N_4553);
nand U5277 (N_5277,N_4633,N_4768);
and U5278 (N_5278,N_4510,N_4272);
xor U5279 (N_5279,N_4750,N_4270);
xnor U5280 (N_5280,N_4261,N_4576);
or U5281 (N_5281,N_4650,N_4388);
nor U5282 (N_5282,N_4593,N_4521);
or U5283 (N_5283,N_4440,N_4595);
nor U5284 (N_5284,N_4710,N_4506);
nor U5285 (N_5285,N_4560,N_4649);
and U5286 (N_5286,N_4541,N_4325);
or U5287 (N_5287,N_4321,N_4205);
xor U5288 (N_5288,N_4761,N_4366);
xnor U5289 (N_5289,N_4495,N_4762);
xnor U5290 (N_5290,N_4361,N_4342);
nand U5291 (N_5291,N_4674,N_4579);
nor U5292 (N_5292,N_4304,N_4585);
or U5293 (N_5293,N_4272,N_4744);
and U5294 (N_5294,N_4491,N_4669);
xnor U5295 (N_5295,N_4344,N_4285);
or U5296 (N_5296,N_4458,N_4406);
nand U5297 (N_5297,N_4452,N_4657);
and U5298 (N_5298,N_4650,N_4707);
and U5299 (N_5299,N_4798,N_4617);
and U5300 (N_5300,N_4462,N_4636);
nand U5301 (N_5301,N_4677,N_4525);
xor U5302 (N_5302,N_4578,N_4238);
nor U5303 (N_5303,N_4540,N_4349);
or U5304 (N_5304,N_4573,N_4232);
or U5305 (N_5305,N_4320,N_4498);
or U5306 (N_5306,N_4707,N_4274);
or U5307 (N_5307,N_4767,N_4472);
xor U5308 (N_5308,N_4232,N_4278);
nor U5309 (N_5309,N_4217,N_4565);
or U5310 (N_5310,N_4609,N_4663);
nand U5311 (N_5311,N_4664,N_4625);
nand U5312 (N_5312,N_4645,N_4648);
nand U5313 (N_5313,N_4250,N_4695);
xnor U5314 (N_5314,N_4545,N_4439);
xnor U5315 (N_5315,N_4781,N_4517);
or U5316 (N_5316,N_4557,N_4629);
and U5317 (N_5317,N_4755,N_4743);
nand U5318 (N_5318,N_4512,N_4524);
nand U5319 (N_5319,N_4571,N_4590);
nand U5320 (N_5320,N_4787,N_4278);
xor U5321 (N_5321,N_4420,N_4754);
or U5322 (N_5322,N_4460,N_4490);
or U5323 (N_5323,N_4256,N_4453);
nor U5324 (N_5324,N_4559,N_4604);
or U5325 (N_5325,N_4615,N_4624);
nor U5326 (N_5326,N_4635,N_4626);
and U5327 (N_5327,N_4285,N_4306);
or U5328 (N_5328,N_4397,N_4334);
nor U5329 (N_5329,N_4609,N_4394);
nand U5330 (N_5330,N_4726,N_4698);
xor U5331 (N_5331,N_4752,N_4651);
nand U5332 (N_5332,N_4380,N_4256);
xor U5333 (N_5333,N_4644,N_4538);
nor U5334 (N_5334,N_4410,N_4766);
nor U5335 (N_5335,N_4422,N_4377);
xnor U5336 (N_5336,N_4580,N_4496);
or U5337 (N_5337,N_4388,N_4581);
nor U5338 (N_5338,N_4449,N_4345);
nor U5339 (N_5339,N_4697,N_4527);
nand U5340 (N_5340,N_4565,N_4215);
nand U5341 (N_5341,N_4247,N_4415);
or U5342 (N_5342,N_4639,N_4404);
xnor U5343 (N_5343,N_4696,N_4589);
nand U5344 (N_5344,N_4382,N_4691);
or U5345 (N_5345,N_4490,N_4553);
nand U5346 (N_5346,N_4362,N_4630);
and U5347 (N_5347,N_4645,N_4664);
nand U5348 (N_5348,N_4555,N_4251);
nand U5349 (N_5349,N_4523,N_4296);
nand U5350 (N_5350,N_4708,N_4225);
nand U5351 (N_5351,N_4414,N_4307);
and U5352 (N_5352,N_4284,N_4395);
xor U5353 (N_5353,N_4221,N_4511);
xnor U5354 (N_5354,N_4356,N_4653);
and U5355 (N_5355,N_4389,N_4742);
nor U5356 (N_5356,N_4222,N_4437);
and U5357 (N_5357,N_4759,N_4646);
nand U5358 (N_5358,N_4357,N_4484);
and U5359 (N_5359,N_4313,N_4375);
or U5360 (N_5360,N_4209,N_4663);
or U5361 (N_5361,N_4397,N_4567);
or U5362 (N_5362,N_4737,N_4710);
nand U5363 (N_5363,N_4642,N_4691);
xor U5364 (N_5364,N_4387,N_4285);
nand U5365 (N_5365,N_4404,N_4258);
or U5366 (N_5366,N_4463,N_4453);
xnor U5367 (N_5367,N_4358,N_4343);
nor U5368 (N_5368,N_4586,N_4355);
and U5369 (N_5369,N_4307,N_4367);
or U5370 (N_5370,N_4418,N_4518);
nor U5371 (N_5371,N_4651,N_4222);
or U5372 (N_5372,N_4489,N_4619);
and U5373 (N_5373,N_4786,N_4330);
nand U5374 (N_5374,N_4486,N_4496);
or U5375 (N_5375,N_4602,N_4255);
xor U5376 (N_5376,N_4687,N_4535);
nor U5377 (N_5377,N_4354,N_4471);
nor U5378 (N_5378,N_4266,N_4249);
and U5379 (N_5379,N_4752,N_4245);
nor U5380 (N_5380,N_4234,N_4501);
xor U5381 (N_5381,N_4740,N_4535);
or U5382 (N_5382,N_4626,N_4698);
and U5383 (N_5383,N_4462,N_4684);
nor U5384 (N_5384,N_4210,N_4627);
nor U5385 (N_5385,N_4534,N_4541);
xnor U5386 (N_5386,N_4572,N_4670);
and U5387 (N_5387,N_4790,N_4372);
nand U5388 (N_5388,N_4383,N_4230);
nand U5389 (N_5389,N_4449,N_4640);
xnor U5390 (N_5390,N_4269,N_4721);
nor U5391 (N_5391,N_4392,N_4295);
xnor U5392 (N_5392,N_4654,N_4603);
or U5393 (N_5393,N_4504,N_4231);
nor U5394 (N_5394,N_4409,N_4233);
and U5395 (N_5395,N_4606,N_4479);
or U5396 (N_5396,N_4254,N_4215);
and U5397 (N_5397,N_4675,N_4732);
nor U5398 (N_5398,N_4249,N_4649);
nand U5399 (N_5399,N_4678,N_4433);
and U5400 (N_5400,N_4943,N_5020);
nor U5401 (N_5401,N_4969,N_5165);
and U5402 (N_5402,N_5102,N_5243);
xor U5403 (N_5403,N_5094,N_5323);
and U5404 (N_5404,N_5191,N_5066);
nand U5405 (N_5405,N_4820,N_5135);
nor U5406 (N_5406,N_5229,N_5247);
or U5407 (N_5407,N_5113,N_5019);
and U5408 (N_5408,N_5070,N_4812);
nor U5409 (N_5409,N_5133,N_5158);
or U5410 (N_5410,N_5272,N_4877);
nor U5411 (N_5411,N_4934,N_4961);
xnor U5412 (N_5412,N_4878,N_5348);
nand U5413 (N_5413,N_5207,N_5117);
and U5414 (N_5414,N_4988,N_4838);
nand U5415 (N_5415,N_5370,N_5076);
xnor U5416 (N_5416,N_5271,N_4976);
and U5417 (N_5417,N_4913,N_4981);
nor U5418 (N_5418,N_5159,N_4870);
nor U5419 (N_5419,N_5236,N_5156);
nor U5420 (N_5420,N_5086,N_5355);
nand U5421 (N_5421,N_4983,N_5262);
and U5422 (N_5422,N_5026,N_5064);
or U5423 (N_5423,N_5208,N_5289);
nor U5424 (N_5424,N_5009,N_4995);
and U5425 (N_5425,N_5365,N_4998);
nor U5426 (N_5426,N_5268,N_5103);
nor U5427 (N_5427,N_4848,N_5153);
or U5428 (N_5428,N_5085,N_4993);
or U5429 (N_5429,N_5163,N_5392);
and U5430 (N_5430,N_4909,N_4922);
nand U5431 (N_5431,N_4999,N_5197);
and U5432 (N_5432,N_5171,N_4886);
or U5433 (N_5433,N_4810,N_4857);
and U5434 (N_5434,N_5280,N_5358);
and U5435 (N_5435,N_4828,N_5288);
and U5436 (N_5436,N_5131,N_5362);
xor U5437 (N_5437,N_4990,N_4971);
or U5438 (N_5438,N_5095,N_5237);
and U5439 (N_5439,N_5169,N_4985);
nand U5440 (N_5440,N_5351,N_4809);
nand U5441 (N_5441,N_5330,N_5250);
xnor U5442 (N_5442,N_5282,N_4826);
nor U5443 (N_5443,N_5279,N_4802);
nand U5444 (N_5444,N_5258,N_5202);
xor U5445 (N_5445,N_4947,N_4949);
or U5446 (N_5446,N_4819,N_4829);
or U5447 (N_5447,N_5188,N_5206);
and U5448 (N_5448,N_5015,N_4973);
or U5449 (N_5449,N_5087,N_4882);
nor U5450 (N_5450,N_4803,N_5230);
xnor U5451 (N_5451,N_5168,N_4950);
or U5452 (N_5452,N_5312,N_5029);
or U5453 (N_5453,N_4929,N_4960);
nand U5454 (N_5454,N_4843,N_5018);
or U5455 (N_5455,N_5075,N_5034);
xor U5456 (N_5456,N_4846,N_4946);
and U5457 (N_5457,N_5195,N_5211);
and U5458 (N_5458,N_5214,N_5345);
xor U5459 (N_5459,N_5264,N_5215);
nand U5460 (N_5460,N_4824,N_5266);
or U5461 (N_5461,N_5028,N_4884);
nand U5462 (N_5462,N_5115,N_5164);
or U5463 (N_5463,N_5007,N_5396);
and U5464 (N_5464,N_5394,N_5297);
xnor U5465 (N_5465,N_5298,N_5201);
xor U5466 (N_5466,N_5128,N_5101);
or U5467 (N_5467,N_4849,N_5361);
xnor U5468 (N_5468,N_4858,N_4924);
nor U5469 (N_5469,N_5056,N_5327);
xnor U5470 (N_5470,N_5142,N_5315);
nor U5471 (N_5471,N_5167,N_5027);
xor U5472 (N_5472,N_5270,N_5353);
xnor U5473 (N_5473,N_5048,N_4875);
nor U5474 (N_5474,N_5154,N_5046);
nor U5475 (N_5475,N_5053,N_4967);
nand U5476 (N_5476,N_4997,N_5317);
nand U5477 (N_5477,N_5308,N_5275);
nand U5478 (N_5478,N_4952,N_4907);
or U5479 (N_5479,N_5319,N_4866);
xnor U5480 (N_5480,N_5013,N_5324);
nor U5481 (N_5481,N_4908,N_5124);
xnor U5482 (N_5482,N_5293,N_4982);
nand U5483 (N_5483,N_5263,N_5233);
xor U5484 (N_5484,N_4987,N_4958);
nor U5485 (N_5485,N_5335,N_5055);
or U5486 (N_5486,N_5210,N_4816);
nand U5487 (N_5487,N_5336,N_4927);
xnor U5488 (N_5488,N_4817,N_4914);
and U5489 (N_5489,N_4885,N_5387);
nor U5490 (N_5490,N_4915,N_5139);
xnor U5491 (N_5491,N_5108,N_5106);
nor U5492 (N_5492,N_5393,N_5363);
or U5493 (N_5493,N_5222,N_4916);
or U5494 (N_5494,N_5097,N_5148);
nor U5495 (N_5495,N_5234,N_5257);
and U5496 (N_5496,N_5132,N_5123);
and U5497 (N_5497,N_5025,N_5054);
and U5498 (N_5498,N_5292,N_5161);
or U5499 (N_5499,N_5294,N_5285);
xnor U5500 (N_5500,N_5241,N_4815);
nand U5501 (N_5501,N_5388,N_5300);
xor U5502 (N_5502,N_4837,N_4984);
xnor U5503 (N_5503,N_4833,N_5039);
or U5504 (N_5504,N_5184,N_4940);
xor U5505 (N_5505,N_5179,N_5339);
xor U5506 (N_5506,N_5231,N_5286);
nor U5507 (N_5507,N_4844,N_5193);
nor U5508 (N_5508,N_5384,N_5160);
and U5509 (N_5509,N_4814,N_4900);
xor U5510 (N_5510,N_4904,N_4956);
nand U5511 (N_5511,N_5024,N_4896);
nor U5512 (N_5512,N_5038,N_4932);
nand U5513 (N_5513,N_5044,N_5313);
nor U5514 (N_5514,N_5252,N_5383);
nor U5515 (N_5515,N_5084,N_4921);
nand U5516 (N_5516,N_5220,N_5374);
nor U5517 (N_5517,N_4941,N_5185);
xor U5518 (N_5518,N_5340,N_4991);
nor U5519 (N_5519,N_5090,N_5379);
nor U5520 (N_5520,N_5138,N_5309);
or U5521 (N_5521,N_4972,N_5256);
nor U5522 (N_5522,N_4948,N_5082);
nand U5523 (N_5523,N_4830,N_4937);
xnor U5524 (N_5524,N_4902,N_5372);
nor U5525 (N_5525,N_5069,N_5259);
xor U5526 (N_5526,N_5314,N_5344);
and U5527 (N_5527,N_5248,N_5307);
nand U5528 (N_5528,N_5040,N_5190);
nor U5529 (N_5529,N_5092,N_5178);
and U5530 (N_5530,N_5091,N_5368);
xnor U5531 (N_5531,N_4897,N_5145);
and U5532 (N_5532,N_5074,N_5342);
nand U5533 (N_5533,N_4847,N_5254);
xnor U5534 (N_5534,N_5032,N_4959);
or U5535 (N_5535,N_5325,N_4890);
nor U5536 (N_5536,N_5350,N_4962);
or U5537 (N_5537,N_4861,N_5352);
nor U5538 (N_5538,N_5045,N_4855);
xor U5539 (N_5539,N_5337,N_4899);
nor U5540 (N_5540,N_5141,N_4888);
xnor U5541 (N_5541,N_5174,N_4994);
or U5542 (N_5542,N_4813,N_5077);
or U5543 (N_5543,N_5320,N_5209);
and U5544 (N_5544,N_5291,N_5283);
nand U5545 (N_5545,N_5112,N_4841);
or U5546 (N_5546,N_4895,N_5036);
xnor U5547 (N_5547,N_5225,N_5110);
xor U5548 (N_5548,N_5037,N_4954);
xnor U5549 (N_5549,N_5006,N_5129);
xnor U5550 (N_5550,N_4965,N_5381);
or U5551 (N_5551,N_4874,N_4917);
nand U5552 (N_5552,N_5043,N_5200);
xor U5553 (N_5553,N_5116,N_5114);
nand U5554 (N_5554,N_4871,N_5093);
nand U5555 (N_5555,N_4951,N_5203);
nor U5556 (N_5556,N_4980,N_5100);
or U5557 (N_5557,N_5192,N_5398);
or U5558 (N_5558,N_5296,N_4898);
nand U5559 (N_5559,N_5239,N_4901);
xor U5560 (N_5560,N_5051,N_5221);
and U5561 (N_5561,N_5079,N_5334);
and U5562 (N_5562,N_4834,N_5251);
or U5563 (N_5563,N_5310,N_5399);
xor U5564 (N_5564,N_5119,N_5157);
nor U5565 (N_5565,N_4905,N_4879);
or U5566 (N_5566,N_5332,N_5014);
or U5567 (N_5567,N_4856,N_5120);
or U5568 (N_5568,N_5261,N_5130);
nor U5569 (N_5569,N_4806,N_5253);
nor U5570 (N_5570,N_5042,N_4808);
and U5571 (N_5571,N_5033,N_5062);
xor U5572 (N_5572,N_5099,N_5078);
and U5573 (N_5573,N_4883,N_4825);
and U5574 (N_5574,N_4989,N_5081);
or U5575 (N_5575,N_4821,N_4872);
xor U5576 (N_5576,N_4807,N_5364);
nand U5577 (N_5577,N_5021,N_4842);
nor U5578 (N_5578,N_5073,N_5311);
nor U5579 (N_5579,N_5284,N_5194);
nor U5580 (N_5580,N_5306,N_5089);
nand U5581 (N_5581,N_4887,N_4918);
or U5582 (N_5582,N_4862,N_5228);
or U5583 (N_5583,N_5390,N_5008);
and U5584 (N_5584,N_5061,N_5299);
and U5585 (N_5585,N_5218,N_5290);
nor U5586 (N_5586,N_5058,N_5003);
nor U5587 (N_5587,N_4869,N_4936);
xor U5588 (N_5588,N_4839,N_5265);
and U5589 (N_5589,N_5052,N_5155);
nand U5590 (N_5590,N_5170,N_5386);
nor U5591 (N_5591,N_4968,N_5223);
nor U5592 (N_5592,N_5240,N_5065);
xor U5593 (N_5593,N_4811,N_4818);
nand U5594 (N_5594,N_5278,N_4867);
nand U5595 (N_5595,N_4860,N_4894);
and U5596 (N_5596,N_4964,N_4978);
or U5597 (N_5597,N_5035,N_5359);
xnor U5598 (N_5598,N_5397,N_5111);
nand U5599 (N_5599,N_4930,N_5151);
xnor U5600 (N_5600,N_4822,N_5172);
xor U5601 (N_5601,N_5244,N_5049);
nor U5602 (N_5602,N_5134,N_4923);
nand U5603 (N_5603,N_4925,N_4979);
xor U5604 (N_5604,N_5002,N_5047);
nand U5605 (N_5605,N_4942,N_5249);
nand U5606 (N_5606,N_5373,N_4801);
xor U5607 (N_5607,N_5071,N_4963);
nand U5608 (N_5608,N_5173,N_4854);
or U5609 (N_5609,N_5176,N_5149);
nand U5610 (N_5610,N_5126,N_4892);
and U5611 (N_5611,N_4992,N_5096);
nand U5612 (N_5612,N_5180,N_4938);
nor U5613 (N_5613,N_5152,N_5219);
or U5614 (N_5614,N_5205,N_4881);
and U5615 (N_5615,N_5137,N_5000);
xnor U5616 (N_5616,N_5162,N_5238);
or U5617 (N_5617,N_4906,N_5212);
nand U5618 (N_5618,N_5166,N_5226);
nor U5619 (N_5619,N_5333,N_5269);
nand U5620 (N_5620,N_4827,N_5107);
or U5621 (N_5621,N_5187,N_4845);
nor U5622 (N_5622,N_5274,N_4831);
nor U5623 (N_5623,N_5063,N_5301);
and U5624 (N_5624,N_5010,N_5357);
nand U5625 (N_5625,N_5098,N_5281);
nand U5626 (N_5626,N_5198,N_4931);
nor U5627 (N_5627,N_4853,N_5341);
or U5628 (N_5628,N_5177,N_4903);
or U5629 (N_5629,N_5175,N_4859);
xnor U5630 (N_5630,N_5088,N_4864);
nor U5631 (N_5631,N_5204,N_5304);
xor U5632 (N_5632,N_5347,N_4868);
nor U5633 (N_5633,N_4823,N_5150);
xor U5634 (N_5634,N_5331,N_5277);
nand U5635 (N_5635,N_5326,N_5377);
and U5636 (N_5636,N_5356,N_5017);
nand U5637 (N_5637,N_5245,N_5023);
nor U5638 (N_5638,N_5216,N_5395);
and U5639 (N_5639,N_5354,N_5182);
nor U5640 (N_5640,N_5224,N_5242);
nand U5641 (N_5641,N_4805,N_5227);
nand U5642 (N_5642,N_4986,N_5183);
xor U5643 (N_5643,N_5217,N_5376);
nor U5644 (N_5644,N_5318,N_5321);
nor U5645 (N_5645,N_5011,N_4945);
and U5646 (N_5646,N_5196,N_5105);
nand U5647 (N_5647,N_5371,N_5060);
or U5648 (N_5648,N_4977,N_5016);
or U5649 (N_5649,N_5147,N_5287);
nand U5650 (N_5650,N_4926,N_4975);
nand U5651 (N_5651,N_5273,N_4800);
xor U5652 (N_5652,N_5022,N_5109);
nor U5653 (N_5653,N_4928,N_5144);
and U5654 (N_5654,N_5246,N_5067);
and U5655 (N_5655,N_5127,N_5316);
nor U5656 (N_5656,N_5255,N_4891);
nor U5657 (N_5657,N_4889,N_5004);
nor U5658 (N_5658,N_5213,N_5146);
and U5659 (N_5659,N_5385,N_5125);
nand U5660 (N_5660,N_5305,N_5303);
nand U5661 (N_5661,N_5080,N_4966);
xnor U5662 (N_5662,N_4832,N_4851);
xor U5663 (N_5663,N_5181,N_5235);
or U5664 (N_5664,N_5232,N_5367);
or U5665 (N_5665,N_4912,N_5041);
nor U5666 (N_5666,N_4876,N_4974);
and U5667 (N_5667,N_5012,N_5360);
nand U5668 (N_5668,N_5031,N_4953);
nor U5669 (N_5669,N_5338,N_4944);
and U5670 (N_5670,N_4880,N_4919);
and U5671 (N_5671,N_5302,N_4835);
and U5672 (N_5672,N_4911,N_4836);
or U5673 (N_5673,N_4920,N_5378);
nand U5674 (N_5674,N_4804,N_4955);
nand U5675 (N_5675,N_5375,N_4840);
nand U5676 (N_5676,N_5140,N_5050);
nand U5677 (N_5677,N_4850,N_5295);
and U5678 (N_5678,N_5389,N_5267);
and U5679 (N_5679,N_4996,N_5083);
xor U5680 (N_5680,N_4935,N_5118);
or U5681 (N_5681,N_5329,N_4910);
or U5682 (N_5682,N_5186,N_5057);
xnor U5683 (N_5683,N_4893,N_5122);
and U5684 (N_5684,N_5391,N_4939);
nand U5685 (N_5685,N_5121,N_5276);
xor U5686 (N_5686,N_5382,N_5059);
xor U5687 (N_5687,N_5366,N_5136);
nand U5688 (N_5688,N_4852,N_5001);
and U5689 (N_5689,N_5104,N_5143);
nor U5690 (N_5690,N_5068,N_5322);
and U5691 (N_5691,N_5199,N_5072);
nand U5692 (N_5692,N_5349,N_4970);
xnor U5693 (N_5693,N_5343,N_4957);
or U5694 (N_5694,N_5030,N_4865);
or U5695 (N_5695,N_5005,N_5346);
nor U5696 (N_5696,N_5328,N_4873);
nor U5697 (N_5697,N_5369,N_5260);
xnor U5698 (N_5698,N_5189,N_4863);
xor U5699 (N_5699,N_5380,N_4933);
nor U5700 (N_5700,N_5007,N_5319);
and U5701 (N_5701,N_5164,N_5123);
xor U5702 (N_5702,N_4854,N_5156);
xor U5703 (N_5703,N_5082,N_5071);
nand U5704 (N_5704,N_5353,N_5066);
and U5705 (N_5705,N_5252,N_4968);
nor U5706 (N_5706,N_4910,N_5269);
nand U5707 (N_5707,N_5379,N_4813);
xor U5708 (N_5708,N_4953,N_5324);
xor U5709 (N_5709,N_5178,N_4943);
nand U5710 (N_5710,N_5325,N_5053);
xnor U5711 (N_5711,N_5241,N_4961);
xor U5712 (N_5712,N_5196,N_5298);
and U5713 (N_5713,N_4851,N_4984);
nor U5714 (N_5714,N_5392,N_4916);
nor U5715 (N_5715,N_4842,N_5001);
and U5716 (N_5716,N_4915,N_5029);
xor U5717 (N_5717,N_4941,N_5308);
nand U5718 (N_5718,N_5396,N_5326);
xor U5719 (N_5719,N_5198,N_4828);
and U5720 (N_5720,N_4963,N_5304);
and U5721 (N_5721,N_5318,N_4947);
or U5722 (N_5722,N_4970,N_4979);
or U5723 (N_5723,N_5252,N_5069);
nor U5724 (N_5724,N_5303,N_5368);
nand U5725 (N_5725,N_5168,N_5007);
nand U5726 (N_5726,N_5258,N_5327);
and U5727 (N_5727,N_5088,N_5026);
xnor U5728 (N_5728,N_5377,N_4988);
and U5729 (N_5729,N_4981,N_5360);
nand U5730 (N_5730,N_4994,N_4888);
xor U5731 (N_5731,N_5263,N_5304);
xnor U5732 (N_5732,N_5215,N_5348);
and U5733 (N_5733,N_5321,N_4896);
and U5734 (N_5734,N_5158,N_5132);
nor U5735 (N_5735,N_5084,N_5310);
xor U5736 (N_5736,N_5036,N_5375);
nand U5737 (N_5737,N_5056,N_5265);
and U5738 (N_5738,N_5056,N_5316);
xnor U5739 (N_5739,N_4873,N_5165);
nand U5740 (N_5740,N_4967,N_5017);
xor U5741 (N_5741,N_5389,N_4968);
and U5742 (N_5742,N_5002,N_4816);
xnor U5743 (N_5743,N_5191,N_5107);
and U5744 (N_5744,N_4824,N_5021);
nand U5745 (N_5745,N_4809,N_4910);
and U5746 (N_5746,N_5134,N_5114);
nor U5747 (N_5747,N_4809,N_5032);
nor U5748 (N_5748,N_5139,N_5011);
xor U5749 (N_5749,N_5252,N_5186);
nor U5750 (N_5750,N_5093,N_4911);
nor U5751 (N_5751,N_5064,N_5272);
nand U5752 (N_5752,N_4987,N_5306);
and U5753 (N_5753,N_4808,N_4826);
nand U5754 (N_5754,N_4904,N_5339);
and U5755 (N_5755,N_5387,N_4826);
and U5756 (N_5756,N_4874,N_4806);
or U5757 (N_5757,N_5284,N_4848);
or U5758 (N_5758,N_5221,N_5347);
nand U5759 (N_5759,N_5333,N_4867);
or U5760 (N_5760,N_5259,N_5209);
or U5761 (N_5761,N_4982,N_5393);
and U5762 (N_5762,N_5070,N_5251);
or U5763 (N_5763,N_5287,N_5021);
nor U5764 (N_5764,N_5019,N_4801);
nand U5765 (N_5765,N_5236,N_4892);
xnor U5766 (N_5766,N_5252,N_5016);
and U5767 (N_5767,N_4916,N_5294);
nor U5768 (N_5768,N_5222,N_5151);
nand U5769 (N_5769,N_5018,N_5250);
and U5770 (N_5770,N_5159,N_5011);
and U5771 (N_5771,N_5253,N_5387);
nand U5772 (N_5772,N_5256,N_5399);
xor U5773 (N_5773,N_5176,N_4989);
and U5774 (N_5774,N_4890,N_5042);
and U5775 (N_5775,N_4973,N_4886);
xnor U5776 (N_5776,N_5392,N_5142);
and U5777 (N_5777,N_5121,N_4812);
nand U5778 (N_5778,N_5008,N_5005);
nand U5779 (N_5779,N_5204,N_5138);
and U5780 (N_5780,N_5166,N_4850);
or U5781 (N_5781,N_4871,N_5126);
and U5782 (N_5782,N_5240,N_5055);
nand U5783 (N_5783,N_5126,N_5114);
nor U5784 (N_5784,N_5350,N_4878);
nand U5785 (N_5785,N_5226,N_4944);
xnor U5786 (N_5786,N_5387,N_5332);
and U5787 (N_5787,N_5117,N_5061);
nor U5788 (N_5788,N_4823,N_5074);
nand U5789 (N_5789,N_5072,N_5219);
nor U5790 (N_5790,N_5082,N_4953);
nor U5791 (N_5791,N_5322,N_5344);
nand U5792 (N_5792,N_5094,N_4960);
nor U5793 (N_5793,N_4960,N_5354);
or U5794 (N_5794,N_5151,N_5155);
nand U5795 (N_5795,N_4900,N_4865);
nor U5796 (N_5796,N_4821,N_5336);
and U5797 (N_5797,N_5183,N_4847);
xnor U5798 (N_5798,N_4910,N_5343);
xnor U5799 (N_5799,N_5084,N_5058);
and U5800 (N_5800,N_4854,N_4839);
or U5801 (N_5801,N_4809,N_4967);
nor U5802 (N_5802,N_4818,N_4977);
and U5803 (N_5803,N_5299,N_5027);
nand U5804 (N_5804,N_5317,N_4892);
and U5805 (N_5805,N_5213,N_4956);
xor U5806 (N_5806,N_5261,N_4959);
and U5807 (N_5807,N_5338,N_5115);
nor U5808 (N_5808,N_5072,N_5242);
or U5809 (N_5809,N_4960,N_4994);
or U5810 (N_5810,N_5113,N_5025);
nor U5811 (N_5811,N_4909,N_5028);
xor U5812 (N_5812,N_4900,N_5271);
nand U5813 (N_5813,N_4988,N_4922);
nor U5814 (N_5814,N_4909,N_5206);
nand U5815 (N_5815,N_4908,N_5016);
or U5816 (N_5816,N_5244,N_5142);
nor U5817 (N_5817,N_4969,N_5051);
nand U5818 (N_5818,N_5102,N_5027);
and U5819 (N_5819,N_4955,N_4934);
xnor U5820 (N_5820,N_5178,N_5004);
xnor U5821 (N_5821,N_5054,N_4901);
nand U5822 (N_5822,N_4927,N_4986);
xnor U5823 (N_5823,N_5377,N_5298);
xnor U5824 (N_5824,N_4933,N_4965);
and U5825 (N_5825,N_5281,N_5212);
or U5826 (N_5826,N_4887,N_4942);
nand U5827 (N_5827,N_5303,N_4850);
nor U5828 (N_5828,N_5001,N_5150);
nand U5829 (N_5829,N_5125,N_4852);
and U5830 (N_5830,N_5019,N_4821);
and U5831 (N_5831,N_5262,N_5315);
and U5832 (N_5832,N_4881,N_5158);
and U5833 (N_5833,N_4956,N_5291);
or U5834 (N_5834,N_5030,N_5340);
xnor U5835 (N_5835,N_4854,N_4913);
and U5836 (N_5836,N_5293,N_5395);
nand U5837 (N_5837,N_5303,N_4918);
and U5838 (N_5838,N_5225,N_5182);
nand U5839 (N_5839,N_5124,N_4993);
and U5840 (N_5840,N_5182,N_4827);
and U5841 (N_5841,N_5250,N_4807);
xor U5842 (N_5842,N_4835,N_5222);
and U5843 (N_5843,N_5287,N_4925);
nor U5844 (N_5844,N_4976,N_5080);
nand U5845 (N_5845,N_5010,N_4974);
and U5846 (N_5846,N_5001,N_5377);
and U5847 (N_5847,N_5371,N_5136);
xnor U5848 (N_5848,N_5328,N_4866);
xnor U5849 (N_5849,N_4887,N_4889);
or U5850 (N_5850,N_4927,N_5146);
xor U5851 (N_5851,N_5203,N_4861);
or U5852 (N_5852,N_5320,N_5208);
xnor U5853 (N_5853,N_4869,N_5299);
nor U5854 (N_5854,N_5353,N_4801);
nand U5855 (N_5855,N_5114,N_5154);
and U5856 (N_5856,N_5330,N_5115);
nand U5857 (N_5857,N_5104,N_5326);
nor U5858 (N_5858,N_4904,N_4935);
xor U5859 (N_5859,N_5013,N_4996);
nor U5860 (N_5860,N_5321,N_5308);
and U5861 (N_5861,N_5001,N_5166);
and U5862 (N_5862,N_5375,N_5099);
xor U5863 (N_5863,N_4819,N_4935);
and U5864 (N_5864,N_4949,N_5116);
nor U5865 (N_5865,N_5051,N_5362);
or U5866 (N_5866,N_5162,N_4944);
or U5867 (N_5867,N_5315,N_4882);
nor U5868 (N_5868,N_5006,N_4979);
xnor U5869 (N_5869,N_5340,N_5376);
or U5870 (N_5870,N_4985,N_5307);
nor U5871 (N_5871,N_5281,N_5156);
and U5872 (N_5872,N_4901,N_5266);
nor U5873 (N_5873,N_4805,N_5172);
xnor U5874 (N_5874,N_4961,N_4960);
and U5875 (N_5875,N_5367,N_5301);
xnor U5876 (N_5876,N_5068,N_4869);
and U5877 (N_5877,N_5136,N_4992);
nand U5878 (N_5878,N_5123,N_5345);
and U5879 (N_5879,N_5004,N_5286);
nor U5880 (N_5880,N_5186,N_5236);
nor U5881 (N_5881,N_5168,N_4815);
nand U5882 (N_5882,N_5173,N_4887);
and U5883 (N_5883,N_5332,N_4850);
and U5884 (N_5884,N_5046,N_5352);
nand U5885 (N_5885,N_5058,N_5389);
nor U5886 (N_5886,N_5351,N_5308);
nor U5887 (N_5887,N_4825,N_5069);
nor U5888 (N_5888,N_4808,N_5252);
or U5889 (N_5889,N_5042,N_5381);
nor U5890 (N_5890,N_5272,N_4915);
and U5891 (N_5891,N_5058,N_5176);
or U5892 (N_5892,N_4894,N_5010);
and U5893 (N_5893,N_5039,N_5105);
nand U5894 (N_5894,N_5276,N_5133);
nand U5895 (N_5895,N_5047,N_5173);
xor U5896 (N_5896,N_4856,N_5396);
nand U5897 (N_5897,N_4836,N_5163);
nor U5898 (N_5898,N_4931,N_5181);
nor U5899 (N_5899,N_5195,N_5115);
nand U5900 (N_5900,N_4852,N_5292);
xnor U5901 (N_5901,N_5164,N_5258);
xor U5902 (N_5902,N_5074,N_4941);
nand U5903 (N_5903,N_5127,N_4873);
and U5904 (N_5904,N_5072,N_4955);
nand U5905 (N_5905,N_4850,N_5228);
and U5906 (N_5906,N_4843,N_4913);
or U5907 (N_5907,N_5209,N_5030);
and U5908 (N_5908,N_5389,N_5059);
nor U5909 (N_5909,N_5122,N_5168);
and U5910 (N_5910,N_4954,N_4998);
and U5911 (N_5911,N_5189,N_4902);
xnor U5912 (N_5912,N_5385,N_5299);
nor U5913 (N_5913,N_4960,N_4992);
nor U5914 (N_5914,N_4982,N_5111);
and U5915 (N_5915,N_5318,N_5219);
or U5916 (N_5916,N_5221,N_5053);
xnor U5917 (N_5917,N_5264,N_5298);
nand U5918 (N_5918,N_5290,N_5084);
and U5919 (N_5919,N_5325,N_5081);
or U5920 (N_5920,N_5006,N_5083);
nand U5921 (N_5921,N_5077,N_5215);
nor U5922 (N_5922,N_5009,N_5067);
xor U5923 (N_5923,N_5197,N_5023);
or U5924 (N_5924,N_5117,N_4961);
nor U5925 (N_5925,N_5202,N_5288);
or U5926 (N_5926,N_4880,N_5133);
and U5927 (N_5927,N_4849,N_4955);
and U5928 (N_5928,N_4869,N_5091);
and U5929 (N_5929,N_5348,N_5301);
nor U5930 (N_5930,N_4908,N_5155);
or U5931 (N_5931,N_4988,N_4968);
or U5932 (N_5932,N_4836,N_4820);
nand U5933 (N_5933,N_5109,N_4926);
xor U5934 (N_5934,N_5159,N_5162);
nor U5935 (N_5935,N_5111,N_5223);
xor U5936 (N_5936,N_5100,N_5230);
nor U5937 (N_5937,N_5234,N_5245);
nor U5938 (N_5938,N_5308,N_4922);
or U5939 (N_5939,N_5101,N_4889);
nor U5940 (N_5940,N_5060,N_5203);
nand U5941 (N_5941,N_5129,N_5152);
nand U5942 (N_5942,N_5105,N_5024);
and U5943 (N_5943,N_4985,N_5155);
xnor U5944 (N_5944,N_5141,N_5273);
xnor U5945 (N_5945,N_5131,N_5175);
or U5946 (N_5946,N_4859,N_4880);
xnor U5947 (N_5947,N_5145,N_5342);
and U5948 (N_5948,N_4863,N_5342);
and U5949 (N_5949,N_5117,N_5080);
or U5950 (N_5950,N_5261,N_4899);
nor U5951 (N_5951,N_5215,N_5282);
xnor U5952 (N_5952,N_5042,N_5204);
nor U5953 (N_5953,N_5043,N_5193);
xnor U5954 (N_5954,N_5106,N_5144);
nand U5955 (N_5955,N_5082,N_5106);
and U5956 (N_5956,N_5266,N_5248);
nor U5957 (N_5957,N_4842,N_4872);
nor U5958 (N_5958,N_4883,N_5164);
and U5959 (N_5959,N_5157,N_5145);
and U5960 (N_5960,N_5214,N_5138);
xor U5961 (N_5961,N_5127,N_4994);
nor U5962 (N_5962,N_4835,N_4803);
xor U5963 (N_5963,N_5314,N_5077);
xnor U5964 (N_5964,N_4918,N_5231);
nor U5965 (N_5965,N_4951,N_4961);
nor U5966 (N_5966,N_4960,N_5329);
xor U5967 (N_5967,N_5247,N_5017);
or U5968 (N_5968,N_5281,N_4879);
xor U5969 (N_5969,N_5307,N_5073);
xor U5970 (N_5970,N_5378,N_5055);
nand U5971 (N_5971,N_5076,N_5354);
nand U5972 (N_5972,N_4933,N_5372);
nor U5973 (N_5973,N_5312,N_4972);
and U5974 (N_5974,N_4891,N_4903);
or U5975 (N_5975,N_4882,N_5384);
and U5976 (N_5976,N_5319,N_5276);
and U5977 (N_5977,N_5009,N_4870);
and U5978 (N_5978,N_5200,N_5183);
nor U5979 (N_5979,N_4823,N_4916);
or U5980 (N_5980,N_4959,N_5030);
xnor U5981 (N_5981,N_5160,N_5275);
nand U5982 (N_5982,N_4833,N_5388);
nor U5983 (N_5983,N_5263,N_5108);
nor U5984 (N_5984,N_5064,N_5179);
xor U5985 (N_5985,N_4808,N_4990);
or U5986 (N_5986,N_5304,N_5006);
or U5987 (N_5987,N_5106,N_4980);
or U5988 (N_5988,N_4859,N_5338);
or U5989 (N_5989,N_5075,N_5146);
or U5990 (N_5990,N_5393,N_5199);
xnor U5991 (N_5991,N_5343,N_5087);
and U5992 (N_5992,N_5148,N_5322);
or U5993 (N_5993,N_5222,N_5068);
nand U5994 (N_5994,N_5369,N_4873);
xor U5995 (N_5995,N_5089,N_5360);
nor U5996 (N_5996,N_5217,N_4868);
and U5997 (N_5997,N_5247,N_5262);
and U5998 (N_5998,N_5099,N_5271);
nand U5999 (N_5999,N_5041,N_5013);
xor U6000 (N_6000,N_5627,N_5447);
xor U6001 (N_6001,N_5963,N_5836);
xor U6002 (N_6002,N_5976,N_5639);
nor U6003 (N_6003,N_5427,N_5949);
nor U6004 (N_6004,N_5665,N_5497);
xnor U6005 (N_6005,N_5944,N_5692);
xor U6006 (N_6006,N_5700,N_5844);
xor U6007 (N_6007,N_5551,N_5955);
nand U6008 (N_6008,N_5673,N_5459);
nor U6009 (N_6009,N_5578,N_5643);
nand U6010 (N_6010,N_5406,N_5542);
xor U6011 (N_6011,N_5464,N_5915);
and U6012 (N_6012,N_5428,N_5531);
nor U6013 (N_6013,N_5908,N_5999);
xnor U6014 (N_6014,N_5481,N_5450);
and U6015 (N_6015,N_5588,N_5859);
nand U6016 (N_6016,N_5806,N_5989);
or U6017 (N_6017,N_5528,N_5581);
nand U6018 (N_6018,N_5852,N_5633);
nor U6019 (N_6019,N_5930,N_5832);
xnor U6020 (N_6020,N_5453,N_5722);
xor U6021 (N_6021,N_5672,N_5443);
or U6022 (N_6022,N_5843,N_5761);
and U6023 (N_6023,N_5462,N_5599);
nor U6024 (N_6024,N_5460,N_5540);
xnor U6025 (N_6025,N_5681,N_5650);
nor U6026 (N_6026,N_5611,N_5765);
xor U6027 (N_6027,N_5417,N_5845);
nand U6028 (N_6028,N_5544,N_5704);
and U6029 (N_6029,N_5757,N_5828);
xor U6030 (N_6030,N_5425,N_5532);
nand U6031 (N_6031,N_5418,N_5966);
or U6032 (N_6032,N_5538,N_5810);
xor U6033 (N_6033,N_5735,N_5726);
xnor U6034 (N_6034,N_5896,N_5719);
nor U6035 (N_6035,N_5543,N_5485);
and U6036 (N_6036,N_5594,N_5880);
xor U6037 (N_6037,N_5632,N_5519);
xor U6038 (N_6038,N_5920,N_5940);
xnor U6039 (N_6039,N_5798,N_5463);
or U6040 (N_6040,N_5925,N_5946);
or U6041 (N_6041,N_5970,N_5756);
or U6042 (N_6042,N_5817,N_5648);
and U6043 (N_6043,N_5939,N_5931);
or U6044 (N_6044,N_5446,N_5960);
nand U6045 (N_6045,N_5723,N_5589);
nor U6046 (N_6046,N_5834,N_5616);
or U6047 (N_6047,N_5951,N_5554);
or U6048 (N_6048,N_5548,N_5789);
nand U6049 (N_6049,N_5786,N_5858);
or U6050 (N_6050,N_5586,N_5559);
or U6051 (N_6051,N_5861,N_5598);
nor U6052 (N_6052,N_5558,N_5449);
and U6053 (N_6053,N_5985,N_5936);
and U6054 (N_6054,N_5779,N_5678);
nand U6055 (N_6055,N_5910,N_5675);
nand U6056 (N_6056,N_5452,N_5855);
xnor U6057 (N_6057,N_5711,N_5833);
nand U6058 (N_6058,N_5465,N_5792);
and U6059 (N_6059,N_5895,N_5630);
xor U6060 (N_6060,N_5827,N_5610);
xor U6061 (N_6061,N_5888,N_5900);
xnor U6062 (N_6062,N_5430,N_5890);
and U6063 (N_6063,N_5432,N_5620);
nand U6064 (N_6064,N_5699,N_5518);
nor U6065 (N_6065,N_5736,N_5902);
and U6066 (N_6066,N_5771,N_5776);
or U6067 (N_6067,N_5794,N_5444);
or U6068 (N_6068,N_5402,N_5635);
and U6069 (N_6069,N_5609,N_5868);
nand U6070 (N_6070,N_5911,N_5937);
nand U6071 (N_6071,N_5929,N_5835);
nor U6072 (N_6072,N_5912,N_5516);
and U6073 (N_6073,N_5893,N_5965);
nand U6074 (N_6074,N_5494,N_5696);
nor U6075 (N_6075,N_5524,N_5873);
and U6076 (N_6076,N_5802,N_5811);
nand U6077 (N_6077,N_5694,N_5793);
and U6078 (N_6078,N_5714,N_5891);
and U6079 (N_6079,N_5987,N_5746);
or U6080 (N_6080,N_5788,N_5731);
or U6081 (N_6081,N_5458,N_5654);
xnor U6082 (N_6082,N_5809,N_5864);
nand U6083 (N_6083,N_5437,N_5964);
nand U6084 (N_6084,N_5472,N_5721);
xor U6085 (N_6085,N_5935,N_5954);
and U6086 (N_6086,N_5766,N_5831);
or U6087 (N_6087,N_5566,N_5928);
nor U6088 (N_6088,N_5480,N_5981);
or U6089 (N_6089,N_5737,N_5667);
xor U6090 (N_6090,N_5943,N_5419);
xnor U6091 (N_6091,N_5805,N_5530);
and U6092 (N_6092,N_5784,N_5884);
and U6093 (N_6093,N_5431,N_5603);
or U6094 (N_6094,N_5770,N_5718);
and U6095 (N_6095,N_5568,N_5569);
xor U6096 (N_6096,N_5872,N_5708);
nor U6097 (N_6097,N_5772,N_5584);
and U6098 (N_6098,N_5555,N_5492);
and U6099 (N_6099,N_5433,N_5663);
nand U6100 (N_6100,N_5838,N_5898);
xor U6101 (N_6101,N_5400,N_5442);
nor U6102 (N_6102,N_5749,N_5822);
xnor U6103 (N_6103,N_5881,N_5514);
and U6104 (N_6104,N_5408,N_5753);
nand U6105 (N_6105,N_5475,N_5968);
nand U6106 (N_6106,N_5661,N_5591);
nor U6107 (N_6107,N_5875,N_5471);
and U6108 (N_6108,N_5580,N_5649);
nand U6109 (N_6109,N_5897,N_5874);
nor U6110 (N_6110,N_5579,N_5682);
and U6111 (N_6111,N_5647,N_5695);
xnor U6112 (N_6112,N_5655,N_5483);
nor U6113 (N_6113,N_5903,N_5560);
or U6114 (N_6114,N_5972,N_5950);
or U6115 (N_6115,N_5992,N_5819);
xor U6116 (N_6116,N_5814,N_5993);
and U6117 (N_6117,N_5886,N_5693);
or U6118 (N_6118,N_5642,N_5644);
nand U6119 (N_6119,N_5619,N_5924);
nor U6120 (N_6120,N_5854,N_5758);
xor U6121 (N_6121,N_5601,N_5407);
nand U6122 (N_6122,N_5501,N_5747);
xnor U6123 (N_6123,N_5550,N_5583);
and U6124 (N_6124,N_5426,N_5973);
nand U6125 (N_6125,N_5984,N_5669);
and U6126 (N_6126,N_5625,N_5489);
and U6127 (N_6127,N_5780,N_5597);
nand U6128 (N_6128,N_5752,N_5813);
or U6129 (N_6129,N_5919,N_5905);
and U6130 (N_6130,N_5961,N_5913);
and U6131 (N_6131,N_5659,N_5680);
or U6132 (N_6132,N_5434,N_5690);
nor U6133 (N_6133,N_5503,N_5743);
xor U6134 (N_6134,N_5640,N_5487);
nor U6135 (N_6135,N_5849,N_5707);
or U6136 (N_6136,N_5552,N_5730);
xor U6137 (N_6137,N_5529,N_5498);
nand U6138 (N_6138,N_5573,N_5688);
and U6139 (N_6139,N_5729,N_5435);
or U6140 (N_6140,N_5674,N_5741);
nand U6141 (N_6141,N_5512,N_5783);
and U6142 (N_6142,N_5710,N_5713);
xnor U6143 (N_6143,N_5851,N_5456);
nand U6144 (N_6144,N_5429,N_5777);
and U6145 (N_6145,N_5523,N_5775);
and U6146 (N_6146,N_5445,N_5755);
nor U6147 (N_6147,N_5816,N_5509);
xor U6148 (N_6148,N_5575,N_5623);
and U6149 (N_6149,N_5926,N_5917);
xnor U6150 (N_6150,N_5797,N_5701);
or U6151 (N_6151,N_5706,N_5799);
xnor U6152 (N_6152,N_5956,N_5837);
and U6153 (N_6153,N_5505,N_5561);
and U6154 (N_6154,N_5488,N_5894);
nor U6155 (N_6155,N_5739,N_5995);
xor U6156 (N_6156,N_5605,N_5942);
or U6157 (N_6157,N_5933,N_5879);
nand U6158 (N_6158,N_5687,N_5994);
nand U6159 (N_6159,N_5909,N_5820);
nand U6160 (N_6160,N_5556,N_5716);
xor U6161 (N_6161,N_5405,N_5764);
nand U6162 (N_6162,N_5732,N_5698);
and U6163 (N_6163,N_5626,N_5439);
xor U6164 (N_6164,N_5998,N_5959);
or U6165 (N_6165,N_5549,N_5495);
nor U6166 (N_6166,N_5490,N_5724);
xor U6167 (N_6167,N_5750,N_5657);
xnor U6168 (N_6168,N_5604,N_5803);
nand U6169 (N_6169,N_5684,N_5638);
nor U6170 (N_6170,N_5593,N_5479);
nor U6171 (N_6171,N_5697,N_5889);
nor U6172 (N_6172,N_5451,N_5829);
xor U6173 (N_6173,N_5997,N_5787);
and U6174 (N_6174,N_5740,N_5602);
nor U6175 (N_6175,N_5742,N_5904);
nand U6176 (N_6176,N_5839,N_5536);
nor U6177 (N_6177,N_5653,N_5424);
or U6178 (N_6178,N_5570,N_5870);
nor U6179 (N_6179,N_5941,N_5751);
xor U6180 (N_6180,N_5971,N_5728);
or U6181 (N_6181,N_5702,N_5582);
xnor U6182 (N_6182,N_5423,N_5745);
nand U6183 (N_6183,N_5470,N_5860);
nor U6184 (N_6184,N_5847,N_5482);
or U6185 (N_6185,N_5507,N_5520);
and U6186 (N_6186,N_5760,N_5795);
xor U6187 (N_6187,N_5823,N_5825);
and U6188 (N_6188,N_5521,N_5991);
or U6189 (N_6189,N_5486,N_5785);
and U6190 (N_6190,N_5945,N_5807);
and U6191 (N_6191,N_5685,N_5414);
nor U6192 (N_6192,N_5767,N_5763);
xnor U6193 (N_6193,N_5754,N_5922);
nand U6194 (N_6194,N_5469,N_5637);
xor U6195 (N_6195,N_5413,N_5508);
xnor U6196 (N_6196,N_5869,N_5476);
xnor U6197 (N_6197,N_5411,N_5666);
and U6198 (N_6198,N_5484,N_5978);
nand U6199 (N_6199,N_5448,N_5914);
xor U6200 (N_6200,N_5422,N_5404);
and U6201 (N_6201,N_5537,N_5618);
nor U6202 (N_6202,N_5867,N_5615);
nand U6203 (N_6203,N_5441,N_5934);
nor U6204 (N_6204,N_5821,N_5790);
or U6205 (N_6205,N_5842,N_5474);
nand U6206 (N_6206,N_5535,N_5907);
nor U6207 (N_6207,N_5656,N_5634);
or U6208 (N_6208,N_5906,N_5982);
xnor U6209 (N_6209,N_5557,N_5545);
or U6210 (N_6210,N_5796,N_5436);
and U6211 (N_6211,N_5502,N_5641);
xnor U6212 (N_6212,N_5467,N_5515);
or U6213 (N_6213,N_5608,N_5988);
and U6214 (N_6214,N_5636,N_5979);
xor U6215 (N_6215,N_5967,N_5720);
or U6216 (N_6216,N_5878,N_5815);
xor U6217 (N_6217,N_5553,N_5607);
nand U6218 (N_6218,N_5613,N_5774);
nor U6219 (N_6219,N_5477,N_5525);
xnor U6220 (N_6220,N_5791,N_5952);
nor U6221 (N_6221,N_5679,N_5500);
nor U6222 (N_6222,N_5725,N_5883);
nand U6223 (N_6223,N_5778,N_5932);
nand U6224 (N_6224,N_5923,N_5671);
xor U6225 (N_6225,N_5969,N_5668);
nor U6226 (N_6226,N_5617,N_5606);
or U6227 (N_6227,N_5662,N_5958);
nor U6228 (N_6228,N_5717,N_5440);
xor U6229 (N_6229,N_5808,N_5782);
and U6230 (N_6230,N_5689,N_5401);
nor U6231 (N_6231,N_5403,N_5534);
nor U6232 (N_6232,N_5415,N_5983);
nor U6233 (N_6233,N_5703,N_5614);
nor U6234 (N_6234,N_5980,N_5840);
and U6235 (N_6235,N_5712,N_5499);
and U6236 (N_6236,N_5748,N_5734);
xor U6237 (N_6237,N_5533,N_5596);
xor U6238 (N_6238,N_5812,N_5562);
and U6239 (N_6239,N_5759,N_5709);
xnor U6240 (N_6240,N_5478,N_5841);
xor U6241 (N_6241,N_5491,N_5801);
nand U6242 (N_6242,N_5975,N_5691);
xor U6243 (N_6243,N_5916,N_5493);
nand U6244 (N_6244,N_5658,N_5866);
or U6245 (N_6245,N_5660,N_5670);
nor U6246 (N_6246,N_5567,N_5585);
or U6247 (N_6247,N_5438,N_5865);
or U6248 (N_6248,N_5574,N_5612);
nand U6249 (N_6249,N_5590,N_5409);
or U6250 (N_6250,N_5738,N_5565);
and U6251 (N_6251,N_5517,N_5526);
and U6252 (N_6252,N_5877,N_5629);
nor U6253 (N_6253,N_5927,N_5546);
xor U6254 (N_6254,N_5563,N_5818);
nor U6255 (N_6255,N_5587,N_5473);
and U6256 (N_6256,N_5921,N_5504);
nor U6257 (N_6257,N_5621,N_5769);
and U6258 (N_6258,N_5899,N_5773);
nand U6259 (N_6259,N_5938,N_5466);
nand U6260 (N_6260,N_5676,N_5974);
or U6261 (N_6261,N_5513,N_5622);
nor U6262 (N_6262,N_5850,N_5876);
or U6263 (N_6263,N_5727,N_5651);
or U6264 (N_6264,N_5600,N_5645);
and U6265 (N_6265,N_5857,N_5901);
xnor U6266 (N_6266,N_5804,N_5768);
or U6267 (N_6267,N_5421,N_5416);
xnor U6268 (N_6268,N_5506,N_5522);
nor U6269 (N_6269,N_5830,N_5628);
xor U6270 (N_6270,N_5592,N_5631);
or U6271 (N_6271,N_5541,N_5457);
xnor U6272 (N_6272,N_5686,N_5576);
nor U6273 (N_6273,N_5420,N_5762);
xor U6274 (N_6274,N_5683,N_5715);
or U6275 (N_6275,N_5595,N_5410);
nor U6276 (N_6276,N_5885,N_5953);
or U6277 (N_6277,N_5948,N_5511);
xnor U6278 (N_6278,N_5957,N_5744);
and U6279 (N_6279,N_5624,N_5527);
nor U6280 (N_6280,N_5800,N_5547);
nor U6281 (N_6281,N_5412,N_5496);
and U6282 (N_6282,N_5781,N_5990);
xor U6283 (N_6283,N_5882,N_5539);
xnor U6284 (N_6284,N_5646,N_5918);
nor U6285 (N_6285,N_5962,N_5846);
xnor U6286 (N_6286,N_5848,N_5824);
nor U6287 (N_6287,N_5862,N_5677);
and U6288 (N_6288,N_5871,N_5947);
and U6289 (N_6289,N_5564,N_5572);
nand U6290 (N_6290,N_5664,N_5510);
or U6291 (N_6291,N_5892,N_5733);
nand U6292 (N_6292,N_5977,N_5571);
xor U6293 (N_6293,N_5856,N_5652);
nand U6294 (N_6294,N_5853,N_5887);
nor U6295 (N_6295,N_5986,N_5455);
xor U6296 (N_6296,N_5468,N_5577);
nor U6297 (N_6297,N_5454,N_5461);
nor U6298 (N_6298,N_5863,N_5996);
nor U6299 (N_6299,N_5826,N_5705);
and U6300 (N_6300,N_5866,N_5796);
and U6301 (N_6301,N_5897,N_5808);
nor U6302 (N_6302,N_5707,N_5770);
nor U6303 (N_6303,N_5890,N_5783);
xnor U6304 (N_6304,N_5798,N_5580);
nor U6305 (N_6305,N_5604,N_5826);
nor U6306 (N_6306,N_5514,N_5554);
or U6307 (N_6307,N_5820,N_5464);
xnor U6308 (N_6308,N_5493,N_5586);
nor U6309 (N_6309,N_5865,N_5993);
and U6310 (N_6310,N_5669,N_5525);
and U6311 (N_6311,N_5500,N_5979);
or U6312 (N_6312,N_5401,N_5725);
nor U6313 (N_6313,N_5957,N_5611);
and U6314 (N_6314,N_5526,N_5780);
nor U6315 (N_6315,N_5456,N_5587);
or U6316 (N_6316,N_5986,N_5440);
xnor U6317 (N_6317,N_5463,N_5445);
nor U6318 (N_6318,N_5889,N_5543);
nand U6319 (N_6319,N_5451,N_5578);
and U6320 (N_6320,N_5900,N_5539);
or U6321 (N_6321,N_5515,N_5998);
nor U6322 (N_6322,N_5754,N_5851);
and U6323 (N_6323,N_5400,N_5499);
or U6324 (N_6324,N_5941,N_5435);
nand U6325 (N_6325,N_5935,N_5882);
xor U6326 (N_6326,N_5437,N_5653);
xor U6327 (N_6327,N_5465,N_5618);
nand U6328 (N_6328,N_5949,N_5579);
and U6329 (N_6329,N_5637,N_5663);
nand U6330 (N_6330,N_5575,N_5647);
or U6331 (N_6331,N_5607,N_5500);
nor U6332 (N_6332,N_5576,N_5508);
xor U6333 (N_6333,N_5745,N_5515);
xnor U6334 (N_6334,N_5929,N_5979);
nand U6335 (N_6335,N_5783,N_5959);
and U6336 (N_6336,N_5922,N_5847);
xnor U6337 (N_6337,N_5478,N_5797);
nand U6338 (N_6338,N_5564,N_5728);
and U6339 (N_6339,N_5474,N_5699);
xor U6340 (N_6340,N_5843,N_5466);
and U6341 (N_6341,N_5991,N_5553);
nor U6342 (N_6342,N_5887,N_5595);
nand U6343 (N_6343,N_5845,N_5674);
nand U6344 (N_6344,N_5735,N_5487);
or U6345 (N_6345,N_5721,N_5772);
xor U6346 (N_6346,N_5662,N_5628);
nand U6347 (N_6347,N_5954,N_5829);
or U6348 (N_6348,N_5444,N_5424);
xnor U6349 (N_6349,N_5560,N_5767);
or U6350 (N_6350,N_5818,N_5997);
xnor U6351 (N_6351,N_5464,N_5899);
xor U6352 (N_6352,N_5752,N_5700);
nand U6353 (N_6353,N_5526,N_5516);
nand U6354 (N_6354,N_5859,N_5616);
xnor U6355 (N_6355,N_5734,N_5770);
and U6356 (N_6356,N_5917,N_5594);
nand U6357 (N_6357,N_5709,N_5649);
or U6358 (N_6358,N_5833,N_5485);
nand U6359 (N_6359,N_5765,N_5460);
or U6360 (N_6360,N_5440,N_5631);
nand U6361 (N_6361,N_5995,N_5638);
and U6362 (N_6362,N_5826,N_5538);
nor U6363 (N_6363,N_5836,N_5663);
and U6364 (N_6364,N_5902,N_5744);
xor U6365 (N_6365,N_5698,N_5886);
nand U6366 (N_6366,N_5984,N_5723);
or U6367 (N_6367,N_5883,N_5795);
nor U6368 (N_6368,N_5624,N_5640);
nand U6369 (N_6369,N_5685,N_5878);
nor U6370 (N_6370,N_5471,N_5641);
xor U6371 (N_6371,N_5764,N_5863);
xor U6372 (N_6372,N_5564,N_5500);
xor U6373 (N_6373,N_5824,N_5693);
nand U6374 (N_6374,N_5472,N_5646);
xor U6375 (N_6375,N_5553,N_5484);
nor U6376 (N_6376,N_5724,N_5644);
and U6377 (N_6377,N_5954,N_5817);
xnor U6378 (N_6378,N_5486,N_5649);
nor U6379 (N_6379,N_5526,N_5721);
or U6380 (N_6380,N_5549,N_5460);
xnor U6381 (N_6381,N_5889,N_5911);
or U6382 (N_6382,N_5813,N_5444);
xnor U6383 (N_6383,N_5723,N_5667);
and U6384 (N_6384,N_5795,N_5877);
nor U6385 (N_6385,N_5599,N_5813);
xor U6386 (N_6386,N_5859,N_5715);
nand U6387 (N_6387,N_5536,N_5478);
xnor U6388 (N_6388,N_5763,N_5593);
nor U6389 (N_6389,N_5894,N_5562);
nand U6390 (N_6390,N_5871,N_5572);
xor U6391 (N_6391,N_5976,N_5468);
xnor U6392 (N_6392,N_5975,N_5822);
nor U6393 (N_6393,N_5808,N_5410);
and U6394 (N_6394,N_5600,N_5652);
or U6395 (N_6395,N_5638,N_5602);
and U6396 (N_6396,N_5717,N_5959);
nand U6397 (N_6397,N_5884,N_5991);
or U6398 (N_6398,N_5483,N_5809);
or U6399 (N_6399,N_5414,N_5795);
xnor U6400 (N_6400,N_5475,N_5670);
nand U6401 (N_6401,N_5441,N_5659);
and U6402 (N_6402,N_5986,N_5464);
xnor U6403 (N_6403,N_5426,N_5971);
or U6404 (N_6404,N_5642,N_5423);
and U6405 (N_6405,N_5683,N_5541);
nand U6406 (N_6406,N_5677,N_5940);
or U6407 (N_6407,N_5955,N_5569);
xnor U6408 (N_6408,N_5654,N_5975);
or U6409 (N_6409,N_5516,N_5523);
nor U6410 (N_6410,N_5614,N_5867);
nor U6411 (N_6411,N_5501,N_5628);
or U6412 (N_6412,N_5409,N_5688);
or U6413 (N_6413,N_5401,N_5617);
nor U6414 (N_6414,N_5991,N_5668);
nor U6415 (N_6415,N_5602,N_5982);
nor U6416 (N_6416,N_5879,N_5556);
nand U6417 (N_6417,N_5767,N_5434);
xnor U6418 (N_6418,N_5480,N_5824);
or U6419 (N_6419,N_5459,N_5752);
and U6420 (N_6420,N_5517,N_5983);
xnor U6421 (N_6421,N_5574,N_5698);
and U6422 (N_6422,N_5595,N_5886);
or U6423 (N_6423,N_5968,N_5681);
nor U6424 (N_6424,N_5492,N_5970);
or U6425 (N_6425,N_5831,N_5422);
nand U6426 (N_6426,N_5796,N_5907);
xnor U6427 (N_6427,N_5498,N_5485);
xnor U6428 (N_6428,N_5530,N_5745);
and U6429 (N_6429,N_5412,N_5750);
or U6430 (N_6430,N_5668,N_5620);
nand U6431 (N_6431,N_5494,N_5458);
xnor U6432 (N_6432,N_5448,N_5618);
nand U6433 (N_6433,N_5892,N_5473);
or U6434 (N_6434,N_5748,N_5896);
or U6435 (N_6435,N_5512,N_5469);
nand U6436 (N_6436,N_5554,N_5431);
nand U6437 (N_6437,N_5673,N_5789);
and U6438 (N_6438,N_5886,N_5502);
or U6439 (N_6439,N_5946,N_5594);
or U6440 (N_6440,N_5848,N_5659);
xor U6441 (N_6441,N_5740,N_5714);
nand U6442 (N_6442,N_5688,N_5497);
or U6443 (N_6443,N_5857,N_5410);
nand U6444 (N_6444,N_5589,N_5772);
xnor U6445 (N_6445,N_5936,N_5729);
or U6446 (N_6446,N_5564,N_5714);
or U6447 (N_6447,N_5478,N_5838);
and U6448 (N_6448,N_5676,N_5912);
nor U6449 (N_6449,N_5982,N_5757);
nand U6450 (N_6450,N_5997,N_5762);
and U6451 (N_6451,N_5872,N_5649);
and U6452 (N_6452,N_5586,N_5480);
nor U6453 (N_6453,N_5967,N_5525);
nand U6454 (N_6454,N_5868,N_5937);
or U6455 (N_6455,N_5878,N_5807);
and U6456 (N_6456,N_5711,N_5650);
xor U6457 (N_6457,N_5809,N_5408);
or U6458 (N_6458,N_5547,N_5504);
and U6459 (N_6459,N_5982,N_5608);
or U6460 (N_6460,N_5623,N_5756);
or U6461 (N_6461,N_5962,N_5980);
nand U6462 (N_6462,N_5404,N_5920);
xnor U6463 (N_6463,N_5964,N_5684);
nor U6464 (N_6464,N_5674,N_5605);
or U6465 (N_6465,N_5759,N_5414);
and U6466 (N_6466,N_5634,N_5803);
nor U6467 (N_6467,N_5402,N_5805);
nand U6468 (N_6468,N_5631,N_5983);
nor U6469 (N_6469,N_5855,N_5781);
nand U6470 (N_6470,N_5469,N_5462);
nand U6471 (N_6471,N_5712,N_5400);
and U6472 (N_6472,N_5981,N_5967);
nor U6473 (N_6473,N_5638,N_5767);
xnor U6474 (N_6474,N_5876,N_5514);
or U6475 (N_6475,N_5686,N_5496);
xor U6476 (N_6476,N_5741,N_5508);
nor U6477 (N_6477,N_5628,N_5947);
nor U6478 (N_6478,N_5983,N_5901);
or U6479 (N_6479,N_5770,N_5939);
xor U6480 (N_6480,N_5525,N_5812);
xor U6481 (N_6481,N_5439,N_5647);
xnor U6482 (N_6482,N_5507,N_5447);
xnor U6483 (N_6483,N_5490,N_5532);
nand U6484 (N_6484,N_5891,N_5565);
and U6485 (N_6485,N_5460,N_5436);
xnor U6486 (N_6486,N_5517,N_5823);
nor U6487 (N_6487,N_5990,N_5980);
or U6488 (N_6488,N_5471,N_5592);
and U6489 (N_6489,N_5900,N_5503);
nor U6490 (N_6490,N_5954,N_5549);
and U6491 (N_6491,N_5455,N_5957);
nor U6492 (N_6492,N_5413,N_5701);
xnor U6493 (N_6493,N_5832,N_5992);
and U6494 (N_6494,N_5586,N_5624);
nor U6495 (N_6495,N_5851,N_5644);
xor U6496 (N_6496,N_5817,N_5484);
xnor U6497 (N_6497,N_5990,N_5814);
nor U6498 (N_6498,N_5766,N_5944);
and U6499 (N_6499,N_5964,N_5966);
nand U6500 (N_6500,N_5743,N_5417);
and U6501 (N_6501,N_5719,N_5591);
and U6502 (N_6502,N_5516,N_5654);
and U6503 (N_6503,N_5816,N_5560);
nor U6504 (N_6504,N_5603,N_5401);
and U6505 (N_6505,N_5551,N_5570);
nand U6506 (N_6506,N_5576,N_5903);
nor U6507 (N_6507,N_5953,N_5632);
and U6508 (N_6508,N_5797,N_5545);
or U6509 (N_6509,N_5691,N_5867);
nor U6510 (N_6510,N_5650,N_5677);
xnor U6511 (N_6511,N_5641,N_5659);
nor U6512 (N_6512,N_5891,N_5661);
and U6513 (N_6513,N_5766,N_5605);
and U6514 (N_6514,N_5849,N_5656);
or U6515 (N_6515,N_5768,N_5787);
nand U6516 (N_6516,N_5629,N_5548);
nor U6517 (N_6517,N_5750,N_5852);
or U6518 (N_6518,N_5801,N_5925);
or U6519 (N_6519,N_5604,N_5521);
and U6520 (N_6520,N_5584,N_5505);
nor U6521 (N_6521,N_5699,N_5471);
and U6522 (N_6522,N_5693,N_5567);
nor U6523 (N_6523,N_5406,N_5987);
or U6524 (N_6524,N_5600,N_5646);
nor U6525 (N_6525,N_5797,N_5441);
or U6526 (N_6526,N_5617,N_5849);
nand U6527 (N_6527,N_5464,N_5642);
and U6528 (N_6528,N_5520,N_5418);
nand U6529 (N_6529,N_5892,N_5687);
xnor U6530 (N_6530,N_5716,N_5738);
and U6531 (N_6531,N_5596,N_5975);
nand U6532 (N_6532,N_5669,N_5693);
xor U6533 (N_6533,N_5784,N_5970);
or U6534 (N_6534,N_5725,N_5666);
and U6535 (N_6535,N_5983,N_5789);
nor U6536 (N_6536,N_5846,N_5853);
or U6537 (N_6537,N_5847,N_5595);
and U6538 (N_6538,N_5787,N_5917);
nand U6539 (N_6539,N_5955,N_5543);
or U6540 (N_6540,N_5942,N_5537);
and U6541 (N_6541,N_5944,N_5574);
nand U6542 (N_6542,N_5973,N_5563);
and U6543 (N_6543,N_5943,N_5665);
nor U6544 (N_6544,N_5849,N_5454);
nand U6545 (N_6545,N_5797,N_5591);
nand U6546 (N_6546,N_5745,N_5813);
and U6547 (N_6547,N_5689,N_5736);
nor U6548 (N_6548,N_5641,N_5933);
and U6549 (N_6549,N_5779,N_5839);
or U6550 (N_6550,N_5419,N_5712);
or U6551 (N_6551,N_5835,N_5940);
xnor U6552 (N_6552,N_5829,N_5516);
or U6553 (N_6553,N_5625,N_5537);
nand U6554 (N_6554,N_5935,N_5428);
nand U6555 (N_6555,N_5808,N_5646);
nand U6556 (N_6556,N_5906,N_5574);
xor U6557 (N_6557,N_5659,N_5966);
nand U6558 (N_6558,N_5862,N_5698);
and U6559 (N_6559,N_5753,N_5804);
or U6560 (N_6560,N_5886,N_5573);
nor U6561 (N_6561,N_5516,N_5977);
nor U6562 (N_6562,N_5458,N_5879);
xnor U6563 (N_6563,N_5740,N_5754);
nand U6564 (N_6564,N_5504,N_5798);
nand U6565 (N_6565,N_5496,N_5443);
nor U6566 (N_6566,N_5403,N_5883);
nor U6567 (N_6567,N_5625,N_5849);
and U6568 (N_6568,N_5868,N_5752);
nor U6569 (N_6569,N_5833,N_5801);
nor U6570 (N_6570,N_5952,N_5680);
and U6571 (N_6571,N_5500,N_5668);
nor U6572 (N_6572,N_5994,N_5543);
nor U6573 (N_6573,N_5438,N_5962);
nor U6574 (N_6574,N_5708,N_5964);
nor U6575 (N_6575,N_5492,N_5627);
nand U6576 (N_6576,N_5411,N_5688);
xnor U6577 (N_6577,N_5787,N_5515);
nand U6578 (N_6578,N_5445,N_5422);
nor U6579 (N_6579,N_5495,N_5857);
xnor U6580 (N_6580,N_5925,N_5750);
nor U6581 (N_6581,N_5502,N_5490);
xor U6582 (N_6582,N_5952,N_5499);
and U6583 (N_6583,N_5996,N_5952);
and U6584 (N_6584,N_5895,N_5580);
xnor U6585 (N_6585,N_5981,N_5552);
or U6586 (N_6586,N_5810,N_5428);
xnor U6587 (N_6587,N_5683,N_5914);
nand U6588 (N_6588,N_5996,N_5942);
nor U6589 (N_6589,N_5460,N_5802);
or U6590 (N_6590,N_5941,N_5936);
xnor U6591 (N_6591,N_5765,N_5572);
xor U6592 (N_6592,N_5401,N_5654);
or U6593 (N_6593,N_5820,N_5615);
and U6594 (N_6594,N_5882,N_5884);
and U6595 (N_6595,N_5663,N_5592);
nand U6596 (N_6596,N_5423,N_5990);
xor U6597 (N_6597,N_5707,N_5734);
nor U6598 (N_6598,N_5656,N_5844);
nor U6599 (N_6599,N_5470,N_5943);
or U6600 (N_6600,N_6429,N_6489);
nor U6601 (N_6601,N_6245,N_6559);
or U6602 (N_6602,N_6537,N_6438);
or U6603 (N_6603,N_6261,N_6169);
xor U6604 (N_6604,N_6433,N_6427);
and U6605 (N_6605,N_6138,N_6431);
or U6606 (N_6606,N_6593,N_6465);
nand U6607 (N_6607,N_6084,N_6592);
nand U6608 (N_6608,N_6225,N_6351);
xor U6609 (N_6609,N_6083,N_6510);
or U6610 (N_6610,N_6029,N_6228);
or U6611 (N_6611,N_6162,N_6403);
xor U6612 (N_6612,N_6184,N_6096);
nand U6613 (N_6613,N_6035,N_6092);
nor U6614 (N_6614,N_6240,N_6252);
or U6615 (N_6615,N_6482,N_6369);
nand U6616 (N_6616,N_6532,N_6250);
nand U6617 (N_6617,N_6397,N_6352);
nand U6618 (N_6618,N_6270,N_6405);
nor U6619 (N_6619,N_6416,N_6584);
nor U6620 (N_6620,N_6268,N_6513);
nor U6621 (N_6621,N_6195,N_6202);
xor U6622 (N_6622,N_6053,N_6082);
and U6623 (N_6623,N_6308,N_6086);
xnor U6624 (N_6624,N_6441,N_6103);
and U6625 (N_6625,N_6199,N_6340);
or U6626 (N_6626,N_6129,N_6469);
xnor U6627 (N_6627,N_6004,N_6186);
and U6628 (N_6628,N_6188,N_6260);
xor U6629 (N_6629,N_6020,N_6002);
nand U6630 (N_6630,N_6568,N_6280);
xnor U6631 (N_6631,N_6139,N_6163);
xor U6632 (N_6632,N_6366,N_6254);
or U6633 (N_6633,N_6374,N_6365);
or U6634 (N_6634,N_6316,N_6201);
or U6635 (N_6635,N_6483,N_6233);
xor U6636 (N_6636,N_6312,N_6271);
xnor U6637 (N_6637,N_6549,N_6432);
and U6638 (N_6638,N_6234,N_6590);
or U6639 (N_6639,N_6231,N_6024);
nor U6640 (N_6640,N_6208,N_6331);
nor U6641 (N_6641,N_6281,N_6575);
nand U6642 (N_6642,N_6309,N_6017);
and U6643 (N_6643,N_6028,N_6119);
and U6644 (N_6644,N_6045,N_6110);
nand U6645 (N_6645,N_6353,N_6302);
nand U6646 (N_6646,N_6522,N_6384);
or U6647 (N_6647,N_6544,N_6533);
xnor U6648 (N_6648,N_6241,N_6126);
nor U6649 (N_6649,N_6015,N_6168);
or U6650 (N_6650,N_6075,N_6344);
nand U6651 (N_6651,N_6026,N_6368);
or U6652 (N_6652,N_6335,N_6196);
and U6653 (N_6653,N_6493,N_6107);
or U6654 (N_6654,N_6450,N_6462);
or U6655 (N_6655,N_6220,N_6599);
nor U6656 (N_6656,N_6137,N_6013);
and U6657 (N_6657,N_6311,N_6371);
or U6658 (N_6658,N_6325,N_6550);
or U6659 (N_6659,N_6387,N_6097);
or U6660 (N_6660,N_6258,N_6226);
or U6661 (N_6661,N_6449,N_6222);
nand U6662 (N_6662,N_6211,N_6580);
xor U6663 (N_6663,N_6583,N_6424);
or U6664 (N_6664,N_6236,N_6059);
nor U6665 (N_6665,N_6117,N_6372);
nor U6666 (N_6666,N_6124,N_6329);
nand U6667 (N_6667,N_6389,N_6190);
or U6668 (N_6668,N_6347,N_6262);
and U6669 (N_6669,N_6338,N_6409);
or U6670 (N_6670,N_6414,N_6069);
and U6671 (N_6671,N_6295,N_6571);
or U6672 (N_6672,N_6033,N_6476);
nor U6673 (N_6673,N_6016,N_6244);
and U6674 (N_6674,N_6385,N_6269);
nand U6675 (N_6675,N_6527,N_6061);
or U6676 (N_6676,N_6051,N_6078);
nor U6677 (N_6677,N_6161,N_6079);
xor U6678 (N_6678,N_6223,N_6349);
or U6679 (N_6679,N_6044,N_6382);
nor U6680 (N_6680,N_6273,N_6412);
nor U6681 (N_6681,N_6535,N_6362);
or U6682 (N_6682,N_6067,N_6597);
or U6683 (N_6683,N_6573,N_6404);
xnor U6684 (N_6684,N_6589,N_6496);
nor U6685 (N_6685,N_6560,N_6282);
and U6686 (N_6686,N_6339,N_6379);
nand U6687 (N_6687,N_6102,N_6388);
and U6688 (N_6688,N_6324,N_6164);
or U6689 (N_6689,N_6422,N_6193);
and U6690 (N_6690,N_6361,N_6232);
xor U6691 (N_6691,N_6494,N_6531);
nand U6692 (N_6692,N_6525,N_6536);
nand U6693 (N_6693,N_6547,N_6507);
or U6694 (N_6694,N_6145,N_6401);
and U6695 (N_6695,N_6562,N_6337);
nand U6696 (N_6696,N_6290,N_6418);
or U6697 (N_6697,N_6395,N_6355);
nor U6698 (N_6698,N_6434,N_6506);
nor U6699 (N_6699,N_6293,N_6009);
xor U6700 (N_6700,N_6360,N_6521);
nor U6701 (N_6701,N_6594,N_6046);
xor U6702 (N_6702,N_6218,N_6392);
or U6703 (N_6703,N_6534,N_6134);
nor U6704 (N_6704,N_6070,N_6194);
nor U6705 (N_6705,N_6031,N_6332);
or U6706 (N_6706,N_6495,N_6185);
and U6707 (N_6707,N_6125,N_6093);
or U6708 (N_6708,N_6296,N_6378);
xnor U6709 (N_6709,N_6221,N_6505);
nor U6710 (N_6710,N_6133,N_6249);
nand U6711 (N_6711,N_6548,N_6094);
or U6712 (N_6712,N_6052,N_6068);
nor U6713 (N_6713,N_6181,N_6512);
xnor U6714 (N_6714,N_6251,N_6010);
and U6715 (N_6715,N_6198,N_6173);
or U6716 (N_6716,N_6071,N_6446);
and U6717 (N_6717,N_6229,N_6034);
or U6718 (N_6718,N_6205,N_6417);
or U6719 (N_6719,N_6049,N_6471);
xor U6720 (N_6720,N_6481,N_6146);
or U6721 (N_6721,N_6514,N_6095);
nor U6722 (N_6722,N_6415,N_6557);
and U6723 (N_6723,N_6087,N_6529);
nand U6724 (N_6724,N_6048,N_6171);
nand U6725 (N_6725,N_6130,N_6598);
and U6726 (N_6726,N_6043,N_6555);
nand U6727 (N_6727,N_6516,N_6041);
nand U6728 (N_6728,N_6354,N_6247);
nand U6729 (N_6729,N_6333,N_6459);
and U6730 (N_6730,N_6025,N_6213);
nor U6731 (N_6731,N_6289,N_6488);
nand U6732 (N_6732,N_6058,N_6530);
or U6733 (N_6733,N_6402,N_6539);
nor U6734 (N_6734,N_6330,N_6178);
or U6735 (N_6735,N_6042,N_6430);
nor U6736 (N_6736,N_6005,N_6237);
xnor U6737 (N_6737,N_6565,N_6285);
nor U6738 (N_6738,N_6108,N_6300);
nand U6739 (N_6739,N_6552,N_6538);
xor U6740 (N_6740,N_6179,N_6158);
xor U6741 (N_6741,N_6206,N_6267);
xor U6742 (N_6742,N_6478,N_6182);
nor U6743 (N_6743,N_6187,N_6177);
nor U6744 (N_6744,N_6497,N_6318);
nor U6745 (N_6745,N_6398,N_6588);
and U6746 (N_6746,N_6047,N_6230);
nor U6747 (N_6747,N_6528,N_6159);
and U6748 (N_6748,N_6176,N_6189);
and U6749 (N_6749,N_6081,N_6141);
xor U6750 (N_6750,N_6111,N_6508);
and U6751 (N_6751,N_6012,N_6406);
nor U6752 (N_6752,N_6200,N_6576);
nand U6753 (N_6753,N_6487,N_6131);
or U6754 (N_6754,N_6170,N_6470);
nand U6755 (N_6755,N_6419,N_6065);
or U6756 (N_6756,N_6595,N_6109);
nand U6757 (N_6757,N_6556,N_6467);
nor U6758 (N_6758,N_6348,N_6106);
xnor U6759 (N_6759,N_6008,N_6021);
and U6760 (N_6760,N_6104,N_6574);
nand U6761 (N_6761,N_6322,N_6456);
nor U6762 (N_6762,N_6003,N_6582);
or U6763 (N_6763,N_6057,N_6357);
and U6764 (N_6764,N_6453,N_6359);
nor U6765 (N_6765,N_6219,N_6390);
nor U6766 (N_6766,N_6570,N_6286);
nor U6767 (N_6767,N_6498,N_6135);
nor U6768 (N_6768,N_6410,N_6408);
nor U6769 (N_6769,N_6100,N_6545);
nor U6770 (N_6770,N_6001,N_6586);
nand U6771 (N_6771,N_6203,N_6259);
or U6772 (N_6772,N_6314,N_6321);
xor U6773 (N_6773,N_6501,N_6328);
nor U6774 (N_6774,N_6114,N_6278);
or U6775 (N_6775,N_6306,N_6153);
nor U6776 (N_6776,N_6553,N_6343);
and U6777 (N_6777,N_6143,N_6386);
nor U6778 (N_6778,N_6120,N_6436);
or U6779 (N_6779,N_6447,N_6172);
nor U6780 (N_6780,N_6500,N_6569);
or U6781 (N_6781,N_6437,N_6376);
nor U6782 (N_6782,N_6101,N_6455);
and U6783 (N_6783,N_6444,N_6591);
nor U6784 (N_6784,N_6085,N_6239);
xnor U6785 (N_6785,N_6342,N_6294);
or U6786 (N_6786,N_6090,N_6413);
or U6787 (N_6787,N_6121,N_6373);
nand U6788 (N_6788,N_6310,N_6377);
or U6789 (N_6789,N_6439,N_6297);
nand U6790 (N_6790,N_6350,N_6546);
nor U6791 (N_6791,N_6383,N_6154);
and U6792 (N_6792,N_6291,N_6396);
nor U6793 (N_6793,N_6393,N_6019);
nor U6794 (N_6794,N_6370,N_6473);
or U6795 (N_6795,N_6000,N_6428);
xnor U6796 (N_6796,N_6011,N_6105);
and U6797 (N_6797,N_6007,N_6400);
nand U6798 (N_6798,N_6326,N_6577);
or U6799 (N_6799,N_6144,N_6266);
or U6800 (N_6800,N_6509,N_6255);
or U6801 (N_6801,N_6578,N_6375);
xnor U6802 (N_6802,N_6056,N_6596);
nor U6803 (N_6803,N_6204,N_6216);
and U6804 (N_6804,N_6217,N_6440);
and U6805 (N_6805,N_6517,N_6080);
nand U6806 (N_6806,N_6472,N_6088);
and U6807 (N_6807,N_6442,N_6364);
and U6808 (N_6808,N_6452,N_6468);
xor U6809 (N_6809,N_6558,N_6463);
nor U6810 (N_6810,N_6175,N_6319);
xor U6811 (N_6811,N_6152,N_6060);
and U6812 (N_6812,N_6394,N_6054);
xor U6813 (N_6813,N_6420,N_6038);
or U6814 (N_6814,N_6275,N_6425);
nor U6815 (N_6815,N_6380,N_6464);
and U6816 (N_6816,N_6127,N_6209);
xnor U6817 (N_6817,N_6457,N_6563);
xnor U6818 (N_6818,N_6484,N_6064);
nand U6819 (N_6819,N_6128,N_6018);
nor U6820 (N_6820,N_6142,N_6567);
nor U6821 (N_6821,N_6027,N_6210);
and U6822 (N_6822,N_6477,N_6227);
and U6823 (N_6823,N_6098,N_6006);
nor U6824 (N_6824,N_6490,N_6299);
and U6825 (N_6825,N_6089,N_6475);
xor U6826 (N_6826,N_6055,N_6150);
and U6827 (N_6827,N_6147,N_6160);
or U6828 (N_6828,N_6148,N_6116);
nor U6829 (N_6829,N_6411,N_6180);
nand U6830 (N_6830,N_6304,N_6037);
xor U6831 (N_6831,N_6391,N_6479);
and U6832 (N_6832,N_6356,N_6358);
nand U6833 (N_6833,N_6246,N_6564);
nand U6834 (N_6834,N_6264,N_6077);
xor U6835 (N_6835,N_6305,N_6151);
nor U6836 (N_6836,N_6174,N_6367);
xor U6837 (N_6837,N_6572,N_6486);
nand U6838 (N_6838,N_6118,N_6073);
or U6839 (N_6839,N_6298,N_6561);
nor U6840 (N_6840,N_6140,N_6445);
and U6841 (N_6841,N_6036,N_6551);
or U6842 (N_6842,N_6242,N_6363);
nand U6843 (N_6843,N_6288,N_6072);
and U6844 (N_6844,N_6518,N_6224);
nand U6845 (N_6845,N_6274,N_6454);
xor U6846 (N_6846,N_6115,N_6136);
nand U6847 (N_6847,N_6435,N_6023);
nand U6848 (N_6848,N_6443,N_6014);
nand U6849 (N_6849,N_6543,N_6256);
nand U6850 (N_6850,N_6327,N_6587);
and U6851 (N_6851,N_6461,N_6341);
nor U6852 (N_6852,N_6334,N_6112);
or U6853 (N_6853,N_6458,N_6276);
nand U6854 (N_6854,N_6499,N_6207);
nor U6855 (N_6855,N_6292,N_6554);
nor U6856 (N_6856,N_6566,N_6579);
and U6857 (N_6857,N_6519,N_6149);
and U6858 (N_6858,N_6491,N_6272);
and U6859 (N_6859,N_6215,N_6155);
and U6860 (N_6860,N_6257,N_6301);
nand U6861 (N_6861,N_6032,N_6248);
nand U6862 (N_6862,N_6313,N_6283);
or U6863 (N_6863,N_6520,N_6399);
xnor U6864 (N_6864,N_6113,N_6277);
nor U6865 (N_6865,N_6346,N_6542);
nand U6866 (N_6866,N_6063,N_6345);
and U6867 (N_6867,N_6076,N_6503);
xor U6868 (N_6868,N_6263,N_6284);
nand U6869 (N_6869,N_6279,N_6451);
or U6870 (N_6870,N_6526,N_6485);
nand U6871 (N_6871,N_6156,N_6460);
or U6872 (N_6872,N_6191,N_6197);
or U6873 (N_6873,N_6466,N_6122);
xor U6874 (N_6874,N_6336,N_6091);
xnor U6875 (N_6875,N_6585,N_6524);
xor U6876 (N_6876,N_6166,N_6123);
xnor U6877 (N_6877,N_6030,N_6235);
nand U6878 (N_6878,N_6381,N_6541);
nand U6879 (N_6879,N_6307,N_6407);
and U6880 (N_6880,N_6480,N_6066);
xnor U6881 (N_6881,N_6540,N_6423);
nor U6882 (N_6882,N_6214,N_6515);
and U6883 (N_6883,N_6421,N_6426);
nand U6884 (N_6884,N_6050,N_6303);
xnor U6885 (N_6885,N_6074,N_6320);
xor U6886 (N_6886,N_6040,N_6317);
nor U6887 (N_6887,N_6287,N_6132);
or U6888 (N_6888,N_6167,N_6323);
xnor U6889 (N_6889,N_6474,N_6039);
xnor U6890 (N_6890,N_6212,N_6523);
or U6891 (N_6891,N_6502,N_6315);
nor U6892 (N_6892,N_6165,N_6504);
or U6893 (N_6893,N_6243,N_6265);
nor U6894 (N_6894,N_6099,N_6448);
and U6895 (N_6895,N_6492,N_6062);
nand U6896 (N_6896,N_6511,N_6238);
nand U6897 (N_6897,N_6183,N_6581);
and U6898 (N_6898,N_6253,N_6022);
and U6899 (N_6899,N_6192,N_6157);
and U6900 (N_6900,N_6453,N_6407);
xor U6901 (N_6901,N_6367,N_6189);
or U6902 (N_6902,N_6315,N_6501);
and U6903 (N_6903,N_6158,N_6366);
nand U6904 (N_6904,N_6538,N_6178);
or U6905 (N_6905,N_6037,N_6237);
or U6906 (N_6906,N_6153,N_6380);
and U6907 (N_6907,N_6148,N_6487);
nand U6908 (N_6908,N_6261,N_6090);
nor U6909 (N_6909,N_6319,N_6307);
and U6910 (N_6910,N_6248,N_6462);
nor U6911 (N_6911,N_6556,N_6549);
and U6912 (N_6912,N_6085,N_6354);
nor U6913 (N_6913,N_6460,N_6553);
nand U6914 (N_6914,N_6025,N_6100);
nor U6915 (N_6915,N_6568,N_6538);
nor U6916 (N_6916,N_6430,N_6534);
or U6917 (N_6917,N_6584,N_6427);
and U6918 (N_6918,N_6433,N_6539);
and U6919 (N_6919,N_6585,N_6500);
nand U6920 (N_6920,N_6190,N_6430);
nor U6921 (N_6921,N_6096,N_6058);
nor U6922 (N_6922,N_6127,N_6149);
xnor U6923 (N_6923,N_6211,N_6577);
or U6924 (N_6924,N_6284,N_6381);
nor U6925 (N_6925,N_6441,N_6427);
nor U6926 (N_6926,N_6362,N_6519);
and U6927 (N_6927,N_6530,N_6233);
nor U6928 (N_6928,N_6356,N_6539);
nor U6929 (N_6929,N_6192,N_6424);
and U6930 (N_6930,N_6029,N_6280);
nor U6931 (N_6931,N_6378,N_6417);
or U6932 (N_6932,N_6006,N_6085);
nand U6933 (N_6933,N_6296,N_6085);
nand U6934 (N_6934,N_6082,N_6158);
and U6935 (N_6935,N_6031,N_6491);
nand U6936 (N_6936,N_6097,N_6137);
nand U6937 (N_6937,N_6244,N_6015);
nand U6938 (N_6938,N_6477,N_6303);
nor U6939 (N_6939,N_6404,N_6513);
and U6940 (N_6940,N_6132,N_6566);
nor U6941 (N_6941,N_6519,N_6245);
xnor U6942 (N_6942,N_6189,N_6305);
and U6943 (N_6943,N_6354,N_6398);
and U6944 (N_6944,N_6331,N_6192);
nor U6945 (N_6945,N_6458,N_6123);
and U6946 (N_6946,N_6532,N_6176);
or U6947 (N_6947,N_6081,N_6280);
or U6948 (N_6948,N_6202,N_6218);
or U6949 (N_6949,N_6162,N_6137);
nand U6950 (N_6950,N_6410,N_6403);
nor U6951 (N_6951,N_6200,N_6109);
xnor U6952 (N_6952,N_6104,N_6559);
xor U6953 (N_6953,N_6384,N_6245);
and U6954 (N_6954,N_6297,N_6436);
nor U6955 (N_6955,N_6163,N_6440);
nand U6956 (N_6956,N_6385,N_6522);
and U6957 (N_6957,N_6199,N_6061);
xnor U6958 (N_6958,N_6181,N_6413);
or U6959 (N_6959,N_6040,N_6499);
and U6960 (N_6960,N_6509,N_6510);
and U6961 (N_6961,N_6068,N_6278);
xor U6962 (N_6962,N_6121,N_6074);
or U6963 (N_6963,N_6060,N_6449);
xnor U6964 (N_6964,N_6593,N_6510);
nand U6965 (N_6965,N_6125,N_6240);
or U6966 (N_6966,N_6165,N_6152);
nor U6967 (N_6967,N_6358,N_6586);
xor U6968 (N_6968,N_6311,N_6100);
nor U6969 (N_6969,N_6539,N_6446);
or U6970 (N_6970,N_6028,N_6205);
nor U6971 (N_6971,N_6560,N_6308);
nor U6972 (N_6972,N_6504,N_6203);
nand U6973 (N_6973,N_6564,N_6386);
nor U6974 (N_6974,N_6092,N_6568);
or U6975 (N_6975,N_6276,N_6274);
nor U6976 (N_6976,N_6128,N_6288);
nand U6977 (N_6977,N_6206,N_6534);
or U6978 (N_6978,N_6466,N_6212);
nand U6979 (N_6979,N_6268,N_6286);
xnor U6980 (N_6980,N_6130,N_6020);
nand U6981 (N_6981,N_6287,N_6265);
nand U6982 (N_6982,N_6505,N_6461);
or U6983 (N_6983,N_6226,N_6125);
nand U6984 (N_6984,N_6442,N_6288);
and U6985 (N_6985,N_6535,N_6163);
nand U6986 (N_6986,N_6303,N_6318);
nor U6987 (N_6987,N_6503,N_6154);
xnor U6988 (N_6988,N_6262,N_6204);
nand U6989 (N_6989,N_6157,N_6258);
nor U6990 (N_6990,N_6129,N_6520);
nand U6991 (N_6991,N_6259,N_6575);
xor U6992 (N_6992,N_6237,N_6254);
xor U6993 (N_6993,N_6168,N_6074);
nand U6994 (N_6994,N_6584,N_6424);
and U6995 (N_6995,N_6077,N_6518);
and U6996 (N_6996,N_6127,N_6527);
or U6997 (N_6997,N_6122,N_6337);
xnor U6998 (N_6998,N_6263,N_6040);
xor U6999 (N_6999,N_6249,N_6308);
nand U7000 (N_7000,N_6226,N_6475);
nor U7001 (N_7001,N_6527,N_6330);
xor U7002 (N_7002,N_6335,N_6360);
or U7003 (N_7003,N_6323,N_6512);
nand U7004 (N_7004,N_6559,N_6549);
nor U7005 (N_7005,N_6424,N_6570);
nor U7006 (N_7006,N_6343,N_6270);
nand U7007 (N_7007,N_6465,N_6447);
nand U7008 (N_7008,N_6358,N_6367);
nand U7009 (N_7009,N_6221,N_6119);
or U7010 (N_7010,N_6498,N_6549);
nor U7011 (N_7011,N_6126,N_6532);
or U7012 (N_7012,N_6305,N_6196);
xnor U7013 (N_7013,N_6073,N_6410);
and U7014 (N_7014,N_6113,N_6450);
nor U7015 (N_7015,N_6204,N_6190);
nand U7016 (N_7016,N_6319,N_6477);
xnor U7017 (N_7017,N_6237,N_6448);
xor U7018 (N_7018,N_6011,N_6131);
or U7019 (N_7019,N_6126,N_6502);
nand U7020 (N_7020,N_6094,N_6461);
nor U7021 (N_7021,N_6021,N_6200);
nand U7022 (N_7022,N_6558,N_6190);
or U7023 (N_7023,N_6566,N_6017);
xor U7024 (N_7024,N_6271,N_6129);
nand U7025 (N_7025,N_6393,N_6049);
and U7026 (N_7026,N_6194,N_6211);
nand U7027 (N_7027,N_6099,N_6033);
and U7028 (N_7028,N_6292,N_6594);
and U7029 (N_7029,N_6095,N_6394);
or U7030 (N_7030,N_6230,N_6076);
and U7031 (N_7031,N_6510,N_6505);
and U7032 (N_7032,N_6587,N_6280);
nor U7033 (N_7033,N_6120,N_6558);
nand U7034 (N_7034,N_6282,N_6082);
and U7035 (N_7035,N_6091,N_6144);
or U7036 (N_7036,N_6126,N_6597);
nor U7037 (N_7037,N_6511,N_6428);
and U7038 (N_7038,N_6284,N_6256);
or U7039 (N_7039,N_6038,N_6138);
nand U7040 (N_7040,N_6560,N_6144);
nor U7041 (N_7041,N_6494,N_6486);
nor U7042 (N_7042,N_6336,N_6274);
xnor U7043 (N_7043,N_6521,N_6599);
nor U7044 (N_7044,N_6368,N_6388);
xnor U7045 (N_7045,N_6389,N_6070);
nor U7046 (N_7046,N_6558,N_6195);
xor U7047 (N_7047,N_6153,N_6263);
nor U7048 (N_7048,N_6216,N_6403);
nand U7049 (N_7049,N_6334,N_6589);
and U7050 (N_7050,N_6072,N_6152);
xor U7051 (N_7051,N_6051,N_6279);
xor U7052 (N_7052,N_6218,N_6042);
or U7053 (N_7053,N_6344,N_6304);
nand U7054 (N_7054,N_6549,N_6061);
or U7055 (N_7055,N_6144,N_6227);
nor U7056 (N_7056,N_6116,N_6585);
and U7057 (N_7057,N_6438,N_6515);
xor U7058 (N_7058,N_6393,N_6573);
or U7059 (N_7059,N_6536,N_6139);
nand U7060 (N_7060,N_6069,N_6074);
nor U7061 (N_7061,N_6265,N_6430);
and U7062 (N_7062,N_6592,N_6087);
or U7063 (N_7063,N_6071,N_6391);
or U7064 (N_7064,N_6598,N_6417);
and U7065 (N_7065,N_6537,N_6596);
nor U7066 (N_7066,N_6498,N_6537);
xor U7067 (N_7067,N_6513,N_6241);
nor U7068 (N_7068,N_6269,N_6162);
and U7069 (N_7069,N_6036,N_6335);
and U7070 (N_7070,N_6242,N_6429);
xor U7071 (N_7071,N_6037,N_6223);
or U7072 (N_7072,N_6406,N_6263);
nor U7073 (N_7073,N_6267,N_6320);
nand U7074 (N_7074,N_6305,N_6348);
nand U7075 (N_7075,N_6064,N_6337);
nor U7076 (N_7076,N_6194,N_6230);
and U7077 (N_7077,N_6238,N_6548);
xnor U7078 (N_7078,N_6137,N_6223);
nor U7079 (N_7079,N_6336,N_6392);
nand U7080 (N_7080,N_6141,N_6364);
xor U7081 (N_7081,N_6558,N_6479);
or U7082 (N_7082,N_6553,N_6201);
and U7083 (N_7083,N_6347,N_6010);
or U7084 (N_7084,N_6338,N_6504);
nand U7085 (N_7085,N_6496,N_6108);
nand U7086 (N_7086,N_6591,N_6598);
nand U7087 (N_7087,N_6444,N_6549);
nor U7088 (N_7088,N_6164,N_6256);
and U7089 (N_7089,N_6143,N_6374);
or U7090 (N_7090,N_6189,N_6053);
nand U7091 (N_7091,N_6494,N_6584);
xnor U7092 (N_7092,N_6509,N_6130);
xor U7093 (N_7093,N_6174,N_6205);
nor U7094 (N_7094,N_6467,N_6071);
xor U7095 (N_7095,N_6509,N_6149);
and U7096 (N_7096,N_6097,N_6467);
and U7097 (N_7097,N_6341,N_6589);
or U7098 (N_7098,N_6188,N_6132);
nor U7099 (N_7099,N_6529,N_6441);
xor U7100 (N_7100,N_6277,N_6024);
or U7101 (N_7101,N_6336,N_6394);
nor U7102 (N_7102,N_6311,N_6152);
and U7103 (N_7103,N_6091,N_6329);
xor U7104 (N_7104,N_6333,N_6008);
and U7105 (N_7105,N_6171,N_6293);
or U7106 (N_7106,N_6426,N_6509);
and U7107 (N_7107,N_6115,N_6152);
xor U7108 (N_7108,N_6143,N_6257);
nor U7109 (N_7109,N_6498,N_6376);
and U7110 (N_7110,N_6329,N_6565);
xor U7111 (N_7111,N_6253,N_6345);
and U7112 (N_7112,N_6161,N_6001);
nor U7113 (N_7113,N_6009,N_6418);
nand U7114 (N_7114,N_6491,N_6500);
and U7115 (N_7115,N_6260,N_6489);
nor U7116 (N_7116,N_6136,N_6523);
nand U7117 (N_7117,N_6046,N_6071);
xnor U7118 (N_7118,N_6285,N_6268);
and U7119 (N_7119,N_6114,N_6281);
nand U7120 (N_7120,N_6558,N_6080);
xnor U7121 (N_7121,N_6211,N_6333);
nand U7122 (N_7122,N_6357,N_6123);
and U7123 (N_7123,N_6130,N_6461);
or U7124 (N_7124,N_6256,N_6561);
nor U7125 (N_7125,N_6381,N_6073);
nor U7126 (N_7126,N_6200,N_6568);
and U7127 (N_7127,N_6587,N_6582);
nor U7128 (N_7128,N_6390,N_6014);
nor U7129 (N_7129,N_6436,N_6469);
xnor U7130 (N_7130,N_6170,N_6145);
or U7131 (N_7131,N_6219,N_6577);
nand U7132 (N_7132,N_6338,N_6585);
nor U7133 (N_7133,N_6242,N_6346);
nor U7134 (N_7134,N_6519,N_6148);
xor U7135 (N_7135,N_6254,N_6115);
nor U7136 (N_7136,N_6333,N_6208);
or U7137 (N_7137,N_6544,N_6271);
nor U7138 (N_7138,N_6568,N_6102);
xnor U7139 (N_7139,N_6526,N_6200);
or U7140 (N_7140,N_6252,N_6426);
nor U7141 (N_7141,N_6158,N_6257);
nor U7142 (N_7142,N_6307,N_6097);
nand U7143 (N_7143,N_6057,N_6583);
nor U7144 (N_7144,N_6392,N_6143);
and U7145 (N_7145,N_6350,N_6524);
xor U7146 (N_7146,N_6321,N_6541);
or U7147 (N_7147,N_6096,N_6402);
xnor U7148 (N_7148,N_6295,N_6268);
nand U7149 (N_7149,N_6322,N_6486);
nor U7150 (N_7150,N_6587,N_6420);
nand U7151 (N_7151,N_6412,N_6219);
nor U7152 (N_7152,N_6459,N_6233);
nand U7153 (N_7153,N_6453,N_6165);
nor U7154 (N_7154,N_6266,N_6027);
or U7155 (N_7155,N_6050,N_6034);
nor U7156 (N_7156,N_6076,N_6197);
nand U7157 (N_7157,N_6366,N_6529);
nor U7158 (N_7158,N_6048,N_6561);
nor U7159 (N_7159,N_6444,N_6550);
nand U7160 (N_7160,N_6164,N_6592);
nor U7161 (N_7161,N_6288,N_6027);
nor U7162 (N_7162,N_6277,N_6282);
or U7163 (N_7163,N_6546,N_6311);
or U7164 (N_7164,N_6031,N_6557);
xor U7165 (N_7165,N_6353,N_6356);
and U7166 (N_7166,N_6181,N_6568);
and U7167 (N_7167,N_6400,N_6131);
and U7168 (N_7168,N_6015,N_6212);
and U7169 (N_7169,N_6571,N_6087);
nand U7170 (N_7170,N_6387,N_6240);
xnor U7171 (N_7171,N_6442,N_6131);
or U7172 (N_7172,N_6069,N_6536);
nand U7173 (N_7173,N_6472,N_6168);
nor U7174 (N_7174,N_6026,N_6014);
or U7175 (N_7175,N_6384,N_6535);
or U7176 (N_7176,N_6003,N_6498);
nand U7177 (N_7177,N_6004,N_6214);
nor U7178 (N_7178,N_6538,N_6196);
nor U7179 (N_7179,N_6427,N_6542);
and U7180 (N_7180,N_6526,N_6202);
nor U7181 (N_7181,N_6200,N_6597);
xnor U7182 (N_7182,N_6268,N_6024);
xor U7183 (N_7183,N_6213,N_6279);
xor U7184 (N_7184,N_6119,N_6251);
or U7185 (N_7185,N_6250,N_6387);
and U7186 (N_7186,N_6089,N_6308);
nand U7187 (N_7187,N_6531,N_6199);
and U7188 (N_7188,N_6316,N_6539);
and U7189 (N_7189,N_6108,N_6493);
and U7190 (N_7190,N_6500,N_6100);
and U7191 (N_7191,N_6520,N_6413);
and U7192 (N_7192,N_6506,N_6356);
or U7193 (N_7193,N_6568,N_6145);
or U7194 (N_7194,N_6470,N_6155);
and U7195 (N_7195,N_6497,N_6011);
nand U7196 (N_7196,N_6187,N_6267);
nor U7197 (N_7197,N_6184,N_6511);
nand U7198 (N_7198,N_6189,N_6571);
nand U7199 (N_7199,N_6445,N_6019);
nor U7200 (N_7200,N_7128,N_6696);
and U7201 (N_7201,N_6804,N_6733);
nor U7202 (N_7202,N_6826,N_6907);
nand U7203 (N_7203,N_7175,N_6673);
nand U7204 (N_7204,N_6742,N_6715);
or U7205 (N_7205,N_7090,N_7185);
xnor U7206 (N_7206,N_6991,N_6848);
or U7207 (N_7207,N_7089,N_6676);
xor U7208 (N_7208,N_6736,N_6921);
xnor U7209 (N_7209,N_6602,N_7037);
nor U7210 (N_7210,N_7174,N_6739);
or U7211 (N_7211,N_6900,N_7066);
nor U7212 (N_7212,N_6915,N_6649);
nand U7213 (N_7213,N_6709,N_7130);
nor U7214 (N_7214,N_7087,N_6849);
nand U7215 (N_7215,N_6722,N_6611);
and U7216 (N_7216,N_7168,N_6997);
xor U7217 (N_7217,N_6843,N_6613);
nor U7218 (N_7218,N_6976,N_6610);
and U7219 (N_7219,N_6953,N_7158);
xor U7220 (N_7220,N_6862,N_6979);
nand U7221 (N_7221,N_7118,N_7040);
or U7222 (N_7222,N_7138,N_6652);
xor U7223 (N_7223,N_6809,N_6732);
nand U7224 (N_7224,N_7141,N_6909);
nand U7225 (N_7225,N_7116,N_6894);
xnor U7226 (N_7226,N_7197,N_6872);
and U7227 (N_7227,N_6799,N_6700);
xnor U7228 (N_7228,N_6825,N_6917);
nand U7229 (N_7229,N_6889,N_7076);
nand U7230 (N_7230,N_6723,N_7190);
xnor U7231 (N_7231,N_7113,N_6945);
and U7232 (N_7232,N_7077,N_7104);
xnor U7233 (N_7233,N_6621,N_6833);
and U7234 (N_7234,N_7189,N_7021);
or U7235 (N_7235,N_7013,N_6614);
nor U7236 (N_7236,N_6725,N_7039);
nor U7237 (N_7237,N_6972,N_7196);
and U7238 (N_7238,N_7065,N_6817);
and U7239 (N_7239,N_6663,N_6746);
nand U7240 (N_7240,N_6697,N_7017);
and U7241 (N_7241,N_6781,N_6939);
or U7242 (N_7242,N_6683,N_7131);
or U7243 (N_7243,N_6957,N_6996);
and U7244 (N_7244,N_6648,N_6787);
or U7245 (N_7245,N_6630,N_6837);
xnor U7246 (N_7246,N_7114,N_7094);
or U7247 (N_7247,N_6650,N_6901);
nor U7248 (N_7248,N_6954,N_6759);
nand U7249 (N_7249,N_7069,N_6857);
nand U7250 (N_7250,N_6960,N_7064);
xor U7251 (N_7251,N_7030,N_6776);
nor U7252 (N_7252,N_7092,N_7059);
nand U7253 (N_7253,N_7019,N_6865);
nand U7254 (N_7254,N_6707,N_7156);
and U7255 (N_7255,N_6919,N_7062);
nor U7256 (N_7256,N_7047,N_6974);
xnor U7257 (N_7257,N_6752,N_6705);
nor U7258 (N_7258,N_6858,N_6765);
nand U7259 (N_7259,N_6779,N_7144);
nor U7260 (N_7260,N_6920,N_6823);
and U7261 (N_7261,N_6923,N_6680);
xnor U7262 (N_7262,N_6924,N_6713);
and U7263 (N_7263,N_7070,N_6688);
xor U7264 (N_7264,N_7097,N_6937);
xor U7265 (N_7265,N_6948,N_6698);
or U7266 (N_7266,N_7000,N_6982);
nand U7267 (N_7267,N_7135,N_6691);
xnor U7268 (N_7268,N_7120,N_7148);
nand U7269 (N_7269,N_6987,N_7176);
xnor U7270 (N_7270,N_6681,N_6757);
xor U7271 (N_7271,N_7126,N_6624);
xor U7272 (N_7272,N_6947,N_6975);
nand U7273 (N_7273,N_6803,N_6646);
and U7274 (N_7274,N_6988,N_7181);
or U7275 (N_7275,N_7053,N_6727);
xor U7276 (N_7276,N_6607,N_6835);
or U7277 (N_7277,N_6912,N_6701);
or U7278 (N_7278,N_6639,N_6962);
nand U7279 (N_7279,N_6854,N_6841);
nand U7280 (N_7280,N_7143,N_7057);
xnor U7281 (N_7281,N_6851,N_6895);
xnor U7282 (N_7282,N_7005,N_6969);
nor U7283 (N_7283,N_7006,N_7107);
nand U7284 (N_7284,N_6932,N_7162);
nor U7285 (N_7285,N_7108,N_7075);
nor U7286 (N_7286,N_7027,N_6632);
nor U7287 (N_7287,N_7056,N_6788);
nand U7288 (N_7288,N_7117,N_6684);
and U7289 (N_7289,N_6970,N_7193);
nand U7290 (N_7290,N_6887,N_7096);
nand U7291 (N_7291,N_6821,N_6605);
or U7292 (N_7292,N_6896,N_7038);
or U7293 (N_7293,N_6694,N_6968);
nor U7294 (N_7294,N_6643,N_6884);
and U7295 (N_7295,N_7187,N_6642);
and U7296 (N_7296,N_6675,N_7045);
nor U7297 (N_7297,N_6628,N_6866);
nor U7298 (N_7298,N_6963,N_7018);
and U7299 (N_7299,N_6772,N_6790);
nand U7300 (N_7300,N_6903,N_6877);
nand U7301 (N_7301,N_6710,N_7054);
and U7302 (N_7302,N_6905,N_7020);
and U7303 (N_7303,N_6638,N_7049);
nor U7304 (N_7304,N_6899,N_7186);
and U7305 (N_7305,N_6879,N_7159);
nand U7306 (N_7306,N_6868,N_7008);
xor U7307 (N_7307,N_7034,N_7171);
or U7308 (N_7308,N_6792,N_6936);
and U7309 (N_7309,N_7083,N_6916);
or U7310 (N_7310,N_6778,N_7127);
and U7311 (N_7311,N_6711,N_6795);
nor U7312 (N_7312,N_6925,N_6906);
nand U7313 (N_7313,N_7180,N_6859);
xnor U7314 (N_7314,N_6885,N_7173);
and U7315 (N_7315,N_7080,N_6964);
and U7316 (N_7316,N_6690,N_6748);
xor U7317 (N_7317,N_6961,N_6967);
or U7318 (N_7318,N_6745,N_6898);
nor U7319 (N_7319,N_6949,N_6706);
nor U7320 (N_7320,N_7015,N_6606);
nor U7321 (N_7321,N_6871,N_6782);
or U7322 (N_7322,N_7195,N_7016);
and U7323 (N_7323,N_7051,N_6780);
or U7324 (N_7324,N_7084,N_6761);
xor U7325 (N_7325,N_6717,N_7007);
nor U7326 (N_7326,N_6760,N_6737);
or U7327 (N_7327,N_7145,N_7155);
and U7328 (N_7328,N_7170,N_7035);
nand U7329 (N_7329,N_6758,N_6687);
xnor U7330 (N_7330,N_6796,N_6820);
xnor U7331 (N_7331,N_6721,N_6831);
nand U7332 (N_7332,N_7160,N_6855);
and U7333 (N_7333,N_7029,N_6811);
nor U7334 (N_7334,N_6813,N_7134);
or U7335 (N_7335,N_7178,N_6863);
nor U7336 (N_7336,N_6834,N_6656);
xnor U7337 (N_7337,N_6822,N_6658);
nor U7338 (N_7338,N_6750,N_6892);
xnor U7339 (N_7339,N_6842,N_7022);
and U7340 (N_7340,N_6929,N_6883);
or U7341 (N_7341,N_6989,N_7061);
and U7342 (N_7342,N_6785,N_6873);
and U7343 (N_7343,N_7154,N_6959);
xor U7344 (N_7344,N_7123,N_6838);
xnor U7345 (N_7345,N_6655,N_6720);
and U7346 (N_7346,N_7111,N_6635);
xor U7347 (N_7347,N_6743,N_6881);
or U7348 (N_7348,N_6754,N_6647);
or U7349 (N_7349,N_6994,N_6928);
xor U7350 (N_7350,N_6616,N_6651);
or U7351 (N_7351,N_6603,N_6850);
xor U7352 (N_7352,N_6631,N_6686);
nand U7353 (N_7353,N_6763,N_7101);
nor U7354 (N_7354,N_7102,N_7121);
nor U7355 (N_7355,N_6702,N_7085);
and U7356 (N_7356,N_6617,N_6818);
and U7357 (N_7357,N_6801,N_6791);
xor U7358 (N_7358,N_6993,N_7115);
nor U7359 (N_7359,N_6966,N_6677);
nor U7360 (N_7360,N_6882,N_6660);
and U7361 (N_7361,N_7009,N_7050);
nand U7362 (N_7362,N_6852,N_6674);
nand U7363 (N_7363,N_6672,N_6807);
or U7364 (N_7364,N_7112,N_6682);
nor U7365 (N_7365,N_6731,N_6756);
nor U7366 (N_7366,N_6926,N_6784);
and U7367 (N_7367,N_6845,N_6990);
nand U7368 (N_7368,N_6671,N_7157);
nor U7369 (N_7369,N_6880,N_6771);
nor U7370 (N_7370,N_6814,N_6914);
nor U7371 (N_7371,N_6922,N_6861);
xor U7372 (N_7372,N_7081,N_7055);
nand U7373 (N_7373,N_6714,N_7088);
xnor U7374 (N_7374,N_7191,N_7072);
nor U7375 (N_7375,N_7014,N_7161);
nand U7376 (N_7376,N_6666,N_7025);
nor U7377 (N_7377,N_6755,N_6918);
xnor U7378 (N_7378,N_6867,N_7188);
or U7379 (N_7379,N_6797,N_6653);
or U7380 (N_7380,N_6744,N_6664);
nand U7381 (N_7381,N_6999,N_7172);
nand U7382 (N_7382,N_6703,N_6995);
or U7383 (N_7383,N_6869,N_6890);
or U7384 (N_7384,N_6693,N_7177);
nand U7385 (N_7385,N_7119,N_7140);
and U7386 (N_7386,N_6913,N_6659);
or U7387 (N_7387,N_6747,N_6740);
or U7388 (N_7388,N_6983,N_6773);
and U7389 (N_7389,N_7106,N_6729);
nand U7390 (N_7390,N_7152,N_6728);
and U7391 (N_7391,N_6847,N_6853);
xnor U7392 (N_7392,N_7060,N_6775);
or U7393 (N_7393,N_6668,N_7098);
xnor U7394 (N_7394,N_6934,N_7151);
xor U7395 (N_7395,N_6965,N_6827);
or U7396 (N_7396,N_6808,N_7169);
nand U7397 (N_7397,N_6927,N_6670);
or U7398 (N_7398,N_7183,N_7010);
nor U7399 (N_7399,N_6824,N_6609);
and U7400 (N_7400,N_6645,N_6958);
or U7401 (N_7401,N_6840,N_7136);
xor U7402 (N_7402,N_6931,N_6860);
or U7403 (N_7403,N_6844,N_6793);
xor U7404 (N_7404,N_6839,N_6640);
nand U7405 (N_7405,N_6810,N_7194);
nor U7406 (N_7406,N_7184,N_6626);
or U7407 (N_7407,N_6973,N_6762);
xor U7408 (N_7408,N_6657,N_6886);
or U7409 (N_7409,N_7042,N_6902);
or U7410 (N_7410,N_7164,N_7093);
nor U7411 (N_7411,N_6662,N_6667);
or U7412 (N_7412,N_6956,N_6685);
xnor U7413 (N_7413,N_6941,N_7099);
nand U7414 (N_7414,N_7058,N_6665);
nand U7415 (N_7415,N_7048,N_7110);
nor U7416 (N_7416,N_6981,N_6769);
and U7417 (N_7417,N_7068,N_7012);
nand U7418 (N_7418,N_6897,N_6741);
nor U7419 (N_7419,N_6985,N_7036);
nor U7420 (N_7420,N_6766,N_7028);
xor U7421 (N_7421,N_6789,N_6716);
nand U7422 (N_7422,N_7067,N_6783);
xor U7423 (N_7423,N_7182,N_6695);
xnor U7424 (N_7424,N_6622,N_6812);
nand U7425 (N_7425,N_6946,N_6619);
or U7426 (N_7426,N_7124,N_7044);
and U7427 (N_7427,N_6802,N_6623);
nand U7428 (N_7428,N_6878,N_6777);
nor U7429 (N_7429,N_6891,N_7001);
nor U7430 (N_7430,N_6601,N_6836);
and U7431 (N_7431,N_7082,N_6940);
nand U7432 (N_7432,N_6641,N_7043);
nor U7433 (N_7433,N_6604,N_7004);
nand U7434 (N_7434,N_7199,N_6726);
and U7435 (N_7435,N_6724,N_7105);
xor U7436 (N_7436,N_7198,N_6832);
and U7437 (N_7437,N_7146,N_6980);
nand U7438 (N_7438,N_7002,N_6800);
nand U7439 (N_7439,N_7153,N_6943);
and U7440 (N_7440,N_6692,N_6816);
nand U7441 (N_7441,N_7024,N_7109);
or U7442 (N_7442,N_7103,N_6719);
nor U7443 (N_7443,N_7139,N_6735);
nor U7444 (N_7444,N_6942,N_6955);
nand U7445 (N_7445,N_6904,N_7031);
xnor U7446 (N_7446,N_6828,N_7142);
and U7447 (N_7447,N_6767,N_7086);
or U7448 (N_7448,N_7073,N_6753);
or U7449 (N_7449,N_6749,N_6911);
or U7450 (N_7450,N_6856,N_7122);
or U7451 (N_7451,N_7011,N_7179);
xor U7452 (N_7452,N_6950,N_6794);
nor U7453 (N_7453,N_7079,N_7078);
and U7454 (N_7454,N_7100,N_6633);
or U7455 (N_7455,N_6669,N_6634);
nor U7456 (N_7456,N_7147,N_6819);
or U7457 (N_7457,N_6608,N_6770);
nand U7458 (N_7458,N_6679,N_6846);
nor U7459 (N_7459,N_7063,N_7166);
xnor U7460 (N_7460,N_6875,N_6600);
nor U7461 (N_7461,N_6764,N_6893);
nand U7462 (N_7462,N_6689,N_7150);
xnor U7463 (N_7463,N_6951,N_6708);
or U7464 (N_7464,N_7026,N_6930);
nand U7465 (N_7465,N_6888,N_7052);
xnor U7466 (N_7466,N_6977,N_6933);
and U7467 (N_7467,N_6986,N_7046);
or U7468 (N_7468,N_7129,N_6615);
nand U7469 (N_7469,N_6798,N_6678);
or U7470 (N_7470,N_6618,N_6984);
nor U7471 (N_7471,N_6637,N_7165);
nor U7472 (N_7472,N_7137,N_7167);
nand U7473 (N_7473,N_6876,N_7041);
xnor U7474 (N_7474,N_7023,N_6738);
xnor U7475 (N_7475,N_7091,N_7074);
and U7476 (N_7476,N_6864,N_6730);
or U7477 (N_7477,N_7149,N_6636);
nor U7478 (N_7478,N_6629,N_6699);
and U7479 (N_7479,N_6998,N_7071);
nor U7480 (N_7480,N_7163,N_6971);
nand U7481 (N_7481,N_6830,N_6768);
and U7482 (N_7482,N_6815,N_6718);
and U7483 (N_7483,N_6908,N_6620);
nand U7484 (N_7484,N_6751,N_6661);
nand U7485 (N_7485,N_6712,N_6870);
or U7486 (N_7486,N_6786,N_6644);
and U7487 (N_7487,N_7003,N_6627);
or U7488 (N_7488,N_6704,N_7033);
or U7489 (N_7489,N_7125,N_6938);
or U7490 (N_7490,N_6952,N_7032);
xnor U7491 (N_7491,N_6805,N_6774);
or U7492 (N_7492,N_6829,N_6625);
xnor U7493 (N_7493,N_7192,N_6910);
and U7494 (N_7494,N_6654,N_6612);
nand U7495 (N_7495,N_6935,N_7133);
and U7496 (N_7496,N_7095,N_6978);
and U7497 (N_7497,N_6992,N_6806);
and U7498 (N_7498,N_7132,N_6944);
nand U7499 (N_7499,N_6734,N_6874);
xor U7500 (N_7500,N_6834,N_7186);
and U7501 (N_7501,N_6849,N_7016);
xnor U7502 (N_7502,N_6846,N_6946);
nand U7503 (N_7503,N_7163,N_6922);
and U7504 (N_7504,N_6942,N_7129);
nand U7505 (N_7505,N_7119,N_6838);
nand U7506 (N_7506,N_6860,N_6694);
nand U7507 (N_7507,N_6900,N_6699);
or U7508 (N_7508,N_6656,N_7197);
nor U7509 (N_7509,N_7020,N_6625);
xnor U7510 (N_7510,N_7144,N_7020);
and U7511 (N_7511,N_7051,N_6709);
and U7512 (N_7512,N_6791,N_6675);
xor U7513 (N_7513,N_6691,N_6606);
xor U7514 (N_7514,N_6814,N_7075);
or U7515 (N_7515,N_6857,N_6722);
or U7516 (N_7516,N_7051,N_6644);
xnor U7517 (N_7517,N_7120,N_6780);
nand U7518 (N_7518,N_6663,N_6712);
xor U7519 (N_7519,N_6874,N_6869);
nor U7520 (N_7520,N_6851,N_7009);
xnor U7521 (N_7521,N_6622,N_6819);
xnor U7522 (N_7522,N_7160,N_6889);
xnor U7523 (N_7523,N_7001,N_6965);
or U7524 (N_7524,N_7131,N_7081);
or U7525 (N_7525,N_6658,N_6627);
or U7526 (N_7526,N_6929,N_6697);
nor U7527 (N_7527,N_6984,N_7069);
and U7528 (N_7528,N_7127,N_6698);
nand U7529 (N_7529,N_6883,N_7018);
and U7530 (N_7530,N_6775,N_7109);
nand U7531 (N_7531,N_6805,N_7064);
or U7532 (N_7532,N_7140,N_7137);
nand U7533 (N_7533,N_6813,N_7049);
xor U7534 (N_7534,N_6804,N_7020);
nand U7535 (N_7535,N_6995,N_7033);
nand U7536 (N_7536,N_6659,N_7002);
xor U7537 (N_7537,N_6810,N_6910);
nor U7538 (N_7538,N_7192,N_6748);
xnor U7539 (N_7539,N_6888,N_6857);
and U7540 (N_7540,N_7036,N_6844);
xor U7541 (N_7541,N_6787,N_6927);
nand U7542 (N_7542,N_6617,N_7022);
nor U7543 (N_7543,N_6759,N_7181);
xor U7544 (N_7544,N_6979,N_7002);
nor U7545 (N_7545,N_6621,N_7163);
xnor U7546 (N_7546,N_7041,N_6655);
nor U7547 (N_7547,N_7142,N_6946);
or U7548 (N_7548,N_6990,N_6697);
xor U7549 (N_7549,N_6771,N_6994);
xnor U7550 (N_7550,N_7028,N_7034);
xor U7551 (N_7551,N_6902,N_6963);
nor U7552 (N_7552,N_6847,N_6663);
and U7553 (N_7553,N_6934,N_6996);
or U7554 (N_7554,N_7179,N_7067);
or U7555 (N_7555,N_6970,N_7170);
nand U7556 (N_7556,N_7106,N_6800);
nor U7557 (N_7557,N_6894,N_6890);
or U7558 (N_7558,N_7169,N_7026);
nor U7559 (N_7559,N_7087,N_7027);
nor U7560 (N_7560,N_6695,N_6846);
and U7561 (N_7561,N_6815,N_6888);
and U7562 (N_7562,N_7172,N_6748);
or U7563 (N_7563,N_6627,N_6892);
and U7564 (N_7564,N_6812,N_7170);
nand U7565 (N_7565,N_6779,N_6866);
and U7566 (N_7566,N_6918,N_6686);
nor U7567 (N_7567,N_7129,N_6660);
and U7568 (N_7568,N_7167,N_6705);
or U7569 (N_7569,N_6856,N_7089);
xor U7570 (N_7570,N_7140,N_7085);
and U7571 (N_7571,N_6857,N_7151);
and U7572 (N_7572,N_6981,N_6692);
nor U7573 (N_7573,N_6858,N_7010);
and U7574 (N_7574,N_7054,N_6734);
or U7575 (N_7575,N_7119,N_7051);
or U7576 (N_7576,N_6975,N_6635);
nor U7577 (N_7577,N_7005,N_6786);
xor U7578 (N_7578,N_7047,N_6796);
or U7579 (N_7579,N_6733,N_6961);
nand U7580 (N_7580,N_6914,N_6601);
nand U7581 (N_7581,N_6623,N_7154);
or U7582 (N_7582,N_6750,N_6981);
or U7583 (N_7583,N_6710,N_6678);
or U7584 (N_7584,N_6664,N_7181);
nand U7585 (N_7585,N_6979,N_7117);
xor U7586 (N_7586,N_6875,N_7113);
nand U7587 (N_7587,N_7075,N_6921);
nand U7588 (N_7588,N_6975,N_6830);
xor U7589 (N_7589,N_6988,N_7133);
xor U7590 (N_7590,N_7169,N_6715);
and U7591 (N_7591,N_6940,N_7152);
nor U7592 (N_7592,N_6706,N_6791);
xnor U7593 (N_7593,N_7048,N_6910);
nor U7594 (N_7594,N_6866,N_7148);
nor U7595 (N_7595,N_6703,N_7160);
nor U7596 (N_7596,N_7127,N_6770);
nand U7597 (N_7597,N_6843,N_6665);
xor U7598 (N_7598,N_6885,N_7089);
xor U7599 (N_7599,N_6833,N_6890);
or U7600 (N_7600,N_7161,N_6985);
xor U7601 (N_7601,N_6795,N_7039);
or U7602 (N_7602,N_7114,N_6831);
and U7603 (N_7603,N_6795,N_6810);
or U7604 (N_7604,N_6683,N_7126);
and U7605 (N_7605,N_6707,N_7011);
nor U7606 (N_7606,N_7175,N_7182);
nor U7607 (N_7607,N_6742,N_6854);
and U7608 (N_7608,N_7123,N_7002);
nor U7609 (N_7609,N_7027,N_6681);
nand U7610 (N_7610,N_7136,N_7027);
xnor U7611 (N_7611,N_6954,N_6911);
or U7612 (N_7612,N_7042,N_7004);
xnor U7613 (N_7613,N_6840,N_6939);
nor U7614 (N_7614,N_7110,N_6822);
xnor U7615 (N_7615,N_6859,N_6767);
xor U7616 (N_7616,N_6937,N_6620);
nand U7617 (N_7617,N_7165,N_7193);
or U7618 (N_7618,N_6732,N_6973);
and U7619 (N_7619,N_7110,N_6843);
or U7620 (N_7620,N_6688,N_7046);
nor U7621 (N_7621,N_7088,N_7118);
nor U7622 (N_7622,N_7004,N_7077);
xnor U7623 (N_7623,N_6806,N_6882);
and U7624 (N_7624,N_6838,N_7145);
nand U7625 (N_7625,N_6740,N_6956);
or U7626 (N_7626,N_6745,N_6653);
or U7627 (N_7627,N_6953,N_6985);
xnor U7628 (N_7628,N_6982,N_6794);
nand U7629 (N_7629,N_6633,N_6996);
nor U7630 (N_7630,N_7063,N_6724);
and U7631 (N_7631,N_6788,N_7101);
nand U7632 (N_7632,N_7093,N_6994);
xor U7633 (N_7633,N_6925,N_6851);
xnor U7634 (N_7634,N_7030,N_7004);
and U7635 (N_7635,N_6858,N_6662);
nand U7636 (N_7636,N_7172,N_7149);
and U7637 (N_7637,N_7060,N_6947);
nand U7638 (N_7638,N_7066,N_7055);
nor U7639 (N_7639,N_7165,N_7117);
or U7640 (N_7640,N_6680,N_6801);
nand U7641 (N_7641,N_7128,N_6800);
xnor U7642 (N_7642,N_6980,N_6693);
and U7643 (N_7643,N_7097,N_7174);
nor U7644 (N_7644,N_7058,N_6892);
or U7645 (N_7645,N_6711,N_6894);
nor U7646 (N_7646,N_6740,N_6687);
or U7647 (N_7647,N_6891,N_7098);
nor U7648 (N_7648,N_7077,N_6992);
and U7649 (N_7649,N_6755,N_6787);
xor U7650 (N_7650,N_6823,N_6602);
nand U7651 (N_7651,N_7141,N_6707);
nor U7652 (N_7652,N_6799,N_6632);
and U7653 (N_7653,N_6850,N_6896);
and U7654 (N_7654,N_6818,N_6658);
or U7655 (N_7655,N_6986,N_7087);
xnor U7656 (N_7656,N_6779,N_6723);
nand U7657 (N_7657,N_6734,N_6600);
or U7658 (N_7658,N_6950,N_7008);
or U7659 (N_7659,N_6837,N_7182);
and U7660 (N_7660,N_6853,N_6600);
nor U7661 (N_7661,N_6956,N_6736);
or U7662 (N_7662,N_6709,N_6657);
nor U7663 (N_7663,N_6724,N_7061);
or U7664 (N_7664,N_7143,N_6912);
nand U7665 (N_7665,N_6851,N_6858);
nor U7666 (N_7666,N_6712,N_6861);
and U7667 (N_7667,N_7184,N_6944);
or U7668 (N_7668,N_6990,N_6996);
or U7669 (N_7669,N_7121,N_6665);
nand U7670 (N_7670,N_6822,N_7174);
nand U7671 (N_7671,N_6610,N_7096);
xor U7672 (N_7672,N_6646,N_7159);
or U7673 (N_7673,N_7099,N_6929);
xnor U7674 (N_7674,N_6647,N_6651);
and U7675 (N_7675,N_6618,N_6734);
nor U7676 (N_7676,N_6699,N_6607);
nand U7677 (N_7677,N_6718,N_6944);
nor U7678 (N_7678,N_6641,N_6967);
nor U7679 (N_7679,N_6663,N_6898);
nor U7680 (N_7680,N_6879,N_6921);
or U7681 (N_7681,N_6662,N_6646);
nand U7682 (N_7682,N_6878,N_7043);
and U7683 (N_7683,N_7193,N_6912);
or U7684 (N_7684,N_6638,N_7129);
or U7685 (N_7685,N_6972,N_6726);
and U7686 (N_7686,N_6870,N_6921);
and U7687 (N_7687,N_6643,N_6850);
or U7688 (N_7688,N_6605,N_6600);
xnor U7689 (N_7689,N_6996,N_7058);
nand U7690 (N_7690,N_6742,N_7155);
nand U7691 (N_7691,N_6985,N_6713);
and U7692 (N_7692,N_6815,N_7154);
and U7693 (N_7693,N_7044,N_6774);
or U7694 (N_7694,N_6694,N_7132);
or U7695 (N_7695,N_7162,N_7190);
xor U7696 (N_7696,N_6664,N_6981);
xor U7697 (N_7697,N_7196,N_6999);
nand U7698 (N_7698,N_6651,N_6802);
or U7699 (N_7699,N_6618,N_7173);
nor U7700 (N_7700,N_6667,N_6672);
or U7701 (N_7701,N_6941,N_6924);
or U7702 (N_7702,N_6844,N_6801);
and U7703 (N_7703,N_6865,N_6830);
nor U7704 (N_7704,N_6797,N_6873);
nor U7705 (N_7705,N_7002,N_6693);
and U7706 (N_7706,N_6806,N_7001);
nand U7707 (N_7707,N_6897,N_6655);
xor U7708 (N_7708,N_6824,N_6761);
and U7709 (N_7709,N_6914,N_7034);
and U7710 (N_7710,N_7044,N_6673);
nand U7711 (N_7711,N_6931,N_6728);
nand U7712 (N_7712,N_7065,N_6729);
nor U7713 (N_7713,N_6799,N_7112);
or U7714 (N_7714,N_6820,N_6776);
and U7715 (N_7715,N_6991,N_7147);
and U7716 (N_7716,N_6768,N_6778);
or U7717 (N_7717,N_7110,N_7198);
nor U7718 (N_7718,N_6602,N_7165);
nor U7719 (N_7719,N_6618,N_6942);
and U7720 (N_7720,N_6928,N_6844);
nand U7721 (N_7721,N_6839,N_7132);
and U7722 (N_7722,N_7062,N_6826);
nor U7723 (N_7723,N_6675,N_7008);
and U7724 (N_7724,N_6970,N_6679);
xnor U7725 (N_7725,N_7062,N_6753);
and U7726 (N_7726,N_7176,N_6768);
or U7727 (N_7727,N_6775,N_7079);
nor U7728 (N_7728,N_6985,N_6942);
xnor U7729 (N_7729,N_6739,N_7193);
and U7730 (N_7730,N_6709,N_6825);
or U7731 (N_7731,N_7155,N_6962);
and U7732 (N_7732,N_6618,N_6601);
xor U7733 (N_7733,N_7025,N_6693);
nor U7734 (N_7734,N_6755,N_6852);
nor U7735 (N_7735,N_6879,N_6748);
nand U7736 (N_7736,N_6845,N_6787);
nand U7737 (N_7737,N_7081,N_6994);
and U7738 (N_7738,N_6768,N_6633);
nor U7739 (N_7739,N_6735,N_6832);
xor U7740 (N_7740,N_6706,N_6880);
nand U7741 (N_7741,N_7002,N_7077);
nor U7742 (N_7742,N_6602,N_7184);
and U7743 (N_7743,N_6786,N_6723);
nand U7744 (N_7744,N_6728,N_7060);
or U7745 (N_7745,N_6882,N_6941);
or U7746 (N_7746,N_7033,N_6805);
and U7747 (N_7747,N_6822,N_6789);
xor U7748 (N_7748,N_6838,N_6667);
and U7749 (N_7749,N_6799,N_7055);
xor U7750 (N_7750,N_6791,N_6664);
nor U7751 (N_7751,N_6688,N_7117);
and U7752 (N_7752,N_7052,N_7095);
xnor U7753 (N_7753,N_7017,N_7098);
or U7754 (N_7754,N_7157,N_6651);
nand U7755 (N_7755,N_6994,N_6999);
and U7756 (N_7756,N_6826,N_6686);
nor U7757 (N_7757,N_7168,N_6632);
and U7758 (N_7758,N_6907,N_6946);
and U7759 (N_7759,N_7163,N_6659);
nor U7760 (N_7760,N_7174,N_6965);
or U7761 (N_7761,N_7119,N_7037);
and U7762 (N_7762,N_6939,N_7050);
nor U7763 (N_7763,N_7124,N_7082);
nand U7764 (N_7764,N_6648,N_6760);
nor U7765 (N_7765,N_6834,N_6667);
nor U7766 (N_7766,N_6778,N_6688);
xor U7767 (N_7767,N_7131,N_6729);
or U7768 (N_7768,N_7020,N_6765);
or U7769 (N_7769,N_6828,N_7130);
and U7770 (N_7770,N_6959,N_6975);
nor U7771 (N_7771,N_6861,N_7126);
nor U7772 (N_7772,N_6914,N_6758);
xor U7773 (N_7773,N_7117,N_6844);
nor U7774 (N_7774,N_7092,N_6622);
xor U7775 (N_7775,N_7155,N_6941);
or U7776 (N_7776,N_7053,N_6903);
or U7777 (N_7777,N_6911,N_6766);
xnor U7778 (N_7778,N_7188,N_6713);
nand U7779 (N_7779,N_6771,N_6755);
nor U7780 (N_7780,N_6847,N_6987);
nand U7781 (N_7781,N_6650,N_7082);
nor U7782 (N_7782,N_6939,N_6886);
xnor U7783 (N_7783,N_6761,N_7130);
xor U7784 (N_7784,N_6993,N_7186);
and U7785 (N_7785,N_6716,N_6712);
nor U7786 (N_7786,N_6876,N_6652);
nor U7787 (N_7787,N_6628,N_7191);
nand U7788 (N_7788,N_7161,N_7041);
nand U7789 (N_7789,N_6658,N_7017);
and U7790 (N_7790,N_7143,N_6802);
and U7791 (N_7791,N_6853,N_7189);
and U7792 (N_7792,N_6917,N_6867);
or U7793 (N_7793,N_6967,N_6989);
nand U7794 (N_7794,N_6912,N_7055);
nor U7795 (N_7795,N_7112,N_7079);
or U7796 (N_7796,N_6928,N_6971);
nand U7797 (N_7797,N_7024,N_6862);
nand U7798 (N_7798,N_6657,N_6880);
and U7799 (N_7799,N_6703,N_6797);
nand U7800 (N_7800,N_7588,N_7309);
xor U7801 (N_7801,N_7536,N_7296);
and U7802 (N_7802,N_7324,N_7649);
xnor U7803 (N_7803,N_7485,N_7250);
nor U7804 (N_7804,N_7446,N_7427);
nand U7805 (N_7805,N_7303,N_7423);
xnor U7806 (N_7806,N_7429,N_7537);
xnor U7807 (N_7807,N_7314,N_7683);
nand U7808 (N_7808,N_7738,N_7664);
nor U7809 (N_7809,N_7601,N_7289);
or U7810 (N_7810,N_7501,N_7668);
or U7811 (N_7811,N_7511,N_7430);
nand U7812 (N_7812,N_7504,N_7294);
nand U7813 (N_7813,N_7237,N_7723);
nor U7814 (N_7814,N_7627,N_7736);
or U7815 (N_7815,N_7365,N_7582);
xnor U7816 (N_7816,N_7713,N_7704);
xnor U7817 (N_7817,N_7573,N_7224);
nand U7818 (N_7818,N_7474,N_7796);
or U7819 (N_7819,N_7482,N_7508);
nor U7820 (N_7820,N_7204,N_7781);
and U7821 (N_7821,N_7280,N_7637);
nor U7822 (N_7822,N_7503,N_7559);
and U7823 (N_7823,N_7753,N_7470);
xor U7824 (N_7824,N_7610,N_7413);
nand U7825 (N_7825,N_7475,N_7789);
xnor U7826 (N_7826,N_7759,N_7549);
nor U7827 (N_7827,N_7632,N_7766);
xor U7828 (N_7828,N_7465,N_7785);
and U7829 (N_7829,N_7732,N_7613);
nor U7830 (N_7830,N_7532,N_7251);
nor U7831 (N_7831,N_7200,N_7360);
or U7832 (N_7832,N_7406,N_7367);
xnor U7833 (N_7833,N_7247,N_7357);
nand U7834 (N_7834,N_7264,N_7374);
xnor U7835 (N_7835,N_7600,N_7513);
nand U7836 (N_7836,N_7748,N_7488);
and U7837 (N_7837,N_7287,N_7716);
or U7838 (N_7838,N_7540,N_7304);
or U7839 (N_7839,N_7414,N_7228);
or U7840 (N_7840,N_7246,N_7418);
and U7841 (N_7841,N_7244,N_7266);
and U7842 (N_7842,N_7350,N_7462);
or U7843 (N_7843,N_7592,N_7516);
or U7844 (N_7844,N_7343,N_7467);
and U7845 (N_7845,N_7609,N_7384);
and U7846 (N_7846,N_7369,N_7459);
nor U7847 (N_7847,N_7415,N_7453);
nor U7848 (N_7848,N_7454,N_7428);
and U7849 (N_7849,N_7373,N_7468);
nand U7850 (N_7850,N_7409,N_7650);
xor U7851 (N_7851,N_7354,N_7694);
nor U7852 (N_7852,N_7286,N_7284);
nand U7853 (N_7853,N_7220,N_7569);
nand U7854 (N_7854,N_7331,N_7295);
and U7855 (N_7855,N_7531,N_7703);
or U7856 (N_7856,N_7741,N_7253);
nor U7857 (N_7857,N_7273,N_7596);
or U7858 (N_7858,N_7265,N_7487);
and U7859 (N_7859,N_7407,N_7466);
nand U7860 (N_7860,N_7509,N_7277);
or U7861 (N_7861,N_7227,N_7307);
and U7862 (N_7862,N_7332,N_7538);
nor U7863 (N_7863,N_7481,N_7290);
nand U7864 (N_7864,N_7447,N_7440);
or U7865 (N_7865,N_7777,N_7589);
nand U7866 (N_7866,N_7546,N_7758);
and U7867 (N_7867,N_7576,N_7497);
or U7868 (N_7868,N_7525,N_7492);
and U7869 (N_7869,N_7708,N_7522);
xor U7870 (N_7870,N_7543,N_7791);
nor U7871 (N_7871,N_7461,N_7658);
nand U7872 (N_7872,N_7729,N_7599);
nand U7873 (N_7873,N_7633,N_7463);
nand U7874 (N_7874,N_7398,N_7222);
and U7875 (N_7875,N_7603,N_7387);
nor U7876 (N_7876,N_7257,N_7225);
or U7877 (N_7877,N_7550,N_7292);
and U7878 (N_7878,N_7368,N_7375);
nand U7879 (N_7879,N_7326,N_7740);
xnor U7880 (N_7880,N_7328,N_7624);
and U7881 (N_7881,N_7334,N_7660);
and U7882 (N_7882,N_7379,N_7707);
and U7883 (N_7883,N_7730,N_7595);
nor U7884 (N_7884,N_7233,N_7389);
or U7885 (N_7885,N_7519,N_7383);
nor U7886 (N_7886,N_7241,N_7578);
nor U7887 (N_7887,N_7604,N_7590);
and U7888 (N_7888,N_7666,N_7226);
nor U7889 (N_7889,N_7419,N_7636);
and U7890 (N_7890,N_7445,N_7763);
nand U7891 (N_7891,N_7333,N_7345);
xor U7892 (N_7892,N_7359,N_7269);
nor U7893 (N_7893,N_7211,N_7702);
xnor U7894 (N_7894,N_7319,N_7230);
or U7895 (N_7895,N_7451,N_7715);
or U7896 (N_7896,N_7362,N_7417);
and U7897 (N_7897,N_7378,N_7219);
nor U7898 (N_7898,N_7518,N_7322);
and U7899 (N_7899,N_7556,N_7719);
nand U7900 (N_7900,N_7439,N_7656);
or U7901 (N_7901,N_7252,N_7450);
and U7902 (N_7902,N_7486,N_7260);
nor U7903 (N_7903,N_7533,N_7281);
and U7904 (N_7904,N_7697,N_7744);
or U7905 (N_7905,N_7506,N_7421);
nor U7906 (N_7906,N_7396,N_7458);
xnor U7907 (N_7907,N_7361,N_7714);
nor U7908 (N_7908,N_7757,N_7259);
and U7909 (N_7909,N_7321,N_7655);
nand U7910 (N_7910,N_7436,N_7499);
or U7911 (N_7911,N_7695,N_7755);
xor U7912 (N_7912,N_7388,N_7641);
nand U7913 (N_7913,N_7443,N_7611);
nand U7914 (N_7914,N_7502,N_7215);
xor U7915 (N_7915,N_7438,N_7344);
or U7916 (N_7916,N_7206,N_7783);
nor U7917 (N_7917,N_7762,N_7572);
or U7918 (N_7918,N_7258,N_7737);
nand U7919 (N_7919,N_7448,N_7529);
or U7920 (N_7920,N_7523,N_7583);
or U7921 (N_7921,N_7764,N_7300);
and U7922 (N_7922,N_7679,N_7238);
nor U7923 (N_7923,N_7431,N_7602);
nand U7924 (N_7924,N_7787,N_7709);
and U7925 (N_7925,N_7248,N_7640);
nor U7926 (N_7926,N_7263,N_7297);
nand U7927 (N_7927,N_7394,N_7285);
nor U7928 (N_7928,N_7437,N_7793);
and U7929 (N_7929,N_7495,N_7434);
and U7930 (N_7930,N_7623,N_7372);
nor U7931 (N_7931,N_7771,N_7647);
or U7932 (N_7932,N_7484,N_7710);
nand U7933 (N_7933,N_7393,N_7693);
or U7934 (N_7934,N_7491,N_7216);
nand U7935 (N_7935,N_7784,N_7691);
xor U7936 (N_7936,N_7268,N_7671);
or U7937 (N_7937,N_7336,N_7735);
nor U7938 (N_7938,N_7689,N_7402);
or U7939 (N_7939,N_7201,N_7567);
nand U7940 (N_7940,N_7790,N_7352);
nor U7941 (N_7941,N_7249,N_7725);
xor U7942 (N_7942,N_7382,N_7311);
nor U7943 (N_7943,N_7420,N_7711);
nor U7944 (N_7944,N_7563,N_7597);
xor U7945 (N_7945,N_7229,N_7335);
nand U7946 (N_7946,N_7218,N_7323);
xor U7947 (N_7947,N_7630,N_7355);
nand U7948 (N_7948,N_7464,N_7455);
or U7949 (N_7949,N_7566,N_7262);
xnor U7950 (N_7950,N_7705,N_7593);
nor U7951 (N_7951,N_7698,N_7392);
nand U7952 (N_7952,N_7712,N_7654);
and U7953 (N_7953,N_7242,N_7621);
nand U7954 (N_7954,N_7399,N_7270);
xnor U7955 (N_7955,N_7254,N_7646);
nand U7956 (N_7956,N_7217,N_7773);
and U7957 (N_7957,N_7617,N_7521);
xor U7958 (N_7958,N_7207,N_7320);
nand U7959 (N_7959,N_7585,N_7391);
nor U7960 (N_7960,N_7457,N_7288);
xor U7961 (N_7961,N_7528,N_7329);
nor U7962 (N_7962,N_7645,N_7386);
nand U7963 (N_7963,N_7203,N_7282);
nor U7964 (N_7964,N_7395,N_7298);
and U7965 (N_7965,N_7515,N_7648);
xnor U7966 (N_7966,N_7653,N_7792);
and U7967 (N_7967,N_7306,N_7291);
nand U7968 (N_7968,N_7261,N_7432);
nor U7969 (N_7969,N_7720,N_7469);
or U7970 (N_7970,N_7728,N_7605);
and U7971 (N_7971,N_7435,N_7626);
xor U7972 (N_7972,N_7239,N_7363);
xor U7973 (N_7973,N_7767,N_7701);
nand U7974 (N_7974,N_7622,N_7586);
xor U7975 (N_7975,N_7587,N_7577);
and U7976 (N_7976,N_7562,N_7786);
or U7977 (N_7977,N_7747,N_7634);
nand U7978 (N_7978,N_7795,N_7490);
and U7979 (N_7979,N_7782,N_7726);
and U7980 (N_7980,N_7456,N_7279);
nor U7981 (N_7981,N_7510,N_7615);
nand U7982 (N_7982,N_7699,N_7635);
xnor U7983 (N_7983,N_7442,N_7558);
and U7984 (N_7984,N_7424,N_7769);
nor U7985 (N_7985,N_7524,N_7441);
or U7986 (N_7986,N_7780,N_7272);
xnor U7987 (N_7987,N_7255,N_7325);
and U7988 (N_7988,N_7798,N_7670);
nor U7989 (N_7989,N_7553,N_7642);
nand U7990 (N_7990,N_7338,N_7305);
or U7991 (N_7991,N_7330,N_7686);
nor U7992 (N_7992,N_7643,N_7631);
nor U7993 (N_7993,N_7337,N_7313);
xor U7994 (N_7994,N_7520,N_7659);
or U7995 (N_7995,N_7571,N_7243);
xor U7996 (N_7996,N_7507,N_7449);
xor U7997 (N_7997,N_7400,N_7534);
nand U7998 (N_7998,N_7731,N_7493);
xor U7999 (N_7999,N_7276,N_7267);
or U8000 (N_8000,N_7797,N_7381);
xor U8001 (N_8001,N_7675,N_7620);
nand U8002 (N_8002,N_7223,N_7756);
xnor U8003 (N_8003,N_7568,N_7256);
and U8004 (N_8004,N_7665,N_7214);
xnor U8005 (N_8005,N_7721,N_7681);
nand U8006 (N_8006,N_7754,N_7416);
nand U8007 (N_8007,N_7358,N_7209);
xnor U8008 (N_8008,N_7278,N_7411);
and U8009 (N_8009,N_7564,N_7772);
nor U8010 (N_8010,N_7351,N_7561);
and U8011 (N_8011,N_7208,N_7682);
nor U8012 (N_8012,N_7212,N_7760);
and U8013 (N_8013,N_7271,N_7380);
nand U8014 (N_8014,N_7213,N_7677);
nand U8015 (N_8015,N_7557,N_7751);
xnor U8016 (N_8016,N_7678,N_7356);
or U8017 (N_8017,N_7745,N_7742);
nand U8018 (N_8018,N_7240,N_7340);
nor U8019 (N_8019,N_7341,N_7310);
nor U8020 (N_8020,N_7530,N_7743);
nor U8021 (N_8021,N_7299,N_7514);
or U8022 (N_8022,N_7652,N_7539);
or U8023 (N_8023,N_7348,N_7552);
or U8024 (N_8024,N_7598,N_7746);
and U8025 (N_8025,N_7669,N_7687);
xor U8026 (N_8026,N_7794,N_7498);
xnor U8027 (N_8027,N_7489,N_7618);
nor U8028 (N_8028,N_7739,N_7776);
or U8029 (N_8029,N_7405,N_7496);
xor U8030 (N_8030,N_7734,N_7535);
nor U8031 (N_8031,N_7706,N_7606);
nand U8032 (N_8032,N_7366,N_7770);
xor U8033 (N_8033,N_7555,N_7512);
and U8034 (N_8034,N_7690,N_7376);
xnor U8035 (N_8035,N_7473,N_7302);
or U8036 (N_8036,N_7283,N_7479);
nand U8037 (N_8037,N_7570,N_7476);
nand U8038 (N_8038,N_7625,N_7733);
nor U8039 (N_8039,N_7575,N_7616);
xor U8040 (N_8040,N_7692,N_7444);
and U8041 (N_8041,N_7327,N_7688);
and U8042 (N_8042,N_7560,N_7527);
xor U8043 (N_8043,N_7661,N_7581);
xnor U8044 (N_8044,N_7346,N_7408);
xnor U8045 (N_8045,N_7231,N_7312);
and U8046 (N_8046,N_7517,N_7412);
nor U8047 (N_8047,N_7422,N_7545);
nor U8048 (N_8048,N_7478,N_7628);
nand U8049 (N_8049,N_7724,N_7500);
xor U8050 (N_8050,N_7644,N_7404);
xnor U8051 (N_8051,N_7477,N_7774);
nand U8052 (N_8052,N_7696,N_7353);
and U8053 (N_8053,N_7579,N_7775);
or U8054 (N_8054,N_7717,N_7544);
and U8055 (N_8055,N_7236,N_7480);
xor U8056 (N_8056,N_7722,N_7371);
and U8057 (N_8057,N_7401,N_7390);
nand U8058 (N_8058,N_7672,N_7403);
nand U8059 (N_8059,N_7370,N_7274);
or U8060 (N_8060,N_7397,N_7317);
nand U8061 (N_8061,N_7779,N_7565);
and U8062 (N_8062,N_7685,N_7799);
nand U8063 (N_8063,N_7483,N_7608);
or U8064 (N_8064,N_7718,N_7275);
or U8065 (N_8065,N_7651,N_7316);
xnor U8066 (N_8066,N_7580,N_7761);
nor U8067 (N_8067,N_7639,N_7542);
and U8068 (N_8068,N_7594,N_7778);
or U8069 (N_8069,N_7667,N_7221);
nand U8070 (N_8070,N_7426,N_7349);
or U8071 (N_8071,N_7526,N_7554);
or U8072 (N_8072,N_7638,N_7548);
or U8073 (N_8073,N_7364,N_7210);
nand U8074 (N_8074,N_7750,N_7584);
nand U8075 (N_8075,N_7505,N_7662);
xor U8076 (N_8076,N_7342,N_7749);
nor U8077 (N_8077,N_7318,N_7612);
nand U8078 (N_8078,N_7205,N_7574);
xnor U8079 (N_8079,N_7607,N_7727);
and U8080 (N_8080,N_7680,N_7541);
xor U8081 (N_8081,N_7410,N_7619);
and U8082 (N_8082,N_7657,N_7460);
nor U8083 (N_8083,N_7377,N_7765);
nand U8084 (N_8084,N_7308,N_7551);
or U8085 (N_8085,N_7293,N_7202);
nor U8086 (N_8086,N_7614,N_7425);
or U8087 (N_8087,N_7494,N_7673);
nand U8088 (N_8088,N_7235,N_7768);
nor U8089 (N_8089,N_7674,N_7547);
nand U8090 (N_8090,N_7591,N_7347);
nand U8091 (N_8091,N_7433,N_7232);
nor U8092 (N_8092,N_7752,N_7234);
nand U8093 (N_8093,N_7684,N_7472);
nor U8094 (N_8094,N_7452,N_7339);
nor U8095 (N_8095,N_7385,N_7471);
or U8096 (N_8096,N_7663,N_7301);
nor U8097 (N_8097,N_7315,N_7629);
or U8098 (N_8098,N_7245,N_7788);
and U8099 (N_8099,N_7676,N_7700);
nor U8100 (N_8100,N_7240,N_7514);
nand U8101 (N_8101,N_7654,N_7633);
xor U8102 (N_8102,N_7629,N_7765);
nand U8103 (N_8103,N_7551,N_7381);
nand U8104 (N_8104,N_7563,N_7352);
xnor U8105 (N_8105,N_7577,N_7245);
and U8106 (N_8106,N_7462,N_7347);
nor U8107 (N_8107,N_7600,N_7368);
or U8108 (N_8108,N_7705,N_7316);
nor U8109 (N_8109,N_7670,N_7461);
or U8110 (N_8110,N_7398,N_7357);
and U8111 (N_8111,N_7795,N_7344);
xnor U8112 (N_8112,N_7555,N_7711);
xor U8113 (N_8113,N_7502,N_7724);
and U8114 (N_8114,N_7713,N_7419);
and U8115 (N_8115,N_7513,N_7289);
and U8116 (N_8116,N_7715,N_7444);
xor U8117 (N_8117,N_7694,N_7616);
nand U8118 (N_8118,N_7794,N_7237);
or U8119 (N_8119,N_7606,N_7473);
and U8120 (N_8120,N_7453,N_7737);
or U8121 (N_8121,N_7614,N_7672);
or U8122 (N_8122,N_7752,N_7308);
and U8123 (N_8123,N_7442,N_7223);
or U8124 (N_8124,N_7551,N_7774);
and U8125 (N_8125,N_7256,N_7724);
or U8126 (N_8126,N_7637,N_7527);
and U8127 (N_8127,N_7310,N_7209);
xnor U8128 (N_8128,N_7542,N_7225);
nand U8129 (N_8129,N_7360,N_7229);
nor U8130 (N_8130,N_7781,N_7755);
or U8131 (N_8131,N_7688,N_7443);
nand U8132 (N_8132,N_7227,N_7282);
nor U8133 (N_8133,N_7639,N_7368);
nand U8134 (N_8134,N_7305,N_7757);
xor U8135 (N_8135,N_7682,N_7620);
xnor U8136 (N_8136,N_7336,N_7408);
nor U8137 (N_8137,N_7590,N_7612);
nor U8138 (N_8138,N_7308,N_7768);
nor U8139 (N_8139,N_7394,N_7406);
xor U8140 (N_8140,N_7677,N_7690);
or U8141 (N_8141,N_7606,N_7370);
or U8142 (N_8142,N_7556,N_7682);
nand U8143 (N_8143,N_7213,N_7476);
xnor U8144 (N_8144,N_7616,N_7394);
xor U8145 (N_8145,N_7629,N_7381);
nand U8146 (N_8146,N_7683,N_7424);
or U8147 (N_8147,N_7744,N_7428);
or U8148 (N_8148,N_7518,N_7341);
or U8149 (N_8149,N_7387,N_7641);
or U8150 (N_8150,N_7479,N_7489);
xor U8151 (N_8151,N_7481,N_7316);
nor U8152 (N_8152,N_7434,N_7626);
or U8153 (N_8153,N_7493,N_7677);
nand U8154 (N_8154,N_7598,N_7465);
nand U8155 (N_8155,N_7395,N_7508);
nor U8156 (N_8156,N_7309,N_7299);
nand U8157 (N_8157,N_7440,N_7265);
or U8158 (N_8158,N_7343,N_7644);
and U8159 (N_8159,N_7553,N_7714);
xnor U8160 (N_8160,N_7390,N_7635);
and U8161 (N_8161,N_7371,N_7439);
nand U8162 (N_8162,N_7636,N_7406);
nand U8163 (N_8163,N_7560,N_7473);
nand U8164 (N_8164,N_7345,N_7405);
and U8165 (N_8165,N_7336,N_7396);
nand U8166 (N_8166,N_7339,N_7628);
xor U8167 (N_8167,N_7773,N_7635);
or U8168 (N_8168,N_7617,N_7541);
nand U8169 (N_8169,N_7360,N_7233);
or U8170 (N_8170,N_7463,N_7462);
nor U8171 (N_8171,N_7465,N_7327);
xor U8172 (N_8172,N_7760,N_7751);
or U8173 (N_8173,N_7724,N_7636);
nand U8174 (N_8174,N_7773,N_7769);
or U8175 (N_8175,N_7295,N_7612);
xnor U8176 (N_8176,N_7711,N_7442);
xor U8177 (N_8177,N_7689,N_7547);
and U8178 (N_8178,N_7498,N_7364);
nand U8179 (N_8179,N_7738,N_7587);
nand U8180 (N_8180,N_7756,N_7632);
xnor U8181 (N_8181,N_7373,N_7658);
or U8182 (N_8182,N_7760,N_7763);
nand U8183 (N_8183,N_7461,N_7615);
nand U8184 (N_8184,N_7674,N_7341);
nor U8185 (N_8185,N_7691,N_7455);
nor U8186 (N_8186,N_7687,N_7461);
xor U8187 (N_8187,N_7608,N_7568);
and U8188 (N_8188,N_7531,N_7363);
and U8189 (N_8189,N_7411,N_7343);
or U8190 (N_8190,N_7628,N_7225);
nand U8191 (N_8191,N_7408,N_7599);
nand U8192 (N_8192,N_7364,N_7303);
nand U8193 (N_8193,N_7214,N_7414);
and U8194 (N_8194,N_7420,N_7501);
or U8195 (N_8195,N_7292,N_7558);
and U8196 (N_8196,N_7337,N_7322);
or U8197 (N_8197,N_7223,N_7214);
or U8198 (N_8198,N_7361,N_7633);
xor U8199 (N_8199,N_7649,N_7228);
and U8200 (N_8200,N_7260,N_7449);
or U8201 (N_8201,N_7349,N_7653);
or U8202 (N_8202,N_7528,N_7642);
or U8203 (N_8203,N_7477,N_7255);
nand U8204 (N_8204,N_7442,N_7687);
xnor U8205 (N_8205,N_7774,N_7673);
nand U8206 (N_8206,N_7610,N_7297);
nand U8207 (N_8207,N_7440,N_7378);
nand U8208 (N_8208,N_7519,N_7686);
nor U8209 (N_8209,N_7383,N_7397);
and U8210 (N_8210,N_7270,N_7391);
nor U8211 (N_8211,N_7751,N_7419);
and U8212 (N_8212,N_7302,N_7592);
or U8213 (N_8213,N_7308,N_7663);
xnor U8214 (N_8214,N_7384,N_7587);
or U8215 (N_8215,N_7428,N_7556);
xnor U8216 (N_8216,N_7718,N_7427);
xor U8217 (N_8217,N_7523,N_7529);
and U8218 (N_8218,N_7244,N_7454);
or U8219 (N_8219,N_7764,N_7682);
or U8220 (N_8220,N_7798,N_7661);
nand U8221 (N_8221,N_7474,N_7424);
xnor U8222 (N_8222,N_7282,N_7285);
or U8223 (N_8223,N_7492,N_7712);
nand U8224 (N_8224,N_7275,N_7787);
nor U8225 (N_8225,N_7673,N_7472);
and U8226 (N_8226,N_7469,N_7230);
and U8227 (N_8227,N_7457,N_7430);
nand U8228 (N_8228,N_7625,N_7587);
or U8229 (N_8229,N_7692,N_7437);
xnor U8230 (N_8230,N_7232,N_7458);
nor U8231 (N_8231,N_7733,N_7699);
nand U8232 (N_8232,N_7312,N_7576);
and U8233 (N_8233,N_7759,N_7724);
nor U8234 (N_8234,N_7708,N_7302);
or U8235 (N_8235,N_7480,N_7354);
nor U8236 (N_8236,N_7294,N_7422);
nor U8237 (N_8237,N_7420,N_7334);
and U8238 (N_8238,N_7252,N_7793);
xor U8239 (N_8239,N_7343,N_7746);
or U8240 (N_8240,N_7488,N_7246);
or U8241 (N_8241,N_7667,N_7381);
or U8242 (N_8242,N_7513,N_7392);
or U8243 (N_8243,N_7721,N_7383);
and U8244 (N_8244,N_7211,N_7726);
xnor U8245 (N_8245,N_7699,N_7545);
nand U8246 (N_8246,N_7359,N_7503);
nor U8247 (N_8247,N_7357,N_7682);
or U8248 (N_8248,N_7321,N_7383);
nand U8249 (N_8249,N_7757,N_7608);
nor U8250 (N_8250,N_7509,N_7368);
or U8251 (N_8251,N_7743,N_7742);
nor U8252 (N_8252,N_7771,N_7663);
nand U8253 (N_8253,N_7640,N_7302);
xor U8254 (N_8254,N_7586,N_7688);
xnor U8255 (N_8255,N_7486,N_7718);
nand U8256 (N_8256,N_7374,N_7700);
xor U8257 (N_8257,N_7389,N_7723);
nor U8258 (N_8258,N_7248,N_7794);
nor U8259 (N_8259,N_7309,N_7469);
xor U8260 (N_8260,N_7673,N_7762);
nand U8261 (N_8261,N_7776,N_7674);
xor U8262 (N_8262,N_7551,N_7670);
nand U8263 (N_8263,N_7663,N_7450);
nor U8264 (N_8264,N_7202,N_7442);
xnor U8265 (N_8265,N_7361,N_7432);
nor U8266 (N_8266,N_7612,N_7790);
xor U8267 (N_8267,N_7296,N_7398);
xnor U8268 (N_8268,N_7221,N_7681);
and U8269 (N_8269,N_7463,N_7344);
or U8270 (N_8270,N_7797,N_7507);
and U8271 (N_8271,N_7541,N_7351);
nor U8272 (N_8272,N_7660,N_7261);
or U8273 (N_8273,N_7549,N_7782);
or U8274 (N_8274,N_7656,N_7673);
or U8275 (N_8275,N_7247,N_7404);
nand U8276 (N_8276,N_7390,N_7347);
xnor U8277 (N_8277,N_7596,N_7710);
and U8278 (N_8278,N_7652,N_7340);
nand U8279 (N_8279,N_7530,N_7362);
and U8280 (N_8280,N_7404,N_7563);
nor U8281 (N_8281,N_7271,N_7536);
xor U8282 (N_8282,N_7257,N_7318);
nor U8283 (N_8283,N_7276,N_7585);
and U8284 (N_8284,N_7779,N_7480);
nor U8285 (N_8285,N_7694,N_7319);
and U8286 (N_8286,N_7276,N_7625);
xnor U8287 (N_8287,N_7506,N_7445);
nand U8288 (N_8288,N_7297,N_7515);
nor U8289 (N_8289,N_7583,N_7729);
xnor U8290 (N_8290,N_7408,N_7785);
or U8291 (N_8291,N_7510,N_7769);
nor U8292 (N_8292,N_7278,N_7545);
nor U8293 (N_8293,N_7451,N_7477);
or U8294 (N_8294,N_7282,N_7547);
or U8295 (N_8295,N_7688,N_7478);
nor U8296 (N_8296,N_7408,N_7355);
xor U8297 (N_8297,N_7718,N_7215);
or U8298 (N_8298,N_7276,N_7330);
and U8299 (N_8299,N_7299,N_7735);
nand U8300 (N_8300,N_7272,N_7624);
and U8301 (N_8301,N_7369,N_7477);
or U8302 (N_8302,N_7698,N_7325);
nand U8303 (N_8303,N_7255,N_7515);
nand U8304 (N_8304,N_7476,N_7544);
xnor U8305 (N_8305,N_7435,N_7372);
nand U8306 (N_8306,N_7323,N_7486);
and U8307 (N_8307,N_7416,N_7409);
nand U8308 (N_8308,N_7456,N_7298);
nor U8309 (N_8309,N_7287,N_7518);
and U8310 (N_8310,N_7616,N_7511);
nand U8311 (N_8311,N_7766,N_7202);
or U8312 (N_8312,N_7796,N_7321);
or U8313 (N_8313,N_7334,N_7763);
or U8314 (N_8314,N_7531,N_7394);
nand U8315 (N_8315,N_7636,N_7671);
nand U8316 (N_8316,N_7470,N_7206);
or U8317 (N_8317,N_7368,N_7359);
nor U8318 (N_8318,N_7302,N_7283);
and U8319 (N_8319,N_7496,N_7695);
and U8320 (N_8320,N_7457,N_7772);
and U8321 (N_8321,N_7342,N_7688);
nor U8322 (N_8322,N_7243,N_7404);
nand U8323 (N_8323,N_7452,N_7354);
xor U8324 (N_8324,N_7569,N_7644);
xor U8325 (N_8325,N_7484,N_7581);
nand U8326 (N_8326,N_7298,N_7447);
and U8327 (N_8327,N_7288,N_7639);
nand U8328 (N_8328,N_7230,N_7417);
or U8329 (N_8329,N_7655,N_7251);
and U8330 (N_8330,N_7588,N_7744);
nand U8331 (N_8331,N_7281,N_7502);
nor U8332 (N_8332,N_7798,N_7338);
xnor U8333 (N_8333,N_7404,N_7478);
and U8334 (N_8334,N_7760,N_7226);
or U8335 (N_8335,N_7616,N_7421);
nand U8336 (N_8336,N_7205,N_7392);
nand U8337 (N_8337,N_7773,N_7752);
nand U8338 (N_8338,N_7574,N_7788);
and U8339 (N_8339,N_7302,N_7246);
nor U8340 (N_8340,N_7360,N_7629);
and U8341 (N_8341,N_7658,N_7762);
or U8342 (N_8342,N_7567,N_7677);
nand U8343 (N_8343,N_7725,N_7700);
nand U8344 (N_8344,N_7725,N_7615);
xnor U8345 (N_8345,N_7529,N_7750);
nor U8346 (N_8346,N_7693,N_7250);
or U8347 (N_8347,N_7734,N_7268);
xor U8348 (N_8348,N_7723,N_7448);
nand U8349 (N_8349,N_7308,N_7566);
nand U8350 (N_8350,N_7406,N_7792);
nor U8351 (N_8351,N_7505,N_7792);
and U8352 (N_8352,N_7675,N_7311);
nand U8353 (N_8353,N_7325,N_7799);
and U8354 (N_8354,N_7243,N_7654);
or U8355 (N_8355,N_7374,N_7736);
or U8356 (N_8356,N_7566,N_7551);
nand U8357 (N_8357,N_7429,N_7796);
xor U8358 (N_8358,N_7355,N_7792);
or U8359 (N_8359,N_7603,N_7669);
xnor U8360 (N_8360,N_7663,N_7550);
or U8361 (N_8361,N_7681,N_7206);
nor U8362 (N_8362,N_7319,N_7316);
nor U8363 (N_8363,N_7251,N_7535);
xnor U8364 (N_8364,N_7369,N_7640);
xor U8365 (N_8365,N_7386,N_7584);
nand U8366 (N_8366,N_7653,N_7752);
and U8367 (N_8367,N_7448,N_7202);
nand U8368 (N_8368,N_7590,N_7469);
nand U8369 (N_8369,N_7628,N_7263);
xnor U8370 (N_8370,N_7227,N_7691);
xor U8371 (N_8371,N_7666,N_7325);
nor U8372 (N_8372,N_7728,N_7508);
nand U8373 (N_8373,N_7604,N_7224);
xor U8374 (N_8374,N_7724,N_7320);
nand U8375 (N_8375,N_7725,N_7709);
or U8376 (N_8376,N_7598,N_7403);
nor U8377 (N_8377,N_7456,N_7653);
nor U8378 (N_8378,N_7234,N_7756);
nand U8379 (N_8379,N_7498,N_7442);
xnor U8380 (N_8380,N_7743,N_7486);
and U8381 (N_8381,N_7793,N_7420);
and U8382 (N_8382,N_7377,N_7742);
xnor U8383 (N_8383,N_7757,N_7614);
nand U8384 (N_8384,N_7700,N_7203);
and U8385 (N_8385,N_7399,N_7721);
nor U8386 (N_8386,N_7576,N_7522);
nand U8387 (N_8387,N_7730,N_7717);
xnor U8388 (N_8388,N_7505,N_7285);
or U8389 (N_8389,N_7664,N_7263);
and U8390 (N_8390,N_7527,N_7434);
nor U8391 (N_8391,N_7354,N_7498);
and U8392 (N_8392,N_7445,N_7496);
xor U8393 (N_8393,N_7316,N_7586);
xor U8394 (N_8394,N_7618,N_7528);
nand U8395 (N_8395,N_7731,N_7582);
or U8396 (N_8396,N_7676,N_7249);
xor U8397 (N_8397,N_7296,N_7508);
nor U8398 (N_8398,N_7655,N_7413);
and U8399 (N_8399,N_7669,N_7648);
and U8400 (N_8400,N_8379,N_8019);
and U8401 (N_8401,N_8268,N_8100);
nor U8402 (N_8402,N_7860,N_7874);
or U8403 (N_8403,N_8378,N_7817);
xor U8404 (N_8404,N_8334,N_7812);
xnor U8405 (N_8405,N_8170,N_8184);
nand U8406 (N_8406,N_8140,N_7925);
xnor U8407 (N_8407,N_8207,N_8258);
or U8408 (N_8408,N_7900,N_8182);
or U8409 (N_8409,N_7983,N_8136);
and U8410 (N_8410,N_7819,N_8283);
or U8411 (N_8411,N_8018,N_8021);
xor U8412 (N_8412,N_7954,N_8394);
nor U8413 (N_8413,N_7978,N_7835);
and U8414 (N_8414,N_7813,N_8034);
nor U8415 (N_8415,N_8373,N_8359);
and U8416 (N_8416,N_8356,N_8104);
nand U8417 (N_8417,N_8004,N_8309);
nand U8418 (N_8418,N_7974,N_7850);
nor U8419 (N_8419,N_7946,N_8386);
nand U8420 (N_8420,N_8069,N_8347);
or U8421 (N_8421,N_8224,N_8270);
and U8422 (N_8422,N_8254,N_8231);
and U8423 (N_8423,N_8219,N_8193);
and U8424 (N_8424,N_7879,N_7887);
or U8425 (N_8425,N_8094,N_7808);
and U8426 (N_8426,N_8246,N_7958);
or U8427 (N_8427,N_8340,N_8062);
xor U8428 (N_8428,N_8250,N_8287);
or U8429 (N_8429,N_8297,N_7915);
xor U8430 (N_8430,N_7890,N_8306);
or U8431 (N_8431,N_8134,N_8054);
nor U8432 (N_8432,N_8383,N_8061);
or U8433 (N_8433,N_8279,N_7964);
xnor U8434 (N_8434,N_8229,N_7837);
nand U8435 (N_8435,N_8262,N_7873);
or U8436 (N_8436,N_8282,N_7800);
xor U8437 (N_8437,N_8113,N_7935);
or U8438 (N_8438,N_8336,N_8260);
xnor U8439 (N_8439,N_8166,N_8328);
nand U8440 (N_8440,N_8044,N_8068);
or U8441 (N_8441,N_7941,N_7895);
nor U8442 (N_8442,N_8233,N_8161);
nand U8443 (N_8443,N_8098,N_7910);
nand U8444 (N_8444,N_8345,N_7933);
xnor U8445 (N_8445,N_8278,N_8001);
and U8446 (N_8446,N_8037,N_7904);
nand U8447 (N_8447,N_8101,N_8056);
nand U8448 (N_8448,N_8105,N_8285);
and U8449 (N_8449,N_7940,N_8311);
or U8450 (N_8450,N_7975,N_7864);
nor U8451 (N_8451,N_7862,N_8075);
or U8452 (N_8452,N_8147,N_7923);
nand U8453 (N_8453,N_8040,N_7820);
nor U8454 (N_8454,N_7806,N_8000);
or U8455 (N_8455,N_8025,N_7909);
and U8456 (N_8456,N_8389,N_8276);
xor U8457 (N_8457,N_7942,N_8200);
nor U8458 (N_8458,N_8058,N_7981);
xnor U8459 (N_8459,N_8244,N_8368);
nand U8460 (N_8460,N_7831,N_8307);
and U8461 (N_8461,N_8365,N_8130);
or U8462 (N_8462,N_8103,N_7830);
and U8463 (N_8463,N_8333,N_8125);
xor U8464 (N_8464,N_8057,N_7986);
nand U8465 (N_8465,N_8141,N_8255);
nand U8466 (N_8466,N_8392,N_8181);
and U8467 (N_8467,N_8060,N_7937);
nand U8468 (N_8468,N_8220,N_7977);
and U8469 (N_8469,N_7970,N_7950);
and U8470 (N_8470,N_8256,N_8177);
nand U8471 (N_8471,N_7955,N_8135);
xor U8472 (N_8472,N_8288,N_7918);
nand U8473 (N_8473,N_7944,N_8324);
nand U8474 (N_8474,N_8301,N_8312);
and U8475 (N_8475,N_8002,N_7982);
and U8476 (N_8476,N_7863,N_7809);
nor U8477 (N_8477,N_8222,N_8208);
or U8478 (N_8478,N_8053,N_7969);
nand U8479 (N_8479,N_8242,N_7908);
nand U8480 (N_8480,N_8149,N_7939);
nor U8481 (N_8481,N_7857,N_7811);
or U8482 (N_8482,N_7885,N_7818);
xor U8483 (N_8483,N_8096,N_7931);
and U8484 (N_8484,N_8015,N_8316);
or U8485 (N_8485,N_8310,N_7948);
or U8486 (N_8486,N_7855,N_8248);
and U8487 (N_8487,N_8206,N_7852);
nor U8488 (N_8488,N_8073,N_8252);
and U8489 (N_8489,N_8067,N_8313);
nand U8490 (N_8490,N_7883,N_8127);
nor U8491 (N_8491,N_7841,N_8302);
or U8492 (N_8492,N_7972,N_7927);
or U8493 (N_8493,N_8171,N_8344);
nand U8494 (N_8494,N_8159,N_8032);
and U8495 (N_8495,N_8366,N_8048);
nor U8496 (N_8496,N_8036,N_7859);
and U8497 (N_8497,N_8013,N_8045);
nor U8498 (N_8498,N_7889,N_8038);
and U8499 (N_8499,N_8305,N_7947);
nor U8500 (N_8500,N_7930,N_8196);
or U8501 (N_8501,N_8150,N_8115);
nor U8502 (N_8502,N_8146,N_8362);
nand U8503 (N_8503,N_8008,N_7878);
nand U8504 (N_8504,N_7851,N_8023);
and U8505 (N_8505,N_7840,N_8369);
and U8506 (N_8506,N_7884,N_7987);
xor U8507 (N_8507,N_7913,N_8275);
nand U8508 (N_8508,N_7976,N_8107);
xor U8509 (N_8509,N_7966,N_7814);
or U8510 (N_8510,N_8128,N_8237);
or U8511 (N_8511,N_8372,N_8160);
nor U8512 (N_8512,N_8076,N_8190);
nand U8513 (N_8513,N_8286,N_8041);
xor U8514 (N_8514,N_8064,N_8042);
or U8515 (N_8515,N_8066,N_8388);
or U8516 (N_8516,N_8086,N_8024);
or U8517 (N_8517,N_7869,N_7844);
xnor U8518 (N_8518,N_8380,N_8257);
xor U8519 (N_8519,N_8031,N_8121);
xor U8520 (N_8520,N_8245,N_8367);
xnor U8521 (N_8521,N_8162,N_8352);
nor U8522 (N_8522,N_8236,N_7880);
or U8523 (N_8523,N_8026,N_8174);
nor U8524 (N_8524,N_8143,N_7833);
nand U8525 (N_8525,N_7843,N_8089);
xor U8526 (N_8526,N_7868,N_7861);
and U8527 (N_8527,N_8361,N_8211);
and U8528 (N_8528,N_7824,N_7829);
or U8529 (N_8529,N_7839,N_8203);
xnor U8530 (N_8530,N_8065,N_8168);
xor U8531 (N_8531,N_7832,N_8133);
nor U8532 (N_8532,N_8271,N_8299);
nand U8533 (N_8533,N_8129,N_7845);
or U8534 (N_8534,N_7898,N_7876);
and U8535 (N_8535,N_8215,N_8191);
or U8536 (N_8536,N_8303,N_8051);
nand U8537 (N_8537,N_8261,N_7993);
nand U8538 (N_8538,N_8346,N_8259);
and U8539 (N_8539,N_8077,N_8320);
nor U8540 (N_8540,N_7865,N_8218);
xor U8541 (N_8541,N_7836,N_8173);
and U8542 (N_8542,N_7929,N_8209);
xnor U8543 (N_8543,N_7922,N_8012);
nand U8544 (N_8544,N_7849,N_8329);
or U8545 (N_8545,N_7881,N_7902);
nor U8546 (N_8546,N_8050,N_7996);
nand U8547 (N_8547,N_8396,N_8337);
and U8548 (N_8548,N_7985,N_8033);
and U8549 (N_8549,N_8108,N_7921);
nand U8550 (N_8550,N_8187,N_7801);
and U8551 (N_8551,N_8079,N_7853);
and U8552 (N_8552,N_8382,N_8376);
nor U8553 (N_8553,N_7979,N_7866);
nand U8554 (N_8554,N_7980,N_7877);
xnor U8555 (N_8555,N_8201,N_7894);
and U8556 (N_8556,N_7846,N_8102);
xnor U8557 (N_8557,N_8081,N_7847);
or U8558 (N_8558,N_7823,N_8323);
xnor U8559 (N_8559,N_8354,N_8213);
xnor U8560 (N_8560,N_8020,N_8280);
and U8561 (N_8561,N_7997,N_7956);
and U8562 (N_8562,N_8348,N_7821);
and U8563 (N_8563,N_8385,N_8006);
nor U8564 (N_8564,N_7805,N_8298);
nor U8565 (N_8565,N_8109,N_8003);
xnor U8566 (N_8566,N_8330,N_7990);
nor U8567 (N_8567,N_8185,N_8249);
or U8568 (N_8568,N_8186,N_8029);
nand U8569 (N_8569,N_8082,N_8189);
or U8570 (N_8570,N_7803,N_8084);
or U8571 (N_8571,N_8335,N_8093);
nand U8572 (N_8572,N_7834,N_7991);
xor U8573 (N_8573,N_8167,N_7870);
and U8574 (N_8574,N_7952,N_7911);
nand U8575 (N_8575,N_8142,N_8074);
nand U8576 (N_8576,N_8381,N_7953);
nand U8577 (N_8577,N_7875,N_8106);
nor U8578 (N_8578,N_7858,N_8355);
xor U8579 (N_8579,N_8092,N_8087);
xor U8580 (N_8580,N_8078,N_8214);
nand U8581 (N_8581,N_8202,N_8172);
nand U8582 (N_8582,N_7962,N_8325);
nor U8583 (N_8583,N_7945,N_8374);
and U8584 (N_8584,N_8228,N_8223);
and U8585 (N_8585,N_8027,N_8014);
and U8586 (N_8586,N_8156,N_7871);
and U8587 (N_8587,N_8070,N_8055);
xnor U8588 (N_8588,N_8308,N_8225);
xnor U8589 (N_8589,N_7916,N_8090);
and U8590 (N_8590,N_7912,N_8217);
xnor U8591 (N_8591,N_8377,N_8295);
nand U8592 (N_8592,N_8253,N_7905);
or U8593 (N_8593,N_8212,N_7968);
or U8594 (N_8594,N_7867,N_8204);
and U8595 (N_8595,N_8272,N_7914);
nand U8596 (N_8596,N_7822,N_8251);
or U8597 (N_8597,N_8110,N_7917);
xor U8598 (N_8598,N_8326,N_8291);
nor U8599 (N_8599,N_8183,N_7936);
and U8600 (N_8600,N_8349,N_7932);
xnor U8601 (N_8601,N_7838,N_8071);
xor U8602 (N_8602,N_8357,N_8210);
xor U8603 (N_8603,N_8005,N_7967);
nand U8604 (N_8604,N_8363,N_8175);
xnor U8605 (N_8605,N_7816,N_8290);
or U8606 (N_8606,N_8148,N_7999);
nor U8607 (N_8607,N_8318,N_7882);
and U8608 (N_8608,N_7920,N_8179);
or U8609 (N_8609,N_7827,N_7828);
nand U8610 (N_8610,N_8132,N_8169);
nand U8611 (N_8611,N_8391,N_8384);
and U8612 (N_8612,N_8011,N_8226);
xor U8613 (N_8613,N_8284,N_8116);
or U8614 (N_8614,N_7896,N_7998);
xnor U8615 (N_8615,N_8327,N_8205);
nor U8616 (N_8616,N_7973,N_7892);
nor U8617 (N_8617,N_8341,N_8331);
nor U8618 (N_8618,N_8046,N_7951);
nor U8619 (N_8619,N_8319,N_8126);
or U8620 (N_8620,N_7928,N_8197);
xnor U8621 (N_8621,N_7810,N_7994);
nor U8622 (N_8622,N_8176,N_8266);
xnor U8623 (N_8623,N_8007,N_7888);
nor U8624 (N_8624,N_8360,N_8216);
nand U8625 (N_8625,N_8072,N_8370);
nor U8626 (N_8626,N_7893,N_8095);
xnor U8627 (N_8627,N_8338,N_8111);
nor U8628 (N_8628,N_8234,N_8274);
nand U8629 (N_8629,N_8243,N_8158);
nor U8630 (N_8630,N_8099,N_7891);
xnor U8631 (N_8631,N_8152,N_8139);
nand U8632 (N_8632,N_8157,N_8294);
and U8633 (N_8633,N_8387,N_8395);
xor U8634 (N_8634,N_8343,N_8049);
nand U8635 (N_8635,N_8332,N_8030);
nand U8636 (N_8636,N_8188,N_8293);
nor U8637 (N_8637,N_8364,N_7949);
nand U8638 (N_8638,N_8350,N_8397);
and U8639 (N_8639,N_8144,N_8080);
or U8640 (N_8640,N_8269,N_8180);
and U8641 (N_8641,N_8300,N_8137);
or U8642 (N_8642,N_8398,N_8235);
xor U8643 (N_8643,N_8317,N_8393);
or U8644 (N_8644,N_8238,N_8114);
nand U8645 (N_8645,N_8194,N_8043);
nor U8646 (N_8646,N_8239,N_8165);
xnor U8647 (N_8647,N_8085,N_8151);
nor U8648 (N_8648,N_8017,N_8353);
and U8649 (N_8649,N_7984,N_7804);
or U8650 (N_8650,N_8117,N_8277);
or U8651 (N_8651,N_7934,N_7897);
and U8652 (N_8652,N_7802,N_7995);
nor U8653 (N_8653,N_7807,N_8163);
or U8654 (N_8654,N_8342,N_8227);
nand U8655 (N_8655,N_8314,N_8088);
nor U8656 (N_8656,N_7842,N_8123);
xor U8657 (N_8657,N_7943,N_8059);
xnor U8658 (N_8658,N_8390,N_8118);
or U8659 (N_8659,N_8289,N_8292);
xor U8660 (N_8660,N_8122,N_8119);
nand U8661 (N_8661,N_8371,N_8375);
nand U8662 (N_8662,N_8153,N_8247);
xor U8663 (N_8663,N_8010,N_8178);
nand U8664 (N_8664,N_8131,N_7965);
nor U8665 (N_8665,N_8039,N_8164);
nand U8666 (N_8666,N_7959,N_7957);
nand U8667 (N_8667,N_8240,N_7989);
nor U8668 (N_8668,N_8022,N_7988);
xnor U8669 (N_8669,N_8241,N_7938);
nor U8670 (N_8670,N_7960,N_8304);
xor U8671 (N_8671,N_8047,N_8221);
and U8672 (N_8672,N_8009,N_8321);
and U8673 (N_8673,N_8155,N_7963);
nand U8674 (N_8674,N_8124,N_8358);
nor U8675 (N_8675,N_8145,N_7924);
or U8676 (N_8676,N_7886,N_7961);
nor U8677 (N_8677,N_7854,N_8112);
or U8678 (N_8678,N_8028,N_7815);
xor U8679 (N_8679,N_8281,N_7907);
or U8680 (N_8680,N_7872,N_7903);
nand U8681 (N_8681,N_8138,N_7906);
or U8682 (N_8682,N_8097,N_8052);
and U8683 (N_8683,N_8232,N_8315);
and U8684 (N_8684,N_8264,N_8265);
xnor U8685 (N_8685,N_7899,N_7926);
or U8686 (N_8686,N_8296,N_8199);
nor U8687 (N_8687,N_8192,N_8322);
nor U8688 (N_8688,N_8399,N_7825);
nand U8689 (N_8689,N_7992,N_7826);
nor U8690 (N_8690,N_8016,N_8339);
nand U8691 (N_8691,N_8154,N_8083);
nand U8692 (N_8692,N_8267,N_8198);
and U8693 (N_8693,N_7901,N_8273);
nand U8694 (N_8694,N_8263,N_8195);
nand U8695 (N_8695,N_8035,N_8351);
nor U8696 (N_8696,N_8091,N_7848);
xor U8697 (N_8697,N_8230,N_8120);
or U8698 (N_8698,N_7919,N_8063);
and U8699 (N_8699,N_7856,N_7971);
nand U8700 (N_8700,N_8107,N_8154);
nor U8701 (N_8701,N_8202,N_8027);
or U8702 (N_8702,N_7855,N_8396);
nand U8703 (N_8703,N_8097,N_7945);
and U8704 (N_8704,N_7901,N_7888);
nor U8705 (N_8705,N_7983,N_7853);
nor U8706 (N_8706,N_8262,N_7927);
nand U8707 (N_8707,N_8323,N_7830);
or U8708 (N_8708,N_7943,N_8366);
nand U8709 (N_8709,N_7891,N_8305);
xnor U8710 (N_8710,N_8168,N_8070);
xor U8711 (N_8711,N_8170,N_8132);
or U8712 (N_8712,N_8197,N_8234);
nor U8713 (N_8713,N_7808,N_8082);
nor U8714 (N_8714,N_8291,N_8170);
nor U8715 (N_8715,N_8129,N_8218);
and U8716 (N_8716,N_7848,N_8220);
nor U8717 (N_8717,N_8196,N_8006);
nand U8718 (N_8718,N_8175,N_7941);
nand U8719 (N_8719,N_7948,N_8210);
and U8720 (N_8720,N_8004,N_8145);
nand U8721 (N_8721,N_8371,N_8288);
and U8722 (N_8722,N_7831,N_7820);
xnor U8723 (N_8723,N_8184,N_8155);
nor U8724 (N_8724,N_7924,N_8259);
nand U8725 (N_8725,N_8094,N_8139);
nand U8726 (N_8726,N_8209,N_7855);
and U8727 (N_8727,N_7847,N_7821);
xor U8728 (N_8728,N_8328,N_8230);
nor U8729 (N_8729,N_8289,N_8062);
xor U8730 (N_8730,N_7890,N_8272);
xnor U8731 (N_8731,N_8254,N_8214);
nand U8732 (N_8732,N_8397,N_8081);
or U8733 (N_8733,N_7902,N_8066);
or U8734 (N_8734,N_8290,N_8398);
nor U8735 (N_8735,N_7864,N_8240);
xnor U8736 (N_8736,N_8006,N_7882);
and U8737 (N_8737,N_8018,N_8295);
and U8738 (N_8738,N_8176,N_8157);
or U8739 (N_8739,N_8211,N_7860);
nor U8740 (N_8740,N_8321,N_8353);
xor U8741 (N_8741,N_8334,N_8362);
or U8742 (N_8742,N_8397,N_8330);
or U8743 (N_8743,N_8120,N_8038);
or U8744 (N_8744,N_7906,N_8224);
or U8745 (N_8745,N_8239,N_8229);
and U8746 (N_8746,N_8357,N_7862);
xor U8747 (N_8747,N_8380,N_8294);
and U8748 (N_8748,N_7890,N_8107);
nor U8749 (N_8749,N_7957,N_7892);
nor U8750 (N_8750,N_8178,N_7959);
and U8751 (N_8751,N_8178,N_7922);
and U8752 (N_8752,N_7889,N_7810);
nor U8753 (N_8753,N_8256,N_8325);
nor U8754 (N_8754,N_8074,N_8345);
or U8755 (N_8755,N_8304,N_8131);
or U8756 (N_8756,N_7921,N_8355);
and U8757 (N_8757,N_8350,N_8019);
and U8758 (N_8758,N_8240,N_8176);
nor U8759 (N_8759,N_7917,N_8072);
or U8760 (N_8760,N_8145,N_8200);
or U8761 (N_8761,N_8313,N_8120);
nor U8762 (N_8762,N_8290,N_8276);
nor U8763 (N_8763,N_7816,N_8028);
xnor U8764 (N_8764,N_7917,N_8115);
nor U8765 (N_8765,N_8175,N_7809);
xnor U8766 (N_8766,N_8293,N_8307);
nor U8767 (N_8767,N_8378,N_8129);
or U8768 (N_8768,N_8066,N_8120);
and U8769 (N_8769,N_8076,N_8330);
nor U8770 (N_8770,N_7919,N_8283);
or U8771 (N_8771,N_8309,N_8025);
or U8772 (N_8772,N_7856,N_8243);
xor U8773 (N_8773,N_8166,N_8240);
or U8774 (N_8774,N_8145,N_8109);
and U8775 (N_8775,N_7864,N_8103);
or U8776 (N_8776,N_8050,N_8172);
nand U8777 (N_8777,N_8170,N_7850);
xor U8778 (N_8778,N_8294,N_7943);
and U8779 (N_8779,N_8157,N_8191);
nor U8780 (N_8780,N_7986,N_8337);
or U8781 (N_8781,N_8142,N_7967);
and U8782 (N_8782,N_8152,N_7984);
and U8783 (N_8783,N_8243,N_8176);
xor U8784 (N_8784,N_8156,N_8293);
or U8785 (N_8785,N_8369,N_8142);
nand U8786 (N_8786,N_8191,N_7895);
xnor U8787 (N_8787,N_8047,N_8285);
nand U8788 (N_8788,N_7859,N_7868);
or U8789 (N_8789,N_8116,N_8253);
nand U8790 (N_8790,N_8232,N_8055);
or U8791 (N_8791,N_8029,N_7880);
or U8792 (N_8792,N_8016,N_8086);
or U8793 (N_8793,N_8129,N_8269);
and U8794 (N_8794,N_8076,N_7996);
xor U8795 (N_8795,N_8314,N_8046);
nand U8796 (N_8796,N_8195,N_8211);
xor U8797 (N_8797,N_7832,N_7920);
xor U8798 (N_8798,N_8318,N_7927);
xnor U8799 (N_8799,N_8074,N_8024);
nand U8800 (N_8800,N_7994,N_8353);
xnor U8801 (N_8801,N_8064,N_7951);
and U8802 (N_8802,N_7885,N_8332);
nor U8803 (N_8803,N_8101,N_8036);
or U8804 (N_8804,N_8088,N_8369);
xor U8805 (N_8805,N_7858,N_7806);
or U8806 (N_8806,N_8185,N_8157);
nand U8807 (N_8807,N_8382,N_8320);
and U8808 (N_8808,N_7868,N_8046);
or U8809 (N_8809,N_8116,N_8285);
nor U8810 (N_8810,N_7982,N_7947);
or U8811 (N_8811,N_8337,N_7832);
and U8812 (N_8812,N_8068,N_7971);
and U8813 (N_8813,N_7939,N_7894);
and U8814 (N_8814,N_8076,N_8201);
or U8815 (N_8815,N_8274,N_8097);
xor U8816 (N_8816,N_8035,N_7997);
xnor U8817 (N_8817,N_7817,N_8323);
nand U8818 (N_8818,N_7842,N_8039);
xnor U8819 (N_8819,N_8272,N_8057);
xnor U8820 (N_8820,N_8068,N_7857);
xnor U8821 (N_8821,N_8035,N_8284);
xor U8822 (N_8822,N_8011,N_8108);
xor U8823 (N_8823,N_8124,N_8122);
xnor U8824 (N_8824,N_8074,N_7989);
or U8825 (N_8825,N_8279,N_7945);
nor U8826 (N_8826,N_8361,N_7997);
and U8827 (N_8827,N_8234,N_7911);
and U8828 (N_8828,N_8062,N_8060);
nor U8829 (N_8829,N_7811,N_7842);
nand U8830 (N_8830,N_7830,N_8242);
or U8831 (N_8831,N_8275,N_7909);
xor U8832 (N_8832,N_8306,N_7920);
xor U8833 (N_8833,N_8363,N_7907);
nand U8834 (N_8834,N_8105,N_7879);
nor U8835 (N_8835,N_8078,N_7883);
and U8836 (N_8836,N_8338,N_8242);
and U8837 (N_8837,N_8009,N_8106);
nand U8838 (N_8838,N_7936,N_7878);
nor U8839 (N_8839,N_7860,N_8148);
and U8840 (N_8840,N_8101,N_7947);
nand U8841 (N_8841,N_7937,N_8325);
nor U8842 (N_8842,N_8053,N_8219);
and U8843 (N_8843,N_8000,N_8381);
nor U8844 (N_8844,N_8376,N_8085);
or U8845 (N_8845,N_8143,N_7867);
nor U8846 (N_8846,N_8263,N_7950);
and U8847 (N_8847,N_8267,N_8268);
nor U8848 (N_8848,N_8173,N_8384);
nand U8849 (N_8849,N_8150,N_8289);
xnor U8850 (N_8850,N_7884,N_8198);
xor U8851 (N_8851,N_8080,N_8043);
or U8852 (N_8852,N_8364,N_8007);
xor U8853 (N_8853,N_7876,N_8092);
or U8854 (N_8854,N_8251,N_7916);
nor U8855 (N_8855,N_7816,N_7824);
or U8856 (N_8856,N_8165,N_8104);
xor U8857 (N_8857,N_8117,N_7965);
nor U8858 (N_8858,N_8255,N_7842);
xnor U8859 (N_8859,N_8200,N_8060);
xnor U8860 (N_8860,N_8091,N_8390);
nand U8861 (N_8861,N_8161,N_7955);
or U8862 (N_8862,N_7940,N_8020);
xor U8863 (N_8863,N_8260,N_8133);
nand U8864 (N_8864,N_8264,N_8170);
nor U8865 (N_8865,N_8323,N_8206);
xor U8866 (N_8866,N_8078,N_7934);
nand U8867 (N_8867,N_8176,N_8187);
and U8868 (N_8868,N_8165,N_8069);
nor U8869 (N_8869,N_8276,N_8199);
and U8870 (N_8870,N_7982,N_7944);
or U8871 (N_8871,N_8299,N_7876);
and U8872 (N_8872,N_7904,N_7856);
xnor U8873 (N_8873,N_8169,N_8260);
nand U8874 (N_8874,N_7939,N_8166);
nor U8875 (N_8875,N_7929,N_8038);
nor U8876 (N_8876,N_7841,N_8115);
nor U8877 (N_8877,N_8095,N_8203);
xnor U8878 (N_8878,N_8177,N_7897);
xnor U8879 (N_8879,N_8040,N_8024);
nor U8880 (N_8880,N_8367,N_8144);
and U8881 (N_8881,N_7855,N_8204);
xnor U8882 (N_8882,N_8317,N_7924);
nand U8883 (N_8883,N_8162,N_7868);
nand U8884 (N_8884,N_8236,N_7812);
nand U8885 (N_8885,N_8316,N_8309);
xnor U8886 (N_8886,N_7984,N_7833);
nor U8887 (N_8887,N_8263,N_8108);
and U8888 (N_8888,N_8187,N_7916);
and U8889 (N_8889,N_8232,N_8236);
xor U8890 (N_8890,N_7813,N_8229);
xor U8891 (N_8891,N_7864,N_7998);
or U8892 (N_8892,N_8250,N_8199);
nor U8893 (N_8893,N_8124,N_7986);
nand U8894 (N_8894,N_7819,N_7951);
or U8895 (N_8895,N_8086,N_8174);
and U8896 (N_8896,N_8214,N_7827);
or U8897 (N_8897,N_8141,N_7924);
nor U8898 (N_8898,N_8245,N_8383);
nand U8899 (N_8899,N_8125,N_8003);
xnor U8900 (N_8900,N_8262,N_7981);
and U8901 (N_8901,N_8240,N_8342);
nor U8902 (N_8902,N_8058,N_7901);
nand U8903 (N_8903,N_8020,N_8351);
and U8904 (N_8904,N_7910,N_8177);
xor U8905 (N_8905,N_8276,N_7929);
or U8906 (N_8906,N_8225,N_8313);
xor U8907 (N_8907,N_8228,N_7939);
nand U8908 (N_8908,N_7901,N_7999);
nor U8909 (N_8909,N_8359,N_7907);
or U8910 (N_8910,N_8096,N_7948);
or U8911 (N_8911,N_8252,N_7955);
nor U8912 (N_8912,N_8109,N_8236);
nor U8913 (N_8913,N_7913,N_8076);
nand U8914 (N_8914,N_8002,N_7957);
xor U8915 (N_8915,N_8187,N_7853);
xnor U8916 (N_8916,N_8221,N_8270);
or U8917 (N_8917,N_8142,N_8003);
nor U8918 (N_8918,N_7936,N_8157);
and U8919 (N_8919,N_8112,N_7870);
xor U8920 (N_8920,N_8188,N_8357);
nor U8921 (N_8921,N_8098,N_7927);
xor U8922 (N_8922,N_7855,N_8184);
or U8923 (N_8923,N_8130,N_8355);
xor U8924 (N_8924,N_7926,N_8115);
or U8925 (N_8925,N_8085,N_7822);
or U8926 (N_8926,N_7907,N_7970);
or U8927 (N_8927,N_8266,N_8111);
nor U8928 (N_8928,N_8319,N_7878);
nor U8929 (N_8929,N_7825,N_8300);
or U8930 (N_8930,N_8043,N_8270);
nand U8931 (N_8931,N_8039,N_8125);
nand U8932 (N_8932,N_8060,N_8013);
or U8933 (N_8933,N_8368,N_8137);
nor U8934 (N_8934,N_8226,N_8155);
or U8935 (N_8935,N_8348,N_8195);
nand U8936 (N_8936,N_7810,N_8208);
and U8937 (N_8937,N_8107,N_7893);
and U8938 (N_8938,N_8356,N_7906);
xnor U8939 (N_8939,N_8154,N_8193);
nand U8940 (N_8940,N_8022,N_7817);
nor U8941 (N_8941,N_8283,N_8294);
and U8942 (N_8942,N_8090,N_7994);
or U8943 (N_8943,N_8148,N_8189);
nor U8944 (N_8944,N_7991,N_8049);
nand U8945 (N_8945,N_8200,N_7969);
nand U8946 (N_8946,N_7870,N_8110);
or U8947 (N_8947,N_8075,N_8338);
nand U8948 (N_8948,N_7870,N_7996);
nor U8949 (N_8949,N_7901,N_8115);
or U8950 (N_8950,N_7823,N_8383);
nor U8951 (N_8951,N_8328,N_7971);
and U8952 (N_8952,N_7923,N_7831);
nor U8953 (N_8953,N_8158,N_8307);
nand U8954 (N_8954,N_8153,N_8024);
nand U8955 (N_8955,N_8069,N_7897);
nand U8956 (N_8956,N_8189,N_8319);
nand U8957 (N_8957,N_8391,N_7806);
and U8958 (N_8958,N_7821,N_8275);
xor U8959 (N_8959,N_8310,N_7977);
or U8960 (N_8960,N_8207,N_7960);
nor U8961 (N_8961,N_8162,N_8275);
nor U8962 (N_8962,N_8303,N_8397);
or U8963 (N_8963,N_8094,N_8361);
or U8964 (N_8964,N_8258,N_8284);
xor U8965 (N_8965,N_8056,N_8371);
and U8966 (N_8966,N_7855,N_7884);
xor U8967 (N_8967,N_8017,N_7983);
nand U8968 (N_8968,N_8158,N_7842);
and U8969 (N_8969,N_8202,N_8045);
and U8970 (N_8970,N_7934,N_8294);
and U8971 (N_8971,N_8154,N_8296);
and U8972 (N_8972,N_7856,N_7969);
nor U8973 (N_8973,N_8036,N_8373);
nor U8974 (N_8974,N_7827,N_7903);
or U8975 (N_8975,N_7973,N_7921);
and U8976 (N_8976,N_7810,N_8026);
xor U8977 (N_8977,N_8107,N_8098);
xor U8978 (N_8978,N_7848,N_8065);
xnor U8979 (N_8979,N_8012,N_8099);
nor U8980 (N_8980,N_7873,N_8017);
and U8981 (N_8981,N_8113,N_8056);
nand U8982 (N_8982,N_8322,N_8399);
and U8983 (N_8983,N_8120,N_8285);
or U8984 (N_8984,N_7971,N_7922);
or U8985 (N_8985,N_7871,N_8190);
xnor U8986 (N_8986,N_8377,N_7953);
or U8987 (N_8987,N_8253,N_8219);
xor U8988 (N_8988,N_7832,N_8266);
and U8989 (N_8989,N_8040,N_8288);
nor U8990 (N_8990,N_8256,N_7947);
nor U8991 (N_8991,N_8183,N_8278);
and U8992 (N_8992,N_7884,N_8186);
nand U8993 (N_8993,N_7979,N_8080);
or U8994 (N_8994,N_8301,N_7893);
nand U8995 (N_8995,N_8062,N_8081);
nand U8996 (N_8996,N_8096,N_7891);
and U8997 (N_8997,N_7847,N_8058);
or U8998 (N_8998,N_8149,N_7870);
nor U8999 (N_8999,N_8288,N_7845);
xor U9000 (N_9000,N_8424,N_8802);
or U9001 (N_9001,N_8736,N_8815);
nor U9002 (N_9002,N_8684,N_8586);
xnor U9003 (N_9003,N_8745,N_8696);
xor U9004 (N_9004,N_8492,N_8969);
or U9005 (N_9005,N_8551,N_8841);
or U9006 (N_9006,N_8606,N_8585);
or U9007 (N_9007,N_8409,N_8865);
or U9008 (N_9008,N_8739,N_8809);
nor U9009 (N_9009,N_8598,N_8703);
nor U9010 (N_9010,N_8646,N_8909);
nand U9011 (N_9011,N_8594,N_8746);
nand U9012 (N_9012,N_8765,N_8843);
xor U9013 (N_9013,N_8818,N_8700);
and U9014 (N_9014,N_8812,N_8737);
and U9015 (N_9015,N_8762,N_8524);
or U9016 (N_9016,N_8845,N_8619);
or U9017 (N_9017,N_8501,N_8853);
and U9018 (N_9018,N_8669,N_8849);
or U9019 (N_9019,N_8611,N_8564);
and U9020 (N_9020,N_8698,N_8472);
or U9021 (N_9021,N_8469,N_8904);
and U9022 (N_9022,N_8774,N_8443);
xnor U9023 (N_9023,N_8780,N_8952);
or U9024 (N_9024,N_8931,N_8692);
and U9025 (N_9025,N_8872,N_8577);
or U9026 (N_9026,N_8824,N_8667);
nand U9027 (N_9027,N_8595,N_8691);
xnor U9028 (N_9028,N_8715,N_8694);
and U9029 (N_9029,N_8814,N_8868);
nand U9030 (N_9030,N_8532,N_8444);
nor U9031 (N_9031,N_8782,N_8572);
nand U9032 (N_9032,N_8593,N_8429);
nand U9033 (N_9033,N_8942,N_8450);
or U9034 (N_9034,N_8857,N_8587);
nor U9035 (N_9035,N_8930,N_8880);
and U9036 (N_9036,N_8555,N_8754);
xnor U9037 (N_9037,N_8597,N_8436);
nor U9038 (N_9038,N_8924,N_8738);
and U9039 (N_9039,N_8773,N_8903);
nand U9040 (N_9040,N_8721,N_8975);
or U9041 (N_9041,N_8453,N_8955);
nand U9042 (N_9042,N_8658,N_8860);
nand U9043 (N_9043,N_8592,N_8954);
xor U9044 (N_9044,N_8478,N_8674);
xor U9045 (N_9045,N_8580,N_8718);
nand U9046 (N_9046,N_8601,N_8428);
or U9047 (N_9047,N_8888,N_8591);
or U9048 (N_9048,N_8596,N_8490);
or U9049 (N_9049,N_8829,N_8822);
xor U9050 (N_9050,N_8751,N_8726);
or U9051 (N_9051,N_8633,N_8590);
and U9052 (N_9052,N_8526,N_8432);
xnor U9053 (N_9053,N_8796,N_8949);
or U9054 (N_9054,N_8455,N_8759);
nor U9055 (N_9055,N_8827,N_8886);
nand U9056 (N_9056,N_8426,N_8621);
nand U9057 (N_9057,N_8533,N_8729);
or U9058 (N_9058,N_8400,N_8471);
xnor U9059 (N_9059,N_8465,N_8987);
nor U9060 (N_9060,N_8850,N_8489);
nor U9061 (N_9061,N_8420,N_8846);
and U9062 (N_9062,N_8407,N_8433);
and U9063 (N_9063,N_8803,N_8764);
nor U9064 (N_9064,N_8410,N_8806);
and U9065 (N_9065,N_8517,N_8463);
or U9066 (N_9066,N_8670,N_8999);
nor U9067 (N_9067,N_8608,N_8913);
nand U9068 (N_9068,N_8892,N_8981);
nor U9069 (N_9069,N_8506,N_8530);
or U9070 (N_9070,N_8705,N_8704);
nand U9071 (N_9071,N_8724,N_8874);
nand U9072 (N_9072,N_8602,N_8638);
nor U9073 (N_9073,N_8588,N_8682);
and U9074 (N_9074,N_8878,N_8933);
and U9075 (N_9075,N_8451,N_8749);
nor U9076 (N_9076,N_8474,N_8786);
or U9077 (N_9077,N_8864,N_8567);
and U9078 (N_9078,N_8722,N_8852);
or U9079 (N_9079,N_8760,N_8421);
xnor U9080 (N_9080,N_8734,N_8997);
or U9081 (N_9081,N_8498,N_8673);
xnor U9082 (N_9082,N_8537,N_8816);
and U9083 (N_9083,N_8542,N_8483);
xnor U9084 (N_9084,N_8640,N_8914);
nand U9085 (N_9085,N_8991,N_8541);
nand U9086 (N_9086,N_8512,N_8578);
nand U9087 (N_9087,N_8877,N_8900);
and U9088 (N_9088,N_8659,N_8702);
and U9089 (N_9089,N_8756,N_8761);
and U9090 (N_9090,N_8891,N_8459);
nor U9091 (N_9091,N_8630,N_8821);
nor U9092 (N_9092,N_8953,N_8730);
or U9093 (N_9093,N_8644,N_8716);
nor U9094 (N_9094,N_8466,N_8811);
xor U9095 (N_9095,N_8844,N_8939);
or U9096 (N_9096,N_8748,N_8847);
xnor U9097 (N_9097,N_8576,N_8476);
nand U9098 (N_9098,N_8923,N_8779);
nor U9099 (N_9099,N_8972,N_8701);
nand U9100 (N_9100,N_8959,N_8916);
and U9101 (N_9101,N_8950,N_8623);
nand U9102 (N_9102,N_8507,N_8518);
or U9103 (N_9103,N_8826,N_8529);
xor U9104 (N_9104,N_8744,N_8495);
nand U9105 (N_9105,N_8538,N_8488);
nand U9106 (N_9106,N_8448,N_8560);
or U9107 (N_9107,N_8414,N_8713);
nand U9108 (N_9108,N_8525,N_8966);
nor U9109 (N_9109,N_8415,N_8856);
and U9110 (N_9110,N_8666,N_8990);
nand U9111 (N_9111,N_8895,N_8614);
nor U9112 (N_9112,N_8493,N_8677);
nand U9113 (N_9113,N_8446,N_8511);
or U9114 (N_9114,N_8743,N_8719);
and U9115 (N_9115,N_8487,N_8554);
and U9116 (N_9116,N_8610,N_8613);
nand U9117 (N_9117,N_8976,N_8766);
and U9118 (N_9118,N_8618,N_8571);
nor U9119 (N_9119,N_8984,N_8968);
nor U9120 (N_9120,N_8550,N_8642);
and U9121 (N_9121,N_8604,N_8676);
and U9122 (N_9122,N_8750,N_8731);
nor U9123 (N_9123,N_8648,N_8652);
nand U9124 (N_9124,N_8481,N_8938);
xnor U9125 (N_9125,N_8600,N_8998);
or U9126 (N_9126,N_8695,N_8767);
and U9127 (N_9127,N_8875,N_8539);
and U9128 (N_9128,N_8902,N_8553);
and U9129 (N_9129,N_8449,N_8427);
or U9130 (N_9130,N_8625,N_8770);
and U9131 (N_9131,N_8484,N_8657);
and U9132 (N_9132,N_8906,N_8645);
nand U9133 (N_9133,N_8830,N_8664);
xor U9134 (N_9134,N_8934,N_8548);
nor U9135 (N_9135,N_8989,N_8438);
nor U9136 (N_9136,N_8480,N_8499);
xor U9137 (N_9137,N_8675,N_8650);
and U9138 (N_9138,N_8919,N_8635);
nand U9139 (N_9139,N_8681,N_8974);
and U9140 (N_9140,N_8800,N_8435);
or U9141 (N_9141,N_8519,N_8521);
and U9142 (N_9142,N_8452,N_8647);
xor U9143 (N_9143,N_8817,N_8653);
nand U9144 (N_9144,N_8883,N_8475);
nand U9145 (N_9145,N_8884,N_8683);
nor U9146 (N_9146,N_8755,N_8651);
xnor U9147 (N_9147,N_8561,N_8851);
and U9148 (N_9148,N_8985,N_8528);
nand U9149 (N_9149,N_8535,N_8928);
xnor U9150 (N_9150,N_8876,N_8970);
nor U9151 (N_9151,N_8497,N_8763);
nor U9152 (N_9152,N_8889,N_8871);
nor U9153 (N_9153,N_8482,N_8791);
or U9154 (N_9154,N_8935,N_8839);
xor U9155 (N_9155,N_8869,N_8707);
nand U9156 (N_9156,N_8562,N_8920);
nand U9157 (N_9157,N_8717,N_8977);
and U9158 (N_9158,N_8982,N_8753);
xnor U9159 (N_9159,N_8907,N_8757);
xnor U9160 (N_9160,N_8842,N_8973);
or U9161 (N_9161,N_8685,N_8788);
xor U9162 (N_9162,N_8747,N_8464);
and U9163 (N_9163,N_8879,N_8958);
and U9164 (N_9164,N_8584,N_8566);
nand U9165 (N_9165,N_8454,N_8494);
nor U9166 (N_9166,N_8711,N_8714);
or U9167 (N_9167,N_8838,N_8881);
and U9168 (N_9168,N_8798,N_8793);
and U9169 (N_9169,N_8956,N_8946);
xnor U9170 (N_9170,N_8565,N_8708);
and U9171 (N_9171,N_8859,N_8855);
nor U9172 (N_9172,N_8544,N_8522);
nand U9173 (N_9173,N_8993,N_8470);
and U9174 (N_9174,N_8403,N_8742);
nand U9175 (N_9175,N_8686,N_8558);
xnor U9176 (N_9176,N_8899,N_8500);
nor U9177 (N_9177,N_8479,N_8922);
xor U9178 (N_9178,N_8948,N_8706);
and U9179 (N_9179,N_8994,N_8992);
nand U9180 (N_9180,N_8911,N_8733);
xnor U9181 (N_9181,N_8790,N_8980);
nand U9182 (N_9182,N_8693,N_8617);
or U9183 (N_9183,N_8486,N_8442);
or U9184 (N_9184,N_8965,N_8837);
xor U9185 (N_9185,N_8575,N_8795);
xor U9186 (N_9186,N_8629,N_8505);
nand U9187 (N_9187,N_8679,N_8527);
xor U9188 (N_9188,N_8835,N_8406);
xor U9189 (N_9189,N_8758,N_8634);
nand U9190 (N_9190,N_8418,N_8569);
or U9191 (N_9191,N_8820,N_8688);
nor U9192 (N_9192,N_8962,N_8456);
or U9193 (N_9193,N_8710,N_8639);
and U9194 (N_9194,N_8785,N_8402);
or U9195 (N_9195,N_8534,N_8712);
nor U9196 (N_9196,N_8515,N_8936);
nor U9197 (N_9197,N_8612,N_8727);
nand U9198 (N_9198,N_8599,N_8740);
or U9199 (N_9199,N_8978,N_8858);
and U9200 (N_9200,N_8825,N_8579);
nand U9201 (N_9201,N_8431,N_8461);
nor U9202 (N_9202,N_8967,N_8508);
and U9203 (N_9203,N_8496,N_8901);
and U9204 (N_9204,N_8627,N_8545);
nor U9205 (N_9205,N_8603,N_8626);
or U9206 (N_9206,N_8416,N_8405);
and U9207 (N_9207,N_8531,N_8460);
or U9208 (N_9208,N_8689,N_8964);
nand U9209 (N_9209,N_8732,N_8661);
nor U9210 (N_9210,N_8915,N_8687);
and U9211 (N_9211,N_8557,N_8583);
or U9212 (N_9212,N_8784,N_8996);
or U9213 (N_9213,N_8932,N_8777);
nor U9214 (N_9214,N_8672,N_8794);
xnor U9215 (N_9215,N_8468,N_8951);
nand U9216 (N_9216,N_8411,N_8771);
and U9217 (N_9217,N_8910,N_8504);
or U9218 (N_9218,N_8979,N_8945);
nor U9219 (N_9219,N_8543,N_8632);
nor U9220 (N_9220,N_8840,N_8917);
nor U9221 (N_9221,N_8775,N_8831);
xor U9222 (N_9222,N_8894,N_8781);
xor U9223 (N_9223,N_8641,N_8656);
xor U9224 (N_9224,N_8417,N_8801);
or U9225 (N_9225,N_8918,N_8813);
nor U9226 (N_9226,N_8441,N_8568);
xor U9227 (N_9227,N_8662,N_8609);
nor U9228 (N_9228,N_8631,N_8473);
and U9229 (N_9229,N_8988,N_8908);
or U9230 (N_9230,N_8408,N_8862);
nor U9231 (N_9231,N_8622,N_8581);
xnor U9232 (N_9232,N_8668,N_8447);
or U9233 (N_9233,N_8804,N_8768);
xnor U9234 (N_9234,N_8921,N_8810);
nor U9235 (N_9235,N_8404,N_8728);
xnor U9236 (N_9236,N_8940,N_8440);
nor U9237 (N_9237,N_8573,N_8772);
nor U9238 (N_9238,N_8422,N_8834);
xnor U9239 (N_9239,N_8983,N_8615);
or U9240 (N_9240,N_8873,N_8905);
or U9241 (N_9241,N_8485,N_8699);
or U9242 (N_9242,N_8546,N_8477);
or U9243 (N_9243,N_8552,N_8735);
nand U9244 (N_9244,N_8467,N_8823);
or U9245 (N_9245,N_8799,N_8655);
nor U9246 (N_9246,N_8509,N_8503);
xor U9247 (N_9247,N_8663,N_8514);
nand U9248 (N_9248,N_8995,N_8890);
or U9249 (N_9249,N_8863,N_8605);
nor U9250 (N_9250,N_8412,N_8723);
nand U9251 (N_9251,N_8783,N_8523);
and U9252 (N_9252,N_8654,N_8971);
xor U9253 (N_9253,N_8836,N_8944);
xor U9254 (N_9254,N_8425,N_8607);
nor U9255 (N_9255,N_8709,N_8963);
or U9256 (N_9256,N_8589,N_8792);
nand U9257 (N_9257,N_8439,N_8559);
nor U9258 (N_9258,N_8925,N_8419);
nand U9259 (N_9259,N_8462,N_8437);
or U9260 (N_9260,N_8805,N_8960);
nand U9261 (N_9261,N_8882,N_8536);
xor U9262 (N_9262,N_8671,N_8616);
nand U9263 (N_9263,N_8516,N_8556);
nand U9264 (N_9264,N_8574,N_8697);
nand U9265 (N_9265,N_8866,N_8636);
or U9266 (N_9266,N_8423,N_8885);
or U9267 (N_9267,N_8725,N_8649);
or U9268 (N_9268,N_8628,N_8458);
and U9269 (N_9269,N_8957,N_8540);
xnor U9270 (N_9270,N_8926,N_8943);
nand U9271 (N_9271,N_8789,N_8867);
or U9272 (N_9272,N_8741,N_8720);
or U9273 (N_9273,N_8870,N_8778);
or U9274 (N_9274,N_8896,N_8912);
xor U9275 (N_9275,N_8752,N_8401);
and U9276 (N_9276,N_8808,N_8833);
and U9277 (N_9277,N_8787,N_8620);
nor U9278 (N_9278,N_8854,N_8961);
nand U9279 (N_9279,N_8819,N_8927);
or U9280 (N_9280,N_8848,N_8430);
and U9281 (N_9281,N_8582,N_8520);
and U9282 (N_9282,N_8861,N_8897);
and U9283 (N_9283,N_8665,N_8549);
xnor U9284 (N_9284,N_8502,N_8513);
nor U9285 (N_9285,N_8947,N_8563);
xnor U9286 (N_9286,N_8457,N_8690);
xnor U9287 (N_9287,N_8680,N_8413);
nor U9288 (N_9288,N_8986,N_8941);
xor U9289 (N_9289,N_8570,N_8491);
nor U9290 (N_9290,N_8547,N_8434);
and U9291 (N_9291,N_8797,N_8807);
nand U9292 (N_9292,N_8445,N_8660);
or U9293 (N_9293,N_8643,N_8678);
and U9294 (N_9294,N_8510,N_8769);
nand U9295 (N_9295,N_8624,N_8832);
and U9296 (N_9296,N_8776,N_8828);
or U9297 (N_9297,N_8929,N_8937);
and U9298 (N_9298,N_8893,N_8898);
xnor U9299 (N_9299,N_8637,N_8887);
or U9300 (N_9300,N_8580,N_8509);
and U9301 (N_9301,N_8892,N_8428);
and U9302 (N_9302,N_8426,N_8553);
and U9303 (N_9303,N_8560,N_8643);
nor U9304 (N_9304,N_8856,N_8736);
nor U9305 (N_9305,N_8541,N_8652);
and U9306 (N_9306,N_8567,N_8950);
and U9307 (N_9307,N_8865,N_8579);
xor U9308 (N_9308,N_8507,N_8749);
or U9309 (N_9309,N_8507,N_8895);
nand U9310 (N_9310,N_8951,N_8661);
and U9311 (N_9311,N_8449,N_8550);
or U9312 (N_9312,N_8853,N_8716);
nor U9313 (N_9313,N_8657,N_8461);
nor U9314 (N_9314,N_8887,N_8955);
nand U9315 (N_9315,N_8631,N_8831);
nand U9316 (N_9316,N_8528,N_8668);
xnor U9317 (N_9317,N_8880,N_8519);
nor U9318 (N_9318,N_8914,N_8916);
or U9319 (N_9319,N_8455,N_8981);
and U9320 (N_9320,N_8647,N_8508);
and U9321 (N_9321,N_8737,N_8667);
nor U9322 (N_9322,N_8737,N_8585);
and U9323 (N_9323,N_8674,N_8856);
nand U9324 (N_9324,N_8692,N_8910);
nor U9325 (N_9325,N_8950,N_8643);
xnor U9326 (N_9326,N_8650,N_8415);
nor U9327 (N_9327,N_8652,N_8876);
and U9328 (N_9328,N_8538,N_8808);
or U9329 (N_9329,N_8798,N_8964);
nand U9330 (N_9330,N_8899,N_8843);
nor U9331 (N_9331,N_8601,N_8530);
nor U9332 (N_9332,N_8875,N_8766);
or U9333 (N_9333,N_8812,N_8703);
or U9334 (N_9334,N_8857,N_8526);
nor U9335 (N_9335,N_8718,N_8814);
and U9336 (N_9336,N_8453,N_8669);
and U9337 (N_9337,N_8571,N_8841);
nand U9338 (N_9338,N_8484,N_8798);
nand U9339 (N_9339,N_8628,N_8883);
nand U9340 (N_9340,N_8932,N_8428);
xor U9341 (N_9341,N_8729,N_8703);
and U9342 (N_9342,N_8513,N_8781);
xnor U9343 (N_9343,N_8521,N_8854);
nand U9344 (N_9344,N_8500,N_8848);
nand U9345 (N_9345,N_8933,N_8527);
xnor U9346 (N_9346,N_8642,N_8469);
or U9347 (N_9347,N_8927,N_8782);
and U9348 (N_9348,N_8557,N_8915);
or U9349 (N_9349,N_8913,N_8833);
and U9350 (N_9350,N_8779,N_8595);
and U9351 (N_9351,N_8965,N_8657);
nor U9352 (N_9352,N_8495,N_8614);
or U9353 (N_9353,N_8976,N_8882);
nor U9354 (N_9354,N_8579,N_8624);
and U9355 (N_9355,N_8695,N_8447);
nand U9356 (N_9356,N_8932,N_8480);
or U9357 (N_9357,N_8552,N_8945);
nor U9358 (N_9358,N_8639,N_8483);
or U9359 (N_9359,N_8711,N_8535);
nor U9360 (N_9360,N_8872,N_8707);
nand U9361 (N_9361,N_8591,N_8706);
xor U9362 (N_9362,N_8782,N_8413);
nor U9363 (N_9363,N_8704,N_8434);
and U9364 (N_9364,N_8712,N_8946);
and U9365 (N_9365,N_8957,N_8405);
nand U9366 (N_9366,N_8976,N_8835);
nand U9367 (N_9367,N_8614,N_8772);
nand U9368 (N_9368,N_8656,N_8670);
nor U9369 (N_9369,N_8952,N_8584);
nand U9370 (N_9370,N_8400,N_8763);
and U9371 (N_9371,N_8951,N_8901);
nor U9372 (N_9372,N_8876,N_8556);
xnor U9373 (N_9373,N_8771,N_8517);
nor U9374 (N_9374,N_8699,N_8971);
or U9375 (N_9375,N_8512,N_8588);
nor U9376 (N_9376,N_8491,N_8433);
and U9377 (N_9377,N_8929,N_8444);
or U9378 (N_9378,N_8693,N_8556);
xor U9379 (N_9379,N_8478,N_8709);
or U9380 (N_9380,N_8928,N_8674);
or U9381 (N_9381,N_8488,N_8626);
nand U9382 (N_9382,N_8463,N_8424);
xnor U9383 (N_9383,N_8527,N_8751);
or U9384 (N_9384,N_8726,N_8534);
nand U9385 (N_9385,N_8612,N_8945);
and U9386 (N_9386,N_8693,N_8429);
nand U9387 (N_9387,N_8813,N_8667);
or U9388 (N_9388,N_8541,N_8771);
xnor U9389 (N_9389,N_8904,N_8931);
xnor U9390 (N_9390,N_8732,N_8488);
or U9391 (N_9391,N_8921,N_8780);
or U9392 (N_9392,N_8837,N_8592);
xor U9393 (N_9393,N_8736,N_8642);
and U9394 (N_9394,N_8567,N_8699);
nand U9395 (N_9395,N_8676,N_8478);
and U9396 (N_9396,N_8934,N_8955);
xnor U9397 (N_9397,N_8501,N_8650);
nand U9398 (N_9398,N_8893,N_8806);
xor U9399 (N_9399,N_8928,N_8793);
or U9400 (N_9400,N_8497,N_8478);
nor U9401 (N_9401,N_8910,N_8682);
and U9402 (N_9402,N_8645,N_8671);
xnor U9403 (N_9403,N_8810,N_8499);
xor U9404 (N_9404,N_8587,N_8739);
and U9405 (N_9405,N_8481,N_8748);
nand U9406 (N_9406,N_8604,N_8625);
or U9407 (N_9407,N_8956,N_8790);
or U9408 (N_9408,N_8581,N_8436);
nor U9409 (N_9409,N_8428,N_8822);
nor U9410 (N_9410,N_8801,N_8650);
and U9411 (N_9411,N_8584,N_8783);
nand U9412 (N_9412,N_8665,N_8494);
or U9413 (N_9413,N_8605,N_8684);
nor U9414 (N_9414,N_8829,N_8947);
xor U9415 (N_9415,N_8476,N_8758);
and U9416 (N_9416,N_8643,N_8771);
nand U9417 (N_9417,N_8543,N_8858);
or U9418 (N_9418,N_8685,N_8888);
and U9419 (N_9419,N_8869,N_8665);
or U9420 (N_9420,N_8957,N_8749);
nand U9421 (N_9421,N_8511,N_8796);
and U9422 (N_9422,N_8820,N_8457);
or U9423 (N_9423,N_8450,N_8846);
and U9424 (N_9424,N_8946,N_8485);
nand U9425 (N_9425,N_8669,N_8904);
nand U9426 (N_9426,N_8701,N_8843);
or U9427 (N_9427,N_8809,N_8730);
nand U9428 (N_9428,N_8766,N_8994);
or U9429 (N_9429,N_8661,N_8470);
nor U9430 (N_9430,N_8618,N_8849);
xnor U9431 (N_9431,N_8622,N_8599);
or U9432 (N_9432,N_8869,N_8473);
nor U9433 (N_9433,N_8834,N_8922);
xnor U9434 (N_9434,N_8506,N_8606);
or U9435 (N_9435,N_8472,N_8577);
nand U9436 (N_9436,N_8701,N_8957);
nor U9437 (N_9437,N_8436,N_8734);
or U9438 (N_9438,N_8418,N_8953);
and U9439 (N_9439,N_8822,N_8680);
xor U9440 (N_9440,N_8644,N_8406);
nand U9441 (N_9441,N_8911,N_8863);
xor U9442 (N_9442,N_8431,N_8577);
or U9443 (N_9443,N_8430,N_8780);
or U9444 (N_9444,N_8416,N_8466);
xor U9445 (N_9445,N_8812,N_8920);
and U9446 (N_9446,N_8674,N_8756);
nor U9447 (N_9447,N_8857,N_8852);
xnor U9448 (N_9448,N_8437,N_8936);
xor U9449 (N_9449,N_8829,N_8669);
nand U9450 (N_9450,N_8646,N_8762);
nand U9451 (N_9451,N_8827,N_8967);
nand U9452 (N_9452,N_8544,N_8604);
or U9453 (N_9453,N_8968,N_8495);
xnor U9454 (N_9454,N_8692,N_8512);
nor U9455 (N_9455,N_8949,N_8651);
nand U9456 (N_9456,N_8707,N_8518);
nand U9457 (N_9457,N_8784,N_8834);
nand U9458 (N_9458,N_8924,N_8744);
nand U9459 (N_9459,N_8754,N_8510);
nand U9460 (N_9460,N_8538,N_8811);
xnor U9461 (N_9461,N_8559,N_8535);
nor U9462 (N_9462,N_8768,N_8609);
nor U9463 (N_9463,N_8892,N_8536);
nor U9464 (N_9464,N_8905,N_8870);
and U9465 (N_9465,N_8559,N_8911);
and U9466 (N_9466,N_8801,N_8723);
nand U9467 (N_9467,N_8430,N_8498);
or U9468 (N_9468,N_8482,N_8937);
and U9469 (N_9469,N_8716,N_8705);
and U9470 (N_9470,N_8536,N_8784);
nor U9471 (N_9471,N_8954,N_8806);
xor U9472 (N_9472,N_8689,N_8791);
nor U9473 (N_9473,N_8647,N_8730);
or U9474 (N_9474,N_8528,N_8499);
nand U9475 (N_9475,N_8977,N_8708);
nor U9476 (N_9476,N_8568,N_8995);
nor U9477 (N_9477,N_8504,N_8434);
and U9478 (N_9478,N_8949,N_8642);
nand U9479 (N_9479,N_8918,N_8561);
nor U9480 (N_9480,N_8666,N_8820);
xnor U9481 (N_9481,N_8710,N_8944);
nand U9482 (N_9482,N_8569,N_8901);
xor U9483 (N_9483,N_8835,N_8937);
nand U9484 (N_9484,N_8836,N_8642);
xnor U9485 (N_9485,N_8946,N_8793);
and U9486 (N_9486,N_8428,N_8422);
xor U9487 (N_9487,N_8927,N_8916);
nor U9488 (N_9488,N_8793,N_8628);
nor U9489 (N_9489,N_8705,N_8831);
nand U9490 (N_9490,N_8577,N_8650);
or U9491 (N_9491,N_8922,N_8613);
xnor U9492 (N_9492,N_8513,N_8645);
xnor U9493 (N_9493,N_8993,N_8889);
and U9494 (N_9494,N_8987,N_8949);
or U9495 (N_9495,N_8847,N_8510);
or U9496 (N_9496,N_8964,N_8643);
nor U9497 (N_9497,N_8648,N_8960);
nor U9498 (N_9498,N_8818,N_8730);
nor U9499 (N_9499,N_8700,N_8641);
xor U9500 (N_9500,N_8777,N_8400);
or U9501 (N_9501,N_8680,N_8605);
nor U9502 (N_9502,N_8770,N_8512);
nand U9503 (N_9503,N_8707,N_8807);
nor U9504 (N_9504,N_8995,N_8740);
and U9505 (N_9505,N_8622,N_8612);
nor U9506 (N_9506,N_8702,N_8468);
nor U9507 (N_9507,N_8828,N_8426);
nand U9508 (N_9508,N_8725,N_8643);
nand U9509 (N_9509,N_8913,N_8810);
xnor U9510 (N_9510,N_8770,N_8618);
xnor U9511 (N_9511,N_8653,N_8513);
or U9512 (N_9512,N_8729,N_8797);
nand U9513 (N_9513,N_8836,N_8545);
nor U9514 (N_9514,N_8838,N_8866);
and U9515 (N_9515,N_8907,N_8624);
xor U9516 (N_9516,N_8939,N_8738);
nand U9517 (N_9517,N_8743,N_8748);
nand U9518 (N_9518,N_8646,N_8442);
nand U9519 (N_9519,N_8911,N_8936);
and U9520 (N_9520,N_8834,N_8950);
nand U9521 (N_9521,N_8631,N_8690);
xnor U9522 (N_9522,N_8520,N_8798);
nor U9523 (N_9523,N_8923,N_8704);
or U9524 (N_9524,N_8502,N_8690);
nor U9525 (N_9525,N_8889,N_8950);
and U9526 (N_9526,N_8880,N_8479);
and U9527 (N_9527,N_8941,N_8859);
nand U9528 (N_9528,N_8402,N_8782);
and U9529 (N_9529,N_8935,N_8655);
nor U9530 (N_9530,N_8517,N_8902);
or U9531 (N_9531,N_8743,N_8874);
nand U9532 (N_9532,N_8950,N_8530);
and U9533 (N_9533,N_8909,N_8503);
or U9534 (N_9534,N_8972,N_8861);
xnor U9535 (N_9535,N_8686,N_8507);
and U9536 (N_9536,N_8480,N_8806);
nor U9537 (N_9537,N_8796,N_8522);
nand U9538 (N_9538,N_8899,N_8675);
nand U9539 (N_9539,N_8993,N_8950);
xnor U9540 (N_9540,N_8739,N_8730);
xor U9541 (N_9541,N_8981,N_8688);
or U9542 (N_9542,N_8814,N_8901);
xor U9543 (N_9543,N_8413,N_8979);
nand U9544 (N_9544,N_8697,N_8493);
and U9545 (N_9545,N_8572,N_8952);
nand U9546 (N_9546,N_8975,N_8693);
or U9547 (N_9547,N_8798,N_8791);
nor U9548 (N_9548,N_8635,N_8842);
nor U9549 (N_9549,N_8864,N_8470);
nor U9550 (N_9550,N_8411,N_8800);
and U9551 (N_9551,N_8997,N_8751);
or U9552 (N_9552,N_8926,N_8758);
and U9553 (N_9553,N_8448,N_8430);
xor U9554 (N_9554,N_8544,N_8674);
and U9555 (N_9555,N_8910,N_8636);
nor U9556 (N_9556,N_8411,N_8663);
nor U9557 (N_9557,N_8481,N_8479);
nor U9558 (N_9558,N_8977,N_8930);
nand U9559 (N_9559,N_8425,N_8839);
nand U9560 (N_9560,N_8822,N_8635);
or U9561 (N_9561,N_8504,N_8822);
and U9562 (N_9562,N_8455,N_8912);
nor U9563 (N_9563,N_8961,N_8789);
nand U9564 (N_9564,N_8899,N_8622);
xor U9565 (N_9565,N_8746,N_8673);
or U9566 (N_9566,N_8715,N_8528);
and U9567 (N_9567,N_8909,N_8995);
and U9568 (N_9568,N_8957,N_8478);
and U9569 (N_9569,N_8650,N_8765);
and U9570 (N_9570,N_8898,N_8692);
or U9571 (N_9571,N_8977,N_8862);
nor U9572 (N_9572,N_8656,N_8615);
or U9573 (N_9573,N_8453,N_8729);
nand U9574 (N_9574,N_8594,N_8611);
or U9575 (N_9575,N_8733,N_8558);
xnor U9576 (N_9576,N_8408,N_8806);
nor U9577 (N_9577,N_8459,N_8948);
nor U9578 (N_9578,N_8615,N_8706);
nand U9579 (N_9579,N_8510,N_8996);
or U9580 (N_9580,N_8506,N_8454);
nor U9581 (N_9581,N_8850,N_8769);
xor U9582 (N_9582,N_8408,N_8895);
or U9583 (N_9583,N_8765,N_8642);
nor U9584 (N_9584,N_8551,N_8741);
xnor U9585 (N_9585,N_8425,N_8713);
or U9586 (N_9586,N_8510,N_8705);
and U9587 (N_9587,N_8813,N_8976);
or U9588 (N_9588,N_8871,N_8733);
nor U9589 (N_9589,N_8587,N_8729);
nor U9590 (N_9590,N_8978,N_8837);
nand U9591 (N_9591,N_8638,N_8795);
nand U9592 (N_9592,N_8740,N_8964);
nor U9593 (N_9593,N_8596,N_8859);
nand U9594 (N_9594,N_8447,N_8752);
nand U9595 (N_9595,N_8515,N_8521);
and U9596 (N_9596,N_8946,N_8803);
nand U9597 (N_9597,N_8873,N_8926);
and U9598 (N_9598,N_8431,N_8700);
xor U9599 (N_9599,N_8653,N_8479);
and U9600 (N_9600,N_9371,N_9157);
nand U9601 (N_9601,N_9067,N_9322);
and U9602 (N_9602,N_9253,N_9425);
nand U9603 (N_9603,N_9208,N_9321);
nor U9604 (N_9604,N_9451,N_9180);
nor U9605 (N_9605,N_9367,N_9364);
xnor U9606 (N_9606,N_9350,N_9158);
nor U9607 (N_9607,N_9375,N_9143);
and U9608 (N_9608,N_9230,N_9051);
nor U9609 (N_9609,N_9217,N_9521);
nand U9610 (N_9610,N_9564,N_9196);
or U9611 (N_9611,N_9565,N_9049);
xnor U9612 (N_9612,N_9290,N_9133);
or U9613 (N_9613,N_9060,N_9566);
nor U9614 (N_9614,N_9282,N_9235);
nor U9615 (N_9615,N_9291,N_9265);
or U9616 (N_9616,N_9188,N_9463);
or U9617 (N_9617,N_9512,N_9091);
xnor U9618 (N_9618,N_9190,N_9439);
and U9619 (N_9619,N_9119,N_9095);
nor U9620 (N_9620,N_9129,N_9457);
nor U9621 (N_9621,N_9433,N_9058);
and U9622 (N_9622,N_9094,N_9527);
nand U9623 (N_9623,N_9422,N_9132);
and U9624 (N_9624,N_9387,N_9427);
and U9625 (N_9625,N_9456,N_9223);
nor U9626 (N_9626,N_9488,N_9168);
or U9627 (N_9627,N_9281,N_9563);
or U9628 (N_9628,N_9409,N_9096);
xor U9629 (N_9629,N_9324,N_9345);
or U9630 (N_9630,N_9428,N_9495);
xor U9631 (N_9631,N_9373,N_9480);
and U9632 (N_9632,N_9105,N_9330);
or U9633 (N_9633,N_9030,N_9502);
and U9634 (N_9634,N_9340,N_9474);
nand U9635 (N_9635,N_9165,N_9070);
and U9636 (N_9636,N_9013,N_9469);
or U9637 (N_9637,N_9580,N_9591);
or U9638 (N_9638,N_9156,N_9336);
or U9639 (N_9639,N_9500,N_9264);
xor U9640 (N_9640,N_9307,N_9108);
and U9641 (N_9641,N_9558,N_9396);
xor U9642 (N_9642,N_9528,N_9333);
xnor U9643 (N_9643,N_9314,N_9526);
xnor U9644 (N_9644,N_9161,N_9532);
and U9645 (N_9645,N_9525,N_9538);
nor U9646 (N_9646,N_9582,N_9115);
and U9647 (N_9647,N_9139,N_9550);
xnor U9648 (N_9648,N_9596,N_9019);
xor U9649 (N_9649,N_9034,N_9455);
and U9650 (N_9650,N_9209,N_9297);
and U9651 (N_9651,N_9032,N_9093);
nand U9652 (N_9652,N_9244,N_9412);
nand U9653 (N_9653,N_9250,N_9181);
and U9654 (N_9654,N_9213,N_9357);
and U9655 (N_9655,N_9126,N_9381);
nor U9656 (N_9656,N_9516,N_9329);
or U9657 (N_9657,N_9179,N_9518);
nor U9658 (N_9658,N_9255,N_9256);
xnor U9659 (N_9659,N_9072,N_9420);
and U9660 (N_9660,N_9355,N_9319);
and U9661 (N_9661,N_9260,N_9379);
nand U9662 (N_9662,N_9182,N_9449);
nand U9663 (N_9663,N_9258,N_9514);
and U9664 (N_9664,N_9542,N_9189);
and U9665 (N_9665,N_9413,N_9028);
nor U9666 (N_9666,N_9083,N_9548);
and U9667 (N_9667,N_9234,N_9112);
nor U9668 (N_9668,N_9193,N_9205);
or U9669 (N_9669,N_9224,N_9577);
or U9670 (N_9670,N_9372,N_9218);
or U9671 (N_9671,N_9537,N_9426);
nor U9672 (N_9672,N_9464,N_9530);
or U9673 (N_9673,N_9517,N_9245);
or U9674 (N_9674,N_9394,N_9277);
and U9675 (N_9675,N_9210,N_9098);
and U9676 (N_9676,N_9380,N_9559);
nand U9677 (N_9677,N_9082,N_9087);
xor U9678 (N_9678,N_9454,N_9164);
and U9679 (N_9679,N_9266,N_9077);
or U9680 (N_9680,N_9339,N_9276);
or U9681 (N_9681,N_9207,N_9254);
or U9682 (N_9682,N_9041,N_9232);
nand U9683 (N_9683,N_9391,N_9279);
nor U9684 (N_9684,N_9239,N_9274);
nor U9685 (N_9685,N_9448,N_9405);
or U9686 (N_9686,N_9555,N_9149);
nand U9687 (N_9687,N_9216,N_9511);
nor U9688 (N_9688,N_9174,N_9150);
or U9689 (N_9689,N_9233,N_9313);
xnor U9690 (N_9690,N_9036,N_9088);
nor U9691 (N_9691,N_9163,N_9572);
nor U9692 (N_9692,N_9106,N_9482);
or U9693 (N_9693,N_9261,N_9348);
and U9694 (N_9694,N_9403,N_9344);
or U9695 (N_9695,N_9444,N_9320);
nor U9696 (N_9696,N_9199,N_9465);
nor U9697 (N_9697,N_9491,N_9300);
or U9698 (N_9698,N_9392,N_9560);
and U9699 (N_9699,N_9123,N_9026);
and U9700 (N_9700,N_9222,N_9323);
nor U9701 (N_9701,N_9368,N_9011);
and U9702 (N_9702,N_9192,N_9583);
and U9703 (N_9703,N_9039,N_9584);
and U9704 (N_9704,N_9442,N_9236);
and U9705 (N_9705,N_9069,N_9153);
or U9706 (N_9706,N_9038,N_9268);
nand U9707 (N_9707,N_9318,N_9298);
nand U9708 (N_9708,N_9206,N_9001);
nor U9709 (N_9709,N_9186,N_9354);
or U9710 (N_9710,N_9021,N_9315);
or U9711 (N_9711,N_9401,N_9508);
or U9712 (N_9712,N_9554,N_9309);
or U9713 (N_9713,N_9341,N_9148);
or U9714 (N_9714,N_9490,N_9086);
nand U9715 (N_9715,N_9599,N_9466);
or U9716 (N_9716,N_9018,N_9306);
nor U9717 (N_9717,N_9184,N_9289);
and U9718 (N_9718,N_9346,N_9044);
nor U9719 (N_9719,N_9598,N_9046);
or U9720 (N_9720,N_9238,N_9293);
xor U9721 (N_9721,N_9472,N_9073);
or U9722 (N_9722,N_9140,N_9513);
and U9723 (N_9723,N_9185,N_9269);
xnor U9724 (N_9724,N_9022,N_9204);
or U9725 (N_9725,N_9576,N_9332);
nor U9726 (N_9726,N_9589,N_9361);
nor U9727 (N_9727,N_9562,N_9316);
or U9728 (N_9728,N_9399,N_9534);
nand U9729 (N_9729,N_9195,N_9221);
and U9730 (N_9730,N_9014,N_9540);
xnor U9731 (N_9731,N_9460,N_9178);
and U9732 (N_9732,N_9203,N_9556);
and U9733 (N_9733,N_9492,N_9363);
nand U9734 (N_9734,N_9522,N_9101);
or U9735 (N_9735,N_9327,N_9447);
and U9736 (N_9736,N_9549,N_9064);
nand U9737 (N_9737,N_9202,N_9510);
and U9738 (N_9738,N_9118,N_9066);
and U9739 (N_9739,N_9107,N_9012);
or U9740 (N_9740,N_9506,N_9225);
nor U9741 (N_9741,N_9169,N_9025);
or U9742 (N_9742,N_9334,N_9446);
and U9743 (N_9743,N_9097,N_9587);
xor U9744 (N_9744,N_9220,N_9331);
or U9745 (N_9745,N_9418,N_9027);
and U9746 (N_9746,N_9145,N_9287);
and U9747 (N_9747,N_9303,N_9588);
and U9748 (N_9748,N_9440,N_9084);
nand U9749 (N_9749,N_9481,N_9081);
or U9750 (N_9750,N_9535,N_9138);
nor U9751 (N_9751,N_9541,N_9503);
or U9752 (N_9752,N_9191,N_9231);
nor U9753 (N_9753,N_9365,N_9103);
nor U9754 (N_9754,N_9408,N_9068);
and U9755 (N_9755,N_9214,N_9187);
nand U9756 (N_9756,N_9407,N_9023);
nand U9757 (N_9757,N_9419,N_9008);
and U9758 (N_9758,N_9043,N_9384);
xnor U9759 (N_9759,N_9015,N_9317);
nor U9760 (N_9760,N_9438,N_9079);
nor U9761 (N_9761,N_9259,N_9047);
and U9762 (N_9762,N_9247,N_9100);
xor U9763 (N_9763,N_9507,N_9286);
or U9764 (N_9764,N_9369,N_9135);
nand U9765 (N_9765,N_9295,N_9531);
or U9766 (N_9766,N_9045,N_9383);
nand U9767 (N_9767,N_9414,N_9573);
and U9768 (N_9768,N_9246,N_9240);
nand U9769 (N_9769,N_9519,N_9048);
or U9770 (N_9770,N_9593,N_9104);
and U9771 (N_9771,N_9486,N_9003);
or U9772 (N_9772,N_9062,N_9342);
xnor U9773 (N_9773,N_9410,N_9547);
nor U9774 (N_9774,N_9142,N_9592);
and U9775 (N_9775,N_9347,N_9056);
nand U9776 (N_9776,N_9505,N_9544);
or U9777 (N_9777,N_9243,N_9567);
nand U9778 (N_9778,N_9523,N_9360);
nand U9779 (N_9779,N_9586,N_9552);
xnor U9780 (N_9780,N_9393,N_9476);
xnor U9781 (N_9781,N_9524,N_9176);
xor U9782 (N_9782,N_9198,N_9432);
nand U9783 (N_9783,N_9325,N_9128);
and U9784 (N_9784,N_9078,N_9037);
or U9785 (N_9785,N_9160,N_9151);
and U9786 (N_9786,N_9125,N_9421);
or U9787 (N_9787,N_9292,N_9484);
and U9788 (N_9788,N_9557,N_9194);
or U9789 (N_9789,N_9183,N_9053);
nand U9790 (N_9790,N_9390,N_9571);
xnor U9791 (N_9791,N_9121,N_9000);
or U9792 (N_9792,N_9400,N_9351);
xnor U9793 (N_9793,N_9366,N_9594);
or U9794 (N_9794,N_9111,N_9595);
xor U9795 (N_9795,N_9052,N_9228);
nor U9796 (N_9796,N_9388,N_9109);
xor U9797 (N_9797,N_9029,N_9002);
and U9798 (N_9798,N_9461,N_9114);
nor U9799 (N_9799,N_9061,N_9010);
or U9800 (N_9800,N_9152,N_9515);
nor U9801 (N_9801,N_9501,N_9326);
nor U9802 (N_9802,N_9411,N_9127);
or U9803 (N_9803,N_9569,N_9120);
nand U9804 (N_9804,N_9561,N_9483);
or U9805 (N_9805,N_9270,N_9020);
or U9806 (N_9806,N_9494,N_9374);
or U9807 (N_9807,N_9434,N_9497);
and U9808 (N_9808,N_9075,N_9050);
and U9809 (N_9809,N_9074,N_9251);
nor U9810 (N_9810,N_9172,N_9417);
or U9811 (N_9811,N_9578,N_9533);
nor U9812 (N_9812,N_9443,N_9288);
nor U9813 (N_9813,N_9136,N_9404);
xor U9814 (N_9814,N_9402,N_9113);
or U9815 (N_9815,N_9590,N_9219);
or U9816 (N_9816,N_9200,N_9328);
and U9817 (N_9817,N_9280,N_9478);
or U9818 (N_9818,N_9241,N_9271);
xnor U9819 (N_9819,N_9147,N_9445);
xor U9820 (N_9820,N_9141,N_9035);
xor U9821 (N_9821,N_9489,N_9585);
and U9822 (N_9822,N_9257,N_9435);
nor U9823 (N_9823,N_9033,N_9509);
xnor U9824 (N_9824,N_9337,N_9175);
nor U9825 (N_9825,N_9273,N_9071);
or U9826 (N_9826,N_9487,N_9272);
xnor U9827 (N_9827,N_9376,N_9252);
nor U9828 (N_9828,N_9579,N_9424);
nand U9829 (N_9829,N_9197,N_9545);
nand U9830 (N_9830,N_9080,N_9177);
or U9831 (N_9831,N_9359,N_9470);
nand U9832 (N_9832,N_9263,N_9076);
nor U9833 (N_9833,N_9283,N_9006);
or U9834 (N_9834,N_9431,N_9016);
and U9835 (N_9835,N_9473,N_9301);
xor U9836 (N_9836,N_9310,N_9397);
and U9837 (N_9837,N_9459,N_9308);
nor U9838 (N_9838,N_9063,N_9146);
or U9839 (N_9839,N_9335,N_9134);
nor U9840 (N_9840,N_9275,N_9009);
or U9841 (N_9841,N_9406,N_9296);
or U9842 (N_9842,N_9551,N_9362);
xnor U9843 (N_9843,N_9597,N_9042);
nor U9844 (N_9844,N_9059,N_9574);
nand U9845 (N_9845,N_9430,N_9553);
or U9846 (N_9846,N_9004,N_9294);
and U9847 (N_9847,N_9570,N_9453);
and U9848 (N_9848,N_9437,N_9416);
or U9849 (N_9849,N_9475,N_9493);
and U9850 (N_9850,N_9154,N_9102);
nor U9851 (N_9851,N_9370,N_9499);
nor U9852 (N_9852,N_9415,N_9568);
nor U9853 (N_9853,N_9377,N_9458);
or U9854 (N_9854,N_9467,N_9159);
xnor U9855 (N_9855,N_9386,N_9130);
and U9856 (N_9856,N_9089,N_9356);
or U9857 (N_9857,N_9212,N_9429);
or U9858 (N_9858,N_9312,N_9005);
nand U9859 (N_9859,N_9055,N_9170);
and U9860 (N_9860,N_9278,N_9504);
or U9861 (N_9861,N_9144,N_9441);
nand U9862 (N_9862,N_9462,N_9520);
or U9863 (N_9863,N_9305,N_9352);
and U9864 (N_9864,N_9173,N_9378);
and U9865 (N_9865,N_9452,N_9358);
and U9866 (N_9866,N_9054,N_9284);
and U9867 (N_9867,N_9285,N_9017);
nand U9868 (N_9868,N_9385,N_9024);
nand U9869 (N_9869,N_9137,N_9226);
xor U9870 (N_9870,N_9299,N_9167);
xor U9871 (N_9871,N_9229,N_9131);
or U9872 (N_9872,N_9099,N_9110);
nor U9873 (N_9873,N_9304,N_9382);
xor U9874 (N_9874,N_9242,N_9581);
nor U9875 (N_9875,N_9468,N_9057);
xnor U9876 (N_9876,N_9543,N_9201);
nor U9877 (N_9877,N_9065,N_9302);
xnor U9878 (N_9878,N_9124,N_9031);
nor U9879 (N_9879,N_9007,N_9237);
nand U9880 (N_9880,N_9575,N_9117);
and U9881 (N_9881,N_9040,N_9485);
nor U9882 (N_9882,N_9436,N_9398);
and U9883 (N_9883,N_9248,N_9227);
or U9884 (N_9884,N_9479,N_9353);
nand U9885 (N_9885,N_9338,N_9349);
and U9886 (N_9886,N_9395,N_9211);
or U9887 (N_9887,N_9546,N_9166);
nor U9888 (N_9888,N_9343,N_9536);
or U9889 (N_9889,N_9155,N_9262);
nor U9890 (N_9890,N_9090,N_9267);
xnor U9891 (N_9891,N_9085,N_9498);
nor U9892 (N_9892,N_9389,N_9122);
nor U9893 (N_9893,N_9477,N_9450);
or U9894 (N_9894,N_9311,N_9471);
and U9895 (N_9895,N_9423,N_9092);
or U9896 (N_9896,N_9116,N_9529);
xnor U9897 (N_9897,N_9215,N_9539);
or U9898 (N_9898,N_9162,N_9171);
and U9899 (N_9899,N_9249,N_9496);
nor U9900 (N_9900,N_9250,N_9336);
xnor U9901 (N_9901,N_9495,N_9268);
nor U9902 (N_9902,N_9501,N_9108);
or U9903 (N_9903,N_9193,N_9543);
nor U9904 (N_9904,N_9388,N_9125);
xnor U9905 (N_9905,N_9046,N_9192);
xor U9906 (N_9906,N_9573,N_9188);
nand U9907 (N_9907,N_9226,N_9473);
xnor U9908 (N_9908,N_9591,N_9047);
nor U9909 (N_9909,N_9243,N_9164);
nor U9910 (N_9910,N_9572,N_9327);
or U9911 (N_9911,N_9425,N_9022);
nand U9912 (N_9912,N_9158,N_9529);
and U9913 (N_9913,N_9412,N_9438);
xor U9914 (N_9914,N_9300,N_9258);
nand U9915 (N_9915,N_9491,N_9025);
and U9916 (N_9916,N_9456,N_9328);
or U9917 (N_9917,N_9540,N_9446);
and U9918 (N_9918,N_9533,N_9493);
xnor U9919 (N_9919,N_9564,N_9073);
nand U9920 (N_9920,N_9484,N_9423);
and U9921 (N_9921,N_9011,N_9049);
xor U9922 (N_9922,N_9444,N_9016);
xor U9923 (N_9923,N_9104,N_9235);
nand U9924 (N_9924,N_9422,N_9144);
or U9925 (N_9925,N_9422,N_9547);
and U9926 (N_9926,N_9001,N_9398);
xor U9927 (N_9927,N_9141,N_9180);
or U9928 (N_9928,N_9399,N_9218);
and U9929 (N_9929,N_9142,N_9025);
or U9930 (N_9930,N_9363,N_9553);
or U9931 (N_9931,N_9591,N_9303);
nor U9932 (N_9932,N_9300,N_9117);
nor U9933 (N_9933,N_9106,N_9049);
nand U9934 (N_9934,N_9524,N_9445);
nand U9935 (N_9935,N_9453,N_9053);
or U9936 (N_9936,N_9349,N_9165);
or U9937 (N_9937,N_9448,N_9087);
or U9938 (N_9938,N_9517,N_9066);
and U9939 (N_9939,N_9360,N_9043);
nand U9940 (N_9940,N_9374,N_9336);
nand U9941 (N_9941,N_9584,N_9184);
xnor U9942 (N_9942,N_9462,N_9304);
or U9943 (N_9943,N_9105,N_9082);
or U9944 (N_9944,N_9131,N_9279);
or U9945 (N_9945,N_9161,N_9577);
nor U9946 (N_9946,N_9495,N_9213);
nor U9947 (N_9947,N_9041,N_9495);
xnor U9948 (N_9948,N_9538,N_9579);
nand U9949 (N_9949,N_9166,N_9549);
nor U9950 (N_9950,N_9008,N_9517);
xnor U9951 (N_9951,N_9229,N_9474);
nor U9952 (N_9952,N_9041,N_9310);
and U9953 (N_9953,N_9586,N_9015);
and U9954 (N_9954,N_9020,N_9062);
xnor U9955 (N_9955,N_9565,N_9557);
and U9956 (N_9956,N_9023,N_9134);
xnor U9957 (N_9957,N_9365,N_9525);
nand U9958 (N_9958,N_9590,N_9160);
nand U9959 (N_9959,N_9090,N_9332);
or U9960 (N_9960,N_9332,N_9273);
or U9961 (N_9961,N_9379,N_9286);
and U9962 (N_9962,N_9305,N_9569);
and U9963 (N_9963,N_9061,N_9544);
xnor U9964 (N_9964,N_9187,N_9563);
and U9965 (N_9965,N_9310,N_9429);
xnor U9966 (N_9966,N_9143,N_9519);
and U9967 (N_9967,N_9206,N_9568);
and U9968 (N_9968,N_9043,N_9548);
nor U9969 (N_9969,N_9365,N_9564);
xnor U9970 (N_9970,N_9270,N_9234);
and U9971 (N_9971,N_9454,N_9422);
xnor U9972 (N_9972,N_9572,N_9537);
nand U9973 (N_9973,N_9151,N_9010);
and U9974 (N_9974,N_9582,N_9272);
xnor U9975 (N_9975,N_9357,N_9405);
or U9976 (N_9976,N_9245,N_9564);
nor U9977 (N_9977,N_9302,N_9316);
or U9978 (N_9978,N_9004,N_9342);
nand U9979 (N_9979,N_9225,N_9249);
xor U9980 (N_9980,N_9563,N_9073);
xor U9981 (N_9981,N_9049,N_9393);
or U9982 (N_9982,N_9018,N_9586);
or U9983 (N_9983,N_9298,N_9014);
xor U9984 (N_9984,N_9098,N_9530);
or U9985 (N_9985,N_9188,N_9385);
and U9986 (N_9986,N_9247,N_9308);
and U9987 (N_9987,N_9158,N_9443);
nand U9988 (N_9988,N_9517,N_9130);
or U9989 (N_9989,N_9182,N_9492);
xor U9990 (N_9990,N_9305,N_9582);
or U9991 (N_9991,N_9569,N_9441);
xor U9992 (N_9992,N_9546,N_9354);
nand U9993 (N_9993,N_9116,N_9521);
nand U9994 (N_9994,N_9169,N_9487);
or U9995 (N_9995,N_9072,N_9427);
nand U9996 (N_9996,N_9377,N_9484);
nor U9997 (N_9997,N_9026,N_9495);
and U9998 (N_9998,N_9462,N_9394);
nor U9999 (N_9999,N_9113,N_9279);
nand U10000 (N_10000,N_9456,N_9351);
nor U10001 (N_10001,N_9172,N_9094);
and U10002 (N_10002,N_9226,N_9383);
or U10003 (N_10003,N_9557,N_9125);
nor U10004 (N_10004,N_9143,N_9283);
or U10005 (N_10005,N_9479,N_9541);
nor U10006 (N_10006,N_9126,N_9471);
nor U10007 (N_10007,N_9543,N_9264);
nand U10008 (N_10008,N_9310,N_9444);
nand U10009 (N_10009,N_9418,N_9458);
nor U10010 (N_10010,N_9356,N_9483);
xor U10011 (N_10011,N_9397,N_9151);
or U10012 (N_10012,N_9297,N_9262);
and U10013 (N_10013,N_9222,N_9263);
nor U10014 (N_10014,N_9011,N_9072);
and U10015 (N_10015,N_9337,N_9073);
nand U10016 (N_10016,N_9094,N_9447);
xnor U10017 (N_10017,N_9076,N_9420);
nor U10018 (N_10018,N_9544,N_9376);
or U10019 (N_10019,N_9488,N_9443);
nor U10020 (N_10020,N_9055,N_9586);
nor U10021 (N_10021,N_9321,N_9095);
and U10022 (N_10022,N_9090,N_9067);
xor U10023 (N_10023,N_9080,N_9595);
and U10024 (N_10024,N_9167,N_9529);
and U10025 (N_10025,N_9073,N_9449);
xor U10026 (N_10026,N_9581,N_9534);
and U10027 (N_10027,N_9285,N_9389);
xnor U10028 (N_10028,N_9537,N_9164);
nor U10029 (N_10029,N_9156,N_9154);
and U10030 (N_10030,N_9135,N_9180);
and U10031 (N_10031,N_9165,N_9407);
nor U10032 (N_10032,N_9515,N_9518);
and U10033 (N_10033,N_9047,N_9375);
xnor U10034 (N_10034,N_9336,N_9137);
and U10035 (N_10035,N_9549,N_9181);
or U10036 (N_10036,N_9558,N_9492);
nand U10037 (N_10037,N_9528,N_9136);
nand U10038 (N_10038,N_9126,N_9498);
or U10039 (N_10039,N_9156,N_9171);
nor U10040 (N_10040,N_9090,N_9317);
xor U10041 (N_10041,N_9304,N_9587);
nor U10042 (N_10042,N_9484,N_9280);
and U10043 (N_10043,N_9218,N_9151);
xor U10044 (N_10044,N_9416,N_9188);
nand U10045 (N_10045,N_9527,N_9277);
xnor U10046 (N_10046,N_9202,N_9274);
nand U10047 (N_10047,N_9361,N_9417);
or U10048 (N_10048,N_9472,N_9429);
or U10049 (N_10049,N_9405,N_9181);
xor U10050 (N_10050,N_9431,N_9049);
nand U10051 (N_10051,N_9398,N_9135);
and U10052 (N_10052,N_9196,N_9589);
or U10053 (N_10053,N_9528,N_9367);
or U10054 (N_10054,N_9107,N_9598);
nor U10055 (N_10055,N_9251,N_9086);
and U10056 (N_10056,N_9444,N_9373);
and U10057 (N_10057,N_9026,N_9130);
or U10058 (N_10058,N_9546,N_9243);
and U10059 (N_10059,N_9432,N_9457);
nor U10060 (N_10060,N_9427,N_9215);
nor U10061 (N_10061,N_9219,N_9530);
and U10062 (N_10062,N_9324,N_9465);
xor U10063 (N_10063,N_9215,N_9134);
and U10064 (N_10064,N_9380,N_9087);
nor U10065 (N_10065,N_9348,N_9561);
and U10066 (N_10066,N_9105,N_9362);
xor U10067 (N_10067,N_9010,N_9482);
nand U10068 (N_10068,N_9231,N_9249);
and U10069 (N_10069,N_9035,N_9066);
xnor U10070 (N_10070,N_9525,N_9058);
nand U10071 (N_10071,N_9401,N_9224);
nor U10072 (N_10072,N_9233,N_9113);
or U10073 (N_10073,N_9517,N_9430);
or U10074 (N_10074,N_9503,N_9355);
xnor U10075 (N_10075,N_9226,N_9546);
nor U10076 (N_10076,N_9466,N_9242);
or U10077 (N_10077,N_9007,N_9335);
xor U10078 (N_10078,N_9230,N_9046);
nor U10079 (N_10079,N_9598,N_9526);
nand U10080 (N_10080,N_9282,N_9530);
nor U10081 (N_10081,N_9501,N_9010);
or U10082 (N_10082,N_9270,N_9432);
xnor U10083 (N_10083,N_9377,N_9072);
nand U10084 (N_10084,N_9533,N_9580);
or U10085 (N_10085,N_9095,N_9092);
and U10086 (N_10086,N_9110,N_9561);
or U10087 (N_10087,N_9122,N_9549);
xor U10088 (N_10088,N_9091,N_9429);
nand U10089 (N_10089,N_9030,N_9146);
xnor U10090 (N_10090,N_9096,N_9147);
and U10091 (N_10091,N_9046,N_9287);
and U10092 (N_10092,N_9580,N_9391);
or U10093 (N_10093,N_9332,N_9027);
nand U10094 (N_10094,N_9414,N_9400);
and U10095 (N_10095,N_9512,N_9150);
nand U10096 (N_10096,N_9557,N_9302);
nand U10097 (N_10097,N_9581,N_9044);
nor U10098 (N_10098,N_9365,N_9069);
and U10099 (N_10099,N_9147,N_9274);
xor U10100 (N_10100,N_9367,N_9464);
and U10101 (N_10101,N_9302,N_9304);
or U10102 (N_10102,N_9489,N_9526);
or U10103 (N_10103,N_9511,N_9457);
nor U10104 (N_10104,N_9567,N_9131);
and U10105 (N_10105,N_9176,N_9194);
or U10106 (N_10106,N_9414,N_9577);
nor U10107 (N_10107,N_9313,N_9536);
nor U10108 (N_10108,N_9034,N_9137);
or U10109 (N_10109,N_9048,N_9450);
and U10110 (N_10110,N_9107,N_9064);
nor U10111 (N_10111,N_9101,N_9355);
nand U10112 (N_10112,N_9192,N_9373);
xnor U10113 (N_10113,N_9007,N_9384);
xnor U10114 (N_10114,N_9399,N_9438);
or U10115 (N_10115,N_9108,N_9515);
xor U10116 (N_10116,N_9327,N_9156);
and U10117 (N_10117,N_9145,N_9040);
nor U10118 (N_10118,N_9484,N_9329);
or U10119 (N_10119,N_9147,N_9543);
nor U10120 (N_10120,N_9061,N_9114);
xnor U10121 (N_10121,N_9455,N_9147);
nor U10122 (N_10122,N_9547,N_9307);
and U10123 (N_10123,N_9561,N_9518);
xnor U10124 (N_10124,N_9402,N_9355);
or U10125 (N_10125,N_9356,N_9017);
and U10126 (N_10126,N_9042,N_9093);
nor U10127 (N_10127,N_9076,N_9060);
xnor U10128 (N_10128,N_9200,N_9544);
or U10129 (N_10129,N_9052,N_9560);
nor U10130 (N_10130,N_9254,N_9431);
nor U10131 (N_10131,N_9263,N_9038);
or U10132 (N_10132,N_9508,N_9355);
xor U10133 (N_10133,N_9217,N_9234);
nand U10134 (N_10134,N_9039,N_9410);
or U10135 (N_10135,N_9321,N_9273);
xor U10136 (N_10136,N_9200,N_9421);
nand U10137 (N_10137,N_9209,N_9292);
nor U10138 (N_10138,N_9057,N_9214);
nand U10139 (N_10139,N_9542,N_9257);
or U10140 (N_10140,N_9472,N_9177);
nand U10141 (N_10141,N_9039,N_9304);
nor U10142 (N_10142,N_9375,N_9247);
nand U10143 (N_10143,N_9144,N_9093);
or U10144 (N_10144,N_9102,N_9070);
and U10145 (N_10145,N_9565,N_9448);
nand U10146 (N_10146,N_9384,N_9311);
xnor U10147 (N_10147,N_9478,N_9039);
or U10148 (N_10148,N_9211,N_9274);
nor U10149 (N_10149,N_9182,N_9177);
and U10150 (N_10150,N_9103,N_9461);
nand U10151 (N_10151,N_9312,N_9390);
nor U10152 (N_10152,N_9082,N_9451);
nand U10153 (N_10153,N_9050,N_9543);
nand U10154 (N_10154,N_9086,N_9384);
nand U10155 (N_10155,N_9441,N_9247);
xor U10156 (N_10156,N_9384,N_9021);
nor U10157 (N_10157,N_9504,N_9075);
and U10158 (N_10158,N_9048,N_9357);
nand U10159 (N_10159,N_9339,N_9448);
and U10160 (N_10160,N_9511,N_9589);
or U10161 (N_10161,N_9410,N_9512);
nor U10162 (N_10162,N_9150,N_9161);
or U10163 (N_10163,N_9165,N_9468);
nand U10164 (N_10164,N_9362,N_9544);
nor U10165 (N_10165,N_9349,N_9476);
nand U10166 (N_10166,N_9359,N_9585);
nor U10167 (N_10167,N_9108,N_9124);
or U10168 (N_10168,N_9239,N_9540);
nor U10169 (N_10169,N_9557,N_9532);
or U10170 (N_10170,N_9143,N_9229);
nor U10171 (N_10171,N_9182,N_9469);
and U10172 (N_10172,N_9335,N_9451);
nand U10173 (N_10173,N_9257,N_9081);
and U10174 (N_10174,N_9284,N_9203);
nor U10175 (N_10175,N_9391,N_9200);
nor U10176 (N_10176,N_9286,N_9162);
nand U10177 (N_10177,N_9493,N_9398);
nand U10178 (N_10178,N_9530,N_9075);
and U10179 (N_10179,N_9205,N_9100);
or U10180 (N_10180,N_9508,N_9316);
nand U10181 (N_10181,N_9424,N_9450);
and U10182 (N_10182,N_9282,N_9115);
and U10183 (N_10183,N_9292,N_9568);
nor U10184 (N_10184,N_9001,N_9566);
nand U10185 (N_10185,N_9093,N_9366);
and U10186 (N_10186,N_9416,N_9135);
or U10187 (N_10187,N_9016,N_9138);
xor U10188 (N_10188,N_9105,N_9156);
nor U10189 (N_10189,N_9465,N_9564);
nor U10190 (N_10190,N_9317,N_9501);
and U10191 (N_10191,N_9142,N_9037);
or U10192 (N_10192,N_9012,N_9346);
and U10193 (N_10193,N_9079,N_9172);
xor U10194 (N_10194,N_9257,N_9276);
nor U10195 (N_10195,N_9203,N_9283);
xnor U10196 (N_10196,N_9095,N_9500);
nor U10197 (N_10197,N_9099,N_9574);
or U10198 (N_10198,N_9371,N_9403);
xnor U10199 (N_10199,N_9527,N_9238);
or U10200 (N_10200,N_9999,N_10099);
nor U10201 (N_10201,N_10186,N_10010);
and U10202 (N_10202,N_9762,N_10123);
or U10203 (N_10203,N_9867,N_10125);
nand U10204 (N_10204,N_10004,N_10030);
or U10205 (N_10205,N_9986,N_9754);
or U10206 (N_10206,N_9953,N_10115);
nand U10207 (N_10207,N_9991,N_9615);
nand U10208 (N_10208,N_9657,N_9702);
or U10209 (N_10209,N_10046,N_9653);
xnor U10210 (N_10210,N_9695,N_9707);
nand U10211 (N_10211,N_9641,N_10053);
nand U10212 (N_10212,N_9728,N_10174);
and U10213 (N_10213,N_9870,N_10071);
and U10214 (N_10214,N_10027,N_9771);
or U10215 (N_10215,N_10088,N_10130);
and U10216 (N_10216,N_9611,N_10181);
nor U10217 (N_10217,N_10137,N_9763);
or U10218 (N_10218,N_9995,N_10034);
and U10219 (N_10219,N_9909,N_10145);
or U10220 (N_10220,N_9791,N_9978);
xnor U10221 (N_10221,N_9673,N_9877);
nand U10222 (N_10222,N_9946,N_9988);
nand U10223 (N_10223,N_9891,N_10043);
or U10224 (N_10224,N_9785,N_9942);
nand U10225 (N_10225,N_10126,N_9983);
nor U10226 (N_10226,N_9747,N_9745);
nor U10227 (N_10227,N_9677,N_9955);
nor U10228 (N_10228,N_9948,N_9743);
xnor U10229 (N_10229,N_9619,N_9742);
or U10230 (N_10230,N_10074,N_9820);
xor U10231 (N_10231,N_10122,N_10169);
and U10232 (N_10232,N_10073,N_10078);
nand U10233 (N_10233,N_10159,N_10166);
nand U10234 (N_10234,N_9956,N_9694);
and U10235 (N_10235,N_10149,N_9700);
nand U10236 (N_10236,N_9618,N_9947);
and U10237 (N_10237,N_10023,N_9902);
nor U10238 (N_10238,N_9847,N_10033);
nor U10239 (N_10239,N_10035,N_10037);
nand U10240 (N_10240,N_9784,N_9913);
xor U10241 (N_10241,N_9976,N_10119);
nand U10242 (N_10242,N_9622,N_10013);
nand U10243 (N_10243,N_9683,N_9912);
nand U10244 (N_10244,N_10050,N_10170);
and U10245 (N_10245,N_9688,N_9701);
or U10246 (N_10246,N_9964,N_9860);
nand U10247 (N_10247,N_10146,N_9923);
nand U10248 (N_10248,N_9925,N_10049);
xor U10249 (N_10249,N_10070,N_9984);
or U10250 (N_10250,N_9646,N_9765);
xnor U10251 (N_10251,N_9918,N_9776);
nor U10252 (N_10252,N_10029,N_9645);
nor U10253 (N_10253,N_9853,N_10048);
xnor U10254 (N_10254,N_10045,N_9890);
nand U10255 (N_10255,N_10185,N_9932);
xnor U10256 (N_10256,N_9644,N_10000);
nor U10257 (N_10257,N_10082,N_9778);
and U10258 (N_10258,N_9604,N_10132);
nor U10259 (N_10259,N_9746,N_10002);
nor U10260 (N_10260,N_10171,N_9719);
nor U10261 (N_10261,N_10183,N_9715);
nand U10262 (N_10262,N_9655,N_9665);
nor U10263 (N_10263,N_9833,N_10114);
or U10264 (N_10264,N_9864,N_9687);
and U10265 (N_10265,N_9669,N_10190);
xnor U10266 (N_10266,N_10117,N_9726);
xor U10267 (N_10267,N_9748,N_9672);
or U10268 (N_10268,N_10124,N_10144);
nor U10269 (N_10269,N_9607,N_10005);
or U10270 (N_10270,N_9717,N_9872);
nor U10271 (N_10271,N_9836,N_10022);
and U10272 (N_10272,N_10152,N_9731);
nand U10273 (N_10273,N_10129,N_10176);
and U10274 (N_10274,N_9710,N_9910);
xor U10275 (N_10275,N_9713,N_9940);
xnor U10276 (N_10276,N_9711,N_9917);
or U10277 (N_10277,N_10069,N_9620);
and U10278 (N_10278,N_10109,N_9967);
nor U10279 (N_10279,N_9623,N_10032);
and U10280 (N_10280,N_9671,N_9851);
nand U10281 (N_10281,N_9679,N_10014);
nor U10282 (N_10282,N_9834,N_9662);
nand U10283 (N_10283,N_10056,N_9608);
nand U10284 (N_10284,N_9706,N_9682);
xnor U10285 (N_10285,N_10020,N_9767);
nand U10286 (N_10286,N_10095,N_9812);
and U10287 (N_10287,N_9996,N_9843);
nand U10288 (N_10288,N_10127,N_9854);
nor U10289 (N_10289,N_10128,N_9613);
nand U10290 (N_10290,N_9642,N_10160);
and U10291 (N_10291,N_10135,N_9939);
nand U10292 (N_10292,N_9721,N_9831);
and U10293 (N_10293,N_9814,N_10021);
xor U10294 (N_10294,N_9862,N_10017);
nand U10295 (N_10295,N_9905,N_10012);
nand U10296 (N_10296,N_10092,N_9969);
nand U10297 (N_10297,N_9690,N_9806);
nor U10298 (N_10298,N_9732,N_9938);
nor U10299 (N_10299,N_10178,N_9749);
nor U10300 (N_10300,N_9633,N_10118);
nor U10301 (N_10301,N_9832,N_9884);
nand U10302 (N_10302,N_10041,N_9936);
nor U10303 (N_10303,N_9850,N_10194);
nor U10304 (N_10304,N_9761,N_9980);
nor U10305 (N_10305,N_9972,N_10085);
xor U10306 (N_10306,N_9739,N_9793);
xor U10307 (N_10307,N_9670,N_9603);
nor U10308 (N_10308,N_9827,N_9987);
xor U10309 (N_10309,N_9857,N_9626);
or U10310 (N_10310,N_9949,N_9686);
xnor U10311 (N_10311,N_10054,N_9954);
and U10312 (N_10312,N_9685,N_9751);
xnor U10313 (N_10313,N_10018,N_9977);
nand U10314 (N_10314,N_9807,N_10090);
nor U10315 (N_10315,N_9600,N_9933);
or U10316 (N_10316,N_9758,N_9930);
nand U10317 (N_10317,N_9926,N_10147);
nor U10318 (N_10318,N_10036,N_10162);
nand U10319 (N_10319,N_9922,N_9674);
xnor U10320 (N_10320,N_10155,N_9651);
xor U10321 (N_10321,N_10016,N_9893);
or U10322 (N_10322,N_10015,N_9759);
nor U10323 (N_10323,N_10062,N_10089);
nor U10324 (N_10324,N_9614,N_10184);
or U10325 (N_10325,N_9654,N_9656);
xnor U10326 (N_10326,N_9664,N_9703);
and U10327 (N_10327,N_10199,N_9801);
and U10328 (N_10328,N_10196,N_9965);
nor U10329 (N_10329,N_9681,N_9889);
nor U10330 (N_10330,N_9640,N_9735);
xor U10331 (N_10331,N_10047,N_9699);
nand U10332 (N_10332,N_10151,N_10042);
or U10333 (N_10333,N_9863,N_9628);
xor U10334 (N_10334,N_10094,N_9753);
and U10335 (N_10335,N_9680,N_10110);
xor U10336 (N_10336,N_9773,N_10121);
or U10337 (N_10337,N_9906,N_9770);
nand U10338 (N_10338,N_10133,N_9601);
nand U10339 (N_10339,N_9838,N_9734);
nor U10340 (N_10340,N_9738,N_9824);
nor U10341 (N_10341,N_10044,N_9835);
nor U10342 (N_10342,N_9868,N_9871);
nand U10343 (N_10343,N_9813,N_9904);
or U10344 (N_10344,N_10120,N_9704);
or U10345 (N_10345,N_9819,N_9632);
or U10346 (N_10346,N_9616,N_10108);
or U10347 (N_10347,N_9733,N_9612);
xor U10348 (N_10348,N_9795,N_9828);
nor U10349 (N_10349,N_10001,N_9896);
nor U10350 (N_10350,N_9606,N_9894);
nor U10351 (N_10351,N_9997,N_10028);
nor U10352 (N_10352,N_9783,N_9915);
nand U10353 (N_10353,N_9990,N_9937);
and U10354 (N_10354,N_10026,N_9941);
xor U10355 (N_10355,N_10076,N_9888);
xor U10356 (N_10356,N_9769,N_9823);
and U10357 (N_10357,N_9989,N_10038);
and U10358 (N_10358,N_9855,N_9944);
nor U10359 (N_10359,N_10091,N_9740);
nand U10360 (N_10360,N_9689,N_9709);
or U10361 (N_10361,N_9803,N_9667);
nand U10362 (N_10362,N_10058,N_9992);
nor U10363 (N_10363,N_9757,N_9798);
and U10364 (N_10364,N_10068,N_9817);
nor U10365 (N_10365,N_9708,N_9880);
and U10366 (N_10366,N_9919,N_9931);
or U10367 (N_10367,N_9729,N_9962);
nor U10368 (N_10368,N_10138,N_9609);
and U10369 (N_10369,N_9666,N_10142);
or U10370 (N_10370,N_9659,N_9705);
xnor U10371 (N_10371,N_9636,N_10154);
or U10372 (N_10372,N_10113,N_9974);
and U10373 (N_10373,N_9885,N_10143);
or U10374 (N_10374,N_10193,N_9970);
and U10375 (N_10375,N_9914,N_9876);
or U10376 (N_10376,N_10140,N_10087);
nand U10377 (N_10377,N_9994,N_9768);
xnor U10378 (N_10378,N_10009,N_10148);
nor U10379 (N_10379,N_10187,N_10191);
nor U10380 (N_10380,N_9892,N_10065);
or U10381 (N_10381,N_10051,N_9924);
and U10382 (N_10382,N_9796,N_9895);
and U10383 (N_10383,N_10075,N_9789);
nor U10384 (N_10384,N_9840,N_9998);
and U10385 (N_10385,N_10060,N_9822);
nand U10386 (N_10386,N_10189,N_9718);
and U10387 (N_10387,N_10116,N_10008);
or U10388 (N_10388,N_9693,N_9815);
nor U10389 (N_10389,N_9625,N_9637);
and U10390 (N_10390,N_9961,N_9934);
nor U10391 (N_10391,N_9774,N_9846);
and U10392 (N_10392,N_9816,N_9663);
nand U10393 (N_10393,N_9945,N_9966);
nor U10394 (N_10394,N_9802,N_10167);
nand U10395 (N_10395,N_10156,N_9951);
xnor U10396 (N_10396,N_10011,N_9777);
nand U10397 (N_10397,N_9805,N_9786);
nand U10398 (N_10398,N_10172,N_9883);
xnor U10399 (N_10399,N_10007,N_10072);
and U10400 (N_10400,N_9958,N_9869);
nor U10401 (N_10401,N_9874,N_9900);
and U10402 (N_10402,N_9764,N_9638);
or U10403 (N_10403,N_10102,N_9676);
xor U10404 (N_10404,N_10059,N_9714);
xor U10405 (N_10405,N_9908,N_9730);
nor U10406 (N_10406,N_10101,N_9993);
nand U10407 (N_10407,N_10024,N_10093);
xor U10408 (N_10408,N_10195,N_9650);
and U10409 (N_10409,N_10081,N_9775);
or U10410 (N_10410,N_9950,N_10019);
nand U10411 (N_10411,N_9856,N_9842);
and U10412 (N_10412,N_9920,N_10139);
nand U10413 (N_10413,N_9921,N_9848);
nor U10414 (N_10414,N_9903,N_9660);
nor U10415 (N_10415,N_9981,N_10107);
and U10416 (N_10416,N_9720,N_10103);
or U10417 (N_10417,N_9968,N_9865);
nand U10418 (N_10418,N_9652,N_9825);
or U10419 (N_10419,N_9643,N_9975);
xnor U10420 (N_10420,N_9692,N_9602);
and U10421 (N_10421,N_9875,N_9830);
nand U10422 (N_10422,N_9957,N_10141);
xnor U10423 (N_10423,N_10100,N_9878);
or U10424 (N_10424,N_10083,N_9627);
nand U10425 (N_10425,N_9866,N_9691);
xnor U10426 (N_10426,N_10084,N_9750);
nand U10427 (N_10427,N_9736,N_9724);
and U10428 (N_10428,N_9907,N_10006);
nand U10429 (N_10429,N_10173,N_9661);
and U10430 (N_10430,N_9799,N_9781);
nand U10431 (N_10431,N_10179,N_9755);
and U10432 (N_10432,N_10055,N_9723);
nand U10433 (N_10433,N_9697,N_10188);
xnor U10434 (N_10434,N_9772,N_10063);
xor U10435 (N_10435,N_9852,N_9861);
nand U10436 (N_10436,N_10066,N_9901);
and U10437 (N_10437,N_9752,N_9760);
xor U10438 (N_10438,N_9725,N_9911);
xor U10439 (N_10439,N_10077,N_10097);
and U10440 (N_10440,N_9826,N_10153);
and U10441 (N_10441,N_9675,N_9658);
and U10442 (N_10442,N_9624,N_9792);
xor U10443 (N_10443,N_9897,N_10040);
xor U10444 (N_10444,N_10112,N_9809);
xor U10445 (N_10445,N_9858,N_10061);
nor U10446 (N_10446,N_9886,N_9952);
xor U10447 (N_10447,N_9844,N_9737);
xor U10448 (N_10448,N_9678,N_10197);
nor U10449 (N_10449,N_9882,N_9716);
nor U10450 (N_10450,N_10098,N_9971);
xnor U10451 (N_10451,N_10163,N_9927);
nor U10452 (N_10452,N_10165,N_9979);
xor U10453 (N_10453,N_9722,N_9810);
nor U10454 (N_10454,N_9899,N_9788);
nand U10455 (N_10455,N_9963,N_9766);
and U10456 (N_10456,N_9727,N_9698);
xnor U10457 (N_10457,N_9605,N_9916);
or U10458 (N_10458,N_9782,N_9811);
or U10459 (N_10459,N_10150,N_10003);
xnor U10460 (N_10460,N_10079,N_9800);
or U10461 (N_10461,N_9982,N_9837);
or U10462 (N_10462,N_9849,N_9985);
and U10463 (N_10463,N_10086,N_9648);
xnor U10464 (N_10464,N_10039,N_10182);
nand U10465 (N_10465,N_9647,N_9780);
xnor U10466 (N_10466,N_9881,N_10131);
nor U10467 (N_10467,N_10175,N_9634);
and U10468 (N_10468,N_9943,N_9859);
and U10469 (N_10469,N_9617,N_10168);
and U10470 (N_10470,N_9610,N_10161);
and U10471 (N_10471,N_9756,N_9668);
xor U10472 (N_10472,N_9741,N_9898);
nand U10473 (N_10473,N_10105,N_9629);
or U10474 (N_10474,N_9841,N_10057);
or U10475 (N_10475,N_9649,N_9696);
or U10476 (N_10476,N_10106,N_10096);
nor U10477 (N_10477,N_9935,N_9808);
and U10478 (N_10478,N_10177,N_9960);
nor U10479 (N_10479,N_9712,N_9631);
and U10480 (N_10480,N_9635,N_9779);
and U10481 (N_10481,N_9804,N_10192);
nand U10482 (N_10482,N_9621,N_9821);
nor U10483 (N_10483,N_9818,N_9790);
or U10484 (N_10484,N_9845,N_9630);
xor U10485 (N_10485,N_10064,N_10164);
xnor U10486 (N_10486,N_9928,N_10198);
nor U10487 (N_10487,N_9787,N_10180);
nand U10488 (N_10488,N_9929,N_10157);
and U10489 (N_10489,N_9794,N_10104);
or U10490 (N_10490,N_10158,N_10080);
xor U10491 (N_10491,N_9797,N_9829);
and U10492 (N_10492,N_10134,N_10052);
xnor U10493 (N_10493,N_10111,N_9959);
xnor U10494 (N_10494,N_9873,N_10025);
or U10495 (N_10495,N_9839,N_9887);
and U10496 (N_10496,N_9973,N_10136);
xor U10497 (N_10497,N_10031,N_9744);
nand U10498 (N_10498,N_9684,N_9639);
and U10499 (N_10499,N_9879,N_10067);
and U10500 (N_10500,N_9948,N_10046);
nand U10501 (N_10501,N_10074,N_9926);
nand U10502 (N_10502,N_9731,N_9804);
and U10503 (N_10503,N_9936,N_9935);
and U10504 (N_10504,N_9984,N_10075);
xor U10505 (N_10505,N_9933,N_9886);
nor U10506 (N_10506,N_9631,N_9835);
nand U10507 (N_10507,N_9922,N_9853);
or U10508 (N_10508,N_10091,N_10121);
nand U10509 (N_10509,N_10019,N_9958);
or U10510 (N_10510,N_9773,N_9942);
nor U10511 (N_10511,N_9831,N_9619);
and U10512 (N_10512,N_9857,N_10068);
and U10513 (N_10513,N_10144,N_10197);
or U10514 (N_10514,N_9765,N_9687);
or U10515 (N_10515,N_9734,N_9972);
nand U10516 (N_10516,N_10000,N_9906);
and U10517 (N_10517,N_9673,N_9680);
xor U10518 (N_10518,N_9965,N_9933);
and U10519 (N_10519,N_9634,N_9704);
and U10520 (N_10520,N_9832,N_9673);
and U10521 (N_10521,N_9671,N_9693);
xor U10522 (N_10522,N_9618,N_9897);
nor U10523 (N_10523,N_10125,N_10190);
or U10524 (N_10524,N_9682,N_9720);
xor U10525 (N_10525,N_9749,N_9981);
nand U10526 (N_10526,N_9985,N_10179);
and U10527 (N_10527,N_9667,N_9925);
or U10528 (N_10528,N_9794,N_9602);
xor U10529 (N_10529,N_9959,N_10008);
or U10530 (N_10530,N_9622,N_10066);
xnor U10531 (N_10531,N_9681,N_9937);
and U10532 (N_10532,N_9625,N_9982);
and U10533 (N_10533,N_10037,N_9891);
xor U10534 (N_10534,N_10199,N_9835);
or U10535 (N_10535,N_9880,N_10076);
or U10536 (N_10536,N_9778,N_9794);
or U10537 (N_10537,N_9851,N_9873);
and U10538 (N_10538,N_9645,N_9975);
xnor U10539 (N_10539,N_9880,N_10140);
nor U10540 (N_10540,N_9971,N_9937);
and U10541 (N_10541,N_9822,N_9751);
and U10542 (N_10542,N_9716,N_9824);
nor U10543 (N_10543,N_9864,N_9660);
and U10544 (N_10544,N_9770,N_9652);
and U10545 (N_10545,N_10073,N_9830);
or U10546 (N_10546,N_9626,N_10020);
or U10547 (N_10547,N_9773,N_9688);
xnor U10548 (N_10548,N_10162,N_9934);
and U10549 (N_10549,N_10176,N_10078);
nand U10550 (N_10550,N_10102,N_9737);
or U10551 (N_10551,N_10107,N_9943);
nor U10552 (N_10552,N_9969,N_9900);
nor U10553 (N_10553,N_9715,N_9758);
nand U10554 (N_10554,N_9950,N_9737);
and U10555 (N_10555,N_9769,N_9922);
and U10556 (N_10556,N_10058,N_9844);
nor U10557 (N_10557,N_10083,N_9920);
nor U10558 (N_10558,N_9712,N_9893);
nand U10559 (N_10559,N_9622,N_9934);
xor U10560 (N_10560,N_10197,N_9676);
xnor U10561 (N_10561,N_9622,N_10194);
xor U10562 (N_10562,N_9987,N_10026);
nand U10563 (N_10563,N_9842,N_9743);
and U10564 (N_10564,N_9824,N_10166);
xnor U10565 (N_10565,N_9652,N_9802);
or U10566 (N_10566,N_9924,N_9948);
nand U10567 (N_10567,N_10033,N_9796);
xor U10568 (N_10568,N_9600,N_10128);
nor U10569 (N_10569,N_10082,N_9703);
nor U10570 (N_10570,N_10185,N_9697);
or U10571 (N_10571,N_10002,N_10162);
nand U10572 (N_10572,N_10040,N_9722);
xnor U10573 (N_10573,N_9687,N_10021);
nor U10574 (N_10574,N_9720,N_10043);
nand U10575 (N_10575,N_9615,N_9826);
xor U10576 (N_10576,N_9757,N_9821);
nor U10577 (N_10577,N_10080,N_10194);
and U10578 (N_10578,N_9743,N_9814);
or U10579 (N_10579,N_9836,N_9855);
nand U10580 (N_10580,N_9951,N_10182);
or U10581 (N_10581,N_10185,N_10157);
xnor U10582 (N_10582,N_10189,N_9828);
nand U10583 (N_10583,N_9990,N_9991);
or U10584 (N_10584,N_10106,N_9936);
and U10585 (N_10585,N_9980,N_10061);
nand U10586 (N_10586,N_9713,N_9859);
nand U10587 (N_10587,N_9924,N_9974);
nor U10588 (N_10588,N_9874,N_9958);
xor U10589 (N_10589,N_10038,N_9668);
and U10590 (N_10590,N_9648,N_9884);
xor U10591 (N_10591,N_9744,N_10128);
nor U10592 (N_10592,N_9816,N_10198);
nand U10593 (N_10593,N_9952,N_10146);
and U10594 (N_10594,N_9856,N_9671);
nand U10595 (N_10595,N_10067,N_9864);
or U10596 (N_10596,N_9770,N_9850);
nand U10597 (N_10597,N_10176,N_9859);
xor U10598 (N_10598,N_10132,N_10076);
xnor U10599 (N_10599,N_9992,N_10092);
or U10600 (N_10600,N_9996,N_9829);
nor U10601 (N_10601,N_9832,N_9800);
and U10602 (N_10602,N_9697,N_10172);
nand U10603 (N_10603,N_9803,N_9631);
and U10604 (N_10604,N_9833,N_9700);
nor U10605 (N_10605,N_10117,N_10095);
and U10606 (N_10606,N_9849,N_10189);
nor U10607 (N_10607,N_10135,N_9628);
nand U10608 (N_10608,N_9926,N_10102);
nand U10609 (N_10609,N_9957,N_9950);
and U10610 (N_10610,N_9690,N_10051);
nand U10611 (N_10611,N_10116,N_9813);
or U10612 (N_10612,N_9759,N_9630);
xnor U10613 (N_10613,N_10024,N_9732);
and U10614 (N_10614,N_9760,N_9882);
nor U10615 (N_10615,N_10170,N_9789);
xor U10616 (N_10616,N_9910,N_10137);
xnor U10617 (N_10617,N_9618,N_10076);
or U10618 (N_10618,N_10196,N_10040);
nor U10619 (N_10619,N_9785,N_10100);
nand U10620 (N_10620,N_10051,N_9882);
or U10621 (N_10621,N_9959,N_9723);
nor U10622 (N_10622,N_9890,N_10049);
xnor U10623 (N_10623,N_9848,N_9839);
or U10624 (N_10624,N_10097,N_9737);
xor U10625 (N_10625,N_10041,N_9925);
and U10626 (N_10626,N_9912,N_10100);
nand U10627 (N_10627,N_10142,N_10099);
and U10628 (N_10628,N_9769,N_9655);
or U10629 (N_10629,N_10096,N_9636);
and U10630 (N_10630,N_10095,N_9664);
nand U10631 (N_10631,N_10179,N_10185);
xnor U10632 (N_10632,N_10171,N_10187);
xor U10633 (N_10633,N_10040,N_9767);
and U10634 (N_10634,N_9841,N_10125);
nor U10635 (N_10635,N_9632,N_9827);
or U10636 (N_10636,N_9987,N_9786);
nand U10637 (N_10637,N_9973,N_9912);
and U10638 (N_10638,N_10162,N_10057);
nor U10639 (N_10639,N_9994,N_9906);
nor U10640 (N_10640,N_9767,N_9872);
nor U10641 (N_10641,N_9611,N_9690);
and U10642 (N_10642,N_9996,N_9913);
nor U10643 (N_10643,N_9925,N_10078);
and U10644 (N_10644,N_9962,N_10157);
nand U10645 (N_10645,N_10118,N_9618);
nand U10646 (N_10646,N_9873,N_10181);
and U10647 (N_10647,N_10064,N_9804);
xor U10648 (N_10648,N_10170,N_10134);
and U10649 (N_10649,N_10086,N_9821);
and U10650 (N_10650,N_9692,N_9824);
xnor U10651 (N_10651,N_9774,N_9787);
and U10652 (N_10652,N_9893,N_10083);
and U10653 (N_10653,N_10013,N_9880);
nand U10654 (N_10654,N_10100,N_10081);
xor U10655 (N_10655,N_9907,N_9625);
xor U10656 (N_10656,N_9607,N_9674);
xor U10657 (N_10657,N_9976,N_9800);
or U10658 (N_10658,N_9932,N_9872);
and U10659 (N_10659,N_9656,N_9831);
and U10660 (N_10660,N_9633,N_10070);
or U10661 (N_10661,N_9850,N_10127);
or U10662 (N_10662,N_9789,N_10059);
and U10663 (N_10663,N_9800,N_10070);
xor U10664 (N_10664,N_10028,N_10104);
and U10665 (N_10665,N_9694,N_9692);
nor U10666 (N_10666,N_10083,N_9949);
nand U10667 (N_10667,N_10028,N_9879);
or U10668 (N_10668,N_9849,N_10005);
nand U10669 (N_10669,N_9976,N_9802);
nor U10670 (N_10670,N_9829,N_10055);
nand U10671 (N_10671,N_9984,N_10141);
and U10672 (N_10672,N_10012,N_10129);
nor U10673 (N_10673,N_10027,N_9681);
and U10674 (N_10674,N_10159,N_9721);
nor U10675 (N_10675,N_9751,N_9787);
or U10676 (N_10676,N_9894,N_9760);
nand U10677 (N_10677,N_9768,N_10161);
xor U10678 (N_10678,N_9635,N_10066);
nor U10679 (N_10679,N_10114,N_10007);
or U10680 (N_10680,N_10004,N_9662);
or U10681 (N_10681,N_9957,N_9652);
xor U10682 (N_10682,N_10101,N_10149);
or U10683 (N_10683,N_9925,N_9711);
nor U10684 (N_10684,N_9658,N_9805);
or U10685 (N_10685,N_9950,N_10155);
and U10686 (N_10686,N_9742,N_9826);
or U10687 (N_10687,N_9837,N_9968);
nand U10688 (N_10688,N_9910,N_9703);
xnor U10689 (N_10689,N_10017,N_9959);
nand U10690 (N_10690,N_9666,N_9797);
xnor U10691 (N_10691,N_9988,N_9758);
xor U10692 (N_10692,N_9667,N_9938);
or U10693 (N_10693,N_9615,N_9718);
nor U10694 (N_10694,N_10043,N_10102);
xnor U10695 (N_10695,N_9953,N_9633);
xnor U10696 (N_10696,N_10181,N_10123);
nor U10697 (N_10697,N_9850,N_9905);
or U10698 (N_10698,N_10083,N_9937);
xnor U10699 (N_10699,N_9837,N_9840);
nand U10700 (N_10700,N_9661,N_9677);
xnor U10701 (N_10701,N_9834,N_9657);
nor U10702 (N_10702,N_9756,N_9874);
or U10703 (N_10703,N_10162,N_9853);
and U10704 (N_10704,N_10075,N_9955);
or U10705 (N_10705,N_10056,N_9734);
and U10706 (N_10706,N_9694,N_9953);
nor U10707 (N_10707,N_9864,N_10035);
nor U10708 (N_10708,N_9808,N_9814);
nand U10709 (N_10709,N_9783,N_10047);
nand U10710 (N_10710,N_9968,N_10178);
and U10711 (N_10711,N_9933,N_9610);
or U10712 (N_10712,N_9711,N_9753);
nand U10713 (N_10713,N_10141,N_10009);
nand U10714 (N_10714,N_9732,N_9974);
xnor U10715 (N_10715,N_9821,N_10094);
and U10716 (N_10716,N_10029,N_9752);
or U10717 (N_10717,N_9942,N_9988);
or U10718 (N_10718,N_9792,N_10156);
nor U10719 (N_10719,N_10025,N_9630);
and U10720 (N_10720,N_9772,N_9749);
or U10721 (N_10721,N_9706,N_10051);
and U10722 (N_10722,N_9928,N_9990);
nand U10723 (N_10723,N_9786,N_10021);
nand U10724 (N_10724,N_9609,N_10180);
xnor U10725 (N_10725,N_9779,N_9637);
nand U10726 (N_10726,N_9958,N_10150);
nand U10727 (N_10727,N_10122,N_9937);
or U10728 (N_10728,N_10163,N_9810);
and U10729 (N_10729,N_9645,N_9861);
nor U10730 (N_10730,N_10022,N_9817);
xnor U10731 (N_10731,N_10102,N_9621);
and U10732 (N_10732,N_9670,N_10088);
nor U10733 (N_10733,N_9617,N_9948);
nor U10734 (N_10734,N_9735,N_10007);
nand U10735 (N_10735,N_9640,N_9861);
or U10736 (N_10736,N_10143,N_9960);
xnor U10737 (N_10737,N_9799,N_9690);
nand U10738 (N_10738,N_9704,N_10018);
or U10739 (N_10739,N_9772,N_9763);
or U10740 (N_10740,N_9832,N_10040);
nor U10741 (N_10741,N_10089,N_9932);
xnor U10742 (N_10742,N_9842,N_9894);
nand U10743 (N_10743,N_10094,N_10035);
nor U10744 (N_10744,N_10129,N_9889);
or U10745 (N_10745,N_9726,N_9734);
nor U10746 (N_10746,N_9903,N_9612);
nand U10747 (N_10747,N_9635,N_9667);
xor U10748 (N_10748,N_9761,N_9653);
xnor U10749 (N_10749,N_10008,N_9909);
xnor U10750 (N_10750,N_9650,N_9977);
nor U10751 (N_10751,N_9916,N_10048);
nand U10752 (N_10752,N_9948,N_10165);
or U10753 (N_10753,N_9671,N_9951);
and U10754 (N_10754,N_9772,N_10013);
or U10755 (N_10755,N_9686,N_9666);
and U10756 (N_10756,N_9938,N_9813);
nor U10757 (N_10757,N_9788,N_10000);
nand U10758 (N_10758,N_9814,N_9671);
xor U10759 (N_10759,N_9724,N_10024);
nor U10760 (N_10760,N_9706,N_10004);
and U10761 (N_10761,N_10087,N_9831);
or U10762 (N_10762,N_9768,N_9790);
nand U10763 (N_10763,N_10102,N_9836);
xnor U10764 (N_10764,N_9912,N_9657);
nor U10765 (N_10765,N_9835,N_9868);
and U10766 (N_10766,N_9606,N_9848);
xnor U10767 (N_10767,N_10169,N_9648);
nand U10768 (N_10768,N_10074,N_10151);
nand U10769 (N_10769,N_10187,N_10009);
and U10770 (N_10770,N_9936,N_9735);
or U10771 (N_10771,N_10035,N_10017);
nor U10772 (N_10772,N_10046,N_10100);
and U10773 (N_10773,N_9786,N_9860);
nor U10774 (N_10774,N_9677,N_9924);
or U10775 (N_10775,N_9608,N_9760);
nand U10776 (N_10776,N_9850,N_10008);
and U10777 (N_10777,N_9896,N_9631);
or U10778 (N_10778,N_9714,N_9864);
xnor U10779 (N_10779,N_10003,N_9779);
and U10780 (N_10780,N_10117,N_10086);
xor U10781 (N_10781,N_10171,N_9864);
xnor U10782 (N_10782,N_9961,N_9950);
or U10783 (N_10783,N_9635,N_10132);
and U10784 (N_10784,N_9726,N_9963);
nor U10785 (N_10785,N_10151,N_10064);
nor U10786 (N_10786,N_10143,N_9661);
nand U10787 (N_10787,N_9971,N_9741);
nor U10788 (N_10788,N_10180,N_10080);
or U10789 (N_10789,N_9759,N_10050);
nor U10790 (N_10790,N_9982,N_10113);
and U10791 (N_10791,N_10078,N_9634);
xnor U10792 (N_10792,N_9720,N_10008);
nor U10793 (N_10793,N_10166,N_9924);
xor U10794 (N_10794,N_9741,N_9979);
or U10795 (N_10795,N_10031,N_9930);
and U10796 (N_10796,N_9975,N_9708);
nor U10797 (N_10797,N_9607,N_10129);
xor U10798 (N_10798,N_10071,N_9623);
nor U10799 (N_10799,N_9922,N_9994);
or U10800 (N_10800,N_10258,N_10681);
xor U10801 (N_10801,N_10492,N_10724);
nand U10802 (N_10802,N_10290,N_10275);
or U10803 (N_10803,N_10443,N_10320);
nor U10804 (N_10804,N_10264,N_10509);
nor U10805 (N_10805,N_10407,N_10607);
nor U10806 (N_10806,N_10340,N_10437);
and U10807 (N_10807,N_10202,N_10248);
xor U10808 (N_10808,N_10250,N_10501);
or U10809 (N_10809,N_10459,N_10759);
nand U10810 (N_10810,N_10757,N_10219);
and U10811 (N_10811,N_10451,N_10302);
nor U10812 (N_10812,N_10548,N_10625);
nand U10813 (N_10813,N_10643,N_10515);
xor U10814 (N_10814,N_10427,N_10400);
xnor U10815 (N_10815,N_10610,N_10424);
xor U10816 (N_10816,N_10305,N_10461);
and U10817 (N_10817,N_10673,N_10413);
nor U10818 (N_10818,N_10620,N_10404);
nor U10819 (N_10819,N_10281,N_10429);
nand U10820 (N_10820,N_10351,N_10700);
or U10821 (N_10821,N_10709,N_10708);
xor U10822 (N_10822,N_10683,N_10630);
nand U10823 (N_10823,N_10375,N_10217);
or U10824 (N_10824,N_10448,N_10265);
xnor U10825 (N_10825,N_10260,N_10535);
nand U10826 (N_10826,N_10784,N_10588);
xnor U10827 (N_10827,N_10203,N_10563);
nand U10828 (N_10828,N_10552,N_10334);
nand U10829 (N_10829,N_10431,N_10476);
nor U10830 (N_10830,N_10790,N_10216);
nand U10831 (N_10831,N_10597,N_10464);
nor U10832 (N_10832,N_10726,N_10371);
nor U10833 (N_10833,N_10692,N_10415);
and U10834 (N_10834,N_10321,N_10355);
or U10835 (N_10835,N_10514,N_10398);
xnor U10836 (N_10836,N_10279,N_10298);
nand U10837 (N_10837,N_10335,N_10496);
xnor U10838 (N_10838,N_10299,N_10566);
or U10839 (N_10839,N_10545,N_10278);
or U10840 (N_10840,N_10756,N_10534);
and U10841 (N_10841,N_10395,N_10731);
xnor U10842 (N_10842,N_10263,N_10704);
nor U10843 (N_10843,N_10468,N_10200);
or U10844 (N_10844,N_10269,N_10750);
nand U10845 (N_10845,N_10417,N_10593);
or U10846 (N_10846,N_10783,N_10270);
nor U10847 (N_10847,N_10256,N_10627);
nand U10848 (N_10848,N_10669,N_10456);
nand U10849 (N_10849,N_10656,N_10676);
xnor U10850 (N_10850,N_10328,N_10358);
xor U10851 (N_10851,N_10658,N_10495);
nor U10852 (N_10852,N_10316,N_10477);
nor U10853 (N_10853,N_10695,N_10490);
xor U10854 (N_10854,N_10293,N_10487);
xor U10855 (N_10855,N_10562,N_10774);
xor U10856 (N_10856,N_10277,N_10699);
nor U10857 (N_10857,N_10767,N_10785);
nor U10858 (N_10858,N_10409,N_10352);
nand U10859 (N_10859,N_10603,N_10636);
or U10860 (N_10860,N_10796,N_10241);
xnor U10861 (N_10861,N_10575,N_10434);
and U10862 (N_10862,N_10576,N_10614);
or U10863 (N_10863,N_10787,N_10201);
nor U10864 (N_10864,N_10380,N_10341);
and U10865 (N_10865,N_10420,N_10520);
and U10866 (N_10866,N_10310,N_10581);
nand U10867 (N_10867,N_10317,N_10444);
xor U10868 (N_10868,N_10403,N_10347);
nor U10869 (N_10869,N_10484,N_10578);
or U10870 (N_10870,N_10247,N_10547);
nor U10871 (N_10871,N_10727,N_10349);
xnor U10872 (N_10872,N_10629,N_10589);
xor U10873 (N_10873,N_10306,N_10272);
and U10874 (N_10874,N_10747,N_10594);
nor U10875 (N_10875,N_10628,N_10686);
nor U10876 (N_10876,N_10554,N_10421);
and U10877 (N_10877,N_10367,N_10579);
and U10878 (N_10878,N_10606,N_10243);
and U10879 (N_10879,N_10214,N_10525);
nand U10880 (N_10880,N_10778,N_10729);
nand U10881 (N_10881,N_10518,N_10753);
and U10882 (N_10882,N_10208,N_10679);
xor U10883 (N_10883,N_10622,N_10204);
and U10884 (N_10884,N_10768,N_10227);
xnor U10885 (N_10885,N_10274,N_10454);
xor U10886 (N_10886,N_10325,N_10745);
nand U10887 (N_10887,N_10261,N_10749);
nor U10888 (N_10888,N_10471,N_10493);
xnor U10889 (N_10889,N_10645,N_10458);
xor U10890 (N_10890,N_10654,N_10780);
nand U10891 (N_10891,N_10229,N_10245);
nand U10892 (N_10892,N_10326,N_10678);
nand U10893 (N_10893,N_10285,N_10440);
nand U10894 (N_10894,N_10311,N_10393);
or U10895 (N_10895,N_10693,N_10324);
and U10896 (N_10896,N_10583,N_10396);
xor U10897 (N_10897,N_10213,N_10430);
nand U10898 (N_10898,N_10297,N_10408);
nor U10899 (N_10899,N_10618,N_10551);
nor U10900 (N_10900,N_10315,N_10602);
nand U10901 (N_10901,N_10540,N_10510);
nand U10902 (N_10902,N_10761,N_10498);
nor U10903 (N_10903,N_10668,N_10604);
xor U10904 (N_10904,N_10337,N_10374);
and U10905 (N_10905,N_10527,N_10432);
xnor U10906 (N_10906,N_10388,N_10379);
and U10907 (N_10907,N_10211,N_10572);
and U10908 (N_10908,N_10730,N_10391);
nor U10909 (N_10909,N_10705,N_10283);
or U10910 (N_10910,N_10303,N_10586);
or U10911 (N_10911,N_10291,N_10600);
xor U10912 (N_10912,N_10333,N_10406);
xor U10913 (N_10913,N_10596,N_10573);
or U10914 (N_10914,N_10598,N_10414);
xor U10915 (N_10915,N_10344,N_10276);
xor U10916 (N_10916,N_10226,N_10240);
nand U10917 (N_10917,N_10376,N_10339);
xor U10918 (N_10918,N_10682,N_10218);
nand U10919 (N_10919,N_10402,N_10253);
or U10920 (N_10920,N_10336,N_10743);
nor U10921 (N_10921,N_10296,N_10671);
nor U10922 (N_10922,N_10499,N_10649);
and U10923 (N_10923,N_10307,N_10238);
nor U10924 (N_10924,N_10762,N_10433);
xnor U10925 (N_10925,N_10266,N_10795);
and U10926 (N_10926,N_10512,N_10652);
and U10927 (N_10927,N_10345,N_10262);
or U10928 (N_10928,N_10733,N_10342);
nand U10929 (N_10929,N_10794,N_10478);
xor U10930 (N_10930,N_10770,N_10300);
and U10931 (N_10931,N_10577,N_10390);
and U10932 (N_10932,N_10752,N_10497);
nand U10933 (N_10933,N_10485,N_10505);
xnor U10934 (N_10934,N_10508,N_10397);
or U10935 (N_10935,N_10687,N_10209);
nor U10936 (N_10936,N_10766,N_10222);
and U10937 (N_10937,N_10234,N_10701);
nand U10938 (N_10938,N_10236,N_10631);
xnor U10939 (N_10939,N_10504,N_10529);
nand U10940 (N_10940,N_10777,N_10613);
or U10941 (N_10941,N_10738,N_10585);
and U10942 (N_10942,N_10530,N_10289);
nand U10943 (N_10943,N_10634,N_10282);
or U10944 (N_10944,N_10480,N_10771);
xor U10945 (N_10945,N_10368,N_10372);
nor U10946 (N_10946,N_10313,N_10482);
or U10947 (N_10947,N_10561,N_10455);
xor U10948 (N_10948,N_10318,N_10775);
and U10949 (N_10949,N_10696,N_10354);
and U10950 (N_10950,N_10582,N_10612);
and U10951 (N_10951,N_10254,N_10472);
or U10952 (N_10952,N_10348,N_10748);
nor U10953 (N_10953,N_10373,N_10387);
nor U10954 (N_10954,N_10793,N_10394);
nand U10955 (N_10955,N_10744,N_10591);
nor U10956 (N_10956,N_10740,N_10633);
nand U10957 (N_10957,N_10419,N_10502);
nor U10958 (N_10958,N_10776,N_10584);
and U10959 (N_10959,N_10723,N_10416);
nor U10960 (N_10960,N_10706,N_10511);
xor U10961 (N_10961,N_10550,N_10257);
nand U10962 (N_10962,N_10327,N_10797);
and U10963 (N_10963,N_10732,N_10736);
nor U10964 (N_10964,N_10428,N_10568);
or U10965 (N_10965,N_10553,N_10765);
nor U10966 (N_10966,N_10688,N_10255);
and U10967 (N_10967,N_10605,N_10644);
nor U10968 (N_10968,N_10647,N_10564);
nor U10969 (N_10969,N_10314,N_10792);
nor U10970 (N_10970,N_10287,N_10242);
nor U10971 (N_10971,N_10663,N_10624);
or U10972 (N_10972,N_10786,N_10370);
nor U10973 (N_10973,N_10383,N_10773);
nand U10974 (N_10974,N_10735,N_10378);
xor U10975 (N_10975,N_10539,N_10779);
xor U10976 (N_10976,N_10533,N_10764);
xor U10977 (N_10977,N_10537,N_10423);
and U10978 (N_10978,N_10788,N_10363);
or U10979 (N_10979,N_10516,N_10667);
and U10980 (N_10980,N_10356,N_10452);
or U10981 (N_10981,N_10401,N_10239);
and U10982 (N_10982,N_10689,N_10488);
xor U10983 (N_10983,N_10332,N_10225);
nand U10984 (N_10984,N_10331,N_10721);
xor U10985 (N_10985,N_10251,N_10312);
and U10986 (N_10986,N_10720,N_10309);
or U10987 (N_10987,N_10651,N_10590);
nor U10988 (N_10988,N_10680,N_10481);
nor U10989 (N_10989,N_10574,N_10445);
and U10990 (N_10990,N_10763,N_10364);
and U10991 (N_10991,N_10691,N_10565);
nand U10992 (N_10992,N_10422,N_10426);
nand U10993 (N_10993,N_10304,N_10690);
xnor U10994 (N_10994,N_10556,N_10343);
and U10995 (N_10995,N_10206,N_10694);
xor U10996 (N_10996,N_10411,N_10205);
nor U10997 (N_10997,N_10546,N_10361);
xor U10998 (N_10998,N_10357,N_10728);
and U10999 (N_10999,N_10781,N_10381);
or U11000 (N_11000,N_10301,N_10715);
and U11001 (N_11001,N_10284,N_10460);
nand U11002 (N_11002,N_10292,N_10491);
nand U11003 (N_11003,N_10685,N_10224);
or U11004 (N_11004,N_10467,N_10369);
or U11005 (N_11005,N_10710,N_10639);
and U11006 (N_11006,N_10507,N_10338);
and U11007 (N_11007,N_10223,N_10555);
or U11008 (N_11008,N_10215,N_10295);
and U11009 (N_11009,N_10592,N_10760);
xnor U11010 (N_11010,N_10523,N_10410);
nand U11011 (N_11011,N_10675,N_10718);
nand U11012 (N_11012,N_10670,N_10362);
nand U11013 (N_11013,N_10385,N_10615);
xor U11014 (N_11014,N_10714,N_10323);
xor U11015 (N_11015,N_10465,N_10538);
nand U11016 (N_11016,N_10623,N_10608);
and U11017 (N_11017,N_10382,N_10541);
and U11018 (N_11018,N_10716,N_10470);
or U11019 (N_11019,N_10436,N_10587);
xnor U11020 (N_11020,N_10221,N_10463);
nor U11021 (N_11021,N_10469,N_10271);
xnor U11022 (N_11022,N_10329,N_10653);
nor U11023 (N_11023,N_10717,N_10637);
nand U11024 (N_11024,N_10799,N_10286);
and U11025 (N_11025,N_10473,N_10599);
nand U11026 (N_11026,N_10711,N_10755);
xor U11027 (N_11027,N_10536,N_10734);
nor U11028 (N_11028,N_10237,N_10570);
nor U11029 (N_11029,N_10462,N_10418);
nand U11030 (N_11030,N_10475,N_10447);
nand U11031 (N_11031,N_10319,N_10640);
and U11032 (N_11032,N_10399,N_10611);
nor U11033 (N_11033,N_10233,N_10713);
nand U11034 (N_11034,N_10280,N_10601);
or U11035 (N_11035,N_10366,N_10609);
and U11036 (N_11036,N_10228,N_10489);
and U11037 (N_11037,N_10405,N_10425);
nand U11038 (N_11038,N_10674,N_10742);
xor U11039 (N_11039,N_10642,N_10494);
or U11040 (N_11040,N_10486,N_10466);
and U11041 (N_11041,N_10531,N_10703);
nand U11042 (N_11042,N_10769,N_10249);
and U11043 (N_11043,N_10549,N_10662);
xor U11044 (N_11044,N_10210,N_10626);
and U11045 (N_11045,N_10360,N_10503);
nand U11046 (N_11046,N_10791,N_10522);
nand U11047 (N_11047,N_10737,N_10751);
xnor U11048 (N_11048,N_10412,N_10619);
nand U11049 (N_11049,N_10660,N_10595);
nor U11050 (N_11050,N_10580,N_10544);
xnor U11051 (N_11051,N_10648,N_10442);
xnor U11052 (N_11052,N_10521,N_10641);
and U11053 (N_11053,N_10230,N_10782);
nor U11054 (N_11054,N_10386,N_10246);
or U11055 (N_11055,N_10632,N_10308);
xnor U11056 (N_11056,N_10702,N_10353);
nand U11057 (N_11057,N_10559,N_10288);
nor U11058 (N_11058,N_10500,N_10513);
nor U11059 (N_11059,N_10268,N_10235);
or U11060 (N_11060,N_10438,N_10677);
xor U11061 (N_11061,N_10543,N_10244);
and U11062 (N_11062,N_10392,N_10621);
nor U11063 (N_11063,N_10772,N_10722);
and U11064 (N_11064,N_10212,N_10567);
and U11065 (N_11065,N_10267,N_10571);
and U11066 (N_11066,N_10558,N_10273);
or U11067 (N_11067,N_10542,N_10446);
nor U11068 (N_11068,N_10389,N_10725);
nand U11069 (N_11069,N_10557,N_10758);
or U11070 (N_11070,N_10479,N_10483);
nor U11071 (N_11071,N_10453,N_10439);
or U11072 (N_11072,N_10754,N_10322);
or U11073 (N_11073,N_10617,N_10569);
xnor U11074 (N_11074,N_10532,N_10655);
xnor U11075 (N_11075,N_10746,N_10207);
or U11076 (N_11076,N_10441,N_10560);
nand U11077 (N_11077,N_10635,N_10798);
xor U11078 (N_11078,N_10789,N_10526);
nand U11079 (N_11079,N_10666,N_10528);
or U11080 (N_11080,N_10524,N_10359);
xor U11081 (N_11081,N_10657,N_10659);
nor U11082 (N_11082,N_10739,N_10232);
nor U11083 (N_11083,N_10697,N_10457);
or U11084 (N_11084,N_10741,N_10664);
nand U11085 (N_11085,N_10377,N_10252);
nor U11086 (N_11086,N_10330,N_10665);
or U11087 (N_11087,N_10707,N_10638);
xnor U11088 (N_11088,N_10684,N_10646);
or U11089 (N_11089,N_10449,N_10616);
or U11090 (N_11090,N_10474,N_10346);
xnor U11091 (N_11091,N_10661,N_10517);
nor U11092 (N_11092,N_10712,N_10698);
and U11093 (N_11093,N_10294,N_10650);
nor U11094 (N_11094,N_10435,N_10672);
nand U11095 (N_11095,N_10384,N_10259);
nand U11096 (N_11096,N_10365,N_10719);
nand U11097 (N_11097,N_10350,N_10231);
xnor U11098 (N_11098,N_10506,N_10519);
nand U11099 (N_11099,N_10220,N_10450);
and U11100 (N_11100,N_10796,N_10644);
nand U11101 (N_11101,N_10658,N_10334);
or U11102 (N_11102,N_10756,N_10323);
nand U11103 (N_11103,N_10343,N_10357);
nor U11104 (N_11104,N_10265,N_10532);
nand U11105 (N_11105,N_10422,N_10756);
nor U11106 (N_11106,N_10607,N_10250);
xnor U11107 (N_11107,N_10449,N_10626);
nand U11108 (N_11108,N_10352,N_10254);
xor U11109 (N_11109,N_10512,N_10265);
xnor U11110 (N_11110,N_10485,N_10490);
and U11111 (N_11111,N_10431,N_10450);
and U11112 (N_11112,N_10223,N_10701);
nor U11113 (N_11113,N_10366,N_10218);
nand U11114 (N_11114,N_10405,N_10522);
and U11115 (N_11115,N_10506,N_10741);
nand U11116 (N_11116,N_10507,N_10367);
nor U11117 (N_11117,N_10522,N_10280);
and U11118 (N_11118,N_10403,N_10223);
and U11119 (N_11119,N_10598,N_10699);
xor U11120 (N_11120,N_10773,N_10762);
nor U11121 (N_11121,N_10213,N_10374);
or U11122 (N_11122,N_10694,N_10261);
nand U11123 (N_11123,N_10329,N_10568);
nand U11124 (N_11124,N_10711,N_10259);
nor U11125 (N_11125,N_10665,N_10583);
or U11126 (N_11126,N_10720,N_10741);
xor U11127 (N_11127,N_10294,N_10713);
or U11128 (N_11128,N_10699,N_10321);
or U11129 (N_11129,N_10543,N_10628);
or U11130 (N_11130,N_10547,N_10748);
and U11131 (N_11131,N_10798,N_10326);
xnor U11132 (N_11132,N_10659,N_10443);
nand U11133 (N_11133,N_10440,N_10600);
nor U11134 (N_11134,N_10721,N_10738);
xnor U11135 (N_11135,N_10252,N_10509);
nor U11136 (N_11136,N_10335,N_10282);
nand U11137 (N_11137,N_10253,N_10455);
nor U11138 (N_11138,N_10286,N_10558);
xor U11139 (N_11139,N_10392,N_10274);
and U11140 (N_11140,N_10789,N_10359);
nor U11141 (N_11141,N_10236,N_10559);
and U11142 (N_11142,N_10605,N_10366);
nand U11143 (N_11143,N_10554,N_10440);
nand U11144 (N_11144,N_10639,N_10213);
and U11145 (N_11145,N_10574,N_10578);
and U11146 (N_11146,N_10505,N_10664);
nand U11147 (N_11147,N_10685,N_10775);
or U11148 (N_11148,N_10310,N_10405);
or U11149 (N_11149,N_10486,N_10759);
and U11150 (N_11150,N_10511,N_10250);
or U11151 (N_11151,N_10311,N_10356);
and U11152 (N_11152,N_10304,N_10586);
and U11153 (N_11153,N_10564,N_10656);
xnor U11154 (N_11154,N_10438,N_10321);
or U11155 (N_11155,N_10570,N_10575);
xnor U11156 (N_11156,N_10394,N_10515);
or U11157 (N_11157,N_10300,N_10413);
or U11158 (N_11158,N_10533,N_10675);
nor U11159 (N_11159,N_10321,N_10591);
nand U11160 (N_11160,N_10664,N_10545);
nor U11161 (N_11161,N_10701,N_10444);
or U11162 (N_11162,N_10642,N_10282);
xnor U11163 (N_11163,N_10698,N_10412);
xor U11164 (N_11164,N_10341,N_10513);
nand U11165 (N_11165,N_10665,N_10732);
nor U11166 (N_11166,N_10409,N_10705);
and U11167 (N_11167,N_10782,N_10747);
nor U11168 (N_11168,N_10766,N_10626);
nor U11169 (N_11169,N_10704,N_10748);
nor U11170 (N_11170,N_10377,N_10793);
nor U11171 (N_11171,N_10510,N_10384);
nor U11172 (N_11172,N_10225,N_10278);
and U11173 (N_11173,N_10389,N_10252);
nand U11174 (N_11174,N_10234,N_10324);
nor U11175 (N_11175,N_10319,N_10726);
nor U11176 (N_11176,N_10582,N_10364);
xor U11177 (N_11177,N_10705,N_10402);
nand U11178 (N_11178,N_10718,N_10622);
or U11179 (N_11179,N_10537,N_10324);
nor U11180 (N_11180,N_10489,N_10314);
xor U11181 (N_11181,N_10532,N_10277);
and U11182 (N_11182,N_10641,N_10540);
nand U11183 (N_11183,N_10252,N_10504);
or U11184 (N_11184,N_10434,N_10437);
or U11185 (N_11185,N_10757,N_10643);
or U11186 (N_11186,N_10534,N_10421);
or U11187 (N_11187,N_10203,N_10388);
nor U11188 (N_11188,N_10614,N_10439);
xnor U11189 (N_11189,N_10612,N_10706);
or U11190 (N_11190,N_10600,N_10217);
nor U11191 (N_11191,N_10660,N_10579);
nor U11192 (N_11192,N_10475,N_10668);
xnor U11193 (N_11193,N_10382,N_10261);
nand U11194 (N_11194,N_10244,N_10275);
and U11195 (N_11195,N_10543,N_10660);
or U11196 (N_11196,N_10601,N_10424);
nand U11197 (N_11197,N_10358,N_10278);
and U11198 (N_11198,N_10589,N_10415);
nor U11199 (N_11199,N_10607,N_10298);
nor U11200 (N_11200,N_10699,N_10317);
nand U11201 (N_11201,N_10664,N_10571);
xnor U11202 (N_11202,N_10616,N_10400);
or U11203 (N_11203,N_10410,N_10735);
nand U11204 (N_11204,N_10534,N_10441);
nand U11205 (N_11205,N_10747,N_10734);
xor U11206 (N_11206,N_10629,N_10320);
xor U11207 (N_11207,N_10661,N_10515);
nand U11208 (N_11208,N_10714,N_10590);
nand U11209 (N_11209,N_10763,N_10350);
nand U11210 (N_11210,N_10328,N_10217);
nand U11211 (N_11211,N_10204,N_10407);
and U11212 (N_11212,N_10357,N_10303);
nor U11213 (N_11213,N_10347,N_10555);
nor U11214 (N_11214,N_10483,N_10524);
and U11215 (N_11215,N_10451,N_10732);
and U11216 (N_11216,N_10336,N_10733);
nand U11217 (N_11217,N_10521,N_10381);
and U11218 (N_11218,N_10348,N_10429);
xor U11219 (N_11219,N_10513,N_10375);
xor U11220 (N_11220,N_10698,N_10789);
nor U11221 (N_11221,N_10787,N_10384);
or U11222 (N_11222,N_10211,N_10625);
or U11223 (N_11223,N_10670,N_10687);
nor U11224 (N_11224,N_10547,N_10369);
xor U11225 (N_11225,N_10359,N_10522);
nor U11226 (N_11226,N_10613,N_10328);
nand U11227 (N_11227,N_10561,N_10750);
xnor U11228 (N_11228,N_10342,N_10732);
nor U11229 (N_11229,N_10561,N_10770);
xnor U11230 (N_11230,N_10797,N_10442);
or U11231 (N_11231,N_10629,N_10362);
xnor U11232 (N_11232,N_10592,N_10497);
or U11233 (N_11233,N_10340,N_10729);
and U11234 (N_11234,N_10285,N_10253);
nor U11235 (N_11235,N_10648,N_10545);
xnor U11236 (N_11236,N_10789,N_10393);
and U11237 (N_11237,N_10763,N_10713);
nor U11238 (N_11238,N_10594,N_10797);
nor U11239 (N_11239,N_10697,N_10710);
and U11240 (N_11240,N_10656,N_10783);
or U11241 (N_11241,N_10755,N_10563);
xnor U11242 (N_11242,N_10222,N_10763);
xor U11243 (N_11243,N_10447,N_10278);
xor U11244 (N_11244,N_10442,N_10765);
and U11245 (N_11245,N_10347,N_10447);
and U11246 (N_11246,N_10709,N_10217);
xnor U11247 (N_11247,N_10418,N_10729);
nand U11248 (N_11248,N_10485,N_10700);
nor U11249 (N_11249,N_10360,N_10293);
nor U11250 (N_11250,N_10270,N_10710);
nor U11251 (N_11251,N_10268,N_10385);
xnor U11252 (N_11252,N_10424,N_10381);
nor U11253 (N_11253,N_10383,N_10418);
nor U11254 (N_11254,N_10522,N_10743);
and U11255 (N_11255,N_10784,N_10393);
xnor U11256 (N_11256,N_10363,N_10701);
and U11257 (N_11257,N_10703,N_10357);
and U11258 (N_11258,N_10343,N_10422);
nor U11259 (N_11259,N_10266,N_10553);
and U11260 (N_11260,N_10535,N_10692);
nand U11261 (N_11261,N_10447,N_10729);
nand U11262 (N_11262,N_10301,N_10619);
and U11263 (N_11263,N_10397,N_10716);
and U11264 (N_11264,N_10313,N_10285);
nand U11265 (N_11265,N_10303,N_10335);
and U11266 (N_11266,N_10545,N_10690);
xor U11267 (N_11267,N_10392,N_10360);
xor U11268 (N_11268,N_10459,N_10785);
nor U11269 (N_11269,N_10623,N_10491);
nand U11270 (N_11270,N_10234,N_10763);
nor U11271 (N_11271,N_10221,N_10201);
nand U11272 (N_11272,N_10236,N_10622);
nand U11273 (N_11273,N_10739,N_10454);
nor U11274 (N_11274,N_10571,N_10789);
or U11275 (N_11275,N_10508,N_10349);
or U11276 (N_11276,N_10408,N_10474);
nand U11277 (N_11277,N_10282,N_10759);
nor U11278 (N_11278,N_10314,N_10720);
nand U11279 (N_11279,N_10408,N_10749);
or U11280 (N_11280,N_10478,N_10256);
nand U11281 (N_11281,N_10385,N_10665);
nand U11282 (N_11282,N_10367,N_10556);
nand U11283 (N_11283,N_10673,N_10247);
nand U11284 (N_11284,N_10494,N_10371);
or U11285 (N_11285,N_10245,N_10372);
nand U11286 (N_11286,N_10642,N_10453);
xnor U11287 (N_11287,N_10415,N_10665);
nor U11288 (N_11288,N_10607,N_10674);
or U11289 (N_11289,N_10601,N_10493);
nor U11290 (N_11290,N_10396,N_10536);
and U11291 (N_11291,N_10544,N_10319);
or U11292 (N_11292,N_10606,N_10369);
xor U11293 (N_11293,N_10650,N_10520);
xnor U11294 (N_11294,N_10613,N_10434);
nor U11295 (N_11295,N_10262,N_10395);
nor U11296 (N_11296,N_10668,N_10628);
and U11297 (N_11297,N_10466,N_10689);
nor U11298 (N_11298,N_10321,N_10755);
xor U11299 (N_11299,N_10375,N_10422);
or U11300 (N_11300,N_10485,N_10533);
or U11301 (N_11301,N_10571,N_10288);
and U11302 (N_11302,N_10306,N_10783);
xnor U11303 (N_11303,N_10505,N_10236);
nand U11304 (N_11304,N_10363,N_10720);
nor U11305 (N_11305,N_10639,N_10305);
or U11306 (N_11306,N_10287,N_10441);
xnor U11307 (N_11307,N_10511,N_10458);
and U11308 (N_11308,N_10740,N_10501);
and U11309 (N_11309,N_10414,N_10468);
and U11310 (N_11310,N_10362,N_10380);
nand U11311 (N_11311,N_10625,N_10703);
or U11312 (N_11312,N_10242,N_10416);
nor U11313 (N_11313,N_10328,N_10319);
nor U11314 (N_11314,N_10634,N_10692);
xor U11315 (N_11315,N_10454,N_10442);
nor U11316 (N_11316,N_10680,N_10225);
or U11317 (N_11317,N_10391,N_10376);
xor U11318 (N_11318,N_10556,N_10549);
nand U11319 (N_11319,N_10495,N_10260);
and U11320 (N_11320,N_10611,N_10367);
xnor U11321 (N_11321,N_10212,N_10374);
or U11322 (N_11322,N_10549,N_10761);
or U11323 (N_11323,N_10700,N_10202);
or U11324 (N_11324,N_10532,N_10761);
nand U11325 (N_11325,N_10416,N_10600);
nand U11326 (N_11326,N_10295,N_10642);
and U11327 (N_11327,N_10770,N_10488);
xor U11328 (N_11328,N_10365,N_10243);
nand U11329 (N_11329,N_10417,N_10358);
xnor U11330 (N_11330,N_10330,N_10670);
xnor U11331 (N_11331,N_10613,N_10402);
xnor U11332 (N_11332,N_10583,N_10514);
nor U11333 (N_11333,N_10790,N_10371);
xor U11334 (N_11334,N_10263,N_10685);
nor U11335 (N_11335,N_10581,N_10746);
nand U11336 (N_11336,N_10286,N_10768);
nand U11337 (N_11337,N_10342,N_10618);
nand U11338 (N_11338,N_10527,N_10423);
and U11339 (N_11339,N_10544,N_10648);
nand U11340 (N_11340,N_10601,N_10309);
nand U11341 (N_11341,N_10416,N_10761);
nor U11342 (N_11342,N_10341,N_10612);
xor U11343 (N_11343,N_10779,N_10270);
and U11344 (N_11344,N_10502,N_10620);
or U11345 (N_11345,N_10298,N_10789);
or U11346 (N_11346,N_10234,N_10729);
nor U11347 (N_11347,N_10264,N_10537);
xor U11348 (N_11348,N_10339,N_10361);
nor U11349 (N_11349,N_10611,N_10619);
and U11350 (N_11350,N_10750,N_10520);
or U11351 (N_11351,N_10259,N_10713);
nor U11352 (N_11352,N_10578,N_10316);
and U11353 (N_11353,N_10554,N_10595);
nor U11354 (N_11354,N_10321,N_10373);
nor U11355 (N_11355,N_10702,N_10355);
and U11356 (N_11356,N_10213,N_10672);
nand U11357 (N_11357,N_10599,N_10239);
nand U11358 (N_11358,N_10328,N_10240);
nor U11359 (N_11359,N_10642,N_10454);
nor U11360 (N_11360,N_10212,N_10635);
nand U11361 (N_11361,N_10708,N_10474);
and U11362 (N_11362,N_10374,N_10527);
and U11363 (N_11363,N_10215,N_10262);
nand U11364 (N_11364,N_10555,N_10546);
xnor U11365 (N_11365,N_10355,N_10450);
and U11366 (N_11366,N_10633,N_10265);
and U11367 (N_11367,N_10233,N_10204);
and U11368 (N_11368,N_10490,N_10435);
nor U11369 (N_11369,N_10745,N_10759);
nor U11370 (N_11370,N_10680,N_10428);
xor U11371 (N_11371,N_10602,N_10732);
nand U11372 (N_11372,N_10318,N_10782);
or U11373 (N_11373,N_10252,N_10640);
nand U11374 (N_11374,N_10478,N_10628);
nand U11375 (N_11375,N_10230,N_10329);
or U11376 (N_11376,N_10538,N_10760);
nor U11377 (N_11377,N_10222,N_10734);
and U11378 (N_11378,N_10682,N_10570);
xnor U11379 (N_11379,N_10204,N_10402);
xor U11380 (N_11380,N_10328,N_10473);
or U11381 (N_11381,N_10255,N_10308);
nand U11382 (N_11382,N_10646,N_10791);
nor U11383 (N_11383,N_10572,N_10682);
or U11384 (N_11384,N_10273,N_10586);
nand U11385 (N_11385,N_10256,N_10549);
and U11386 (N_11386,N_10515,N_10766);
xnor U11387 (N_11387,N_10548,N_10701);
and U11388 (N_11388,N_10784,N_10301);
nand U11389 (N_11389,N_10599,N_10455);
nor U11390 (N_11390,N_10429,N_10261);
and U11391 (N_11391,N_10510,N_10344);
or U11392 (N_11392,N_10672,N_10233);
xnor U11393 (N_11393,N_10528,N_10720);
nand U11394 (N_11394,N_10475,N_10336);
or U11395 (N_11395,N_10673,N_10569);
nor U11396 (N_11396,N_10778,N_10340);
and U11397 (N_11397,N_10328,N_10294);
and U11398 (N_11398,N_10268,N_10779);
nor U11399 (N_11399,N_10784,N_10778);
nand U11400 (N_11400,N_11297,N_10926);
nand U11401 (N_11401,N_11253,N_10852);
nand U11402 (N_11402,N_10827,N_10813);
and U11403 (N_11403,N_11160,N_10989);
nor U11404 (N_11404,N_11063,N_11113);
or U11405 (N_11405,N_10885,N_11201);
and U11406 (N_11406,N_10940,N_11101);
or U11407 (N_11407,N_10875,N_11048);
and U11408 (N_11408,N_10973,N_11339);
xnor U11409 (N_11409,N_11270,N_10917);
nand U11410 (N_11410,N_11143,N_10945);
nor U11411 (N_11411,N_11138,N_10980);
nand U11412 (N_11412,N_11250,N_11040);
xnor U11413 (N_11413,N_10888,N_11019);
nand U11414 (N_11414,N_10892,N_11249);
nor U11415 (N_11415,N_11075,N_10893);
nor U11416 (N_11416,N_11089,N_11306);
nor U11417 (N_11417,N_11151,N_10990);
xnor U11418 (N_11418,N_11059,N_11193);
nor U11419 (N_11419,N_11009,N_10804);
nand U11420 (N_11420,N_11294,N_11285);
nand U11421 (N_11421,N_11357,N_10933);
nand U11422 (N_11422,N_11218,N_11343);
and U11423 (N_11423,N_11240,N_10809);
or U11424 (N_11424,N_11200,N_10992);
nand U11425 (N_11425,N_10877,N_11356);
or U11426 (N_11426,N_11196,N_11399);
xor U11427 (N_11427,N_10821,N_10944);
nor U11428 (N_11428,N_10899,N_10906);
nor U11429 (N_11429,N_11037,N_11368);
and U11430 (N_11430,N_11332,N_11102);
and U11431 (N_11431,N_11100,N_10812);
and U11432 (N_11432,N_11382,N_11152);
and U11433 (N_11433,N_11271,N_11024);
xor U11434 (N_11434,N_11360,N_10900);
or U11435 (N_11435,N_11128,N_10842);
nand U11436 (N_11436,N_11350,N_10865);
and U11437 (N_11437,N_11117,N_10832);
and U11438 (N_11438,N_10960,N_11094);
nor U11439 (N_11439,N_10864,N_10919);
xor U11440 (N_11440,N_10853,N_11182);
nor U11441 (N_11441,N_10898,N_11067);
or U11442 (N_11442,N_10830,N_11066);
or U11443 (N_11443,N_11081,N_11302);
or U11444 (N_11444,N_11351,N_11046);
nor U11445 (N_11445,N_11324,N_10946);
nor U11446 (N_11446,N_11349,N_11011);
and U11447 (N_11447,N_11247,N_10996);
nand U11448 (N_11448,N_10897,N_11261);
xnor U11449 (N_11449,N_10984,N_10907);
nor U11450 (N_11450,N_10987,N_11042);
or U11451 (N_11451,N_10856,N_10835);
nor U11452 (N_11452,N_10872,N_10878);
nand U11453 (N_11453,N_10924,N_11062);
nor U11454 (N_11454,N_10905,N_11124);
and U11455 (N_11455,N_10998,N_10948);
nand U11456 (N_11456,N_11251,N_11219);
or U11457 (N_11457,N_11252,N_11105);
or U11458 (N_11458,N_11029,N_10951);
and U11459 (N_11459,N_10814,N_11224);
nand U11460 (N_11460,N_10895,N_11359);
or U11461 (N_11461,N_10970,N_10894);
nor U11462 (N_11462,N_11340,N_11053);
xor U11463 (N_11463,N_11018,N_11006);
and U11464 (N_11464,N_11178,N_11111);
or U11465 (N_11465,N_11181,N_11173);
xnor U11466 (N_11466,N_10965,N_11312);
nor U11467 (N_11467,N_10995,N_11300);
nor U11468 (N_11468,N_11090,N_10811);
or U11469 (N_11469,N_11236,N_11192);
or U11470 (N_11470,N_10824,N_11103);
or U11471 (N_11471,N_11217,N_11171);
nor U11472 (N_11472,N_11311,N_11303);
xor U11473 (N_11473,N_11381,N_10857);
xnor U11474 (N_11474,N_11309,N_11329);
or U11475 (N_11475,N_11248,N_11284);
and U11476 (N_11476,N_10845,N_11327);
and U11477 (N_11477,N_11167,N_10890);
nand U11478 (N_11478,N_10803,N_11195);
and U11479 (N_11479,N_10927,N_11266);
or U11480 (N_11480,N_11330,N_11206);
and U11481 (N_11481,N_10818,N_11183);
or U11482 (N_11482,N_10952,N_11384);
or U11483 (N_11483,N_11280,N_11320);
or U11484 (N_11484,N_11121,N_10939);
nand U11485 (N_11485,N_11083,N_10870);
xnor U11486 (N_11486,N_10855,N_11374);
xnor U11487 (N_11487,N_11142,N_11108);
and U11488 (N_11488,N_11077,N_11198);
and U11489 (N_11489,N_10836,N_11234);
or U11490 (N_11490,N_11353,N_11185);
nand U11491 (N_11491,N_11354,N_11134);
nand U11492 (N_11492,N_10964,N_11216);
xor U11493 (N_11493,N_11383,N_11220);
or U11494 (N_11494,N_11110,N_11197);
and U11495 (N_11495,N_11323,N_10993);
and U11496 (N_11496,N_11060,N_11025);
nand U11497 (N_11497,N_10896,N_11325);
or U11498 (N_11498,N_11267,N_11375);
xor U11499 (N_11499,N_11237,N_11337);
nor U11500 (N_11500,N_11050,N_11052);
or U11501 (N_11501,N_11047,N_11398);
nor U11502 (N_11502,N_11127,N_11289);
nor U11503 (N_11503,N_10977,N_10873);
or U11504 (N_11504,N_11378,N_11049);
nor U11505 (N_11505,N_10982,N_10807);
nor U11506 (N_11506,N_11145,N_11211);
nand U11507 (N_11507,N_10909,N_11363);
nor U11508 (N_11508,N_11209,N_10916);
nand U11509 (N_11509,N_10859,N_11308);
and U11510 (N_11510,N_11273,N_10861);
or U11511 (N_11511,N_11076,N_11393);
nor U11512 (N_11512,N_11369,N_10912);
xnor U11513 (N_11513,N_11017,N_11336);
and U11514 (N_11514,N_11345,N_11085);
and U11515 (N_11515,N_11346,N_11118);
and U11516 (N_11516,N_11022,N_11086);
nand U11517 (N_11517,N_11222,N_11045);
nor U11518 (N_11518,N_10962,N_11057);
xor U11519 (N_11519,N_11115,N_10954);
and U11520 (N_11520,N_10886,N_11159);
nand U11521 (N_11521,N_11321,N_11304);
nor U11522 (N_11522,N_11314,N_11287);
and U11523 (N_11523,N_10860,N_11109);
or U11524 (N_11524,N_11079,N_11116);
or U11525 (N_11525,N_11044,N_10808);
and U11526 (N_11526,N_11051,N_10866);
nor U11527 (N_11527,N_11188,N_10806);
nor U11528 (N_11528,N_11317,N_11227);
and U11529 (N_11529,N_10887,N_11335);
nand U11530 (N_11530,N_11093,N_11348);
or U11531 (N_11531,N_11352,N_11032);
nor U11532 (N_11532,N_11361,N_11379);
nor U11533 (N_11533,N_10915,N_10834);
xor U11534 (N_11534,N_11290,N_11260);
nand U11535 (N_11535,N_11184,N_11283);
nor U11536 (N_11536,N_10957,N_11041);
nor U11537 (N_11537,N_10959,N_11164);
nor U11538 (N_11538,N_10949,N_11131);
nand U11539 (N_11539,N_11269,N_10863);
or U11540 (N_11540,N_11010,N_10972);
xor U11541 (N_11541,N_10941,N_11301);
nand U11542 (N_11542,N_11136,N_10953);
xnor U11543 (N_11543,N_10978,N_11072);
nand U11544 (N_11544,N_11265,N_11043);
xor U11545 (N_11545,N_11229,N_11038);
nor U11546 (N_11546,N_11278,N_11396);
or U11547 (N_11547,N_11364,N_10958);
xnor U11548 (N_11548,N_11245,N_10801);
and U11549 (N_11549,N_11141,N_11214);
xnor U11550 (N_11550,N_10891,N_11228);
or U11551 (N_11551,N_11298,N_10843);
or U11552 (N_11552,N_11007,N_11186);
or U11553 (N_11553,N_11146,N_11333);
and U11554 (N_11554,N_11023,N_11122);
or U11555 (N_11555,N_10911,N_11084);
nor U11556 (N_11556,N_11373,N_10874);
nand U11557 (N_11557,N_11395,N_11069);
or U11558 (N_11558,N_11114,N_11068);
and U11559 (N_11559,N_11231,N_11254);
and U11560 (N_11560,N_11291,N_10928);
xnor U11561 (N_11561,N_11190,N_11215);
and U11562 (N_11562,N_11326,N_11039);
xor U11563 (N_11563,N_11262,N_10823);
nand U11564 (N_11564,N_11238,N_11177);
and U11565 (N_11565,N_11119,N_11073);
nand U11566 (N_11566,N_10826,N_11169);
xnor U11567 (N_11567,N_11061,N_11056);
or U11568 (N_11568,N_10994,N_10947);
nor U11569 (N_11569,N_11233,N_11034);
or U11570 (N_11570,N_10828,N_10844);
xor U11571 (N_11571,N_11288,N_10838);
xnor U11572 (N_11572,N_11358,N_11002);
nand U11573 (N_11573,N_10901,N_11213);
or U11574 (N_11574,N_11104,N_10950);
nor U11575 (N_11575,N_11021,N_10902);
or U11576 (N_11576,N_10983,N_10985);
xor U11577 (N_11577,N_10846,N_11355);
nor U11578 (N_11578,N_10932,N_10816);
nand U11579 (N_11579,N_11055,N_10805);
nand U11580 (N_11580,N_11133,N_10903);
nand U11581 (N_11581,N_11033,N_11126);
xnor U11582 (N_11582,N_11276,N_11344);
nor U11583 (N_11583,N_11386,N_10943);
and U11584 (N_11584,N_11054,N_10997);
xnor U11585 (N_11585,N_11135,N_11307);
nand U11586 (N_11586,N_11070,N_10867);
xor U11587 (N_11587,N_10868,N_10815);
nand U11588 (N_11588,N_11322,N_10862);
or U11589 (N_11589,N_11390,N_10931);
nand U11590 (N_11590,N_10937,N_11275);
xnor U11591 (N_11591,N_11315,N_10968);
nor U11592 (N_11592,N_11129,N_11362);
or U11593 (N_11593,N_11334,N_10882);
nand U11594 (N_11594,N_11099,N_11153);
nand U11595 (N_11595,N_11207,N_11005);
nor U11596 (N_11596,N_11028,N_10918);
nand U11597 (N_11597,N_10961,N_11095);
or U11598 (N_11598,N_11163,N_11392);
nand U11599 (N_11599,N_11221,N_11258);
xnor U11600 (N_11600,N_10871,N_11365);
or U11601 (N_11601,N_11203,N_11071);
and U11602 (N_11602,N_11154,N_11080);
nor U11603 (N_11603,N_10921,N_11263);
xor U11604 (N_11604,N_11140,N_10956);
xor U11605 (N_11605,N_11031,N_11205);
nand U11606 (N_11606,N_11004,N_10839);
and U11607 (N_11607,N_11305,N_10854);
xnor U11608 (N_11608,N_11328,N_10934);
nand U11609 (N_11609,N_11150,N_11157);
and U11610 (N_11610,N_11020,N_11014);
nand U11611 (N_11611,N_11397,N_11235);
nor U11612 (N_11612,N_11008,N_11242);
or U11613 (N_11613,N_11012,N_11030);
or U11614 (N_11614,N_11170,N_11161);
nor U11615 (N_11615,N_10879,N_11096);
or U11616 (N_11616,N_10914,N_10966);
nor U11617 (N_11617,N_11058,N_11367);
nor U11618 (N_11618,N_11264,N_11149);
nand U11619 (N_11619,N_11168,N_10935);
or U11620 (N_11620,N_11387,N_11064);
nor U11621 (N_11621,N_10999,N_10876);
xnor U11622 (N_11622,N_11179,N_10922);
nor U11623 (N_11623,N_11204,N_11166);
and U11624 (N_11624,N_11091,N_11123);
xnor U11625 (N_11625,N_10820,N_10889);
xnor U11626 (N_11626,N_11331,N_11027);
or U11627 (N_11627,N_10991,N_11013);
and U11628 (N_11628,N_10849,N_11313);
nand U11629 (N_11629,N_11293,N_10810);
or U11630 (N_11630,N_11036,N_11098);
xnor U11631 (N_11631,N_11246,N_11394);
or U11632 (N_11632,N_11180,N_11274);
nand U11633 (N_11633,N_11226,N_10847);
and U11634 (N_11634,N_10904,N_11174);
nor U11635 (N_11635,N_11156,N_11165);
xor U11636 (N_11636,N_11241,N_10920);
or U11637 (N_11637,N_11162,N_11389);
nor U11638 (N_11638,N_11388,N_10979);
nand U11639 (N_11639,N_10848,N_11316);
nor U11640 (N_11640,N_11176,N_11268);
nand U11641 (N_11641,N_11155,N_11255);
xor U11642 (N_11642,N_11282,N_10831);
nor U11643 (N_11643,N_10975,N_10913);
and U11644 (N_11644,N_10833,N_11286);
nand U11645 (N_11645,N_11191,N_11230);
nor U11646 (N_11646,N_10851,N_10981);
or U11647 (N_11647,N_11347,N_10923);
nor U11648 (N_11648,N_10880,N_10930);
xnor U11649 (N_11649,N_11016,N_11158);
and U11650 (N_11650,N_10837,N_10936);
nor U11651 (N_11651,N_10822,N_11310);
xnor U11652 (N_11652,N_11106,N_10955);
and U11653 (N_11653,N_11257,N_10800);
or U11654 (N_11654,N_11074,N_10976);
nor U11655 (N_11655,N_11130,N_10908);
or U11656 (N_11656,N_11026,N_11239);
nand U11657 (N_11657,N_11194,N_11377);
nand U11658 (N_11658,N_11199,N_11015);
or U11659 (N_11659,N_11338,N_10910);
and U11660 (N_11660,N_11202,N_10817);
xor U11661 (N_11661,N_11078,N_11292);
xor U11662 (N_11662,N_10881,N_11097);
nand U11663 (N_11663,N_11281,N_11187);
xor U11664 (N_11664,N_11244,N_11147);
and U11665 (N_11665,N_10971,N_10986);
and U11666 (N_11666,N_11277,N_11259);
nand U11667 (N_11667,N_11371,N_11223);
and U11668 (N_11668,N_11112,N_10969);
and U11669 (N_11669,N_11296,N_11189);
or U11670 (N_11670,N_11299,N_11380);
or U11671 (N_11671,N_10858,N_11318);
nand U11672 (N_11672,N_10840,N_10819);
or U11673 (N_11673,N_11341,N_11225);
xnor U11674 (N_11674,N_11087,N_11137);
xor U11675 (N_11675,N_11172,N_10942);
nor U11676 (N_11676,N_11125,N_10802);
or U11677 (N_11677,N_11082,N_11391);
nor U11678 (N_11678,N_11175,N_10850);
or U11679 (N_11679,N_10988,N_11372);
xor U11680 (N_11680,N_11065,N_10829);
nand U11681 (N_11681,N_11144,N_11272);
nand U11682 (N_11682,N_11000,N_11210);
or U11683 (N_11683,N_11120,N_11243);
or U11684 (N_11684,N_10883,N_11212);
nand U11685 (N_11685,N_11319,N_10925);
xnor U11686 (N_11686,N_10841,N_11385);
and U11687 (N_11687,N_11132,N_11256);
and U11688 (N_11688,N_11035,N_11148);
and U11689 (N_11689,N_10825,N_11139);
nor U11690 (N_11690,N_10974,N_11232);
xnor U11691 (N_11691,N_11366,N_11342);
xnor U11692 (N_11692,N_11088,N_11295);
nor U11693 (N_11693,N_10938,N_11107);
nand U11694 (N_11694,N_10869,N_11376);
nor U11695 (N_11695,N_10963,N_10884);
and U11696 (N_11696,N_10967,N_11003);
xnor U11697 (N_11697,N_11370,N_11279);
nor U11698 (N_11698,N_10929,N_11001);
xor U11699 (N_11699,N_11208,N_11092);
or U11700 (N_11700,N_11065,N_10814);
nor U11701 (N_11701,N_11254,N_11377);
nand U11702 (N_11702,N_10979,N_11156);
and U11703 (N_11703,N_11206,N_10984);
nand U11704 (N_11704,N_10846,N_11331);
xnor U11705 (N_11705,N_10906,N_11308);
nor U11706 (N_11706,N_10987,N_11109);
nand U11707 (N_11707,N_11342,N_10947);
nor U11708 (N_11708,N_11161,N_11151);
or U11709 (N_11709,N_11107,N_11099);
xor U11710 (N_11710,N_10904,N_11044);
and U11711 (N_11711,N_11000,N_11026);
nand U11712 (N_11712,N_11354,N_11048);
xnor U11713 (N_11713,N_11020,N_10993);
nor U11714 (N_11714,N_11069,N_10926);
nand U11715 (N_11715,N_11108,N_11168);
and U11716 (N_11716,N_11350,N_10975);
nand U11717 (N_11717,N_11306,N_11032);
xor U11718 (N_11718,N_11275,N_11379);
nand U11719 (N_11719,N_11308,N_11210);
and U11720 (N_11720,N_11213,N_11097);
or U11721 (N_11721,N_11261,N_11271);
and U11722 (N_11722,N_11280,N_11334);
xor U11723 (N_11723,N_11243,N_11296);
nand U11724 (N_11724,N_11259,N_11340);
nand U11725 (N_11725,N_11117,N_11235);
and U11726 (N_11726,N_10857,N_10982);
nand U11727 (N_11727,N_11250,N_11090);
or U11728 (N_11728,N_11091,N_11219);
nand U11729 (N_11729,N_11389,N_11221);
or U11730 (N_11730,N_10893,N_11242);
and U11731 (N_11731,N_10914,N_11172);
xnor U11732 (N_11732,N_11196,N_10889);
xnor U11733 (N_11733,N_11375,N_10860);
or U11734 (N_11734,N_11052,N_11313);
and U11735 (N_11735,N_11096,N_11200);
and U11736 (N_11736,N_11000,N_11079);
xnor U11737 (N_11737,N_11212,N_10902);
or U11738 (N_11738,N_11070,N_11098);
nor U11739 (N_11739,N_11126,N_10856);
and U11740 (N_11740,N_11386,N_11344);
xor U11741 (N_11741,N_10942,N_11179);
or U11742 (N_11742,N_10974,N_11030);
and U11743 (N_11743,N_11096,N_11347);
and U11744 (N_11744,N_11137,N_11188);
nand U11745 (N_11745,N_11122,N_11010);
nand U11746 (N_11746,N_10953,N_11233);
or U11747 (N_11747,N_10809,N_11122);
nand U11748 (N_11748,N_11190,N_11094);
nand U11749 (N_11749,N_11154,N_11305);
nand U11750 (N_11750,N_11194,N_11150);
nor U11751 (N_11751,N_10970,N_10865);
and U11752 (N_11752,N_10937,N_10889);
nand U11753 (N_11753,N_11291,N_11330);
nor U11754 (N_11754,N_10900,N_10902);
or U11755 (N_11755,N_11356,N_11242);
nand U11756 (N_11756,N_11181,N_11388);
or U11757 (N_11757,N_10885,N_10902);
or U11758 (N_11758,N_11232,N_11034);
and U11759 (N_11759,N_11258,N_11091);
or U11760 (N_11760,N_11187,N_11061);
or U11761 (N_11761,N_11252,N_11112);
nor U11762 (N_11762,N_11336,N_11060);
nand U11763 (N_11763,N_11100,N_10985);
nand U11764 (N_11764,N_11120,N_11206);
and U11765 (N_11765,N_11263,N_11179);
or U11766 (N_11766,N_11049,N_10931);
nor U11767 (N_11767,N_11169,N_10892);
nand U11768 (N_11768,N_10855,N_11164);
xnor U11769 (N_11769,N_10991,N_11291);
nor U11770 (N_11770,N_11154,N_11208);
or U11771 (N_11771,N_11040,N_11363);
xnor U11772 (N_11772,N_10878,N_10999);
or U11773 (N_11773,N_10898,N_11399);
and U11774 (N_11774,N_10988,N_11289);
nor U11775 (N_11775,N_11370,N_10907);
and U11776 (N_11776,N_10844,N_10938);
and U11777 (N_11777,N_11267,N_11049);
or U11778 (N_11778,N_11015,N_11333);
xor U11779 (N_11779,N_11148,N_10953);
nor U11780 (N_11780,N_10983,N_11099);
xnor U11781 (N_11781,N_11388,N_11047);
nand U11782 (N_11782,N_11184,N_10846);
nor U11783 (N_11783,N_11209,N_10830);
xor U11784 (N_11784,N_11290,N_11295);
nand U11785 (N_11785,N_10889,N_10855);
and U11786 (N_11786,N_10849,N_11302);
or U11787 (N_11787,N_10829,N_11357);
or U11788 (N_11788,N_10998,N_11366);
nor U11789 (N_11789,N_10994,N_11271);
nand U11790 (N_11790,N_11110,N_10953);
nand U11791 (N_11791,N_11033,N_11203);
xnor U11792 (N_11792,N_10960,N_10859);
or U11793 (N_11793,N_10882,N_11211);
or U11794 (N_11794,N_11143,N_10833);
and U11795 (N_11795,N_10888,N_11092);
and U11796 (N_11796,N_11053,N_11146);
nand U11797 (N_11797,N_11099,N_11132);
xor U11798 (N_11798,N_10983,N_10930);
nand U11799 (N_11799,N_11134,N_10996);
xor U11800 (N_11800,N_10814,N_11245);
xor U11801 (N_11801,N_11166,N_10843);
nand U11802 (N_11802,N_11073,N_11142);
nor U11803 (N_11803,N_11329,N_11303);
xor U11804 (N_11804,N_11364,N_10941);
nor U11805 (N_11805,N_11311,N_11230);
and U11806 (N_11806,N_11125,N_11337);
nor U11807 (N_11807,N_11303,N_10832);
or U11808 (N_11808,N_11140,N_11278);
nand U11809 (N_11809,N_11390,N_10912);
and U11810 (N_11810,N_10811,N_11389);
nor U11811 (N_11811,N_10840,N_11026);
nor U11812 (N_11812,N_11085,N_10923);
xnor U11813 (N_11813,N_11172,N_11164);
nand U11814 (N_11814,N_10871,N_11288);
or U11815 (N_11815,N_10818,N_11287);
and U11816 (N_11816,N_11266,N_11281);
nand U11817 (N_11817,N_11236,N_10849);
nor U11818 (N_11818,N_10942,N_11275);
and U11819 (N_11819,N_11204,N_11133);
nor U11820 (N_11820,N_11121,N_11026);
xnor U11821 (N_11821,N_10923,N_11250);
nand U11822 (N_11822,N_11024,N_11392);
and U11823 (N_11823,N_11307,N_11154);
xnor U11824 (N_11824,N_10805,N_10816);
nand U11825 (N_11825,N_11298,N_10989);
nand U11826 (N_11826,N_11058,N_11285);
nand U11827 (N_11827,N_10816,N_10920);
nand U11828 (N_11828,N_11110,N_11320);
and U11829 (N_11829,N_11237,N_10822);
nand U11830 (N_11830,N_11076,N_11003);
or U11831 (N_11831,N_10963,N_11120);
nand U11832 (N_11832,N_11049,N_10885);
nor U11833 (N_11833,N_10903,N_11377);
xnor U11834 (N_11834,N_11306,N_11023);
or U11835 (N_11835,N_10882,N_11020);
xnor U11836 (N_11836,N_10890,N_11018);
and U11837 (N_11837,N_11355,N_11050);
xnor U11838 (N_11838,N_10883,N_10870);
and U11839 (N_11839,N_10928,N_10897);
and U11840 (N_11840,N_11100,N_10972);
nand U11841 (N_11841,N_10852,N_11188);
or U11842 (N_11842,N_10829,N_11291);
nor U11843 (N_11843,N_10893,N_10843);
xnor U11844 (N_11844,N_11021,N_11183);
and U11845 (N_11845,N_10890,N_11184);
and U11846 (N_11846,N_11008,N_11138);
nor U11847 (N_11847,N_11139,N_11340);
nor U11848 (N_11848,N_10814,N_10934);
and U11849 (N_11849,N_10991,N_10899);
or U11850 (N_11850,N_10943,N_10821);
and U11851 (N_11851,N_11166,N_11031);
nand U11852 (N_11852,N_10818,N_11209);
xnor U11853 (N_11853,N_11119,N_11080);
nor U11854 (N_11854,N_10812,N_11278);
nor U11855 (N_11855,N_10897,N_11162);
nand U11856 (N_11856,N_11152,N_11256);
nand U11857 (N_11857,N_11353,N_10922);
nand U11858 (N_11858,N_11011,N_11147);
nor U11859 (N_11859,N_11100,N_10980);
or U11860 (N_11860,N_11142,N_10813);
or U11861 (N_11861,N_11395,N_11140);
nand U11862 (N_11862,N_11268,N_10912);
xor U11863 (N_11863,N_10919,N_11223);
or U11864 (N_11864,N_10894,N_10810);
and U11865 (N_11865,N_10992,N_10899);
nor U11866 (N_11866,N_10840,N_10927);
xnor U11867 (N_11867,N_11212,N_11216);
and U11868 (N_11868,N_11151,N_11322);
or U11869 (N_11869,N_11328,N_11388);
and U11870 (N_11870,N_11298,N_11006);
and U11871 (N_11871,N_11279,N_11376);
nand U11872 (N_11872,N_10968,N_10964);
nand U11873 (N_11873,N_10825,N_11147);
and U11874 (N_11874,N_11136,N_10952);
and U11875 (N_11875,N_10879,N_11229);
and U11876 (N_11876,N_11022,N_10998);
nand U11877 (N_11877,N_10948,N_11013);
xnor U11878 (N_11878,N_10926,N_10966);
or U11879 (N_11879,N_11384,N_11023);
nor U11880 (N_11880,N_10890,N_10972);
nand U11881 (N_11881,N_11129,N_11054);
and U11882 (N_11882,N_11188,N_11146);
or U11883 (N_11883,N_11340,N_11378);
and U11884 (N_11884,N_10872,N_10932);
xnor U11885 (N_11885,N_10948,N_11257);
and U11886 (N_11886,N_11257,N_10828);
nor U11887 (N_11887,N_11284,N_10868);
nand U11888 (N_11888,N_11226,N_10893);
nor U11889 (N_11889,N_11188,N_11281);
nand U11890 (N_11890,N_11234,N_11150);
xnor U11891 (N_11891,N_11000,N_10831);
nor U11892 (N_11892,N_11052,N_11356);
or U11893 (N_11893,N_11286,N_11273);
xnor U11894 (N_11894,N_10917,N_11331);
nor U11895 (N_11895,N_11239,N_11340);
nor U11896 (N_11896,N_11007,N_11299);
or U11897 (N_11897,N_11356,N_11272);
nor U11898 (N_11898,N_11131,N_11004);
and U11899 (N_11899,N_11133,N_10876);
and U11900 (N_11900,N_10994,N_10911);
nor U11901 (N_11901,N_10887,N_11004);
or U11902 (N_11902,N_11049,N_11311);
nand U11903 (N_11903,N_11038,N_11179);
xor U11904 (N_11904,N_11188,N_11147);
xor U11905 (N_11905,N_10984,N_11042);
xor U11906 (N_11906,N_11030,N_11219);
and U11907 (N_11907,N_11344,N_11054);
and U11908 (N_11908,N_11245,N_11121);
nor U11909 (N_11909,N_10835,N_11237);
nor U11910 (N_11910,N_11064,N_11190);
nor U11911 (N_11911,N_11022,N_10866);
and U11912 (N_11912,N_11015,N_11232);
or U11913 (N_11913,N_10805,N_11136);
and U11914 (N_11914,N_11189,N_11040);
nor U11915 (N_11915,N_11399,N_11374);
nand U11916 (N_11916,N_11095,N_10917);
xnor U11917 (N_11917,N_11315,N_11299);
xnor U11918 (N_11918,N_11114,N_10903);
and U11919 (N_11919,N_11121,N_10912);
nor U11920 (N_11920,N_10813,N_11384);
or U11921 (N_11921,N_11258,N_10890);
nand U11922 (N_11922,N_10852,N_11279);
or U11923 (N_11923,N_11030,N_11337);
nor U11924 (N_11924,N_10989,N_11393);
or U11925 (N_11925,N_10989,N_11276);
nor U11926 (N_11926,N_10878,N_10833);
xor U11927 (N_11927,N_10994,N_11342);
xnor U11928 (N_11928,N_10914,N_11175);
or U11929 (N_11929,N_11147,N_11065);
or U11930 (N_11930,N_10873,N_11017);
or U11931 (N_11931,N_11145,N_11225);
and U11932 (N_11932,N_11068,N_11116);
or U11933 (N_11933,N_11012,N_11140);
nor U11934 (N_11934,N_11247,N_11397);
xnor U11935 (N_11935,N_11057,N_11246);
xor U11936 (N_11936,N_10876,N_10968);
nand U11937 (N_11937,N_10877,N_10806);
nor U11938 (N_11938,N_10941,N_11231);
or U11939 (N_11939,N_11210,N_10987);
nor U11940 (N_11940,N_10967,N_11253);
nand U11941 (N_11941,N_11163,N_11158);
and U11942 (N_11942,N_11203,N_11252);
nor U11943 (N_11943,N_11241,N_11369);
or U11944 (N_11944,N_10900,N_11323);
nand U11945 (N_11945,N_11038,N_10812);
xnor U11946 (N_11946,N_11333,N_11027);
nand U11947 (N_11947,N_11237,N_11227);
nor U11948 (N_11948,N_10814,N_11187);
and U11949 (N_11949,N_10811,N_11384);
xor U11950 (N_11950,N_10958,N_10875);
and U11951 (N_11951,N_11022,N_11180);
and U11952 (N_11952,N_11211,N_10859);
nor U11953 (N_11953,N_11010,N_11111);
or U11954 (N_11954,N_11293,N_11016);
or U11955 (N_11955,N_10822,N_11086);
nand U11956 (N_11956,N_11192,N_10823);
xor U11957 (N_11957,N_10980,N_11047);
nand U11958 (N_11958,N_10923,N_11387);
nand U11959 (N_11959,N_11355,N_10873);
or U11960 (N_11960,N_11123,N_10916);
nor U11961 (N_11961,N_10909,N_11007);
and U11962 (N_11962,N_10864,N_11125);
or U11963 (N_11963,N_11361,N_10809);
and U11964 (N_11964,N_10940,N_11267);
nand U11965 (N_11965,N_10992,N_11279);
nand U11966 (N_11966,N_10845,N_11142);
xor U11967 (N_11967,N_11396,N_11133);
and U11968 (N_11968,N_10819,N_10981);
nand U11969 (N_11969,N_10851,N_10945);
and U11970 (N_11970,N_11160,N_11075);
and U11971 (N_11971,N_10897,N_11393);
xnor U11972 (N_11972,N_10943,N_11219);
xor U11973 (N_11973,N_10900,N_10896);
or U11974 (N_11974,N_11018,N_11285);
xnor U11975 (N_11975,N_10807,N_10873);
nand U11976 (N_11976,N_11073,N_10992);
nor U11977 (N_11977,N_11371,N_11121);
and U11978 (N_11978,N_11051,N_11273);
nor U11979 (N_11979,N_10821,N_11130);
nand U11980 (N_11980,N_10978,N_11029);
and U11981 (N_11981,N_11057,N_11068);
nor U11982 (N_11982,N_11212,N_10897);
or U11983 (N_11983,N_11107,N_10825);
and U11984 (N_11984,N_10917,N_11220);
nor U11985 (N_11985,N_11081,N_11216);
and U11986 (N_11986,N_11007,N_11330);
nor U11987 (N_11987,N_10821,N_11187);
and U11988 (N_11988,N_10964,N_11342);
xor U11989 (N_11989,N_11365,N_10804);
nor U11990 (N_11990,N_11121,N_11356);
xnor U11991 (N_11991,N_11109,N_11183);
and U11992 (N_11992,N_11289,N_10861);
nand U11993 (N_11993,N_10817,N_11307);
and U11994 (N_11994,N_11166,N_11289);
and U11995 (N_11995,N_11217,N_10984);
or U11996 (N_11996,N_11240,N_11166);
and U11997 (N_11997,N_11122,N_10963);
nor U11998 (N_11998,N_10885,N_11279);
and U11999 (N_11999,N_11258,N_10963);
or U12000 (N_12000,N_11452,N_11613);
or U12001 (N_12001,N_11717,N_11701);
or U12002 (N_12002,N_11818,N_11893);
xor U12003 (N_12003,N_11736,N_11415);
or U12004 (N_12004,N_11669,N_11885);
xnor U12005 (N_12005,N_11878,N_11605);
nor U12006 (N_12006,N_11460,N_11611);
nor U12007 (N_12007,N_11903,N_11985);
or U12008 (N_12008,N_11989,N_11779);
or U12009 (N_12009,N_11775,N_11913);
nand U12010 (N_12010,N_11550,N_11483);
nor U12011 (N_12011,N_11479,N_11868);
xnor U12012 (N_12012,N_11651,N_11525);
nand U12013 (N_12013,N_11936,N_11750);
xor U12014 (N_12014,N_11951,N_11658);
and U12015 (N_12015,N_11730,N_11741);
and U12016 (N_12016,N_11875,N_11752);
or U12017 (N_12017,N_11497,N_11964);
or U12018 (N_12018,N_11558,N_11708);
nand U12019 (N_12019,N_11765,N_11599);
nor U12020 (N_12020,N_11512,N_11952);
or U12021 (N_12021,N_11932,N_11542);
and U12022 (N_12022,N_11766,N_11592);
or U12023 (N_12023,N_11958,N_11480);
or U12024 (N_12024,N_11482,N_11748);
and U12025 (N_12025,N_11873,N_11762);
nor U12026 (N_12026,N_11834,N_11530);
xor U12027 (N_12027,N_11824,N_11821);
xnor U12028 (N_12028,N_11612,N_11674);
nand U12029 (N_12029,N_11901,N_11724);
nor U12030 (N_12030,N_11865,N_11880);
nand U12031 (N_12031,N_11648,N_11683);
xnor U12032 (N_12032,N_11891,N_11892);
nand U12033 (N_12033,N_11496,N_11929);
xnor U12034 (N_12034,N_11538,N_11641);
or U12035 (N_12035,N_11581,N_11511);
nor U12036 (N_12036,N_11737,N_11809);
and U12037 (N_12037,N_11950,N_11709);
and U12038 (N_12038,N_11907,N_11746);
xnor U12039 (N_12039,N_11793,N_11478);
or U12040 (N_12040,N_11920,N_11516);
or U12041 (N_12041,N_11532,N_11491);
nor U12042 (N_12042,N_11976,N_11505);
xor U12043 (N_12043,N_11606,N_11998);
nor U12044 (N_12044,N_11947,N_11515);
nand U12045 (N_12045,N_11797,N_11799);
and U12046 (N_12046,N_11690,N_11441);
or U12047 (N_12047,N_11977,N_11785);
nor U12048 (N_12048,N_11859,N_11796);
nand U12049 (N_12049,N_11753,N_11722);
nor U12050 (N_12050,N_11575,N_11484);
and U12051 (N_12051,N_11853,N_11771);
or U12052 (N_12052,N_11840,N_11904);
or U12053 (N_12053,N_11405,N_11414);
xor U12054 (N_12054,N_11798,N_11548);
and U12055 (N_12055,N_11992,N_11576);
xor U12056 (N_12056,N_11691,N_11634);
or U12057 (N_12057,N_11468,N_11996);
xor U12058 (N_12058,N_11774,N_11833);
nand U12059 (N_12059,N_11828,N_11778);
nand U12060 (N_12060,N_11896,N_11434);
nor U12061 (N_12061,N_11650,N_11458);
and U12062 (N_12062,N_11430,N_11973);
and U12063 (N_12063,N_11409,N_11697);
xnor U12064 (N_12064,N_11849,N_11623);
nand U12065 (N_12065,N_11805,N_11566);
nand U12066 (N_12066,N_11624,N_11935);
xnor U12067 (N_12067,N_11573,N_11933);
or U12068 (N_12068,N_11732,N_11693);
xor U12069 (N_12069,N_11858,N_11463);
and U12070 (N_12070,N_11960,N_11584);
and U12071 (N_12071,N_11789,N_11703);
or U12072 (N_12072,N_11632,N_11751);
and U12073 (N_12073,N_11604,N_11467);
nand U12074 (N_12074,N_11676,N_11991);
and U12075 (N_12075,N_11879,N_11817);
nand U12076 (N_12076,N_11617,N_11871);
or U12077 (N_12077,N_11881,N_11787);
or U12078 (N_12078,N_11686,N_11403);
and U12079 (N_12079,N_11546,N_11522);
or U12080 (N_12080,N_11735,N_11850);
and U12081 (N_12081,N_11924,N_11614);
nand U12082 (N_12082,N_11493,N_11551);
or U12083 (N_12083,N_11547,N_11925);
and U12084 (N_12084,N_11439,N_11602);
and U12085 (N_12085,N_11677,N_11969);
or U12086 (N_12086,N_11743,N_11968);
nor U12087 (N_12087,N_11541,N_11580);
nand U12088 (N_12088,N_11569,N_11436);
nor U12089 (N_12089,N_11510,N_11930);
nand U12090 (N_12090,N_11984,N_11459);
xnor U12091 (N_12091,N_11595,N_11823);
and U12092 (N_12092,N_11812,N_11464);
or U12093 (N_12093,N_11927,N_11715);
or U12094 (N_12094,N_11504,N_11555);
xor U12095 (N_12095,N_11666,N_11656);
nand U12096 (N_12096,N_11433,N_11781);
xor U12097 (N_12097,N_11987,N_11419);
nand U12098 (N_12098,N_11861,N_11431);
nand U12099 (N_12099,N_11937,N_11682);
nand U12100 (N_12100,N_11445,N_11972);
and U12101 (N_12101,N_11627,N_11931);
or U12102 (N_12102,N_11589,N_11685);
or U12103 (N_12103,N_11745,N_11792);
xor U12104 (N_12104,N_11727,N_11601);
nand U12105 (N_12105,N_11842,N_11990);
nor U12106 (N_12106,N_11596,N_11600);
nand U12107 (N_12107,N_11928,N_11883);
nand U12108 (N_12108,N_11640,N_11456);
nand U12109 (N_12109,N_11945,N_11501);
nand U12110 (N_12110,N_11450,N_11738);
nor U12111 (N_12111,N_11417,N_11832);
and U12112 (N_12112,N_11477,N_11628);
xor U12113 (N_12113,N_11609,N_11747);
xor U12114 (N_12114,N_11435,N_11837);
xnor U12115 (N_12115,N_11949,N_11923);
and U12116 (N_12116,N_11487,N_11572);
nor U12117 (N_12117,N_11783,N_11938);
xor U12118 (N_12118,N_11437,N_11876);
nor U12119 (N_12119,N_11588,N_11440);
or U12120 (N_12120,N_11673,N_11570);
or U12121 (N_12121,N_11653,N_11788);
and U12122 (N_12122,N_11618,N_11702);
xor U12123 (N_12123,N_11506,N_11919);
nor U12124 (N_12124,N_11637,N_11654);
or U12125 (N_12125,N_11536,N_11803);
xnor U12126 (N_12126,N_11744,N_11442);
and U12127 (N_12127,N_11723,N_11784);
and U12128 (N_12128,N_11585,N_11946);
and U12129 (N_12129,N_11539,N_11975);
and U12130 (N_12130,N_11999,N_11769);
nor U12131 (N_12131,N_11644,N_11524);
xnor U12132 (N_12132,N_11986,N_11594);
xor U12133 (N_12133,N_11528,N_11866);
or U12134 (N_12134,N_11942,N_11791);
and U12135 (N_12135,N_11995,N_11438);
or U12136 (N_12136,N_11465,N_11616);
or U12137 (N_12137,N_11782,N_11647);
and U12138 (N_12138,N_11767,N_11763);
nand U12139 (N_12139,N_11667,N_11869);
nor U12140 (N_12140,N_11508,N_11894);
xor U12141 (N_12141,N_11681,N_11704);
nand U12142 (N_12142,N_11802,N_11513);
xor U12143 (N_12143,N_11423,N_11944);
xnor U12144 (N_12144,N_11527,N_11485);
nand U12145 (N_12145,N_11620,N_11714);
xor U12146 (N_12146,N_11490,N_11526);
nor U12147 (N_12147,N_11655,N_11446);
and U12148 (N_12148,N_11979,N_11926);
or U12149 (N_12149,N_11954,N_11461);
nor U12150 (N_12150,N_11489,N_11915);
and U12151 (N_12151,N_11671,N_11448);
or U12152 (N_12152,N_11810,N_11672);
and U12153 (N_12153,N_11475,N_11696);
nand U12154 (N_12154,N_11549,N_11529);
xnor U12155 (N_12155,N_11565,N_11670);
nand U12156 (N_12156,N_11854,N_11401);
or U12157 (N_12157,N_11642,N_11556);
nor U12158 (N_12158,N_11710,N_11568);
nand U12159 (N_12159,N_11827,N_11728);
nand U12160 (N_12160,N_11740,N_11684);
nor U12161 (N_12161,N_11971,N_11662);
nor U12162 (N_12162,N_11811,N_11520);
xnor U12163 (N_12163,N_11564,N_11813);
nor U12164 (N_12164,N_11453,N_11786);
xnor U12165 (N_12165,N_11416,N_11909);
nor U12166 (N_12166,N_11980,N_11961);
and U12167 (N_12167,N_11498,N_11957);
or U12168 (N_12168,N_11940,N_11941);
or U12169 (N_12169,N_11836,N_11993);
nand U12170 (N_12170,N_11918,N_11561);
xor U12171 (N_12171,N_11590,N_11507);
xor U12172 (N_12172,N_11706,N_11841);
or U12173 (N_12173,N_11820,N_11848);
xor U12174 (N_12174,N_11424,N_11872);
nand U12175 (N_12175,N_11754,N_11852);
xor U12176 (N_12176,N_11906,N_11649);
and U12177 (N_12177,N_11462,N_11553);
or U12178 (N_12178,N_11804,N_11695);
xor U12179 (N_12179,N_11898,N_11910);
and U12180 (N_12180,N_11959,N_11713);
or U12181 (N_12181,N_11420,N_11598);
and U12182 (N_12182,N_11429,N_11579);
xnor U12183 (N_12183,N_11877,N_11502);
and U12184 (N_12184,N_11406,N_11646);
nor U12185 (N_12185,N_11899,N_11408);
xnor U12186 (N_12186,N_11692,N_11659);
nor U12187 (N_12187,N_11770,N_11582);
and U12188 (N_12188,N_11567,N_11629);
nor U12189 (N_12189,N_11720,N_11756);
or U12190 (N_12190,N_11889,N_11800);
xnor U12191 (N_12191,N_11578,N_11657);
xnor U12192 (N_12192,N_11402,N_11794);
and U12193 (N_12193,N_11886,N_11470);
or U12194 (N_12194,N_11425,N_11939);
xor U12195 (N_12195,N_11608,N_11533);
nand U12196 (N_12196,N_11764,N_11523);
and U12197 (N_12197,N_11997,N_11635);
nand U12198 (N_12198,N_11801,N_11486);
or U12199 (N_12199,N_11739,N_11761);
nor U12200 (N_12200,N_11963,N_11822);
or U12201 (N_12201,N_11887,N_11807);
and U12202 (N_12202,N_11610,N_11413);
nand U12203 (N_12203,N_11543,N_11863);
xnor U12204 (N_12204,N_11689,N_11587);
xnor U12205 (N_12205,N_11934,N_11825);
and U12206 (N_12206,N_11457,N_11678);
or U12207 (N_12207,N_11661,N_11698);
nor U12208 (N_12208,N_11410,N_11521);
and U12209 (N_12209,N_11500,N_11772);
nand U12210 (N_12210,N_11687,N_11830);
nand U12211 (N_12211,N_11780,N_11535);
and U12212 (N_12212,N_11631,N_11922);
nor U12213 (N_12213,N_11711,N_11831);
nor U12214 (N_12214,N_11776,N_11974);
and U12215 (N_12215,N_11773,N_11843);
or U12216 (N_12216,N_11679,N_11574);
nor U12217 (N_12217,N_11994,N_11731);
xnor U12218 (N_12218,N_11897,N_11777);
nor U12219 (N_12219,N_11469,N_11603);
or U12220 (N_12220,N_11421,N_11426);
nand U12221 (N_12221,N_11943,N_11867);
xnor U12222 (N_12222,N_11829,N_11422);
and U12223 (N_12223,N_11492,N_11545);
or U12224 (N_12224,N_11912,N_11638);
nor U12225 (N_12225,N_11495,N_11953);
and U12226 (N_12226,N_11734,N_11808);
xnor U12227 (N_12227,N_11494,N_11680);
nand U12228 (N_12228,N_11760,N_11481);
and U12229 (N_12229,N_11514,N_11699);
nor U12230 (N_12230,N_11552,N_11956);
nand U12231 (N_12231,N_11844,N_11476);
or U12232 (N_12232,N_11725,N_11404);
nor U12233 (N_12233,N_11888,N_11726);
or U12234 (N_12234,N_11411,N_11643);
or U12235 (N_12235,N_11563,N_11583);
and U12236 (N_12236,N_11948,N_11607);
nor U12237 (N_12237,N_11597,N_11855);
or U12238 (N_12238,N_11593,N_11664);
xnor U12239 (N_12239,N_11428,N_11712);
or U12240 (N_12240,N_11472,N_11826);
nand U12241 (N_12241,N_11921,N_11874);
xnor U12242 (N_12242,N_11636,N_11839);
nand U12243 (N_12243,N_11729,N_11864);
xor U12244 (N_12244,N_11917,N_11432);
and U12245 (N_12245,N_11705,N_11845);
nor U12246 (N_12246,N_11733,N_11499);
xor U12247 (N_12247,N_11443,N_11718);
nor U12248 (N_12248,N_11619,N_11534);
nand U12249 (N_12249,N_11540,N_11455);
or U12250 (N_12250,N_11645,N_11652);
nor U12251 (N_12251,N_11882,N_11466);
or U12252 (N_12252,N_11795,N_11707);
nand U12253 (N_12253,N_11755,N_11815);
and U12254 (N_12254,N_11626,N_11473);
nor U12255 (N_12255,N_11970,N_11895);
and U12256 (N_12256,N_11471,N_11721);
nor U12257 (N_12257,N_11916,N_11966);
nand U12258 (N_12258,N_11571,N_11742);
nor U12259 (N_12259,N_11665,N_11838);
and U12260 (N_12260,N_11503,N_11562);
and U12261 (N_12261,N_11983,N_11819);
nor U12262 (N_12262,N_11517,N_11544);
nand U12263 (N_12263,N_11694,N_11860);
nand U12264 (N_12264,N_11625,N_11400);
nand U12265 (N_12265,N_11890,N_11790);
nor U12266 (N_12266,N_11630,N_11531);
xnor U12267 (N_12267,N_11768,N_11474);
or U12268 (N_12268,N_11757,N_11965);
nor U12269 (N_12269,N_11615,N_11719);
xor U12270 (N_12270,N_11978,N_11900);
xor U12271 (N_12271,N_11758,N_11700);
or U12272 (N_12272,N_11668,N_11908);
and U12273 (N_12273,N_11560,N_11982);
and U12274 (N_12274,N_11559,N_11519);
nand U12275 (N_12275,N_11577,N_11688);
and U12276 (N_12276,N_11988,N_11816);
or U12277 (N_12277,N_11902,N_11557);
nand U12278 (N_12278,N_11591,N_11884);
xor U12279 (N_12279,N_11835,N_11412);
or U12280 (N_12280,N_11454,N_11967);
nand U12281 (N_12281,N_11749,N_11846);
nand U12282 (N_12282,N_11862,N_11554);
nor U12283 (N_12283,N_11911,N_11814);
and U12284 (N_12284,N_11444,N_11451);
xnor U12285 (N_12285,N_11716,N_11806);
xor U12286 (N_12286,N_11488,N_11962);
or U12287 (N_12287,N_11639,N_11537);
nor U12288 (N_12288,N_11914,N_11981);
nand U12289 (N_12289,N_11759,N_11447);
nor U12290 (N_12290,N_11586,N_11857);
nor U12291 (N_12291,N_11622,N_11418);
xnor U12292 (N_12292,N_11621,N_11905);
and U12293 (N_12293,N_11870,N_11660);
nand U12294 (N_12294,N_11633,N_11675);
nand U12295 (N_12295,N_11955,N_11663);
or U12296 (N_12296,N_11518,N_11851);
and U12297 (N_12297,N_11427,N_11407);
or U12298 (N_12298,N_11847,N_11509);
xor U12299 (N_12299,N_11449,N_11856);
nor U12300 (N_12300,N_11769,N_11684);
xor U12301 (N_12301,N_11532,N_11626);
nor U12302 (N_12302,N_11544,N_11705);
and U12303 (N_12303,N_11535,N_11649);
and U12304 (N_12304,N_11925,N_11594);
and U12305 (N_12305,N_11699,N_11516);
xnor U12306 (N_12306,N_11847,N_11468);
and U12307 (N_12307,N_11839,N_11459);
or U12308 (N_12308,N_11498,N_11779);
or U12309 (N_12309,N_11685,N_11603);
nand U12310 (N_12310,N_11574,N_11618);
and U12311 (N_12311,N_11621,N_11408);
and U12312 (N_12312,N_11925,N_11619);
nand U12313 (N_12313,N_11843,N_11805);
xnor U12314 (N_12314,N_11961,N_11635);
nand U12315 (N_12315,N_11906,N_11606);
nand U12316 (N_12316,N_11456,N_11707);
nor U12317 (N_12317,N_11883,N_11984);
and U12318 (N_12318,N_11523,N_11732);
xor U12319 (N_12319,N_11679,N_11882);
xnor U12320 (N_12320,N_11852,N_11950);
xor U12321 (N_12321,N_11659,N_11857);
nand U12322 (N_12322,N_11589,N_11541);
and U12323 (N_12323,N_11664,N_11432);
or U12324 (N_12324,N_11842,N_11602);
nor U12325 (N_12325,N_11710,N_11964);
xnor U12326 (N_12326,N_11540,N_11429);
xnor U12327 (N_12327,N_11971,N_11899);
or U12328 (N_12328,N_11943,N_11524);
nor U12329 (N_12329,N_11959,N_11654);
xor U12330 (N_12330,N_11719,N_11729);
nor U12331 (N_12331,N_11892,N_11482);
nand U12332 (N_12332,N_11903,N_11887);
nor U12333 (N_12333,N_11843,N_11842);
or U12334 (N_12334,N_11547,N_11557);
xnor U12335 (N_12335,N_11726,N_11873);
or U12336 (N_12336,N_11504,N_11693);
and U12337 (N_12337,N_11981,N_11537);
nand U12338 (N_12338,N_11503,N_11974);
nor U12339 (N_12339,N_11953,N_11472);
and U12340 (N_12340,N_11443,N_11925);
or U12341 (N_12341,N_11984,N_11865);
nand U12342 (N_12342,N_11593,N_11522);
nor U12343 (N_12343,N_11428,N_11566);
nand U12344 (N_12344,N_11728,N_11701);
or U12345 (N_12345,N_11905,N_11700);
nor U12346 (N_12346,N_11440,N_11511);
or U12347 (N_12347,N_11926,N_11694);
nand U12348 (N_12348,N_11623,N_11511);
nor U12349 (N_12349,N_11445,N_11965);
or U12350 (N_12350,N_11960,N_11527);
and U12351 (N_12351,N_11701,N_11403);
and U12352 (N_12352,N_11893,N_11449);
and U12353 (N_12353,N_11616,N_11568);
nand U12354 (N_12354,N_11430,N_11998);
nand U12355 (N_12355,N_11517,N_11996);
nor U12356 (N_12356,N_11552,N_11610);
nor U12357 (N_12357,N_11750,N_11803);
and U12358 (N_12358,N_11473,N_11919);
or U12359 (N_12359,N_11405,N_11811);
and U12360 (N_12360,N_11831,N_11851);
nand U12361 (N_12361,N_11989,N_11922);
or U12362 (N_12362,N_11929,N_11623);
nand U12363 (N_12363,N_11584,N_11760);
and U12364 (N_12364,N_11873,N_11806);
or U12365 (N_12365,N_11869,N_11426);
or U12366 (N_12366,N_11408,N_11637);
nand U12367 (N_12367,N_11985,N_11423);
nor U12368 (N_12368,N_11639,N_11778);
or U12369 (N_12369,N_11656,N_11728);
and U12370 (N_12370,N_11974,N_11474);
nand U12371 (N_12371,N_11805,N_11841);
and U12372 (N_12372,N_11889,N_11408);
nand U12373 (N_12373,N_11592,N_11467);
nor U12374 (N_12374,N_11761,N_11695);
nor U12375 (N_12375,N_11671,N_11453);
xnor U12376 (N_12376,N_11412,N_11413);
nor U12377 (N_12377,N_11643,N_11873);
nor U12378 (N_12378,N_11460,N_11589);
nand U12379 (N_12379,N_11547,N_11745);
xor U12380 (N_12380,N_11751,N_11438);
xnor U12381 (N_12381,N_11429,N_11869);
and U12382 (N_12382,N_11873,N_11810);
or U12383 (N_12383,N_11689,N_11761);
nand U12384 (N_12384,N_11571,N_11812);
or U12385 (N_12385,N_11454,N_11549);
nand U12386 (N_12386,N_11719,N_11488);
xnor U12387 (N_12387,N_11900,N_11669);
and U12388 (N_12388,N_11778,N_11630);
and U12389 (N_12389,N_11905,N_11417);
nor U12390 (N_12390,N_11644,N_11527);
and U12391 (N_12391,N_11822,N_11749);
and U12392 (N_12392,N_11808,N_11971);
and U12393 (N_12393,N_11538,N_11920);
or U12394 (N_12394,N_11562,N_11526);
nor U12395 (N_12395,N_11695,N_11489);
xnor U12396 (N_12396,N_11470,N_11500);
nand U12397 (N_12397,N_11701,N_11707);
or U12398 (N_12398,N_11713,N_11684);
and U12399 (N_12399,N_11896,N_11573);
nand U12400 (N_12400,N_11765,N_11778);
nor U12401 (N_12401,N_11918,N_11448);
or U12402 (N_12402,N_11781,N_11587);
nor U12403 (N_12403,N_11423,N_11899);
and U12404 (N_12404,N_11707,N_11738);
xor U12405 (N_12405,N_11411,N_11829);
nand U12406 (N_12406,N_11796,N_11738);
or U12407 (N_12407,N_11423,N_11721);
xnor U12408 (N_12408,N_11749,N_11949);
or U12409 (N_12409,N_11599,N_11689);
or U12410 (N_12410,N_11448,N_11929);
and U12411 (N_12411,N_11576,N_11936);
or U12412 (N_12412,N_11676,N_11848);
or U12413 (N_12413,N_11732,N_11950);
nand U12414 (N_12414,N_11767,N_11755);
xor U12415 (N_12415,N_11932,N_11914);
nor U12416 (N_12416,N_11489,N_11921);
or U12417 (N_12417,N_11834,N_11950);
nand U12418 (N_12418,N_11822,N_11443);
or U12419 (N_12419,N_11486,N_11650);
nand U12420 (N_12420,N_11791,N_11433);
or U12421 (N_12421,N_11994,N_11414);
nand U12422 (N_12422,N_11826,N_11628);
or U12423 (N_12423,N_11613,N_11727);
xnor U12424 (N_12424,N_11833,N_11506);
nor U12425 (N_12425,N_11749,N_11479);
xnor U12426 (N_12426,N_11510,N_11683);
and U12427 (N_12427,N_11423,N_11412);
nand U12428 (N_12428,N_11489,N_11417);
xor U12429 (N_12429,N_11506,N_11964);
and U12430 (N_12430,N_11682,N_11508);
xnor U12431 (N_12431,N_11706,N_11744);
and U12432 (N_12432,N_11656,N_11480);
nor U12433 (N_12433,N_11632,N_11840);
nand U12434 (N_12434,N_11874,N_11803);
nor U12435 (N_12435,N_11591,N_11787);
xnor U12436 (N_12436,N_11670,N_11409);
nor U12437 (N_12437,N_11767,N_11489);
and U12438 (N_12438,N_11742,N_11757);
and U12439 (N_12439,N_11868,N_11960);
and U12440 (N_12440,N_11974,N_11466);
nor U12441 (N_12441,N_11429,N_11860);
nor U12442 (N_12442,N_11701,N_11438);
nor U12443 (N_12443,N_11736,N_11935);
and U12444 (N_12444,N_11629,N_11428);
nand U12445 (N_12445,N_11720,N_11877);
and U12446 (N_12446,N_11895,N_11652);
and U12447 (N_12447,N_11911,N_11436);
nor U12448 (N_12448,N_11667,N_11540);
or U12449 (N_12449,N_11406,N_11944);
xor U12450 (N_12450,N_11809,N_11502);
nor U12451 (N_12451,N_11911,N_11921);
or U12452 (N_12452,N_11470,N_11614);
or U12453 (N_12453,N_11460,N_11941);
nand U12454 (N_12454,N_11452,N_11955);
nor U12455 (N_12455,N_11772,N_11760);
nand U12456 (N_12456,N_11451,N_11995);
or U12457 (N_12457,N_11455,N_11935);
xor U12458 (N_12458,N_11791,N_11757);
nand U12459 (N_12459,N_11517,N_11639);
nand U12460 (N_12460,N_11440,N_11586);
nand U12461 (N_12461,N_11920,N_11438);
or U12462 (N_12462,N_11809,N_11637);
nor U12463 (N_12463,N_11516,N_11847);
xnor U12464 (N_12464,N_11486,N_11590);
nand U12465 (N_12465,N_11772,N_11931);
nand U12466 (N_12466,N_11578,N_11787);
xor U12467 (N_12467,N_11767,N_11909);
or U12468 (N_12468,N_11930,N_11773);
nand U12469 (N_12469,N_11986,N_11657);
or U12470 (N_12470,N_11730,N_11561);
or U12471 (N_12471,N_11646,N_11859);
xor U12472 (N_12472,N_11757,N_11940);
xor U12473 (N_12473,N_11702,N_11640);
xnor U12474 (N_12474,N_11562,N_11673);
xor U12475 (N_12475,N_11621,N_11958);
and U12476 (N_12476,N_11438,N_11404);
nor U12477 (N_12477,N_11414,N_11539);
nand U12478 (N_12478,N_11578,N_11934);
or U12479 (N_12479,N_11974,N_11978);
nand U12480 (N_12480,N_11716,N_11560);
nand U12481 (N_12481,N_11506,N_11815);
xnor U12482 (N_12482,N_11575,N_11429);
and U12483 (N_12483,N_11906,N_11645);
xnor U12484 (N_12484,N_11838,N_11804);
or U12485 (N_12485,N_11657,N_11753);
nor U12486 (N_12486,N_11707,N_11484);
nor U12487 (N_12487,N_11694,N_11606);
xor U12488 (N_12488,N_11736,N_11817);
or U12489 (N_12489,N_11815,N_11880);
xor U12490 (N_12490,N_11993,N_11752);
xnor U12491 (N_12491,N_11732,N_11737);
and U12492 (N_12492,N_11473,N_11660);
and U12493 (N_12493,N_11673,N_11430);
or U12494 (N_12494,N_11489,N_11667);
and U12495 (N_12495,N_11440,N_11551);
nand U12496 (N_12496,N_11906,N_11659);
and U12497 (N_12497,N_11749,N_11484);
xnor U12498 (N_12498,N_11625,N_11612);
and U12499 (N_12499,N_11534,N_11472);
nor U12500 (N_12500,N_11413,N_11936);
or U12501 (N_12501,N_11809,N_11615);
and U12502 (N_12502,N_11564,N_11515);
and U12503 (N_12503,N_11456,N_11785);
nor U12504 (N_12504,N_11556,N_11413);
nor U12505 (N_12505,N_11920,N_11739);
nand U12506 (N_12506,N_11517,N_11524);
nor U12507 (N_12507,N_11575,N_11519);
xnor U12508 (N_12508,N_11638,N_11601);
nor U12509 (N_12509,N_11410,N_11555);
nand U12510 (N_12510,N_11732,N_11776);
xor U12511 (N_12511,N_11533,N_11559);
nand U12512 (N_12512,N_11456,N_11878);
nand U12513 (N_12513,N_11768,N_11949);
xnor U12514 (N_12514,N_11615,N_11437);
xor U12515 (N_12515,N_11649,N_11458);
nor U12516 (N_12516,N_11536,N_11662);
nor U12517 (N_12517,N_11976,N_11503);
and U12518 (N_12518,N_11864,N_11884);
nor U12519 (N_12519,N_11448,N_11902);
or U12520 (N_12520,N_11495,N_11581);
nor U12521 (N_12521,N_11839,N_11651);
nand U12522 (N_12522,N_11952,N_11890);
or U12523 (N_12523,N_11402,N_11740);
nor U12524 (N_12524,N_11530,N_11551);
or U12525 (N_12525,N_11938,N_11478);
nor U12526 (N_12526,N_11708,N_11949);
nor U12527 (N_12527,N_11910,N_11650);
xor U12528 (N_12528,N_11992,N_11861);
nor U12529 (N_12529,N_11472,N_11979);
nand U12530 (N_12530,N_11643,N_11421);
xnor U12531 (N_12531,N_11650,N_11534);
nor U12532 (N_12532,N_11963,N_11979);
nand U12533 (N_12533,N_11480,N_11603);
xor U12534 (N_12534,N_11996,N_11644);
xnor U12535 (N_12535,N_11526,N_11710);
nand U12536 (N_12536,N_11846,N_11454);
or U12537 (N_12537,N_11642,N_11958);
xnor U12538 (N_12538,N_11766,N_11497);
nand U12539 (N_12539,N_11672,N_11456);
nand U12540 (N_12540,N_11768,N_11529);
or U12541 (N_12541,N_11967,N_11469);
nor U12542 (N_12542,N_11811,N_11583);
nor U12543 (N_12543,N_11761,N_11450);
or U12544 (N_12544,N_11965,N_11876);
and U12545 (N_12545,N_11631,N_11648);
nor U12546 (N_12546,N_11725,N_11556);
and U12547 (N_12547,N_11870,N_11610);
nand U12548 (N_12548,N_11814,N_11925);
and U12549 (N_12549,N_11788,N_11433);
xor U12550 (N_12550,N_11970,N_11416);
and U12551 (N_12551,N_11924,N_11762);
xor U12552 (N_12552,N_11436,N_11494);
or U12553 (N_12553,N_11797,N_11968);
and U12554 (N_12554,N_11939,N_11584);
and U12555 (N_12555,N_11560,N_11401);
nor U12556 (N_12556,N_11642,N_11869);
nor U12557 (N_12557,N_11443,N_11807);
nand U12558 (N_12558,N_11684,N_11894);
nand U12559 (N_12559,N_11718,N_11714);
and U12560 (N_12560,N_11917,N_11878);
xor U12561 (N_12561,N_11999,N_11445);
xnor U12562 (N_12562,N_11614,N_11699);
or U12563 (N_12563,N_11433,N_11560);
nand U12564 (N_12564,N_11704,N_11893);
xor U12565 (N_12565,N_11593,N_11540);
xnor U12566 (N_12566,N_11405,N_11603);
or U12567 (N_12567,N_11757,N_11852);
nand U12568 (N_12568,N_11801,N_11664);
or U12569 (N_12569,N_11847,N_11798);
and U12570 (N_12570,N_11475,N_11824);
or U12571 (N_12571,N_11777,N_11965);
nor U12572 (N_12572,N_11628,N_11430);
nor U12573 (N_12573,N_11626,N_11474);
xnor U12574 (N_12574,N_11975,N_11633);
nand U12575 (N_12575,N_11952,N_11558);
nand U12576 (N_12576,N_11486,N_11642);
or U12577 (N_12577,N_11405,N_11821);
xor U12578 (N_12578,N_11504,N_11819);
xor U12579 (N_12579,N_11476,N_11561);
or U12580 (N_12580,N_11544,N_11506);
and U12581 (N_12581,N_11799,N_11469);
or U12582 (N_12582,N_11908,N_11713);
and U12583 (N_12583,N_11763,N_11956);
xnor U12584 (N_12584,N_11457,N_11721);
and U12585 (N_12585,N_11673,N_11589);
nor U12586 (N_12586,N_11908,N_11823);
xor U12587 (N_12587,N_11559,N_11514);
or U12588 (N_12588,N_11426,N_11976);
and U12589 (N_12589,N_11907,N_11452);
nor U12590 (N_12590,N_11838,N_11900);
xor U12591 (N_12591,N_11640,N_11493);
xor U12592 (N_12592,N_11454,N_11507);
nor U12593 (N_12593,N_11421,N_11524);
or U12594 (N_12594,N_11929,N_11889);
and U12595 (N_12595,N_11718,N_11517);
nor U12596 (N_12596,N_11775,N_11675);
nand U12597 (N_12597,N_11667,N_11722);
xnor U12598 (N_12598,N_11817,N_11940);
or U12599 (N_12599,N_11921,N_11445);
and U12600 (N_12600,N_12448,N_12097);
and U12601 (N_12601,N_12539,N_12236);
or U12602 (N_12602,N_12359,N_12307);
and U12603 (N_12603,N_12257,N_12244);
xnor U12604 (N_12604,N_12194,N_12521);
xor U12605 (N_12605,N_12163,N_12082);
nor U12606 (N_12606,N_12078,N_12021);
or U12607 (N_12607,N_12351,N_12000);
nand U12608 (N_12608,N_12306,N_12496);
xnor U12609 (N_12609,N_12535,N_12027);
and U12610 (N_12610,N_12446,N_12435);
or U12611 (N_12611,N_12129,N_12550);
xnor U12612 (N_12612,N_12003,N_12484);
nand U12613 (N_12613,N_12554,N_12059);
nor U12614 (N_12614,N_12478,N_12256);
and U12615 (N_12615,N_12210,N_12486);
xnor U12616 (N_12616,N_12282,N_12471);
or U12617 (N_12617,N_12443,N_12442);
or U12618 (N_12618,N_12090,N_12036);
and U12619 (N_12619,N_12066,N_12353);
nor U12620 (N_12620,N_12406,N_12531);
xor U12621 (N_12621,N_12118,N_12017);
and U12622 (N_12622,N_12470,N_12575);
xnor U12623 (N_12623,N_12513,N_12170);
nand U12624 (N_12624,N_12056,N_12425);
nand U12625 (N_12625,N_12157,N_12193);
nand U12626 (N_12626,N_12290,N_12124);
and U12627 (N_12627,N_12105,N_12213);
nand U12628 (N_12628,N_12143,N_12196);
and U12629 (N_12629,N_12560,N_12012);
and U12630 (N_12630,N_12107,N_12084);
nor U12631 (N_12631,N_12291,N_12127);
nor U12632 (N_12632,N_12552,N_12054);
nand U12633 (N_12633,N_12596,N_12152);
nor U12634 (N_12634,N_12266,N_12315);
nor U12635 (N_12635,N_12172,N_12134);
or U12636 (N_12636,N_12009,N_12508);
nor U12637 (N_12637,N_12460,N_12312);
xor U12638 (N_12638,N_12038,N_12489);
xnor U12639 (N_12639,N_12275,N_12474);
nand U12640 (N_12640,N_12298,N_12372);
and U12641 (N_12641,N_12179,N_12039);
xnor U12642 (N_12642,N_12265,N_12006);
nor U12643 (N_12643,N_12354,N_12013);
and U12644 (N_12644,N_12375,N_12243);
and U12645 (N_12645,N_12431,N_12562);
or U12646 (N_12646,N_12419,N_12240);
or U12647 (N_12647,N_12360,N_12412);
and U12648 (N_12648,N_12304,N_12438);
or U12649 (N_12649,N_12379,N_12204);
xnor U12650 (N_12650,N_12183,N_12577);
and U12651 (N_12651,N_12102,N_12181);
nand U12652 (N_12652,N_12010,N_12004);
nand U12653 (N_12653,N_12449,N_12592);
nor U12654 (N_12654,N_12215,N_12480);
nor U12655 (N_12655,N_12093,N_12355);
or U12656 (N_12656,N_12258,N_12281);
or U12657 (N_12657,N_12395,N_12219);
xor U12658 (N_12658,N_12116,N_12033);
and U12659 (N_12659,N_12051,N_12020);
nand U12660 (N_12660,N_12579,N_12416);
nand U12661 (N_12661,N_12585,N_12436);
xnor U12662 (N_12662,N_12547,N_12482);
nand U12663 (N_12663,N_12561,N_12593);
nor U12664 (N_12664,N_12061,N_12566);
or U12665 (N_12665,N_12008,N_12404);
nand U12666 (N_12666,N_12524,N_12378);
and U12667 (N_12667,N_12267,N_12289);
nand U12668 (N_12668,N_12103,N_12072);
xnor U12669 (N_12669,N_12148,N_12408);
or U12670 (N_12670,N_12405,N_12316);
nand U12671 (N_12671,N_12221,N_12299);
nor U12672 (N_12672,N_12024,N_12487);
nor U12673 (N_12673,N_12171,N_12195);
xnor U12674 (N_12674,N_12297,N_12330);
nand U12675 (N_12675,N_12300,N_12384);
nand U12676 (N_12676,N_12321,N_12136);
xnor U12677 (N_12677,N_12162,N_12301);
or U12678 (N_12678,N_12277,N_12514);
nand U12679 (N_12679,N_12346,N_12160);
xnor U12680 (N_12680,N_12386,N_12510);
xor U12681 (N_12681,N_12132,N_12542);
xnor U12682 (N_12682,N_12518,N_12590);
and U12683 (N_12683,N_12106,N_12400);
nand U12684 (N_12684,N_12037,N_12279);
xor U12685 (N_12685,N_12546,N_12516);
nand U12686 (N_12686,N_12182,N_12523);
or U12687 (N_12687,N_12490,N_12340);
nor U12688 (N_12688,N_12035,N_12276);
xor U12689 (N_12689,N_12032,N_12366);
nor U12690 (N_12690,N_12526,N_12198);
and U12691 (N_12691,N_12156,N_12085);
or U12692 (N_12692,N_12326,N_12147);
and U12693 (N_12693,N_12248,N_12041);
nor U12694 (N_12694,N_12533,N_12507);
or U12695 (N_12695,N_12166,N_12371);
xor U12696 (N_12696,N_12070,N_12357);
nand U12697 (N_12697,N_12403,N_12580);
nand U12698 (N_12698,N_12511,N_12427);
nand U12699 (N_12699,N_12069,N_12383);
xor U12700 (N_12700,N_12374,N_12123);
nor U12701 (N_12701,N_12466,N_12071);
nand U12702 (N_12702,N_12356,N_12168);
nor U12703 (N_12703,N_12045,N_12463);
or U12704 (N_12704,N_12492,N_12043);
nand U12705 (N_12705,N_12563,N_12441);
or U12706 (N_12706,N_12556,N_12188);
and U12707 (N_12707,N_12016,N_12104);
nand U12708 (N_12708,N_12002,N_12122);
and U12709 (N_12709,N_12216,N_12454);
and U12710 (N_12710,N_12376,N_12241);
and U12711 (N_12711,N_12459,N_12119);
nor U12712 (N_12712,N_12100,N_12462);
nor U12713 (N_12713,N_12421,N_12325);
nand U12714 (N_12714,N_12109,N_12467);
and U12715 (N_12715,N_12394,N_12284);
and U12716 (N_12716,N_12174,N_12440);
or U12717 (N_12717,N_12567,N_12578);
and U12718 (N_12718,N_12083,N_12031);
xor U12719 (N_12719,N_12161,N_12073);
nand U12720 (N_12720,N_12135,N_12381);
or U12721 (N_12721,N_12541,N_12365);
xor U12722 (N_12722,N_12005,N_12225);
and U12723 (N_12723,N_12452,N_12030);
nor U12724 (N_12724,N_12227,N_12551);
xor U12725 (N_12725,N_12397,N_12058);
xnor U12726 (N_12726,N_12238,N_12268);
xor U12727 (N_12727,N_12506,N_12150);
xor U12728 (N_12728,N_12029,N_12544);
nand U12729 (N_12729,N_12559,N_12461);
and U12730 (N_12730,N_12209,N_12251);
and U12731 (N_12731,N_12586,N_12253);
and U12732 (N_12732,N_12450,N_12197);
xor U12733 (N_12733,N_12303,N_12588);
nor U12734 (N_12734,N_12469,N_12223);
xor U12735 (N_12735,N_12271,N_12331);
xnor U12736 (N_12736,N_12433,N_12332);
nor U12737 (N_12737,N_12347,N_12153);
nand U12738 (N_12738,N_12293,N_12324);
xnor U12739 (N_12739,N_12595,N_12140);
xor U12740 (N_12740,N_12473,N_12234);
or U12741 (N_12741,N_12553,N_12120);
nor U12742 (N_12742,N_12110,N_12396);
xor U12743 (N_12743,N_12191,N_12437);
xor U12744 (N_12744,N_12349,N_12529);
and U12745 (N_12745,N_12111,N_12545);
and U12746 (N_12746,N_12011,N_12414);
or U12747 (N_12747,N_12040,N_12398);
xnor U12748 (N_12748,N_12060,N_12399);
or U12749 (N_12749,N_12336,N_12068);
nand U12750 (N_12750,N_12475,N_12247);
or U12751 (N_12751,N_12565,N_12491);
xor U12752 (N_12752,N_12228,N_12587);
nand U12753 (N_12753,N_12505,N_12497);
or U12754 (N_12754,N_12549,N_12048);
nor U12755 (N_12755,N_12570,N_12087);
or U12756 (N_12756,N_12426,N_12101);
and U12757 (N_12757,N_12028,N_12310);
nor U12758 (N_12758,N_12364,N_12014);
xnor U12759 (N_12759,N_12285,N_12173);
nor U12760 (N_12760,N_12576,N_12389);
xnor U12761 (N_12761,N_12065,N_12503);
xor U12762 (N_12762,N_12447,N_12025);
nor U12763 (N_12763,N_12472,N_12226);
and U12764 (N_12764,N_12167,N_12339);
and U12765 (N_12765,N_12259,N_12237);
xor U12766 (N_12766,N_12117,N_12274);
or U12767 (N_12767,N_12249,N_12308);
xor U12768 (N_12768,N_12515,N_12528);
nand U12769 (N_12769,N_12125,N_12320);
xnor U12770 (N_12770,N_12338,N_12242);
xnor U12771 (N_12771,N_12314,N_12094);
nor U12772 (N_12772,N_12569,N_12222);
nor U12773 (N_12773,N_12214,N_12262);
xnor U12774 (N_12774,N_12113,N_12062);
or U12775 (N_12775,N_12430,N_12512);
and U12776 (N_12776,N_12534,N_12597);
nor U12777 (N_12777,N_12458,N_12273);
and U12778 (N_12778,N_12574,N_12538);
or U12779 (N_12779,N_12380,N_12335);
nand U12780 (N_12780,N_12434,N_12067);
xnor U12781 (N_12781,N_12149,N_12283);
nor U12782 (N_12782,N_12589,N_12422);
and U12783 (N_12783,N_12114,N_12131);
and U12784 (N_12784,N_12192,N_12233);
nand U12785 (N_12785,N_12525,N_12250);
and U12786 (N_12786,N_12230,N_12342);
nor U12787 (N_12787,N_12270,N_12571);
xor U12788 (N_12788,N_12115,N_12184);
nor U12789 (N_12789,N_12558,N_12245);
nor U12790 (N_12790,N_12096,N_12327);
and U12791 (N_12791,N_12481,N_12420);
nand U12792 (N_12792,N_12260,N_12564);
or U12793 (N_12793,N_12211,N_12246);
and U12794 (N_12794,N_12158,N_12345);
and U12795 (N_12795,N_12278,N_12089);
nand U12796 (N_12796,N_12137,N_12296);
nor U12797 (N_12797,N_12205,N_12317);
nand U12798 (N_12798,N_12456,N_12146);
nand U12799 (N_12799,N_12599,N_12465);
and U12800 (N_12800,N_12064,N_12333);
or U12801 (N_12801,N_12254,N_12178);
or U12802 (N_12802,N_12477,N_12361);
nor U12803 (N_12803,N_12231,N_12369);
or U12804 (N_12804,N_12502,N_12189);
nand U12805 (N_12805,N_12530,N_12220);
and U12806 (N_12806,N_12392,N_12206);
nand U12807 (N_12807,N_12207,N_12536);
and U12808 (N_12808,N_12583,N_12232);
and U12809 (N_12809,N_12318,N_12522);
xor U12810 (N_12810,N_12328,N_12201);
and U12811 (N_12811,N_12520,N_12057);
or U12812 (N_12812,N_12287,N_12572);
and U12813 (N_12813,N_12130,N_12509);
nor U12814 (N_12814,N_12418,N_12432);
xnor U12815 (N_12815,N_12165,N_12074);
or U12816 (N_12816,N_12428,N_12185);
xor U12817 (N_12817,N_12417,N_12142);
nand U12818 (N_12818,N_12264,N_12363);
nor U12819 (N_12819,N_12092,N_12501);
and U12820 (N_12820,N_12410,N_12540);
xnor U12821 (N_12821,N_12464,N_12527);
nor U12822 (N_12822,N_12164,N_12429);
xor U12823 (N_12823,N_12555,N_12341);
nand U12824 (N_12824,N_12145,N_12483);
or U12825 (N_12825,N_12007,N_12079);
xor U12826 (N_12826,N_12019,N_12292);
and U12827 (N_12827,N_12385,N_12411);
xnor U12828 (N_12828,N_12517,N_12272);
nor U12829 (N_12829,N_12343,N_12500);
or U12830 (N_12830,N_12387,N_12023);
xor U12831 (N_12831,N_12362,N_12370);
nand U12832 (N_12832,N_12413,N_12532);
nor U12833 (N_12833,N_12015,N_12439);
or U12834 (N_12834,N_12295,N_12288);
nor U12835 (N_12835,N_12423,N_12088);
or U12836 (N_12836,N_12075,N_12455);
xnor U12837 (N_12837,N_12108,N_12269);
xor U12838 (N_12838,N_12488,N_12144);
and U12839 (N_12839,N_12373,N_12046);
xor U12840 (N_12840,N_12537,N_12519);
nand U12841 (N_12841,N_12255,N_12190);
and U12842 (N_12842,N_12176,N_12485);
nand U12843 (N_12843,N_12573,N_12445);
nand U12844 (N_12844,N_12239,N_12063);
or U12845 (N_12845,N_12095,N_12294);
xnor U12846 (N_12846,N_12368,N_12080);
nor U12847 (N_12847,N_12493,N_12598);
nand U12848 (N_12848,N_12382,N_12001);
nor U12849 (N_12849,N_12584,N_12350);
xor U12850 (N_12850,N_12098,N_12044);
nand U12851 (N_12851,N_12581,N_12453);
nor U12852 (N_12852,N_12479,N_12263);
or U12853 (N_12853,N_12591,N_12138);
xor U12854 (N_12854,N_12208,N_12077);
nor U12855 (N_12855,N_12022,N_12309);
or U12856 (N_12856,N_12081,N_12543);
and U12857 (N_12857,N_12568,N_12177);
nand U12858 (N_12858,N_12367,N_12034);
nand U12859 (N_12859,N_12159,N_12224);
nor U12860 (N_12860,N_12286,N_12217);
xnor U12861 (N_12861,N_12390,N_12494);
or U12862 (N_12862,N_12169,N_12393);
nand U12863 (N_12863,N_12313,N_12086);
xor U12864 (N_12864,N_12126,N_12557);
nand U12865 (N_12865,N_12305,N_12141);
xor U12866 (N_12866,N_12391,N_12052);
nand U12867 (N_12867,N_12076,N_12235);
nor U12868 (N_12868,N_12334,N_12388);
and U12869 (N_12869,N_12498,N_12329);
and U12870 (N_12870,N_12348,N_12199);
or U12871 (N_12871,N_12409,N_12175);
nor U12872 (N_12872,N_12026,N_12337);
or U12873 (N_12873,N_12154,N_12050);
xnor U12874 (N_12874,N_12047,N_12200);
nor U12875 (N_12875,N_12133,N_12499);
xor U12876 (N_12876,N_12186,N_12457);
and U12877 (N_12877,N_12407,N_12139);
and U12878 (N_12878,N_12468,N_12322);
nand U12879 (N_12879,N_12444,N_12424);
nand U12880 (N_12880,N_12402,N_12495);
nor U12881 (N_12881,N_12202,N_12212);
nand U12882 (N_12882,N_12302,N_12112);
nor U12883 (N_12883,N_12180,N_12252);
nor U12884 (N_12884,N_12053,N_12187);
and U12885 (N_12885,N_12401,N_12261);
nand U12886 (N_12886,N_12229,N_12091);
nand U12887 (N_12887,N_12358,N_12476);
and U12888 (N_12888,N_12504,N_12203);
or U12889 (N_12889,N_12548,N_12018);
xor U12890 (N_12890,N_12594,N_12128);
and U12891 (N_12891,N_12377,N_12121);
xnor U12892 (N_12892,N_12344,N_12049);
nand U12893 (N_12893,N_12451,N_12352);
xnor U12894 (N_12894,N_12055,N_12582);
or U12895 (N_12895,N_12099,N_12415);
xor U12896 (N_12896,N_12042,N_12280);
nand U12897 (N_12897,N_12151,N_12323);
xor U12898 (N_12898,N_12218,N_12319);
and U12899 (N_12899,N_12155,N_12311);
nand U12900 (N_12900,N_12324,N_12116);
or U12901 (N_12901,N_12096,N_12453);
or U12902 (N_12902,N_12029,N_12478);
nor U12903 (N_12903,N_12553,N_12376);
nand U12904 (N_12904,N_12308,N_12013);
or U12905 (N_12905,N_12394,N_12280);
and U12906 (N_12906,N_12450,N_12206);
nand U12907 (N_12907,N_12507,N_12133);
or U12908 (N_12908,N_12189,N_12222);
nand U12909 (N_12909,N_12385,N_12349);
nor U12910 (N_12910,N_12586,N_12577);
nand U12911 (N_12911,N_12565,N_12100);
xnor U12912 (N_12912,N_12517,N_12301);
or U12913 (N_12913,N_12077,N_12470);
nor U12914 (N_12914,N_12078,N_12224);
nand U12915 (N_12915,N_12208,N_12505);
nand U12916 (N_12916,N_12078,N_12449);
nor U12917 (N_12917,N_12184,N_12000);
and U12918 (N_12918,N_12139,N_12598);
xor U12919 (N_12919,N_12307,N_12364);
and U12920 (N_12920,N_12329,N_12344);
or U12921 (N_12921,N_12409,N_12139);
nand U12922 (N_12922,N_12121,N_12576);
nor U12923 (N_12923,N_12577,N_12236);
xor U12924 (N_12924,N_12575,N_12326);
and U12925 (N_12925,N_12503,N_12375);
nor U12926 (N_12926,N_12191,N_12498);
and U12927 (N_12927,N_12080,N_12174);
nor U12928 (N_12928,N_12140,N_12582);
nor U12929 (N_12929,N_12404,N_12437);
or U12930 (N_12930,N_12077,N_12036);
nor U12931 (N_12931,N_12183,N_12036);
xnor U12932 (N_12932,N_12401,N_12277);
and U12933 (N_12933,N_12265,N_12125);
or U12934 (N_12934,N_12589,N_12285);
nand U12935 (N_12935,N_12551,N_12514);
and U12936 (N_12936,N_12212,N_12385);
nor U12937 (N_12937,N_12113,N_12324);
nor U12938 (N_12938,N_12564,N_12295);
nand U12939 (N_12939,N_12547,N_12567);
nand U12940 (N_12940,N_12225,N_12194);
nor U12941 (N_12941,N_12558,N_12130);
or U12942 (N_12942,N_12372,N_12386);
and U12943 (N_12943,N_12232,N_12031);
or U12944 (N_12944,N_12119,N_12283);
xor U12945 (N_12945,N_12382,N_12264);
nor U12946 (N_12946,N_12030,N_12199);
and U12947 (N_12947,N_12573,N_12583);
xnor U12948 (N_12948,N_12407,N_12266);
xor U12949 (N_12949,N_12434,N_12135);
nand U12950 (N_12950,N_12318,N_12043);
xor U12951 (N_12951,N_12364,N_12298);
or U12952 (N_12952,N_12554,N_12065);
and U12953 (N_12953,N_12097,N_12248);
and U12954 (N_12954,N_12436,N_12395);
and U12955 (N_12955,N_12564,N_12381);
nor U12956 (N_12956,N_12500,N_12539);
and U12957 (N_12957,N_12067,N_12415);
xor U12958 (N_12958,N_12344,N_12417);
or U12959 (N_12959,N_12242,N_12268);
nand U12960 (N_12960,N_12250,N_12283);
or U12961 (N_12961,N_12067,N_12551);
xnor U12962 (N_12962,N_12347,N_12279);
nand U12963 (N_12963,N_12396,N_12016);
and U12964 (N_12964,N_12215,N_12416);
or U12965 (N_12965,N_12191,N_12455);
and U12966 (N_12966,N_12419,N_12009);
nor U12967 (N_12967,N_12587,N_12023);
or U12968 (N_12968,N_12297,N_12435);
and U12969 (N_12969,N_12444,N_12479);
xor U12970 (N_12970,N_12208,N_12594);
xnor U12971 (N_12971,N_12395,N_12545);
nor U12972 (N_12972,N_12114,N_12193);
and U12973 (N_12973,N_12080,N_12521);
nor U12974 (N_12974,N_12541,N_12406);
or U12975 (N_12975,N_12341,N_12443);
nor U12976 (N_12976,N_12435,N_12271);
and U12977 (N_12977,N_12073,N_12592);
nor U12978 (N_12978,N_12089,N_12337);
nor U12979 (N_12979,N_12171,N_12289);
and U12980 (N_12980,N_12107,N_12446);
or U12981 (N_12981,N_12033,N_12013);
nor U12982 (N_12982,N_12009,N_12034);
or U12983 (N_12983,N_12499,N_12095);
xor U12984 (N_12984,N_12535,N_12240);
nor U12985 (N_12985,N_12514,N_12079);
or U12986 (N_12986,N_12445,N_12063);
nor U12987 (N_12987,N_12098,N_12450);
and U12988 (N_12988,N_12035,N_12246);
nand U12989 (N_12989,N_12342,N_12484);
or U12990 (N_12990,N_12233,N_12285);
and U12991 (N_12991,N_12057,N_12215);
and U12992 (N_12992,N_12271,N_12584);
and U12993 (N_12993,N_12232,N_12468);
or U12994 (N_12994,N_12536,N_12038);
nand U12995 (N_12995,N_12591,N_12293);
xnor U12996 (N_12996,N_12453,N_12501);
and U12997 (N_12997,N_12202,N_12338);
nand U12998 (N_12998,N_12589,N_12101);
nor U12999 (N_12999,N_12525,N_12404);
nand U13000 (N_13000,N_12573,N_12073);
nand U13001 (N_13001,N_12127,N_12247);
nand U13002 (N_13002,N_12373,N_12087);
xnor U13003 (N_13003,N_12525,N_12209);
nor U13004 (N_13004,N_12227,N_12073);
and U13005 (N_13005,N_12595,N_12347);
or U13006 (N_13006,N_12415,N_12518);
nand U13007 (N_13007,N_12284,N_12195);
and U13008 (N_13008,N_12549,N_12521);
or U13009 (N_13009,N_12556,N_12053);
nor U13010 (N_13010,N_12412,N_12380);
and U13011 (N_13011,N_12059,N_12249);
and U13012 (N_13012,N_12161,N_12278);
nor U13013 (N_13013,N_12351,N_12022);
nand U13014 (N_13014,N_12243,N_12381);
xor U13015 (N_13015,N_12182,N_12136);
xor U13016 (N_13016,N_12424,N_12014);
nand U13017 (N_13017,N_12321,N_12151);
nand U13018 (N_13018,N_12071,N_12238);
xnor U13019 (N_13019,N_12212,N_12419);
xor U13020 (N_13020,N_12288,N_12422);
and U13021 (N_13021,N_12424,N_12199);
or U13022 (N_13022,N_12563,N_12399);
and U13023 (N_13023,N_12178,N_12228);
nand U13024 (N_13024,N_12192,N_12074);
or U13025 (N_13025,N_12449,N_12390);
nor U13026 (N_13026,N_12231,N_12026);
and U13027 (N_13027,N_12488,N_12487);
nor U13028 (N_13028,N_12003,N_12522);
nor U13029 (N_13029,N_12217,N_12456);
or U13030 (N_13030,N_12237,N_12566);
nor U13031 (N_13031,N_12335,N_12122);
xnor U13032 (N_13032,N_12157,N_12150);
and U13033 (N_13033,N_12035,N_12323);
xnor U13034 (N_13034,N_12061,N_12312);
xnor U13035 (N_13035,N_12368,N_12587);
xnor U13036 (N_13036,N_12112,N_12521);
or U13037 (N_13037,N_12582,N_12340);
and U13038 (N_13038,N_12150,N_12026);
xor U13039 (N_13039,N_12496,N_12579);
and U13040 (N_13040,N_12321,N_12111);
and U13041 (N_13041,N_12348,N_12415);
or U13042 (N_13042,N_12206,N_12309);
xnor U13043 (N_13043,N_12099,N_12131);
or U13044 (N_13044,N_12025,N_12220);
nor U13045 (N_13045,N_12588,N_12015);
nor U13046 (N_13046,N_12060,N_12056);
and U13047 (N_13047,N_12000,N_12355);
nor U13048 (N_13048,N_12547,N_12564);
and U13049 (N_13049,N_12580,N_12444);
nand U13050 (N_13050,N_12229,N_12315);
and U13051 (N_13051,N_12430,N_12435);
nor U13052 (N_13052,N_12030,N_12590);
or U13053 (N_13053,N_12237,N_12465);
nand U13054 (N_13054,N_12231,N_12427);
and U13055 (N_13055,N_12472,N_12006);
and U13056 (N_13056,N_12054,N_12046);
or U13057 (N_13057,N_12516,N_12396);
and U13058 (N_13058,N_12274,N_12430);
xnor U13059 (N_13059,N_12224,N_12128);
and U13060 (N_13060,N_12131,N_12280);
nor U13061 (N_13061,N_12276,N_12352);
nand U13062 (N_13062,N_12088,N_12256);
or U13063 (N_13063,N_12223,N_12360);
xor U13064 (N_13064,N_12075,N_12314);
or U13065 (N_13065,N_12560,N_12004);
nor U13066 (N_13066,N_12391,N_12016);
nor U13067 (N_13067,N_12535,N_12356);
or U13068 (N_13068,N_12086,N_12134);
nand U13069 (N_13069,N_12506,N_12227);
nand U13070 (N_13070,N_12258,N_12017);
nor U13071 (N_13071,N_12127,N_12319);
or U13072 (N_13072,N_12393,N_12256);
xnor U13073 (N_13073,N_12003,N_12143);
nand U13074 (N_13074,N_12488,N_12235);
nand U13075 (N_13075,N_12562,N_12201);
xnor U13076 (N_13076,N_12266,N_12511);
xnor U13077 (N_13077,N_12503,N_12447);
nor U13078 (N_13078,N_12564,N_12222);
nor U13079 (N_13079,N_12036,N_12170);
or U13080 (N_13080,N_12059,N_12161);
nor U13081 (N_13081,N_12372,N_12147);
and U13082 (N_13082,N_12325,N_12281);
nor U13083 (N_13083,N_12023,N_12360);
or U13084 (N_13084,N_12108,N_12514);
nor U13085 (N_13085,N_12116,N_12501);
xnor U13086 (N_13086,N_12147,N_12486);
nand U13087 (N_13087,N_12119,N_12528);
nor U13088 (N_13088,N_12157,N_12094);
and U13089 (N_13089,N_12300,N_12254);
nor U13090 (N_13090,N_12361,N_12402);
nand U13091 (N_13091,N_12490,N_12021);
nor U13092 (N_13092,N_12080,N_12028);
or U13093 (N_13093,N_12430,N_12047);
nor U13094 (N_13094,N_12461,N_12575);
nor U13095 (N_13095,N_12096,N_12234);
nand U13096 (N_13096,N_12148,N_12544);
nor U13097 (N_13097,N_12507,N_12344);
and U13098 (N_13098,N_12225,N_12092);
and U13099 (N_13099,N_12417,N_12306);
nor U13100 (N_13100,N_12184,N_12230);
nor U13101 (N_13101,N_12416,N_12143);
or U13102 (N_13102,N_12069,N_12040);
nor U13103 (N_13103,N_12093,N_12402);
nor U13104 (N_13104,N_12036,N_12056);
and U13105 (N_13105,N_12416,N_12432);
or U13106 (N_13106,N_12300,N_12296);
nand U13107 (N_13107,N_12137,N_12431);
or U13108 (N_13108,N_12221,N_12293);
nor U13109 (N_13109,N_12264,N_12288);
xor U13110 (N_13110,N_12175,N_12388);
nor U13111 (N_13111,N_12356,N_12302);
xor U13112 (N_13112,N_12267,N_12398);
nor U13113 (N_13113,N_12551,N_12077);
nor U13114 (N_13114,N_12469,N_12348);
nand U13115 (N_13115,N_12509,N_12275);
nor U13116 (N_13116,N_12248,N_12549);
xnor U13117 (N_13117,N_12134,N_12025);
and U13118 (N_13118,N_12555,N_12502);
and U13119 (N_13119,N_12219,N_12281);
xor U13120 (N_13120,N_12190,N_12128);
or U13121 (N_13121,N_12261,N_12304);
or U13122 (N_13122,N_12313,N_12258);
or U13123 (N_13123,N_12075,N_12055);
nand U13124 (N_13124,N_12469,N_12250);
or U13125 (N_13125,N_12460,N_12097);
xnor U13126 (N_13126,N_12048,N_12360);
and U13127 (N_13127,N_12005,N_12512);
or U13128 (N_13128,N_12359,N_12504);
xnor U13129 (N_13129,N_12145,N_12337);
or U13130 (N_13130,N_12346,N_12110);
and U13131 (N_13131,N_12491,N_12025);
and U13132 (N_13132,N_12260,N_12382);
nor U13133 (N_13133,N_12036,N_12092);
nand U13134 (N_13134,N_12237,N_12005);
xnor U13135 (N_13135,N_12120,N_12109);
xnor U13136 (N_13136,N_12486,N_12511);
and U13137 (N_13137,N_12478,N_12559);
xor U13138 (N_13138,N_12101,N_12058);
nor U13139 (N_13139,N_12119,N_12368);
nand U13140 (N_13140,N_12471,N_12504);
nand U13141 (N_13141,N_12129,N_12538);
or U13142 (N_13142,N_12468,N_12273);
nand U13143 (N_13143,N_12163,N_12275);
nor U13144 (N_13144,N_12256,N_12313);
nor U13145 (N_13145,N_12480,N_12500);
nand U13146 (N_13146,N_12194,N_12141);
and U13147 (N_13147,N_12393,N_12087);
xor U13148 (N_13148,N_12344,N_12597);
nand U13149 (N_13149,N_12412,N_12134);
xnor U13150 (N_13150,N_12475,N_12356);
or U13151 (N_13151,N_12592,N_12426);
nand U13152 (N_13152,N_12312,N_12494);
nor U13153 (N_13153,N_12571,N_12193);
and U13154 (N_13154,N_12022,N_12397);
and U13155 (N_13155,N_12132,N_12410);
nor U13156 (N_13156,N_12192,N_12105);
nor U13157 (N_13157,N_12249,N_12292);
xor U13158 (N_13158,N_12220,N_12356);
xor U13159 (N_13159,N_12229,N_12121);
and U13160 (N_13160,N_12529,N_12376);
xor U13161 (N_13161,N_12266,N_12557);
nor U13162 (N_13162,N_12383,N_12203);
xnor U13163 (N_13163,N_12528,N_12364);
or U13164 (N_13164,N_12097,N_12251);
xnor U13165 (N_13165,N_12116,N_12311);
xor U13166 (N_13166,N_12478,N_12356);
and U13167 (N_13167,N_12539,N_12025);
and U13168 (N_13168,N_12386,N_12598);
or U13169 (N_13169,N_12195,N_12235);
or U13170 (N_13170,N_12549,N_12119);
nor U13171 (N_13171,N_12243,N_12121);
nand U13172 (N_13172,N_12566,N_12249);
and U13173 (N_13173,N_12467,N_12168);
nand U13174 (N_13174,N_12361,N_12024);
or U13175 (N_13175,N_12092,N_12363);
xnor U13176 (N_13176,N_12206,N_12085);
and U13177 (N_13177,N_12062,N_12584);
nand U13178 (N_13178,N_12498,N_12383);
nand U13179 (N_13179,N_12133,N_12417);
xnor U13180 (N_13180,N_12310,N_12034);
and U13181 (N_13181,N_12402,N_12165);
nand U13182 (N_13182,N_12456,N_12228);
nand U13183 (N_13183,N_12058,N_12160);
and U13184 (N_13184,N_12566,N_12295);
or U13185 (N_13185,N_12031,N_12474);
nand U13186 (N_13186,N_12597,N_12280);
or U13187 (N_13187,N_12430,N_12411);
nand U13188 (N_13188,N_12027,N_12461);
and U13189 (N_13189,N_12009,N_12199);
and U13190 (N_13190,N_12330,N_12120);
xnor U13191 (N_13191,N_12348,N_12577);
xor U13192 (N_13192,N_12303,N_12222);
nor U13193 (N_13193,N_12290,N_12335);
xor U13194 (N_13194,N_12140,N_12421);
and U13195 (N_13195,N_12074,N_12484);
xor U13196 (N_13196,N_12137,N_12236);
or U13197 (N_13197,N_12366,N_12523);
xor U13198 (N_13198,N_12366,N_12068);
or U13199 (N_13199,N_12447,N_12406);
and U13200 (N_13200,N_12646,N_12706);
nand U13201 (N_13201,N_12639,N_12687);
and U13202 (N_13202,N_13144,N_13152);
and U13203 (N_13203,N_13067,N_12975);
nand U13204 (N_13204,N_12952,N_12732);
nand U13205 (N_13205,N_13062,N_13155);
xnor U13206 (N_13206,N_12962,N_13079);
nor U13207 (N_13207,N_12722,N_13118);
xor U13208 (N_13208,N_12818,N_12878);
or U13209 (N_13209,N_12977,N_12634);
xnor U13210 (N_13210,N_12872,N_13158);
nor U13211 (N_13211,N_12815,N_12883);
and U13212 (N_13212,N_13128,N_12990);
nand U13213 (N_13213,N_12955,N_12623);
xor U13214 (N_13214,N_12672,N_12868);
nor U13215 (N_13215,N_12823,N_12617);
and U13216 (N_13216,N_13187,N_13153);
or U13217 (N_13217,N_13149,N_12663);
nor U13218 (N_13218,N_12629,N_12921);
nor U13219 (N_13219,N_12717,N_12744);
nor U13220 (N_13220,N_12814,N_13107);
nor U13221 (N_13221,N_13094,N_12835);
nor U13222 (N_13222,N_12601,N_12602);
or U13223 (N_13223,N_12802,N_13073);
and U13224 (N_13224,N_12754,N_12898);
nor U13225 (N_13225,N_12656,N_12607);
nand U13226 (N_13226,N_12766,N_13189);
nand U13227 (N_13227,N_12979,N_12632);
and U13228 (N_13228,N_13151,N_12905);
or U13229 (N_13229,N_13035,N_13085);
nor U13230 (N_13230,N_13096,N_12807);
nor U13231 (N_13231,N_12963,N_12782);
nand U13232 (N_13232,N_13197,N_12831);
or U13233 (N_13233,N_12861,N_13059);
nor U13234 (N_13234,N_12929,N_12606);
or U13235 (N_13235,N_12635,N_12772);
and U13236 (N_13236,N_12638,N_12981);
xnor U13237 (N_13237,N_12703,N_13044);
or U13238 (N_13238,N_12956,N_13184);
xnor U13239 (N_13239,N_12851,N_12763);
or U13240 (N_13240,N_13164,N_12705);
and U13241 (N_13241,N_12696,N_13194);
nor U13242 (N_13242,N_12641,N_12985);
and U13243 (N_13243,N_12912,N_12933);
or U13244 (N_13244,N_12746,N_12695);
xor U13245 (N_13245,N_13100,N_12715);
and U13246 (N_13246,N_12890,N_12885);
or U13247 (N_13247,N_12992,N_12865);
nor U13248 (N_13248,N_12904,N_13078);
xor U13249 (N_13249,N_12832,N_12725);
and U13250 (N_13250,N_12935,N_12896);
xor U13251 (N_13251,N_13072,N_12858);
or U13252 (N_13252,N_12742,N_13193);
and U13253 (N_13253,N_12704,N_12988);
nand U13254 (N_13254,N_12936,N_12828);
nor U13255 (N_13255,N_12893,N_13143);
xnor U13256 (N_13256,N_13023,N_12651);
nor U13257 (N_13257,N_13051,N_13003);
and U13258 (N_13258,N_12825,N_12771);
xor U13259 (N_13259,N_12863,N_12674);
or U13260 (N_13260,N_13137,N_12738);
and U13261 (N_13261,N_12873,N_13070);
and U13262 (N_13262,N_13131,N_12655);
xnor U13263 (N_13263,N_12932,N_12862);
or U13264 (N_13264,N_13002,N_12681);
xnor U13265 (N_13265,N_12650,N_12809);
nor U13266 (N_13266,N_13126,N_12892);
and U13267 (N_13267,N_12743,N_13154);
nand U13268 (N_13268,N_12781,N_12653);
or U13269 (N_13269,N_13016,N_12874);
nand U13270 (N_13270,N_13123,N_13117);
xnor U13271 (N_13271,N_13093,N_12694);
or U13272 (N_13272,N_12751,N_12877);
nor U13273 (N_13273,N_12652,N_13139);
nand U13274 (N_13274,N_12608,N_13156);
nor U13275 (N_13275,N_13007,N_12958);
or U13276 (N_13276,N_12881,N_12942);
xnor U13277 (N_13277,N_12791,N_12849);
nor U13278 (N_13278,N_12884,N_12662);
xnor U13279 (N_13279,N_13160,N_12856);
or U13280 (N_13280,N_12978,N_12908);
nand U13281 (N_13281,N_12848,N_12900);
xor U13282 (N_13282,N_13091,N_12661);
and U13283 (N_13283,N_12622,N_12909);
nor U13284 (N_13284,N_12643,N_12668);
nor U13285 (N_13285,N_12991,N_12768);
nand U13286 (N_13286,N_12691,N_12750);
nand U13287 (N_13287,N_13077,N_12899);
or U13288 (N_13288,N_13081,N_12923);
and U13289 (N_13289,N_13052,N_12930);
or U13290 (N_13290,N_12774,N_13146);
and U13291 (N_13291,N_12779,N_13025);
nand U13292 (N_13292,N_12647,N_13064);
and U13293 (N_13293,N_13112,N_12792);
nand U13294 (N_13294,N_12973,N_12755);
nor U13295 (N_13295,N_12969,N_12723);
nand U13296 (N_13296,N_12800,N_13054);
nor U13297 (N_13297,N_12943,N_13068);
nor U13298 (N_13298,N_12918,N_13020);
or U13299 (N_13299,N_13090,N_13110);
nand U13300 (N_13300,N_12659,N_12735);
nand U13301 (N_13301,N_13017,N_12716);
xor U13302 (N_13302,N_12836,N_13161);
nor U13303 (N_13303,N_13142,N_12951);
and U13304 (N_13304,N_13180,N_13125);
nand U13305 (N_13305,N_12971,N_12619);
or U13306 (N_13306,N_13005,N_13106);
or U13307 (N_13307,N_13089,N_12852);
and U13308 (N_13308,N_12948,N_12631);
nand U13309 (N_13309,N_13047,N_13133);
nor U13310 (N_13310,N_12702,N_12678);
nor U13311 (N_13311,N_13098,N_12924);
nor U13312 (N_13312,N_13022,N_12821);
nand U13313 (N_13313,N_12820,N_12897);
xnor U13314 (N_13314,N_12927,N_13182);
or U13315 (N_13315,N_12701,N_12726);
nor U13316 (N_13316,N_12710,N_12645);
and U13317 (N_13317,N_12871,N_13055);
and U13318 (N_13318,N_12997,N_12867);
or U13319 (N_13319,N_13141,N_12983);
nand U13320 (N_13320,N_12670,N_12829);
or U13321 (N_13321,N_12960,N_12688);
nor U13322 (N_13322,N_12685,N_13175);
nand U13323 (N_13323,N_12959,N_13039);
nand U13324 (N_13324,N_12915,N_12797);
or U13325 (N_13325,N_12759,N_12803);
nor U13326 (N_13326,N_13033,N_13173);
nor U13327 (N_13327,N_12986,N_13115);
xnor U13328 (N_13328,N_12838,N_12667);
or U13329 (N_13329,N_13008,N_13080);
and U13330 (N_13330,N_12998,N_12840);
or U13331 (N_13331,N_12712,N_12677);
or U13332 (N_13332,N_12785,N_12749);
and U13333 (N_13333,N_13119,N_12664);
or U13334 (N_13334,N_12972,N_13046);
or U13335 (N_13335,N_12679,N_12767);
nor U13336 (N_13336,N_13087,N_12680);
nor U13337 (N_13337,N_12798,N_13066);
nand U13338 (N_13338,N_13157,N_12786);
and U13339 (N_13339,N_13147,N_13138);
nand U13340 (N_13340,N_12733,N_12644);
xor U13341 (N_13341,N_12922,N_12628);
nor U13342 (N_13342,N_13043,N_12669);
or U13343 (N_13343,N_12762,N_12709);
or U13344 (N_13344,N_13140,N_13050);
and U13345 (N_13345,N_13006,N_13104);
nand U13346 (N_13346,N_13038,N_13012);
xor U13347 (N_13347,N_12658,N_12843);
nor U13348 (N_13348,N_12813,N_12699);
nand U13349 (N_13349,N_12689,N_13037);
nand U13350 (N_13350,N_12938,N_12752);
or U13351 (N_13351,N_12757,N_12925);
nor U13352 (N_13352,N_12911,N_13063);
nand U13353 (N_13353,N_13060,N_12673);
or U13354 (N_13354,N_12618,N_12614);
and U13355 (N_13355,N_12724,N_12919);
or U13356 (N_13356,N_12736,N_12642);
or U13357 (N_13357,N_12914,N_12693);
nand U13358 (N_13358,N_12708,N_13083);
nor U13359 (N_13359,N_12966,N_13127);
xor U13360 (N_13360,N_13191,N_13045);
or U13361 (N_13361,N_13092,N_12944);
nand U13362 (N_13362,N_12995,N_12799);
nand U13363 (N_13363,N_12875,N_12698);
xor U13364 (N_13364,N_12889,N_13188);
xnor U13365 (N_13365,N_13178,N_13082);
and U13366 (N_13366,N_12739,N_12700);
xor U13367 (N_13367,N_12690,N_13074);
and U13368 (N_13368,N_12682,N_12740);
nand U13369 (N_13369,N_12996,N_13136);
or U13370 (N_13370,N_13053,N_12769);
nor U13371 (N_13371,N_12764,N_12713);
or U13372 (N_13372,N_12753,N_12854);
or U13373 (N_13373,N_12649,N_12824);
nor U13374 (N_13374,N_13027,N_13088);
nand U13375 (N_13375,N_12993,N_13105);
nor U13376 (N_13376,N_12615,N_13185);
or U13377 (N_13377,N_13076,N_12660);
xor U13378 (N_13378,N_12857,N_13192);
nor U13379 (N_13379,N_12654,N_12734);
and U13380 (N_13380,N_12866,N_12964);
or U13381 (N_13381,N_13024,N_12837);
xor U13382 (N_13382,N_13165,N_12826);
nor U13383 (N_13383,N_13010,N_12741);
nor U13384 (N_13384,N_13120,N_12834);
or U13385 (N_13385,N_13186,N_12666);
and U13386 (N_13386,N_13111,N_12603);
or U13387 (N_13387,N_13145,N_12609);
xnor U13388 (N_13388,N_12793,N_12633);
nand U13389 (N_13389,N_12817,N_12737);
nor U13390 (N_13390,N_13198,N_12665);
or U13391 (N_13391,N_13114,N_13122);
xnor U13392 (N_13392,N_13028,N_13166);
xnor U13393 (N_13393,N_12940,N_13172);
and U13394 (N_13394,N_12946,N_13199);
nor U13395 (N_13395,N_13001,N_13162);
and U13396 (N_13396,N_12999,N_12637);
nand U13397 (N_13397,N_12711,N_12675);
xor U13398 (N_13398,N_12928,N_13075);
and U13399 (N_13399,N_12676,N_13169);
or U13400 (N_13400,N_12855,N_12913);
xor U13401 (N_13401,N_13103,N_13109);
nor U13402 (N_13402,N_12920,N_12683);
xnor U13403 (N_13403,N_12901,N_13097);
or U13404 (N_13404,N_12748,N_12967);
and U13405 (N_13405,N_12845,N_12810);
nand U13406 (N_13406,N_12630,N_13168);
nor U13407 (N_13407,N_13084,N_12621);
xor U13408 (N_13408,N_12787,N_13034);
xnor U13409 (N_13409,N_12949,N_12806);
and U13410 (N_13410,N_12613,N_12895);
and U13411 (N_13411,N_12758,N_12954);
xor U13412 (N_13412,N_12729,N_12745);
and U13413 (N_13413,N_12879,N_12945);
nor U13414 (N_13414,N_12794,N_13134);
nand U13415 (N_13415,N_12788,N_12937);
nor U13416 (N_13416,N_13113,N_13021);
and U13417 (N_13417,N_12808,N_13056);
xor U13418 (N_13418,N_12728,N_12853);
xor U13419 (N_13419,N_12605,N_13031);
and U13420 (N_13420,N_13061,N_12869);
or U13421 (N_13421,N_13004,N_12616);
nand U13422 (N_13422,N_12902,N_12620);
or U13423 (N_13423,N_12894,N_13167);
nand U13424 (N_13424,N_12917,N_12839);
and U13425 (N_13425,N_13040,N_13057);
or U13426 (N_13426,N_13171,N_12720);
xnor U13427 (N_13427,N_13015,N_13048);
nor U13428 (N_13428,N_12625,N_12714);
nand U13429 (N_13429,N_13086,N_12859);
xnor U13430 (N_13430,N_12941,N_13019);
nor U13431 (N_13431,N_12789,N_12844);
nand U13432 (N_13432,N_13177,N_12627);
nand U13433 (N_13433,N_12805,N_12657);
nor U13434 (N_13434,N_12790,N_12795);
or U13435 (N_13435,N_13069,N_12776);
nor U13436 (N_13436,N_13042,N_13026);
and U13437 (N_13437,N_13101,N_12721);
and U13438 (N_13438,N_12957,N_12801);
nand U13439 (N_13439,N_12989,N_12718);
and U13440 (N_13440,N_13135,N_12982);
or U13441 (N_13441,N_12600,N_13121);
nand U13442 (N_13442,N_12626,N_13095);
xnor U13443 (N_13443,N_12850,N_13195);
xor U13444 (N_13444,N_12624,N_13009);
or U13445 (N_13445,N_12907,N_13014);
nor U13446 (N_13446,N_12611,N_13032);
nand U13447 (N_13447,N_12640,N_12864);
nor U13448 (N_13448,N_12916,N_12830);
and U13449 (N_13449,N_12761,N_13041);
and U13450 (N_13450,N_12819,N_13183);
nand U13451 (N_13451,N_13148,N_13190);
or U13452 (N_13452,N_12610,N_12968);
nand U13453 (N_13453,N_13196,N_12970);
nor U13454 (N_13454,N_12939,N_12812);
and U13455 (N_13455,N_13116,N_12976);
nor U13456 (N_13456,N_12648,N_13058);
and U13457 (N_13457,N_12934,N_13036);
xnor U13458 (N_13458,N_12947,N_12686);
nand U13459 (N_13459,N_12730,N_13011);
nand U13460 (N_13460,N_13179,N_12980);
and U13461 (N_13461,N_13049,N_13176);
or U13462 (N_13462,N_12775,N_12903);
and U13463 (N_13463,N_12887,N_12876);
or U13464 (N_13464,N_12926,N_13065);
nand U13465 (N_13465,N_12891,N_12780);
xor U13466 (N_13466,N_13150,N_13000);
or U13467 (N_13467,N_13174,N_12684);
nor U13468 (N_13468,N_12671,N_12950);
or U13469 (N_13469,N_12994,N_13102);
nor U13470 (N_13470,N_12965,N_13132);
xor U13471 (N_13471,N_12847,N_12636);
xnor U13472 (N_13472,N_12756,N_12953);
nand U13473 (N_13473,N_12870,N_12784);
xor U13474 (N_13474,N_12961,N_12727);
nand U13475 (N_13475,N_13099,N_12841);
and U13476 (N_13476,N_12846,N_12777);
and U13477 (N_13477,N_13129,N_13071);
or U13478 (N_13478,N_12612,N_12811);
xnor U13479 (N_13479,N_12773,N_13108);
or U13480 (N_13480,N_13029,N_12697);
and U13481 (N_13481,N_12731,N_13159);
and U13482 (N_13482,N_13030,N_12783);
or U13483 (N_13483,N_12747,N_12827);
and U13484 (N_13484,N_12796,N_12974);
and U13485 (N_13485,N_13170,N_12882);
and U13486 (N_13486,N_12833,N_12906);
and U13487 (N_13487,N_12886,N_12842);
and U13488 (N_13488,N_12707,N_12984);
nor U13489 (N_13489,N_12778,N_12910);
and U13490 (N_13490,N_13124,N_12692);
and U13491 (N_13491,N_12931,N_13181);
nand U13492 (N_13492,N_12816,N_12770);
or U13493 (N_13493,N_13018,N_12804);
nand U13494 (N_13494,N_12604,N_12760);
xor U13495 (N_13495,N_12822,N_13163);
or U13496 (N_13496,N_12860,N_13130);
nor U13497 (N_13497,N_12765,N_12987);
nor U13498 (N_13498,N_13013,N_12880);
or U13499 (N_13499,N_12719,N_12888);
and U13500 (N_13500,N_12974,N_12801);
or U13501 (N_13501,N_12722,N_12662);
nand U13502 (N_13502,N_13068,N_13034);
nand U13503 (N_13503,N_12923,N_13090);
nand U13504 (N_13504,N_12721,N_12895);
nand U13505 (N_13505,N_13111,N_13191);
nor U13506 (N_13506,N_12753,N_12714);
nor U13507 (N_13507,N_13071,N_12944);
xnor U13508 (N_13508,N_12838,N_13087);
xor U13509 (N_13509,N_12787,N_13074);
and U13510 (N_13510,N_12907,N_13099);
nor U13511 (N_13511,N_12763,N_12759);
and U13512 (N_13512,N_12668,N_13152);
nand U13513 (N_13513,N_12964,N_13143);
or U13514 (N_13514,N_12754,N_12806);
and U13515 (N_13515,N_12925,N_12950);
nor U13516 (N_13516,N_12798,N_12890);
nand U13517 (N_13517,N_12835,N_13093);
and U13518 (N_13518,N_13009,N_13066);
or U13519 (N_13519,N_12985,N_12768);
nor U13520 (N_13520,N_12684,N_12876);
nor U13521 (N_13521,N_12781,N_13025);
and U13522 (N_13522,N_12978,N_13159);
nor U13523 (N_13523,N_12619,N_12936);
or U13524 (N_13524,N_12975,N_12896);
nand U13525 (N_13525,N_13172,N_13030);
nor U13526 (N_13526,N_12913,N_13155);
xor U13527 (N_13527,N_12938,N_13096);
or U13528 (N_13528,N_12697,N_12907);
and U13529 (N_13529,N_13075,N_12675);
nor U13530 (N_13530,N_12900,N_12873);
and U13531 (N_13531,N_13048,N_12762);
and U13532 (N_13532,N_12923,N_12692);
nor U13533 (N_13533,N_12964,N_13140);
xnor U13534 (N_13534,N_12692,N_12887);
and U13535 (N_13535,N_12887,N_12798);
nand U13536 (N_13536,N_12888,N_13091);
or U13537 (N_13537,N_13018,N_13040);
or U13538 (N_13538,N_13033,N_13089);
nor U13539 (N_13539,N_13141,N_13199);
nand U13540 (N_13540,N_12888,N_12808);
xnor U13541 (N_13541,N_13143,N_12679);
and U13542 (N_13542,N_13053,N_13109);
nand U13543 (N_13543,N_12931,N_13064);
xnor U13544 (N_13544,N_12908,N_13144);
nor U13545 (N_13545,N_12769,N_12662);
nor U13546 (N_13546,N_12879,N_13118);
xor U13547 (N_13547,N_12950,N_13021);
and U13548 (N_13548,N_12893,N_12897);
nand U13549 (N_13549,N_12769,N_13117);
xor U13550 (N_13550,N_12623,N_12851);
or U13551 (N_13551,N_13056,N_12741);
or U13552 (N_13552,N_12927,N_12833);
xnor U13553 (N_13553,N_12651,N_12654);
and U13554 (N_13554,N_12820,N_13039);
nand U13555 (N_13555,N_12640,N_12923);
or U13556 (N_13556,N_12983,N_12764);
xnor U13557 (N_13557,N_12880,N_13046);
xor U13558 (N_13558,N_12802,N_13111);
xor U13559 (N_13559,N_12715,N_12834);
and U13560 (N_13560,N_13182,N_13067);
nand U13561 (N_13561,N_12808,N_12839);
xnor U13562 (N_13562,N_12601,N_13109);
or U13563 (N_13563,N_13016,N_12712);
nor U13564 (N_13564,N_12637,N_12938);
or U13565 (N_13565,N_13114,N_12838);
and U13566 (N_13566,N_12801,N_12642);
xor U13567 (N_13567,N_12706,N_12850);
xor U13568 (N_13568,N_12964,N_13017);
or U13569 (N_13569,N_12772,N_12868);
xnor U13570 (N_13570,N_13157,N_13021);
nor U13571 (N_13571,N_12787,N_13197);
nand U13572 (N_13572,N_12854,N_12781);
or U13573 (N_13573,N_12849,N_12955);
or U13574 (N_13574,N_13108,N_13033);
or U13575 (N_13575,N_13144,N_13194);
nand U13576 (N_13576,N_12819,N_13163);
nand U13577 (N_13577,N_12966,N_12786);
nor U13578 (N_13578,N_12710,N_12855);
nor U13579 (N_13579,N_12697,N_12747);
and U13580 (N_13580,N_12793,N_12982);
nand U13581 (N_13581,N_12638,N_13158);
and U13582 (N_13582,N_12662,N_12898);
and U13583 (N_13583,N_12737,N_12852);
or U13584 (N_13584,N_13143,N_13193);
nand U13585 (N_13585,N_12817,N_12883);
nor U13586 (N_13586,N_13138,N_13000);
nand U13587 (N_13587,N_13130,N_13117);
and U13588 (N_13588,N_12624,N_13042);
nand U13589 (N_13589,N_12960,N_12833);
or U13590 (N_13590,N_12866,N_12854);
or U13591 (N_13591,N_12672,N_12883);
or U13592 (N_13592,N_12806,N_13138);
and U13593 (N_13593,N_12626,N_13098);
and U13594 (N_13594,N_12604,N_12910);
or U13595 (N_13595,N_13001,N_12617);
nor U13596 (N_13596,N_13194,N_12832);
or U13597 (N_13597,N_13162,N_12995);
nor U13598 (N_13598,N_12997,N_12730);
xnor U13599 (N_13599,N_12735,N_13016);
and U13600 (N_13600,N_12870,N_12788);
xnor U13601 (N_13601,N_12691,N_13157);
xor U13602 (N_13602,N_13102,N_12885);
and U13603 (N_13603,N_12945,N_12932);
nor U13604 (N_13604,N_12712,N_12961);
and U13605 (N_13605,N_12873,N_12898);
nand U13606 (N_13606,N_12723,N_13079);
nor U13607 (N_13607,N_12683,N_12628);
or U13608 (N_13608,N_12847,N_12987);
and U13609 (N_13609,N_12646,N_13058);
and U13610 (N_13610,N_12826,N_12642);
xor U13611 (N_13611,N_12850,N_12767);
or U13612 (N_13612,N_12838,N_13079);
nand U13613 (N_13613,N_12791,N_13008);
or U13614 (N_13614,N_13085,N_12742);
nand U13615 (N_13615,N_13198,N_12811);
nand U13616 (N_13616,N_12695,N_12889);
nor U13617 (N_13617,N_12984,N_12628);
nor U13618 (N_13618,N_12713,N_12779);
nor U13619 (N_13619,N_13068,N_12772);
or U13620 (N_13620,N_12614,N_12885);
xnor U13621 (N_13621,N_12666,N_13111);
or U13622 (N_13622,N_12873,N_13143);
nand U13623 (N_13623,N_13159,N_13039);
nor U13624 (N_13624,N_12635,N_12628);
xnor U13625 (N_13625,N_12791,N_13099);
or U13626 (N_13626,N_12812,N_12645);
and U13627 (N_13627,N_12897,N_12927);
nor U13628 (N_13628,N_12754,N_12739);
nand U13629 (N_13629,N_13096,N_12959);
nor U13630 (N_13630,N_12838,N_12660);
and U13631 (N_13631,N_13196,N_12903);
or U13632 (N_13632,N_13033,N_12767);
nand U13633 (N_13633,N_13177,N_13123);
xnor U13634 (N_13634,N_12681,N_12971);
nand U13635 (N_13635,N_12724,N_13017);
xor U13636 (N_13636,N_12898,N_12736);
and U13637 (N_13637,N_13072,N_13197);
and U13638 (N_13638,N_12710,N_13044);
or U13639 (N_13639,N_13028,N_12862);
nand U13640 (N_13640,N_12907,N_12822);
xor U13641 (N_13641,N_12804,N_12644);
xnor U13642 (N_13642,N_12738,N_12882);
xor U13643 (N_13643,N_13131,N_12644);
and U13644 (N_13644,N_12676,N_13082);
or U13645 (N_13645,N_13041,N_12927);
or U13646 (N_13646,N_12860,N_12679);
xnor U13647 (N_13647,N_12834,N_13095);
nor U13648 (N_13648,N_13191,N_12910);
nor U13649 (N_13649,N_13163,N_12707);
nand U13650 (N_13650,N_12947,N_12633);
nand U13651 (N_13651,N_12670,N_12768);
xor U13652 (N_13652,N_13055,N_12757);
or U13653 (N_13653,N_13061,N_12913);
nor U13654 (N_13654,N_12680,N_12991);
xor U13655 (N_13655,N_12901,N_12603);
nor U13656 (N_13656,N_12950,N_12908);
nand U13657 (N_13657,N_13181,N_13024);
or U13658 (N_13658,N_13001,N_12672);
or U13659 (N_13659,N_12901,N_12643);
nand U13660 (N_13660,N_12963,N_12985);
xor U13661 (N_13661,N_12888,N_12885);
xnor U13662 (N_13662,N_12668,N_13097);
and U13663 (N_13663,N_13034,N_13197);
nand U13664 (N_13664,N_12884,N_12907);
xnor U13665 (N_13665,N_12905,N_13086);
xnor U13666 (N_13666,N_12870,N_12996);
and U13667 (N_13667,N_13007,N_12709);
and U13668 (N_13668,N_12816,N_12715);
xnor U13669 (N_13669,N_12962,N_12625);
nand U13670 (N_13670,N_12734,N_12815);
xor U13671 (N_13671,N_12886,N_12721);
xnor U13672 (N_13672,N_12786,N_12722);
and U13673 (N_13673,N_13000,N_13070);
nor U13674 (N_13674,N_12986,N_13156);
or U13675 (N_13675,N_12833,N_12793);
and U13676 (N_13676,N_12705,N_12995);
nor U13677 (N_13677,N_12955,N_12689);
xnor U13678 (N_13678,N_13134,N_13029);
xor U13679 (N_13679,N_12950,N_12975);
nand U13680 (N_13680,N_12727,N_12895);
nor U13681 (N_13681,N_12802,N_12612);
nand U13682 (N_13682,N_12753,N_13183);
nor U13683 (N_13683,N_13085,N_12847);
nand U13684 (N_13684,N_12808,N_12636);
nand U13685 (N_13685,N_12731,N_13119);
nand U13686 (N_13686,N_13192,N_12713);
nand U13687 (N_13687,N_13161,N_12990);
nand U13688 (N_13688,N_13083,N_12731);
xor U13689 (N_13689,N_13003,N_12677);
xnor U13690 (N_13690,N_13077,N_13149);
and U13691 (N_13691,N_12737,N_12611);
xor U13692 (N_13692,N_12945,N_12848);
nor U13693 (N_13693,N_12678,N_12859);
nand U13694 (N_13694,N_12934,N_12618);
and U13695 (N_13695,N_13107,N_12999);
or U13696 (N_13696,N_13089,N_13195);
nor U13697 (N_13697,N_12725,N_12669);
and U13698 (N_13698,N_12929,N_13162);
or U13699 (N_13699,N_13189,N_13168);
xor U13700 (N_13700,N_12958,N_13146);
nand U13701 (N_13701,N_12891,N_12610);
nor U13702 (N_13702,N_12970,N_12683);
and U13703 (N_13703,N_13009,N_12772);
nor U13704 (N_13704,N_12965,N_13069);
xnor U13705 (N_13705,N_12765,N_13001);
xnor U13706 (N_13706,N_12718,N_13117);
or U13707 (N_13707,N_12815,N_12773);
and U13708 (N_13708,N_12629,N_12855);
xor U13709 (N_13709,N_12767,N_12772);
xnor U13710 (N_13710,N_12769,N_12821);
nor U13711 (N_13711,N_12793,N_12937);
and U13712 (N_13712,N_12874,N_12959);
or U13713 (N_13713,N_13108,N_13092);
nor U13714 (N_13714,N_12795,N_12840);
and U13715 (N_13715,N_13188,N_12739);
and U13716 (N_13716,N_12961,N_12988);
xor U13717 (N_13717,N_12608,N_13067);
and U13718 (N_13718,N_12648,N_12890);
xor U13719 (N_13719,N_12888,N_12647);
nand U13720 (N_13720,N_13082,N_12945);
or U13721 (N_13721,N_12991,N_12681);
nor U13722 (N_13722,N_13143,N_12623);
and U13723 (N_13723,N_13084,N_13042);
and U13724 (N_13724,N_13107,N_12926);
nand U13725 (N_13725,N_13043,N_13147);
nand U13726 (N_13726,N_12886,N_13083);
nor U13727 (N_13727,N_13142,N_13066);
or U13728 (N_13728,N_13172,N_13018);
xor U13729 (N_13729,N_12992,N_12820);
xnor U13730 (N_13730,N_12657,N_12633);
and U13731 (N_13731,N_13110,N_13128);
xor U13732 (N_13732,N_12995,N_12732);
and U13733 (N_13733,N_12609,N_12779);
nand U13734 (N_13734,N_12626,N_12937);
nand U13735 (N_13735,N_12739,N_12924);
nand U13736 (N_13736,N_12714,N_13042);
nor U13737 (N_13737,N_13041,N_13061);
nor U13738 (N_13738,N_13141,N_13063);
and U13739 (N_13739,N_12751,N_12872);
nor U13740 (N_13740,N_12839,N_12976);
xor U13741 (N_13741,N_12967,N_13021);
and U13742 (N_13742,N_12665,N_12967);
or U13743 (N_13743,N_12682,N_13126);
and U13744 (N_13744,N_13179,N_12790);
and U13745 (N_13745,N_12660,N_12622);
or U13746 (N_13746,N_12708,N_12929);
or U13747 (N_13747,N_12973,N_12928);
xnor U13748 (N_13748,N_13191,N_12668);
nand U13749 (N_13749,N_12986,N_12794);
or U13750 (N_13750,N_13098,N_13005);
nor U13751 (N_13751,N_13185,N_12773);
and U13752 (N_13752,N_13054,N_12863);
or U13753 (N_13753,N_13060,N_12629);
nor U13754 (N_13754,N_13009,N_12926);
nor U13755 (N_13755,N_12936,N_13037);
or U13756 (N_13756,N_12735,N_12973);
nor U13757 (N_13757,N_13108,N_13172);
nor U13758 (N_13758,N_13081,N_12870);
nand U13759 (N_13759,N_12792,N_13094);
nor U13760 (N_13760,N_12846,N_12767);
or U13761 (N_13761,N_13043,N_12785);
nand U13762 (N_13762,N_13166,N_12780);
or U13763 (N_13763,N_13080,N_13055);
or U13764 (N_13764,N_13182,N_12728);
xor U13765 (N_13765,N_13089,N_13123);
and U13766 (N_13766,N_12913,N_12716);
nand U13767 (N_13767,N_12934,N_13021);
xor U13768 (N_13768,N_12738,N_12745);
and U13769 (N_13769,N_12830,N_13099);
and U13770 (N_13770,N_12754,N_13040);
nand U13771 (N_13771,N_12663,N_13043);
nor U13772 (N_13772,N_12929,N_13110);
or U13773 (N_13773,N_12984,N_13177);
and U13774 (N_13774,N_12873,N_12791);
nor U13775 (N_13775,N_12732,N_13030);
or U13776 (N_13776,N_12670,N_13062);
nand U13777 (N_13777,N_12675,N_12672);
nor U13778 (N_13778,N_12721,N_12711);
or U13779 (N_13779,N_13041,N_12915);
xor U13780 (N_13780,N_13057,N_12965);
nand U13781 (N_13781,N_12755,N_13037);
or U13782 (N_13782,N_12689,N_12940);
xor U13783 (N_13783,N_12888,N_12722);
nor U13784 (N_13784,N_12702,N_12987);
xnor U13785 (N_13785,N_12767,N_12798);
nor U13786 (N_13786,N_12777,N_12613);
and U13787 (N_13787,N_13053,N_12689);
nand U13788 (N_13788,N_12765,N_12841);
and U13789 (N_13789,N_13048,N_12894);
and U13790 (N_13790,N_12854,N_12698);
or U13791 (N_13791,N_12891,N_12719);
or U13792 (N_13792,N_12687,N_12877);
nand U13793 (N_13793,N_12936,N_12919);
and U13794 (N_13794,N_12711,N_12939);
nand U13795 (N_13795,N_12628,N_13143);
and U13796 (N_13796,N_13123,N_12739);
and U13797 (N_13797,N_13115,N_12884);
nand U13798 (N_13798,N_13049,N_12602);
nand U13799 (N_13799,N_12659,N_13013);
and U13800 (N_13800,N_13659,N_13287);
nor U13801 (N_13801,N_13793,N_13467);
or U13802 (N_13802,N_13343,N_13402);
and U13803 (N_13803,N_13585,N_13388);
or U13804 (N_13804,N_13645,N_13376);
nor U13805 (N_13805,N_13705,N_13258);
nand U13806 (N_13806,N_13590,N_13517);
or U13807 (N_13807,N_13259,N_13533);
or U13808 (N_13808,N_13309,N_13480);
nor U13809 (N_13809,N_13752,N_13294);
or U13810 (N_13810,N_13320,N_13534);
or U13811 (N_13811,N_13211,N_13505);
or U13812 (N_13812,N_13262,N_13694);
xnor U13813 (N_13813,N_13638,N_13246);
or U13814 (N_13814,N_13663,N_13269);
xnor U13815 (N_13815,N_13639,N_13564);
and U13816 (N_13816,N_13243,N_13536);
xnor U13817 (N_13817,N_13518,N_13510);
nand U13818 (N_13818,N_13702,N_13687);
and U13819 (N_13819,N_13722,N_13756);
or U13820 (N_13820,N_13568,N_13677);
nand U13821 (N_13821,N_13425,N_13263);
or U13822 (N_13822,N_13511,N_13597);
and U13823 (N_13823,N_13535,N_13474);
nor U13824 (N_13824,N_13653,N_13557);
and U13825 (N_13825,N_13278,N_13339);
xor U13826 (N_13826,N_13734,N_13767);
or U13827 (N_13827,N_13633,N_13202);
nand U13828 (N_13828,N_13247,N_13443);
nand U13829 (N_13829,N_13283,N_13553);
or U13830 (N_13830,N_13319,N_13224);
nand U13831 (N_13831,N_13304,N_13365);
nor U13832 (N_13832,N_13241,N_13556);
and U13833 (N_13833,N_13234,N_13798);
nand U13834 (N_13834,N_13631,N_13759);
nand U13835 (N_13835,N_13378,N_13623);
and U13836 (N_13836,N_13682,N_13476);
or U13837 (N_13837,N_13695,N_13377);
or U13838 (N_13838,N_13448,N_13544);
and U13839 (N_13839,N_13451,N_13383);
nand U13840 (N_13840,N_13504,N_13289);
or U13841 (N_13841,N_13223,N_13417);
or U13842 (N_13842,N_13348,N_13628);
nand U13843 (N_13843,N_13362,N_13358);
and U13844 (N_13844,N_13455,N_13254);
nor U13845 (N_13845,N_13543,N_13416);
and U13846 (N_13846,N_13469,N_13424);
nand U13847 (N_13847,N_13708,N_13747);
or U13848 (N_13848,N_13710,N_13739);
xnor U13849 (N_13849,N_13356,N_13303);
and U13850 (N_13850,N_13444,N_13665);
and U13851 (N_13851,N_13586,N_13554);
nand U13852 (N_13852,N_13714,N_13599);
xnor U13853 (N_13853,N_13494,N_13342);
and U13854 (N_13854,N_13650,N_13324);
xnor U13855 (N_13855,N_13531,N_13546);
or U13856 (N_13856,N_13668,N_13613);
nor U13857 (N_13857,N_13770,N_13693);
and U13858 (N_13858,N_13366,N_13244);
or U13859 (N_13859,N_13379,N_13338);
nand U13860 (N_13860,N_13351,N_13288);
xor U13861 (N_13861,N_13589,N_13565);
or U13862 (N_13862,N_13499,N_13403);
nand U13863 (N_13863,N_13606,N_13225);
nor U13864 (N_13864,N_13352,N_13523);
or U13865 (N_13865,N_13232,N_13251);
or U13866 (N_13866,N_13592,N_13472);
or U13867 (N_13867,N_13354,N_13560);
xnor U13868 (N_13868,N_13215,N_13736);
and U13869 (N_13869,N_13760,N_13295);
nor U13870 (N_13870,N_13249,N_13331);
and U13871 (N_13871,N_13337,N_13373);
and U13872 (N_13872,N_13541,N_13781);
nor U13873 (N_13873,N_13239,N_13521);
nand U13874 (N_13874,N_13399,N_13780);
xor U13875 (N_13875,N_13522,N_13284);
and U13876 (N_13876,N_13790,N_13216);
or U13877 (N_13877,N_13408,N_13484);
or U13878 (N_13878,N_13618,N_13754);
nor U13879 (N_13879,N_13411,N_13669);
xnor U13880 (N_13880,N_13250,N_13570);
nand U13881 (N_13881,N_13741,N_13488);
and U13882 (N_13882,N_13656,N_13430);
nand U13883 (N_13883,N_13374,N_13611);
or U13884 (N_13884,N_13271,N_13502);
nor U13885 (N_13885,N_13773,N_13612);
or U13886 (N_13886,N_13328,N_13290);
nand U13887 (N_13887,N_13367,N_13248);
xnor U13888 (N_13888,N_13532,N_13579);
nand U13889 (N_13889,N_13266,N_13561);
or U13890 (N_13890,N_13470,N_13575);
nor U13891 (N_13891,N_13762,N_13721);
or U13892 (N_13892,N_13349,N_13280);
nand U13893 (N_13893,N_13203,N_13406);
nor U13894 (N_13894,N_13626,N_13418);
or U13895 (N_13895,N_13587,N_13607);
or U13896 (N_13896,N_13456,N_13256);
and U13897 (N_13897,N_13768,N_13396);
nand U13898 (N_13898,N_13621,N_13363);
nand U13899 (N_13899,N_13226,N_13577);
and U13900 (N_13900,N_13359,N_13686);
xnor U13901 (N_13901,N_13765,N_13222);
nand U13902 (N_13902,N_13753,N_13576);
xnor U13903 (N_13903,N_13322,N_13779);
nand U13904 (N_13904,N_13397,N_13784);
and U13905 (N_13905,N_13206,N_13654);
or U13906 (N_13906,N_13620,N_13441);
xor U13907 (N_13907,N_13421,N_13335);
or U13908 (N_13908,N_13699,N_13412);
nor U13909 (N_13909,N_13582,N_13387);
xor U13910 (N_13910,N_13624,N_13240);
or U13911 (N_13911,N_13644,N_13748);
xor U13912 (N_13912,N_13371,N_13700);
xnor U13913 (N_13913,N_13300,N_13242);
nor U13914 (N_13914,N_13219,N_13709);
nand U13915 (N_13915,N_13208,N_13477);
and U13916 (N_13916,N_13459,N_13527);
xnor U13917 (N_13917,N_13483,N_13272);
or U13918 (N_13918,N_13245,N_13666);
or U13919 (N_13919,N_13433,N_13528);
and U13920 (N_13920,N_13725,N_13398);
xor U13921 (N_13921,N_13370,N_13487);
xor U13922 (N_13922,N_13720,N_13310);
or U13923 (N_13923,N_13588,N_13641);
nand U13924 (N_13924,N_13566,N_13675);
nand U13925 (N_13925,N_13299,N_13479);
xnor U13926 (N_13926,N_13347,N_13436);
nand U13927 (N_13927,N_13706,N_13719);
nor U13928 (N_13928,N_13391,N_13593);
xor U13929 (N_13929,N_13419,N_13563);
xor U13930 (N_13930,N_13672,N_13345);
nor U13931 (N_13931,N_13540,N_13750);
xnor U13932 (N_13932,N_13594,N_13707);
or U13933 (N_13933,N_13423,N_13799);
nand U13934 (N_13934,N_13210,N_13268);
and U13935 (N_13935,N_13415,N_13450);
nor U13936 (N_13936,N_13745,N_13385);
xor U13937 (N_13937,N_13260,N_13610);
nand U13938 (N_13938,N_13233,N_13746);
and U13939 (N_13939,N_13698,N_13490);
nor U13940 (N_13940,N_13662,N_13434);
nor U13941 (N_13941,N_13212,N_13787);
xor U13942 (N_13942,N_13596,N_13237);
nand U13943 (N_13943,N_13583,N_13395);
nor U13944 (N_13944,N_13697,N_13350);
nor U13945 (N_13945,N_13205,N_13273);
xnor U13946 (N_13946,N_13530,N_13652);
nand U13947 (N_13947,N_13489,N_13440);
xnor U13948 (N_13948,N_13696,N_13730);
nor U13949 (N_13949,N_13547,N_13794);
xor U13950 (N_13950,N_13325,N_13316);
nand U13951 (N_13951,N_13600,N_13390);
nor U13952 (N_13952,N_13204,N_13384);
and U13953 (N_13953,N_13313,N_13427);
nand U13954 (N_13954,N_13758,N_13726);
xnor U13955 (N_13955,N_13314,N_13495);
nor U13956 (N_13956,N_13293,N_13252);
nor U13957 (N_13957,N_13270,N_13603);
xor U13958 (N_13958,N_13764,N_13584);
nand U13959 (N_13959,N_13545,N_13506);
nand U13960 (N_13960,N_13711,N_13619);
xnor U13961 (N_13961,N_13305,N_13307);
nand U13962 (N_13962,N_13292,N_13636);
and U13963 (N_13963,N_13218,N_13353);
xor U13964 (N_13964,N_13743,N_13513);
nor U13965 (N_13965,N_13389,N_13524);
nor U13966 (N_13966,N_13716,N_13286);
or U13967 (N_13967,N_13516,N_13712);
xor U13968 (N_13968,N_13414,N_13431);
or U13969 (N_13969,N_13704,N_13267);
xor U13970 (N_13970,N_13327,N_13605);
nand U13971 (N_13971,N_13311,N_13783);
nor U13972 (N_13972,N_13786,N_13723);
xor U13973 (N_13973,N_13209,N_13382);
or U13974 (N_13974,N_13360,N_13514);
nand U13975 (N_13975,N_13742,N_13775);
and U13976 (N_13976,N_13785,N_13789);
nor U13977 (N_13977,N_13567,N_13318);
nand U13978 (N_13978,N_13729,N_13296);
and U13979 (N_13979,N_13630,N_13410);
and U13980 (N_13980,N_13622,N_13392);
or U13981 (N_13981,N_13475,N_13372);
nor U13982 (N_13982,N_13769,N_13717);
or U13983 (N_13983,N_13330,N_13409);
nand U13984 (N_13984,N_13369,N_13478);
nor U13985 (N_13985,N_13637,N_13526);
nand U13986 (N_13986,N_13649,N_13558);
or U13987 (N_13987,N_13674,N_13458);
nand U13988 (N_13988,N_13615,N_13333);
or U13989 (N_13989,N_13598,N_13386);
nor U13990 (N_13990,N_13548,N_13580);
xnor U13991 (N_13991,N_13275,N_13673);
nor U13992 (N_13992,N_13461,N_13407);
nor U13993 (N_13993,N_13255,N_13380);
nand U13994 (N_13994,N_13643,N_13713);
nand U13995 (N_13995,N_13670,N_13449);
or U13996 (N_13996,N_13221,N_13685);
or U13997 (N_13997,N_13617,N_13651);
or U13998 (N_13998,N_13572,N_13749);
xnor U13999 (N_13999,N_13400,N_13733);
nor U14000 (N_14000,N_13782,N_13657);
xnor U14001 (N_14001,N_13508,N_13446);
and U14002 (N_14002,N_13276,N_13432);
nor U14003 (N_14003,N_13229,N_13261);
and U14004 (N_14004,N_13774,N_13393);
xnor U14005 (N_14005,N_13236,N_13394);
and U14006 (N_14006,N_13520,N_13253);
nand U14007 (N_14007,N_13442,N_13660);
and U14008 (N_14008,N_13689,N_13552);
nor U14009 (N_14009,N_13681,N_13285);
or U14010 (N_14010,N_13452,N_13306);
or U14011 (N_14011,N_13381,N_13559);
nor U14012 (N_14012,N_13691,N_13315);
nor U14013 (N_14013,N_13632,N_13515);
or U14014 (N_14014,N_13496,N_13491);
nor U14015 (N_14015,N_13703,N_13627);
xor U14016 (N_14016,N_13493,N_13321);
nor U14017 (N_14017,N_13336,N_13757);
xor U14018 (N_14018,N_13683,N_13634);
or U14019 (N_14019,N_13667,N_13602);
or U14020 (N_14020,N_13507,N_13792);
or U14021 (N_14021,N_13437,N_13529);
nand U14022 (N_14022,N_13364,N_13308);
or U14023 (N_14023,N_13238,N_13728);
or U14024 (N_14024,N_13265,N_13701);
or U14025 (N_14025,N_13550,N_13738);
xor U14026 (N_14026,N_13569,N_13578);
nand U14027 (N_14027,N_13684,N_13473);
nor U14028 (N_14028,N_13281,N_13227);
nor U14029 (N_14029,N_13763,N_13573);
xnor U14030 (N_14030,N_13332,N_13646);
nor U14031 (N_14031,N_13466,N_13405);
or U14032 (N_14032,N_13201,N_13549);
or U14033 (N_14033,N_13778,N_13420);
nand U14034 (N_14034,N_13482,N_13772);
and U14035 (N_14035,N_13542,N_13581);
and U14036 (N_14036,N_13788,N_13795);
nand U14037 (N_14037,N_13676,N_13655);
or U14038 (N_14038,N_13539,N_13481);
nand U14039 (N_14039,N_13642,N_13571);
nand U14040 (N_14040,N_13608,N_13731);
or U14041 (N_14041,N_13498,N_13766);
and U14042 (N_14042,N_13401,N_13447);
nor U14043 (N_14043,N_13438,N_13344);
or U14044 (N_14044,N_13301,N_13797);
nand U14045 (N_14045,N_13346,N_13274);
nand U14046 (N_14046,N_13404,N_13796);
nor U14047 (N_14047,N_13340,N_13361);
nor U14048 (N_14048,N_13228,N_13616);
and U14049 (N_14049,N_13740,N_13312);
xnor U14050 (N_14050,N_13323,N_13678);
and U14051 (N_14051,N_13429,N_13688);
and U14052 (N_14052,N_13718,N_13679);
or U14053 (N_14053,N_13551,N_13230);
or U14054 (N_14054,N_13355,N_13485);
xor U14055 (N_14055,N_13454,N_13279);
xnor U14056 (N_14056,N_13680,N_13329);
xnor U14057 (N_14057,N_13214,N_13690);
and U14058 (N_14058,N_13519,N_13334);
nor U14059 (N_14059,N_13213,N_13375);
or U14060 (N_14060,N_13435,N_13422);
nand U14061 (N_14061,N_13471,N_13724);
nand U14062 (N_14062,N_13291,N_13595);
nand U14063 (N_14063,N_13648,N_13509);
or U14064 (N_14064,N_13257,N_13264);
nand U14065 (N_14065,N_13357,N_13562);
nand U14066 (N_14066,N_13755,N_13468);
or U14067 (N_14067,N_13326,N_13200);
and U14068 (N_14068,N_13302,N_13625);
and U14069 (N_14069,N_13462,N_13537);
and U14070 (N_14070,N_13465,N_13777);
or U14071 (N_14071,N_13715,N_13604);
or U14072 (N_14072,N_13503,N_13463);
xnor U14073 (N_14073,N_13614,N_13658);
xnor U14074 (N_14074,N_13671,N_13235);
nor U14075 (N_14075,N_13207,N_13497);
nand U14076 (N_14076,N_13692,N_13297);
or U14077 (N_14077,N_13661,N_13220);
xor U14078 (N_14078,N_13555,N_13282);
nand U14079 (N_14079,N_13727,N_13601);
nand U14080 (N_14080,N_13486,N_13635);
xnor U14081 (N_14081,N_13776,N_13737);
and U14082 (N_14082,N_13457,N_13492);
nand U14083 (N_14083,N_13647,N_13368);
or U14084 (N_14084,N_13426,N_13445);
and U14085 (N_14085,N_13439,N_13500);
xnor U14086 (N_14086,N_13525,N_13501);
nand U14087 (N_14087,N_13277,N_13341);
and U14088 (N_14088,N_13664,N_13629);
nor U14089 (N_14089,N_13761,N_13732);
and U14090 (N_14090,N_13217,N_13298);
or U14091 (N_14091,N_13771,N_13751);
nor U14092 (N_14092,N_13428,N_13453);
or U14093 (N_14093,N_13744,N_13735);
nor U14094 (N_14094,N_13231,N_13317);
nand U14095 (N_14095,N_13464,N_13591);
and U14096 (N_14096,N_13574,N_13538);
or U14097 (N_14097,N_13791,N_13460);
xor U14098 (N_14098,N_13640,N_13413);
nand U14099 (N_14099,N_13512,N_13609);
and U14100 (N_14100,N_13400,N_13353);
and U14101 (N_14101,N_13621,N_13642);
and U14102 (N_14102,N_13694,N_13494);
and U14103 (N_14103,N_13760,N_13700);
nor U14104 (N_14104,N_13223,N_13460);
or U14105 (N_14105,N_13535,N_13530);
and U14106 (N_14106,N_13719,N_13303);
nor U14107 (N_14107,N_13280,N_13338);
nand U14108 (N_14108,N_13449,N_13361);
nor U14109 (N_14109,N_13391,N_13600);
nor U14110 (N_14110,N_13742,N_13688);
xor U14111 (N_14111,N_13705,N_13285);
or U14112 (N_14112,N_13481,N_13548);
nand U14113 (N_14113,N_13536,N_13443);
xor U14114 (N_14114,N_13261,N_13634);
and U14115 (N_14115,N_13408,N_13593);
nand U14116 (N_14116,N_13233,N_13451);
or U14117 (N_14117,N_13509,N_13405);
or U14118 (N_14118,N_13377,N_13473);
nor U14119 (N_14119,N_13765,N_13240);
or U14120 (N_14120,N_13541,N_13737);
xor U14121 (N_14121,N_13394,N_13588);
and U14122 (N_14122,N_13784,N_13584);
nor U14123 (N_14123,N_13314,N_13661);
xnor U14124 (N_14124,N_13528,N_13651);
and U14125 (N_14125,N_13636,N_13512);
and U14126 (N_14126,N_13699,N_13314);
nor U14127 (N_14127,N_13681,N_13486);
and U14128 (N_14128,N_13337,N_13581);
nand U14129 (N_14129,N_13686,N_13362);
nor U14130 (N_14130,N_13569,N_13761);
or U14131 (N_14131,N_13437,N_13626);
and U14132 (N_14132,N_13344,N_13284);
and U14133 (N_14133,N_13712,N_13438);
nor U14134 (N_14134,N_13254,N_13788);
xor U14135 (N_14135,N_13452,N_13747);
nor U14136 (N_14136,N_13499,N_13703);
xor U14137 (N_14137,N_13620,N_13332);
and U14138 (N_14138,N_13575,N_13351);
and U14139 (N_14139,N_13341,N_13446);
nor U14140 (N_14140,N_13620,N_13785);
xor U14141 (N_14141,N_13541,N_13744);
xor U14142 (N_14142,N_13662,N_13592);
or U14143 (N_14143,N_13582,N_13618);
xor U14144 (N_14144,N_13311,N_13378);
nand U14145 (N_14145,N_13398,N_13324);
nand U14146 (N_14146,N_13701,N_13385);
nor U14147 (N_14147,N_13249,N_13318);
and U14148 (N_14148,N_13513,N_13488);
xor U14149 (N_14149,N_13496,N_13224);
xor U14150 (N_14150,N_13283,N_13528);
nor U14151 (N_14151,N_13326,N_13554);
xnor U14152 (N_14152,N_13202,N_13730);
nor U14153 (N_14153,N_13289,N_13284);
nand U14154 (N_14154,N_13430,N_13621);
xor U14155 (N_14155,N_13748,N_13583);
and U14156 (N_14156,N_13356,N_13468);
xnor U14157 (N_14157,N_13658,N_13683);
nand U14158 (N_14158,N_13552,N_13720);
and U14159 (N_14159,N_13686,N_13681);
nand U14160 (N_14160,N_13661,N_13436);
nor U14161 (N_14161,N_13370,N_13649);
and U14162 (N_14162,N_13413,N_13333);
nand U14163 (N_14163,N_13600,N_13254);
xor U14164 (N_14164,N_13557,N_13467);
nand U14165 (N_14165,N_13230,N_13426);
xor U14166 (N_14166,N_13355,N_13525);
and U14167 (N_14167,N_13791,N_13228);
and U14168 (N_14168,N_13525,N_13634);
nor U14169 (N_14169,N_13212,N_13245);
nor U14170 (N_14170,N_13614,N_13420);
nor U14171 (N_14171,N_13694,N_13317);
nor U14172 (N_14172,N_13456,N_13372);
nor U14173 (N_14173,N_13328,N_13404);
and U14174 (N_14174,N_13524,N_13253);
and U14175 (N_14175,N_13233,N_13436);
xor U14176 (N_14176,N_13467,N_13283);
or U14177 (N_14177,N_13538,N_13685);
nor U14178 (N_14178,N_13654,N_13791);
and U14179 (N_14179,N_13758,N_13662);
xnor U14180 (N_14180,N_13665,N_13262);
or U14181 (N_14181,N_13346,N_13241);
nor U14182 (N_14182,N_13743,N_13216);
xnor U14183 (N_14183,N_13763,N_13307);
nor U14184 (N_14184,N_13389,N_13605);
and U14185 (N_14185,N_13208,N_13469);
and U14186 (N_14186,N_13537,N_13745);
nand U14187 (N_14187,N_13542,N_13294);
xnor U14188 (N_14188,N_13644,N_13569);
xnor U14189 (N_14189,N_13499,N_13700);
or U14190 (N_14190,N_13637,N_13261);
xnor U14191 (N_14191,N_13646,N_13530);
nand U14192 (N_14192,N_13478,N_13567);
and U14193 (N_14193,N_13454,N_13304);
xor U14194 (N_14194,N_13206,N_13317);
nor U14195 (N_14195,N_13453,N_13267);
xor U14196 (N_14196,N_13532,N_13584);
or U14197 (N_14197,N_13376,N_13426);
nand U14198 (N_14198,N_13384,N_13674);
nor U14199 (N_14199,N_13318,N_13278);
nand U14200 (N_14200,N_13701,N_13560);
nor U14201 (N_14201,N_13444,N_13246);
nand U14202 (N_14202,N_13739,N_13260);
and U14203 (N_14203,N_13608,N_13432);
nand U14204 (N_14204,N_13599,N_13372);
and U14205 (N_14205,N_13255,N_13427);
nor U14206 (N_14206,N_13782,N_13756);
nor U14207 (N_14207,N_13528,N_13449);
nand U14208 (N_14208,N_13201,N_13511);
or U14209 (N_14209,N_13234,N_13520);
nand U14210 (N_14210,N_13228,N_13756);
xnor U14211 (N_14211,N_13321,N_13713);
nand U14212 (N_14212,N_13781,N_13585);
nand U14213 (N_14213,N_13380,N_13335);
or U14214 (N_14214,N_13373,N_13456);
or U14215 (N_14215,N_13595,N_13642);
nor U14216 (N_14216,N_13329,N_13728);
xor U14217 (N_14217,N_13541,N_13724);
or U14218 (N_14218,N_13555,N_13733);
and U14219 (N_14219,N_13308,N_13530);
xor U14220 (N_14220,N_13311,N_13712);
xnor U14221 (N_14221,N_13211,N_13257);
xnor U14222 (N_14222,N_13592,N_13733);
nand U14223 (N_14223,N_13728,N_13316);
nand U14224 (N_14224,N_13776,N_13576);
xnor U14225 (N_14225,N_13410,N_13346);
or U14226 (N_14226,N_13232,N_13718);
and U14227 (N_14227,N_13649,N_13482);
or U14228 (N_14228,N_13489,N_13607);
nand U14229 (N_14229,N_13793,N_13322);
or U14230 (N_14230,N_13282,N_13220);
nand U14231 (N_14231,N_13774,N_13305);
nand U14232 (N_14232,N_13536,N_13460);
xor U14233 (N_14233,N_13303,N_13471);
or U14234 (N_14234,N_13531,N_13205);
nand U14235 (N_14235,N_13448,N_13462);
or U14236 (N_14236,N_13505,N_13301);
xor U14237 (N_14237,N_13451,N_13509);
nand U14238 (N_14238,N_13787,N_13369);
and U14239 (N_14239,N_13264,N_13610);
or U14240 (N_14240,N_13602,N_13786);
xor U14241 (N_14241,N_13566,N_13533);
or U14242 (N_14242,N_13536,N_13295);
nand U14243 (N_14243,N_13363,N_13676);
or U14244 (N_14244,N_13204,N_13205);
nand U14245 (N_14245,N_13520,N_13547);
and U14246 (N_14246,N_13455,N_13573);
xnor U14247 (N_14247,N_13402,N_13653);
xor U14248 (N_14248,N_13660,N_13303);
nor U14249 (N_14249,N_13470,N_13403);
and U14250 (N_14250,N_13654,N_13498);
nand U14251 (N_14251,N_13483,N_13405);
nand U14252 (N_14252,N_13421,N_13672);
nor U14253 (N_14253,N_13621,N_13442);
nor U14254 (N_14254,N_13500,N_13299);
and U14255 (N_14255,N_13603,N_13589);
or U14256 (N_14256,N_13209,N_13275);
and U14257 (N_14257,N_13694,N_13764);
xnor U14258 (N_14258,N_13233,N_13356);
or U14259 (N_14259,N_13586,N_13346);
nor U14260 (N_14260,N_13453,N_13559);
xnor U14261 (N_14261,N_13705,N_13461);
xnor U14262 (N_14262,N_13339,N_13675);
xnor U14263 (N_14263,N_13205,N_13450);
xor U14264 (N_14264,N_13356,N_13261);
nor U14265 (N_14265,N_13411,N_13712);
nand U14266 (N_14266,N_13604,N_13514);
nor U14267 (N_14267,N_13362,N_13717);
nand U14268 (N_14268,N_13634,N_13451);
and U14269 (N_14269,N_13349,N_13311);
or U14270 (N_14270,N_13759,N_13440);
nand U14271 (N_14271,N_13782,N_13404);
or U14272 (N_14272,N_13230,N_13780);
xnor U14273 (N_14273,N_13757,N_13466);
xnor U14274 (N_14274,N_13414,N_13701);
xnor U14275 (N_14275,N_13437,N_13658);
xor U14276 (N_14276,N_13732,N_13567);
nand U14277 (N_14277,N_13376,N_13307);
nor U14278 (N_14278,N_13546,N_13408);
or U14279 (N_14279,N_13452,N_13587);
or U14280 (N_14280,N_13643,N_13790);
nor U14281 (N_14281,N_13522,N_13245);
nor U14282 (N_14282,N_13657,N_13222);
and U14283 (N_14283,N_13729,N_13607);
nor U14284 (N_14284,N_13313,N_13473);
nor U14285 (N_14285,N_13757,N_13714);
xor U14286 (N_14286,N_13436,N_13497);
or U14287 (N_14287,N_13457,N_13795);
xnor U14288 (N_14288,N_13313,N_13297);
xor U14289 (N_14289,N_13792,N_13528);
xor U14290 (N_14290,N_13641,N_13435);
or U14291 (N_14291,N_13298,N_13206);
and U14292 (N_14292,N_13673,N_13697);
and U14293 (N_14293,N_13209,N_13676);
and U14294 (N_14294,N_13266,N_13443);
nand U14295 (N_14295,N_13647,N_13227);
and U14296 (N_14296,N_13504,N_13256);
xnor U14297 (N_14297,N_13299,N_13510);
nor U14298 (N_14298,N_13744,N_13222);
nor U14299 (N_14299,N_13589,N_13261);
nor U14300 (N_14300,N_13752,N_13585);
or U14301 (N_14301,N_13303,N_13663);
xnor U14302 (N_14302,N_13443,N_13497);
nor U14303 (N_14303,N_13694,N_13427);
nand U14304 (N_14304,N_13493,N_13613);
nand U14305 (N_14305,N_13555,N_13642);
or U14306 (N_14306,N_13574,N_13495);
and U14307 (N_14307,N_13662,N_13485);
and U14308 (N_14308,N_13386,N_13762);
nor U14309 (N_14309,N_13630,N_13368);
xnor U14310 (N_14310,N_13545,N_13535);
or U14311 (N_14311,N_13401,N_13265);
or U14312 (N_14312,N_13290,N_13734);
nor U14313 (N_14313,N_13371,N_13521);
xor U14314 (N_14314,N_13547,N_13643);
and U14315 (N_14315,N_13266,N_13355);
and U14316 (N_14316,N_13229,N_13776);
nand U14317 (N_14317,N_13700,N_13609);
nand U14318 (N_14318,N_13505,N_13280);
nor U14319 (N_14319,N_13513,N_13716);
and U14320 (N_14320,N_13795,N_13760);
nand U14321 (N_14321,N_13309,N_13243);
nand U14322 (N_14322,N_13600,N_13436);
nor U14323 (N_14323,N_13711,N_13273);
xor U14324 (N_14324,N_13227,N_13285);
xnor U14325 (N_14325,N_13562,N_13288);
xor U14326 (N_14326,N_13675,N_13669);
and U14327 (N_14327,N_13309,N_13717);
and U14328 (N_14328,N_13549,N_13772);
and U14329 (N_14329,N_13528,N_13262);
nand U14330 (N_14330,N_13375,N_13771);
nand U14331 (N_14331,N_13714,N_13467);
or U14332 (N_14332,N_13512,N_13211);
xnor U14333 (N_14333,N_13487,N_13355);
nand U14334 (N_14334,N_13338,N_13240);
and U14335 (N_14335,N_13760,N_13329);
nand U14336 (N_14336,N_13406,N_13555);
or U14337 (N_14337,N_13748,N_13431);
or U14338 (N_14338,N_13563,N_13604);
nand U14339 (N_14339,N_13714,N_13742);
nor U14340 (N_14340,N_13761,N_13519);
or U14341 (N_14341,N_13728,N_13287);
nand U14342 (N_14342,N_13604,N_13208);
and U14343 (N_14343,N_13748,N_13312);
nor U14344 (N_14344,N_13697,N_13451);
xor U14345 (N_14345,N_13694,N_13337);
xor U14346 (N_14346,N_13368,N_13269);
nor U14347 (N_14347,N_13461,N_13515);
and U14348 (N_14348,N_13735,N_13248);
xor U14349 (N_14349,N_13724,N_13514);
nor U14350 (N_14350,N_13249,N_13596);
xor U14351 (N_14351,N_13726,N_13461);
xor U14352 (N_14352,N_13221,N_13520);
and U14353 (N_14353,N_13461,N_13660);
nand U14354 (N_14354,N_13657,N_13757);
nand U14355 (N_14355,N_13765,N_13583);
and U14356 (N_14356,N_13741,N_13491);
nor U14357 (N_14357,N_13613,N_13702);
and U14358 (N_14358,N_13503,N_13575);
and U14359 (N_14359,N_13522,N_13482);
xor U14360 (N_14360,N_13321,N_13733);
and U14361 (N_14361,N_13360,N_13264);
nor U14362 (N_14362,N_13355,N_13683);
xor U14363 (N_14363,N_13536,N_13710);
and U14364 (N_14364,N_13702,N_13227);
xnor U14365 (N_14365,N_13795,N_13301);
xor U14366 (N_14366,N_13652,N_13597);
or U14367 (N_14367,N_13647,N_13646);
nor U14368 (N_14368,N_13568,N_13472);
or U14369 (N_14369,N_13326,N_13211);
or U14370 (N_14370,N_13213,N_13314);
xnor U14371 (N_14371,N_13317,N_13505);
nand U14372 (N_14372,N_13594,N_13456);
xor U14373 (N_14373,N_13201,N_13764);
and U14374 (N_14374,N_13247,N_13251);
xnor U14375 (N_14375,N_13734,N_13497);
and U14376 (N_14376,N_13332,N_13626);
and U14377 (N_14377,N_13580,N_13552);
and U14378 (N_14378,N_13648,N_13482);
nor U14379 (N_14379,N_13349,N_13279);
and U14380 (N_14380,N_13729,N_13341);
or U14381 (N_14381,N_13498,N_13247);
xor U14382 (N_14382,N_13339,N_13327);
nor U14383 (N_14383,N_13207,N_13452);
nand U14384 (N_14384,N_13764,N_13333);
nand U14385 (N_14385,N_13314,N_13257);
or U14386 (N_14386,N_13461,N_13588);
xor U14387 (N_14387,N_13496,N_13618);
nor U14388 (N_14388,N_13204,N_13254);
and U14389 (N_14389,N_13392,N_13613);
xnor U14390 (N_14390,N_13595,N_13603);
and U14391 (N_14391,N_13509,N_13659);
nand U14392 (N_14392,N_13261,N_13210);
or U14393 (N_14393,N_13735,N_13318);
nand U14394 (N_14394,N_13313,N_13713);
and U14395 (N_14395,N_13747,N_13520);
nor U14396 (N_14396,N_13643,N_13688);
nand U14397 (N_14397,N_13436,N_13396);
xor U14398 (N_14398,N_13475,N_13424);
or U14399 (N_14399,N_13779,N_13255);
xor U14400 (N_14400,N_13834,N_14204);
or U14401 (N_14401,N_13896,N_13883);
nor U14402 (N_14402,N_14148,N_14058);
nor U14403 (N_14403,N_14340,N_14364);
and U14404 (N_14404,N_13993,N_14033);
nor U14405 (N_14405,N_14296,N_13940);
nor U14406 (N_14406,N_13962,N_14381);
xor U14407 (N_14407,N_14036,N_14317);
xnor U14408 (N_14408,N_14182,N_14277);
nor U14409 (N_14409,N_14184,N_14162);
xor U14410 (N_14410,N_14374,N_14105);
or U14411 (N_14411,N_13835,N_13821);
nor U14412 (N_14412,N_14074,N_14301);
nand U14413 (N_14413,N_14055,N_14202);
xor U14414 (N_14414,N_14150,N_14208);
xnor U14415 (N_14415,N_14152,N_14091);
or U14416 (N_14416,N_13840,N_14328);
nor U14417 (N_14417,N_14028,N_13944);
xor U14418 (N_14418,N_13863,N_13911);
nor U14419 (N_14419,N_14051,N_14021);
xor U14420 (N_14420,N_13918,N_13870);
nand U14421 (N_14421,N_14332,N_14156);
or U14422 (N_14422,N_14329,N_14026);
xor U14423 (N_14423,N_14214,N_14285);
xor U14424 (N_14424,N_14002,N_13963);
xnor U14425 (N_14425,N_13864,N_14312);
xor U14426 (N_14426,N_14327,N_13809);
or U14427 (N_14427,N_13984,N_13819);
nand U14428 (N_14428,N_13897,N_14271);
nor U14429 (N_14429,N_13965,N_13887);
or U14430 (N_14430,N_13970,N_13989);
xor U14431 (N_14431,N_13894,N_13941);
or U14432 (N_14432,N_14313,N_14183);
and U14433 (N_14433,N_14205,N_13899);
nor U14434 (N_14434,N_13842,N_14016);
nor U14435 (N_14435,N_13853,N_14009);
xor U14436 (N_14436,N_14114,N_14196);
nor U14437 (N_14437,N_14174,N_14286);
nor U14438 (N_14438,N_14392,N_13966);
and U14439 (N_14439,N_14001,N_14255);
nor U14440 (N_14440,N_13841,N_14014);
nand U14441 (N_14441,N_14127,N_13979);
nand U14442 (N_14442,N_14115,N_13826);
xor U14443 (N_14443,N_14319,N_14056);
and U14444 (N_14444,N_14044,N_14297);
xor U14445 (N_14445,N_13959,N_13855);
or U14446 (N_14446,N_14294,N_14275);
nor U14447 (N_14447,N_14380,N_13927);
nor U14448 (N_14448,N_13983,N_13866);
and U14449 (N_14449,N_14195,N_14180);
nor U14450 (N_14450,N_14092,N_13806);
nand U14451 (N_14451,N_14300,N_13831);
or U14452 (N_14452,N_14308,N_14052);
nand U14453 (N_14453,N_14269,N_13987);
xnor U14454 (N_14454,N_14015,N_14065);
nor U14455 (N_14455,N_14358,N_14295);
or U14456 (N_14456,N_14139,N_14355);
nor U14457 (N_14457,N_13800,N_13933);
and U14458 (N_14458,N_14071,N_13914);
nor U14459 (N_14459,N_14024,N_14228);
xor U14460 (N_14460,N_14124,N_13872);
or U14461 (N_14461,N_14304,N_14389);
or U14462 (N_14462,N_13923,N_14087);
nand U14463 (N_14463,N_13907,N_13937);
and U14464 (N_14464,N_14034,N_13879);
xor U14465 (N_14465,N_13801,N_14059);
or U14466 (N_14466,N_14060,N_14216);
xor U14467 (N_14467,N_13902,N_14106);
xnor U14468 (N_14468,N_13884,N_14070);
xnor U14469 (N_14469,N_13804,N_14351);
or U14470 (N_14470,N_14006,N_14047);
and U14471 (N_14471,N_14226,N_14221);
xor U14472 (N_14472,N_14081,N_13868);
and U14473 (N_14473,N_14191,N_13985);
or U14474 (N_14474,N_14102,N_14238);
or U14475 (N_14475,N_14069,N_13816);
xnor U14476 (N_14476,N_14222,N_13992);
nor U14477 (N_14477,N_13869,N_14395);
nand U14478 (N_14478,N_14235,N_13968);
xor U14479 (N_14479,N_14266,N_13846);
and U14480 (N_14480,N_13981,N_14223);
xnor U14481 (N_14481,N_14012,N_14163);
xor U14482 (N_14482,N_13848,N_13890);
or U14483 (N_14483,N_13861,N_13891);
and U14484 (N_14484,N_14258,N_13917);
xnor U14485 (N_14485,N_14200,N_14210);
or U14486 (N_14486,N_14085,N_13932);
nand U14487 (N_14487,N_14019,N_14178);
or U14488 (N_14488,N_14213,N_13935);
nor U14489 (N_14489,N_14372,N_14306);
nand U14490 (N_14490,N_14324,N_13929);
or U14491 (N_14491,N_14347,N_14027);
nor U14492 (N_14492,N_13916,N_14384);
xor U14493 (N_14493,N_14383,N_14088);
nand U14494 (N_14494,N_14370,N_13910);
nor U14495 (N_14495,N_14030,N_14145);
nand U14496 (N_14496,N_14382,N_14177);
and U14497 (N_14497,N_14288,N_14113);
or U14498 (N_14498,N_13847,N_13971);
or U14499 (N_14499,N_14118,N_13900);
or U14500 (N_14500,N_14217,N_14067);
nand U14501 (N_14501,N_13924,N_13943);
nor U14502 (N_14502,N_14144,N_13808);
nand U14503 (N_14503,N_13871,N_14337);
and U14504 (N_14504,N_14349,N_13803);
and U14505 (N_14505,N_14246,N_14008);
and U14506 (N_14506,N_14134,N_14287);
or U14507 (N_14507,N_14397,N_14320);
xor U14508 (N_14508,N_13920,N_14338);
or U14509 (N_14509,N_14146,N_14289);
nand U14510 (N_14510,N_13969,N_14042);
and U14511 (N_14511,N_14326,N_13998);
nand U14512 (N_14512,N_13892,N_13986);
nand U14513 (N_14513,N_14140,N_13901);
nor U14514 (N_14514,N_14386,N_13844);
or U14515 (N_14515,N_14053,N_14315);
xnor U14516 (N_14516,N_13827,N_14101);
and U14517 (N_14517,N_14108,N_14399);
nand U14518 (N_14518,N_13812,N_14198);
nand U14519 (N_14519,N_14242,N_14171);
xor U14520 (N_14520,N_13905,N_14083);
and U14521 (N_14521,N_13909,N_13802);
and U14522 (N_14522,N_14378,N_13825);
and U14523 (N_14523,N_14187,N_13858);
or U14524 (N_14524,N_13849,N_14166);
nor U14525 (N_14525,N_14253,N_13865);
and U14526 (N_14526,N_13805,N_14283);
xnor U14527 (N_14527,N_14048,N_14076);
and U14528 (N_14528,N_14369,N_13996);
nand U14529 (N_14529,N_14181,N_14151);
nor U14530 (N_14530,N_14393,N_14125);
or U14531 (N_14531,N_14259,N_13851);
or U14532 (N_14532,N_14398,N_14316);
nor U14533 (N_14533,N_13975,N_14066);
nor U14534 (N_14534,N_14190,N_14194);
nor U14535 (N_14535,N_14330,N_14334);
xor U14536 (N_14536,N_14079,N_14149);
nand U14537 (N_14537,N_13814,N_13915);
and U14538 (N_14538,N_13953,N_14078);
xnor U14539 (N_14539,N_14090,N_14251);
nand U14540 (N_14540,N_13836,N_14230);
nor U14541 (N_14541,N_14038,N_13955);
and U14542 (N_14542,N_13921,N_13919);
nor U14543 (N_14543,N_14179,N_14031);
nor U14544 (N_14544,N_14385,N_13823);
nand U14545 (N_14545,N_14344,N_13936);
nand U14546 (N_14546,N_13876,N_14335);
nor U14547 (N_14547,N_14169,N_14075);
nand U14548 (N_14548,N_13889,N_13854);
or U14549 (N_14549,N_14303,N_14023);
or U14550 (N_14550,N_13845,N_13999);
or U14551 (N_14551,N_14201,N_14314);
xnor U14552 (N_14552,N_14160,N_14360);
nand U14553 (N_14553,N_14096,N_14121);
nor U14554 (N_14554,N_14284,N_14310);
and U14555 (N_14555,N_14131,N_14130);
or U14556 (N_14556,N_14159,N_13991);
nor U14557 (N_14557,N_13873,N_14062);
or U14558 (N_14558,N_14260,N_14143);
or U14559 (N_14559,N_13925,N_14017);
nor U14560 (N_14560,N_14043,N_14290);
and U14561 (N_14561,N_13967,N_14197);
nor U14562 (N_14562,N_14274,N_14270);
and U14563 (N_14563,N_14233,N_14396);
or U14564 (N_14564,N_14354,N_13949);
nand U14565 (N_14565,N_14186,N_14005);
nand U14566 (N_14566,N_14292,N_14132);
xnor U14567 (N_14567,N_14359,N_14098);
nor U14568 (N_14568,N_13839,N_14170);
nor U14569 (N_14569,N_14388,N_14095);
and U14570 (N_14570,N_14129,N_14367);
nor U14571 (N_14571,N_13833,N_14211);
xnor U14572 (N_14572,N_13928,N_13995);
and U14573 (N_14573,N_13880,N_14199);
and U14574 (N_14574,N_14050,N_14264);
and U14575 (N_14575,N_13922,N_14352);
nor U14576 (N_14576,N_14215,N_14077);
or U14577 (N_14577,N_14120,N_14072);
nand U14578 (N_14578,N_13945,N_14248);
or U14579 (N_14579,N_14164,N_14321);
and U14580 (N_14580,N_14390,N_14080);
and U14581 (N_14581,N_14133,N_13964);
nand U14582 (N_14582,N_13973,N_14040);
xor U14583 (N_14583,N_13982,N_14203);
or U14584 (N_14584,N_13958,N_13980);
or U14585 (N_14585,N_14141,N_13837);
nor U14586 (N_14586,N_14362,N_14035);
nand U14587 (N_14587,N_14192,N_14110);
nor U14588 (N_14588,N_14346,N_14045);
xor U14589 (N_14589,N_13824,N_14161);
and U14590 (N_14590,N_13947,N_14004);
nor U14591 (N_14591,N_14020,N_13939);
and U14592 (N_14592,N_14342,N_14366);
xnor U14593 (N_14593,N_14007,N_13811);
nand U14594 (N_14594,N_14206,N_13807);
and U14595 (N_14595,N_13882,N_14307);
nor U14596 (N_14596,N_14084,N_13938);
and U14597 (N_14597,N_14176,N_14137);
and U14598 (N_14598,N_14054,N_13857);
nor U14599 (N_14599,N_14229,N_14273);
nor U14600 (N_14600,N_14231,N_13829);
xnor U14601 (N_14601,N_14357,N_14268);
or U14602 (N_14602,N_14094,N_13862);
or U14603 (N_14603,N_14138,N_13843);
nand U14604 (N_14604,N_14112,N_13926);
nor U14605 (N_14605,N_14325,N_14086);
or U14606 (N_14606,N_13815,N_14368);
and U14607 (N_14607,N_14247,N_14135);
or U14608 (N_14608,N_14291,N_14227);
or U14609 (N_14609,N_14158,N_13912);
or U14610 (N_14610,N_14254,N_13850);
and U14611 (N_14611,N_14013,N_14082);
or U14612 (N_14612,N_14039,N_14391);
and U14613 (N_14613,N_14239,N_14363);
xnor U14614 (N_14614,N_14103,N_13931);
nand U14615 (N_14615,N_14175,N_14157);
nor U14616 (N_14616,N_14123,N_13972);
nand U14617 (N_14617,N_13874,N_14350);
or U14618 (N_14618,N_14099,N_13994);
nand U14619 (N_14619,N_13978,N_13828);
nor U14620 (N_14620,N_14298,N_13852);
nor U14621 (N_14621,N_13988,N_14063);
xnor U14622 (N_14622,N_13822,N_14220);
nor U14623 (N_14623,N_14376,N_14185);
nand U14624 (N_14624,N_14377,N_13913);
and U14625 (N_14625,N_13934,N_14155);
nor U14626 (N_14626,N_13930,N_14282);
nand U14627 (N_14627,N_14100,N_14263);
xnor U14628 (N_14628,N_14212,N_14061);
or U14629 (N_14629,N_14341,N_14237);
nor U14630 (N_14630,N_14265,N_14064);
or U14631 (N_14631,N_13948,N_13952);
nand U14632 (N_14632,N_14049,N_14373);
nand U14633 (N_14633,N_14046,N_14336);
nand U14634 (N_14634,N_14029,N_13903);
xor U14635 (N_14635,N_13977,N_14257);
and U14636 (N_14636,N_13888,N_14003);
or U14637 (N_14637,N_13820,N_14224);
nor U14638 (N_14638,N_13904,N_14107);
xor U14639 (N_14639,N_14387,N_14281);
and U14640 (N_14640,N_13877,N_13898);
or U14641 (N_14641,N_13942,N_14219);
nor U14642 (N_14642,N_13867,N_14097);
and U14643 (N_14643,N_14188,N_14122);
nand U14644 (N_14644,N_14168,N_14371);
nor U14645 (N_14645,N_14037,N_13832);
or U14646 (N_14646,N_14172,N_14278);
nand U14647 (N_14647,N_14207,N_14375);
or U14648 (N_14648,N_14218,N_13908);
and U14649 (N_14649,N_14165,N_13976);
or U14650 (N_14650,N_13950,N_13878);
or U14651 (N_14651,N_13956,N_13817);
or U14652 (N_14652,N_14032,N_14331);
xnor U14653 (N_14653,N_14272,N_13946);
or U14654 (N_14654,N_13856,N_14240);
nor U14655 (N_14655,N_14142,N_14057);
and U14656 (N_14656,N_13813,N_14356);
nor U14657 (N_14657,N_13875,N_14345);
and U14658 (N_14658,N_14267,N_14116);
and U14659 (N_14659,N_14189,N_14243);
and U14660 (N_14660,N_14068,N_14153);
or U14661 (N_14661,N_14343,N_14305);
xor U14662 (N_14662,N_13886,N_13810);
xnor U14663 (N_14663,N_14323,N_14394);
or U14664 (N_14664,N_14302,N_14128);
and U14665 (N_14665,N_14348,N_13893);
nor U14666 (N_14666,N_14073,N_14109);
nand U14667 (N_14667,N_14241,N_14261);
xnor U14668 (N_14668,N_13838,N_14353);
nor U14669 (N_14669,N_14173,N_13960);
nor U14670 (N_14670,N_14322,N_14041);
xnor U14671 (N_14671,N_14147,N_13974);
and U14672 (N_14672,N_14000,N_13957);
xor U14673 (N_14673,N_13990,N_14256);
nor U14674 (N_14674,N_14311,N_14089);
or U14675 (N_14675,N_14252,N_14244);
or U14676 (N_14676,N_14293,N_14209);
and U14677 (N_14677,N_14339,N_14154);
nand U14678 (N_14678,N_14234,N_13997);
xor U14679 (N_14679,N_14361,N_14236);
xor U14680 (N_14680,N_14025,N_14119);
or U14681 (N_14681,N_14117,N_14276);
nor U14682 (N_14682,N_13895,N_14193);
and U14683 (N_14683,N_13961,N_14250);
nor U14684 (N_14684,N_14232,N_14167);
nand U14685 (N_14685,N_14379,N_14018);
or U14686 (N_14686,N_14225,N_13885);
nand U14687 (N_14687,N_13881,N_14318);
nand U14688 (N_14688,N_13954,N_14104);
xnor U14689 (N_14689,N_14111,N_13906);
nor U14690 (N_14690,N_13860,N_14333);
nand U14691 (N_14691,N_14249,N_14245);
nor U14692 (N_14692,N_14136,N_14262);
xor U14693 (N_14693,N_14279,N_14093);
xnor U14694 (N_14694,N_14365,N_13951);
and U14695 (N_14695,N_14299,N_13818);
nor U14696 (N_14696,N_14309,N_14126);
and U14697 (N_14697,N_14010,N_13830);
nand U14698 (N_14698,N_14011,N_13859);
xor U14699 (N_14699,N_14022,N_14280);
nand U14700 (N_14700,N_14064,N_14246);
nand U14701 (N_14701,N_14047,N_14108);
or U14702 (N_14702,N_13902,N_14217);
nor U14703 (N_14703,N_13855,N_14382);
and U14704 (N_14704,N_14066,N_14251);
nor U14705 (N_14705,N_14006,N_14204);
nand U14706 (N_14706,N_14077,N_14367);
xnor U14707 (N_14707,N_14206,N_14128);
nor U14708 (N_14708,N_14247,N_14215);
nand U14709 (N_14709,N_14117,N_14024);
nand U14710 (N_14710,N_14074,N_13922);
and U14711 (N_14711,N_13822,N_13900);
xor U14712 (N_14712,N_14184,N_14094);
and U14713 (N_14713,N_14294,N_14311);
nor U14714 (N_14714,N_14186,N_14105);
xor U14715 (N_14715,N_14125,N_14056);
and U14716 (N_14716,N_14316,N_14184);
and U14717 (N_14717,N_13925,N_13811);
and U14718 (N_14718,N_13804,N_13924);
nor U14719 (N_14719,N_13805,N_14266);
and U14720 (N_14720,N_13901,N_14096);
or U14721 (N_14721,N_14314,N_14039);
nand U14722 (N_14722,N_13855,N_13928);
or U14723 (N_14723,N_14276,N_13854);
nand U14724 (N_14724,N_13832,N_14345);
nor U14725 (N_14725,N_13972,N_14023);
and U14726 (N_14726,N_14084,N_13953);
nand U14727 (N_14727,N_14033,N_13882);
nand U14728 (N_14728,N_14037,N_14035);
or U14729 (N_14729,N_14229,N_14383);
xnor U14730 (N_14730,N_14137,N_14239);
nor U14731 (N_14731,N_14084,N_14203);
and U14732 (N_14732,N_14136,N_14204);
xor U14733 (N_14733,N_13817,N_14198);
nor U14734 (N_14734,N_14230,N_13834);
nand U14735 (N_14735,N_14235,N_14281);
nor U14736 (N_14736,N_13805,N_14267);
xor U14737 (N_14737,N_14352,N_13834);
nand U14738 (N_14738,N_13931,N_14086);
and U14739 (N_14739,N_14313,N_14121);
nand U14740 (N_14740,N_14270,N_14096);
and U14741 (N_14741,N_14127,N_13803);
and U14742 (N_14742,N_14232,N_14087);
nand U14743 (N_14743,N_14203,N_14108);
or U14744 (N_14744,N_13818,N_14193);
or U14745 (N_14745,N_14049,N_14208);
xnor U14746 (N_14746,N_14267,N_14106);
nand U14747 (N_14747,N_13960,N_14187);
and U14748 (N_14748,N_14187,N_14256);
and U14749 (N_14749,N_14029,N_14044);
or U14750 (N_14750,N_13981,N_13804);
xor U14751 (N_14751,N_14242,N_14005);
xor U14752 (N_14752,N_14390,N_13955);
nor U14753 (N_14753,N_13842,N_14217);
nand U14754 (N_14754,N_13833,N_14108);
and U14755 (N_14755,N_13806,N_14062);
nand U14756 (N_14756,N_14246,N_13921);
or U14757 (N_14757,N_13886,N_14294);
nand U14758 (N_14758,N_14344,N_14087);
nand U14759 (N_14759,N_13936,N_13997);
nand U14760 (N_14760,N_14367,N_14025);
xnor U14761 (N_14761,N_14190,N_13924);
nor U14762 (N_14762,N_13960,N_13992);
or U14763 (N_14763,N_14356,N_13867);
xor U14764 (N_14764,N_14110,N_14181);
and U14765 (N_14765,N_14081,N_14328);
nor U14766 (N_14766,N_13876,N_14250);
or U14767 (N_14767,N_13927,N_13853);
and U14768 (N_14768,N_13946,N_14167);
xnor U14769 (N_14769,N_14123,N_14058);
or U14770 (N_14770,N_13904,N_14377);
or U14771 (N_14771,N_14021,N_13989);
nor U14772 (N_14772,N_14115,N_14104);
xnor U14773 (N_14773,N_13854,N_13864);
and U14774 (N_14774,N_14016,N_14056);
nand U14775 (N_14775,N_14067,N_14071);
or U14776 (N_14776,N_14230,N_14012);
nand U14777 (N_14777,N_13917,N_13935);
or U14778 (N_14778,N_13806,N_13887);
or U14779 (N_14779,N_14375,N_13990);
or U14780 (N_14780,N_14118,N_14083);
xor U14781 (N_14781,N_14133,N_14384);
nand U14782 (N_14782,N_13836,N_14112);
or U14783 (N_14783,N_13812,N_13839);
and U14784 (N_14784,N_14070,N_14032);
and U14785 (N_14785,N_14135,N_14363);
xor U14786 (N_14786,N_14177,N_14179);
nand U14787 (N_14787,N_14356,N_14234);
or U14788 (N_14788,N_14223,N_13813);
nand U14789 (N_14789,N_14317,N_14216);
nor U14790 (N_14790,N_14387,N_13988);
or U14791 (N_14791,N_14114,N_14246);
xnor U14792 (N_14792,N_14071,N_14059);
xor U14793 (N_14793,N_14132,N_14157);
nor U14794 (N_14794,N_14039,N_13904);
or U14795 (N_14795,N_14294,N_14062);
or U14796 (N_14796,N_13866,N_14225);
or U14797 (N_14797,N_14217,N_13916);
and U14798 (N_14798,N_14091,N_14131);
nand U14799 (N_14799,N_14281,N_13857);
or U14800 (N_14800,N_14394,N_14041);
xnor U14801 (N_14801,N_14058,N_14121);
or U14802 (N_14802,N_14064,N_14387);
and U14803 (N_14803,N_14163,N_14197);
and U14804 (N_14804,N_14306,N_13900);
and U14805 (N_14805,N_14024,N_13849);
and U14806 (N_14806,N_13893,N_13917);
and U14807 (N_14807,N_14325,N_13850);
nor U14808 (N_14808,N_14007,N_13923);
and U14809 (N_14809,N_14365,N_14257);
xor U14810 (N_14810,N_14292,N_14375);
nor U14811 (N_14811,N_14231,N_14100);
xnor U14812 (N_14812,N_13827,N_14029);
and U14813 (N_14813,N_14334,N_13911);
nand U14814 (N_14814,N_13813,N_13884);
nor U14815 (N_14815,N_13875,N_14121);
and U14816 (N_14816,N_13962,N_14290);
or U14817 (N_14817,N_13971,N_14308);
nand U14818 (N_14818,N_14341,N_14221);
nand U14819 (N_14819,N_14075,N_13901);
nor U14820 (N_14820,N_14198,N_14389);
nor U14821 (N_14821,N_13824,N_14056);
nor U14822 (N_14822,N_14266,N_14338);
nand U14823 (N_14823,N_14351,N_14205);
and U14824 (N_14824,N_14199,N_14316);
nor U14825 (N_14825,N_14266,N_14138);
or U14826 (N_14826,N_13988,N_13931);
or U14827 (N_14827,N_14293,N_14141);
nor U14828 (N_14828,N_13987,N_14103);
or U14829 (N_14829,N_13838,N_14093);
and U14830 (N_14830,N_13836,N_14131);
nand U14831 (N_14831,N_13833,N_14188);
nand U14832 (N_14832,N_14374,N_13908);
nand U14833 (N_14833,N_14151,N_13965);
and U14834 (N_14834,N_14221,N_13964);
or U14835 (N_14835,N_14372,N_14309);
and U14836 (N_14836,N_14027,N_14254);
and U14837 (N_14837,N_13820,N_13804);
or U14838 (N_14838,N_14189,N_14370);
xor U14839 (N_14839,N_13939,N_13972);
nand U14840 (N_14840,N_13968,N_14373);
xnor U14841 (N_14841,N_14336,N_13899);
nand U14842 (N_14842,N_14359,N_14101);
nand U14843 (N_14843,N_14041,N_14091);
xor U14844 (N_14844,N_14387,N_13967);
nand U14845 (N_14845,N_14382,N_14267);
or U14846 (N_14846,N_14338,N_13927);
nor U14847 (N_14847,N_14100,N_13809);
and U14848 (N_14848,N_14310,N_14045);
or U14849 (N_14849,N_13988,N_14090);
and U14850 (N_14850,N_13864,N_14028);
nand U14851 (N_14851,N_14389,N_13915);
and U14852 (N_14852,N_13822,N_14107);
or U14853 (N_14853,N_14245,N_14151);
xor U14854 (N_14854,N_14181,N_13822);
xnor U14855 (N_14855,N_13890,N_14218);
nor U14856 (N_14856,N_13853,N_13826);
nand U14857 (N_14857,N_14302,N_13967);
xor U14858 (N_14858,N_13817,N_14130);
xor U14859 (N_14859,N_13996,N_13908);
and U14860 (N_14860,N_14300,N_13819);
nand U14861 (N_14861,N_14020,N_13981);
or U14862 (N_14862,N_13927,N_13847);
nor U14863 (N_14863,N_14302,N_13952);
nand U14864 (N_14864,N_14211,N_14034);
nand U14865 (N_14865,N_14299,N_13812);
and U14866 (N_14866,N_14350,N_13851);
or U14867 (N_14867,N_14035,N_14077);
and U14868 (N_14868,N_13832,N_14060);
nand U14869 (N_14869,N_14246,N_14134);
and U14870 (N_14870,N_14153,N_13945);
nand U14871 (N_14871,N_14039,N_13853);
nand U14872 (N_14872,N_14138,N_14374);
nor U14873 (N_14873,N_13843,N_14224);
and U14874 (N_14874,N_14188,N_14372);
nand U14875 (N_14875,N_13962,N_14065);
nor U14876 (N_14876,N_14326,N_13955);
xor U14877 (N_14877,N_14140,N_13944);
xor U14878 (N_14878,N_14070,N_14084);
xor U14879 (N_14879,N_13914,N_14357);
nor U14880 (N_14880,N_14015,N_13960);
nand U14881 (N_14881,N_14234,N_14073);
nor U14882 (N_14882,N_14011,N_14277);
nand U14883 (N_14883,N_14305,N_14023);
nor U14884 (N_14884,N_14144,N_13901);
nand U14885 (N_14885,N_13860,N_14019);
and U14886 (N_14886,N_13831,N_14308);
xnor U14887 (N_14887,N_13892,N_14045);
xor U14888 (N_14888,N_13894,N_14095);
nor U14889 (N_14889,N_13969,N_14276);
xor U14890 (N_14890,N_14354,N_13866);
and U14891 (N_14891,N_14267,N_13817);
nor U14892 (N_14892,N_14276,N_14359);
nand U14893 (N_14893,N_13958,N_14338);
nor U14894 (N_14894,N_14053,N_14312);
nor U14895 (N_14895,N_13808,N_14126);
or U14896 (N_14896,N_13923,N_14387);
nand U14897 (N_14897,N_14082,N_14107);
and U14898 (N_14898,N_13839,N_13817);
or U14899 (N_14899,N_13800,N_14357);
nand U14900 (N_14900,N_14160,N_14184);
or U14901 (N_14901,N_14041,N_14071);
or U14902 (N_14902,N_13849,N_14089);
xnor U14903 (N_14903,N_14123,N_14292);
xnor U14904 (N_14904,N_13999,N_14057);
and U14905 (N_14905,N_14368,N_14242);
or U14906 (N_14906,N_14231,N_13964);
and U14907 (N_14907,N_14383,N_14040);
nor U14908 (N_14908,N_14241,N_14113);
xor U14909 (N_14909,N_14397,N_13961);
nor U14910 (N_14910,N_14393,N_13992);
or U14911 (N_14911,N_13980,N_14107);
or U14912 (N_14912,N_13955,N_14334);
and U14913 (N_14913,N_14364,N_14366);
xor U14914 (N_14914,N_14309,N_13857);
xor U14915 (N_14915,N_14170,N_14075);
or U14916 (N_14916,N_13929,N_13943);
nand U14917 (N_14917,N_14136,N_14396);
nor U14918 (N_14918,N_14061,N_13866);
or U14919 (N_14919,N_14190,N_14180);
xor U14920 (N_14920,N_13820,N_14011);
and U14921 (N_14921,N_13944,N_14258);
nand U14922 (N_14922,N_13890,N_13904);
and U14923 (N_14923,N_13811,N_13924);
nand U14924 (N_14924,N_14160,N_14059);
and U14925 (N_14925,N_13968,N_14144);
nand U14926 (N_14926,N_14084,N_14360);
and U14927 (N_14927,N_14367,N_14187);
xnor U14928 (N_14928,N_13867,N_14209);
xor U14929 (N_14929,N_14359,N_13919);
xnor U14930 (N_14930,N_14258,N_14173);
and U14931 (N_14931,N_14162,N_14000);
nand U14932 (N_14932,N_14065,N_14183);
and U14933 (N_14933,N_14204,N_13917);
nand U14934 (N_14934,N_14206,N_13823);
nor U14935 (N_14935,N_14238,N_14209);
or U14936 (N_14936,N_13870,N_14284);
xor U14937 (N_14937,N_14317,N_13999);
and U14938 (N_14938,N_13927,N_13951);
nor U14939 (N_14939,N_13867,N_13850);
xnor U14940 (N_14940,N_14304,N_13945);
or U14941 (N_14941,N_14101,N_14122);
nor U14942 (N_14942,N_14054,N_14230);
nand U14943 (N_14943,N_13831,N_14223);
and U14944 (N_14944,N_14300,N_13859);
nor U14945 (N_14945,N_14191,N_13997);
nor U14946 (N_14946,N_14330,N_14076);
or U14947 (N_14947,N_13943,N_13816);
or U14948 (N_14948,N_14238,N_13953);
and U14949 (N_14949,N_14023,N_14229);
nor U14950 (N_14950,N_13847,N_14226);
and U14951 (N_14951,N_14344,N_14047);
nand U14952 (N_14952,N_14246,N_14378);
and U14953 (N_14953,N_13991,N_14078);
and U14954 (N_14954,N_13945,N_13833);
and U14955 (N_14955,N_13876,N_13893);
nand U14956 (N_14956,N_14036,N_14048);
nor U14957 (N_14957,N_13916,N_13804);
or U14958 (N_14958,N_14213,N_14209);
or U14959 (N_14959,N_14285,N_14181);
nor U14960 (N_14960,N_14168,N_14227);
nand U14961 (N_14961,N_13836,N_14243);
nand U14962 (N_14962,N_14098,N_13945);
nand U14963 (N_14963,N_13955,N_13958);
and U14964 (N_14964,N_14233,N_14039);
nor U14965 (N_14965,N_14317,N_14024);
nor U14966 (N_14966,N_14220,N_13926);
or U14967 (N_14967,N_13900,N_14244);
xnor U14968 (N_14968,N_14079,N_13829);
xnor U14969 (N_14969,N_14339,N_14025);
nand U14970 (N_14970,N_14022,N_14101);
xnor U14971 (N_14971,N_13927,N_14244);
nor U14972 (N_14972,N_14079,N_14262);
xor U14973 (N_14973,N_14011,N_14368);
nor U14974 (N_14974,N_14205,N_13969);
xor U14975 (N_14975,N_13946,N_14221);
nand U14976 (N_14976,N_13806,N_13872);
nand U14977 (N_14977,N_14086,N_14031);
xnor U14978 (N_14978,N_14291,N_14059);
xor U14979 (N_14979,N_13834,N_14041);
or U14980 (N_14980,N_14018,N_13818);
nand U14981 (N_14981,N_13901,N_14247);
nand U14982 (N_14982,N_14220,N_14286);
nor U14983 (N_14983,N_14109,N_13911);
nor U14984 (N_14984,N_14332,N_13811);
and U14985 (N_14985,N_13907,N_13908);
or U14986 (N_14986,N_14351,N_13961);
nor U14987 (N_14987,N_13964,N_13891);
or U14988 (N_14988,N_14093,N_14108);
and U14989 (N_14989,N_14138,N_13871);
nand U14990 (N_14990,N_14264,N_14143);
and U14991 (N_14991,N_14076,N_13911);
nand U14992 (N_14992,N_14131,N_14066);
and U14993 (N_14993,N_14081,N_14259);
nand U14994 (N_14994,N_14095,N_14009);
and U14995 (N_14995,N_14068,N_14125);
or U14996 (N_14996,N_14179,N_13970);
and U14997 (N_14997,N_14068,N_14026);
nor U14998 (N_14998,N_14047,N_14011);
xnor U14999 (N_14999,N_14222,N_13892);
xor U15000 (N_15000,N_14934,N_14938);
nor U15001 (N_15001,N_14536,N_14486);
xor U15002 (N_15002,N_14549,N_14501);
or U15003 (N_15003,N_14421,N_14449);
or U15004 (N_15004,N_14492,N_14961);
nor U15005 (N_15005,N_14940,N_14650);
nor U15006 (N_15006,N_14956,N_14516);
or U15007 (N_15007,N_14822,N_14728);
or U15008 (N_15008,N_14812,N_14519);
nor U15009 (N_15009,N_14455,N_14733);
or U15010 (N_15010,N_14607,N_14580);
xor U15011 (N_15011,N_14844,N_14847);
nor U15012 (N_15012,N_14843,N_14887);
nor U15013 (N_15013,N_14852,N_14727);
xor U15014 (N_15014,N_14703,N_14625);
and U15015 (N_15015,N_14986,N_14929);
or U15016 (N_15016,N_14636,N_14765);
nor U15017 (N_15017,N_14442,N_14484);
or U15018 (N_15018,N_14820,N_14846);
and U15019 (N_15019,N_14634,N_14572);
and U15020 (N_15020,N_14534,N_14706);
xor U15021 (N_15021,N_14711,N_14584);
nand U15022 (N_15022,N_14712,N_14689);
nor U15023 (N_15023,N_14759,N_14893);
nor U15024 (N_15024,N_14813,N_14988);
or U15025 (N_15025,N_14952,N_14563);
xnor U15026 (N_15026,N_14818,N_14444);
or U15027 (N_15027,N_14408,N_14792);
or U15028 (N_15028,N_14609,N_14453);
nand U15029 (N_15029,N_14987,N_14973);
nor U15030 (N_15030,N_14983,N_14799);
and U15031 (N_15031,N_14806,N_14640);
nor U15032 (N_15032,N_14658,N_14856);
xnor U15033 (N_15033,N_14862,N_14611);
or U15034 (N_15034,N_14979,N_14530);
nor U15035 (N_15035,N_14981,N_14466);
and U15036 (N_15036,N_14606,N_14838);
nand U15037 (N_15037,N_14477,N_14702);
or U15038 (N_15038,N_14890,N_14997);
nor U15039 (N_15039,N_14507,N_14815);
nand U15040 (N_15040,N_14608,N_14425);
xnor U15041 (N_15041,N_14655,N_14430);
and U15042 (N_15042,N_14747,N_14674);
nor U15043 (N_15043,N_14701,N_14744);
nand U15044 (N_15044,N_14600,N_14539);
and U15045 (N_15045,N_14896,N_14676);
nor U15046 (N_15046,N_14552,N_14837);
nor U15047 (N_15047,N_14889,N_14564);
xor U15048 (N_15048,N_14497,N_14710);
nand U15049 (N_15049,N_14402,N_14863);
xor U15050 (N_15050,N_14808,N_14443);
nor U15051 (N_15051,N_14908,N_14754);
or U15052 (N_15052,N_14433,N_14472);
and U15053 (N_15053,N_14639,N_14831);
and U15054 (N_15054,N_14631,N_14581);
or U15055 (N_15055,N_14502,N_14735);
nand U15056 (N_15056,N_14827,N_14500);
nand U15057 (N_15057,N_14478,N_14594);
and U15058 (N_15058,N_14692,N_14816);
xnor U15059 (N_15059,N_14599,N_14664);
and U15060 (N_15060,N_14616,N_14883);
xor U15061 (N_15061,N_14811,N_14546);
nor U15062 (N_15062,N_14524,N_14912);
xor U15063 (N_15063,N_14510,N_14752);
nor U15064 (N_15064,N_14437,N_14750);
and U15065 (N_15065,N_14753,N_14766);
or U15066 (N_15066,N_14420,N_14659);
nand U15067 (N_15067,N_14434,N_14723);
nand U15068 (N_15068,N_14762,N_14669);
nor U15069 (N_15069,N_14646,N_14993);
nand U15070 (N_15070,N_14736,N_14790);
nor U15071 (N_15071,N_14622,N_14508);
nand U15072 (N_15072,N_14869,N_14638);
nor U15073 (N_15073,N_14892,N_14468);
xnor U15074 (N_15074,N_14605,N_14457);
and U15075 (N_15075,N_14708,N_14517);
and U15076 (N_15076,N_14469,N_14568);
or U15077 (N_15077,N_14514,N_14737);
nor U15078 (N_15078,N_14629,N_14794);
xor U15079 (N_15079,N_14906,N_14476);
nand U15080 (N_15080,N_14699,N_14675);
nand U15081 (N_15081,N_14910,N_14898);
nand U15082 (N_15082,N_14569,N_14967);
or U15083 (N_15083,N_14884,N_14968);
or U15084 (N_15084,N_14464,N_14984);
or U15085 (N_15085,N_14496,N_14819);
and U15086 (N_15086,N_14795,N_14465);
and U15087 (N_15087,N_14757,N_14459);
xor U15088 (N_15088,N_14770,N_14949);
xor U15089 (N_15089,N_14401,N_14784);
nor U15090 (N_15090,N_14687,N_14876);
xnor U15091 (N_15091,N_14858,N_14541);
and U15092 (N_15092,N_14579,N_14738);
xnor U15093 (N_15093,N_14920,N_14917);
xor U15094 (N_15094,N_14974,N_14695);
nand U15095 (N_15095,N_14543,N_14957);
or U15096 (N_15096,N_14978,N_14644);
nor U15097 (N_15097,N_14416,N_14592);
and U15098 (N_15098,N_14999,N_14996);
or U15099 (N_15099,N_14963,N_14542);
and U15100 (N_15100,N_14722,N_14427);
nor U15101 (N_15101,N_14960,N_14495);
xor U15102 (N_15102,N_14840,N_14589);
nand U15103 (N_15103,N_14716,N_14897);
or U15104 (N_15104,N_14781,N_14405);
and U15105 (N_15105,N_14797,N_14485);
xnor U15106 (N_15106,N_14732,N_14900);
xnor U15107 (N_15107,N_14774,N_14587);
xnor U15108 (N_15108,N_14585,N_14947);
or U15109 (N_15109,N_14918,N_14551);
and U15110 (N_15110,N_14678,N_14943);
or U15111 (N_15111,N_14407,N_14936);
nand U15112 (N_15112,N_14554,N_14414);
nand U15113 (N_15113,N_14796,N_14419);
xor U15114 (N_15114,N_14870,N_14595);
or U15115 (N_15115,N_14432,N_14426);
xnor U15116 (N_15116,N_14707,N_14801);
nand U15117 (N_15117,N_14868,N_14654);
nor U15118 (N_15118,N_14962,N_14673);
nand U15119 (N_15119,N_14612,N_14730);
nor U15120 (N_15120,N_14901,N_14959);
or U15121 (N_15121,N_14866,N_14994);
nand U15122 (N_15122,N_14793,N_14621);
nand U15123 (N_15123,N_14851,N_14691);
xor U15124 (N_15124,N_14891,N_14470);
nand U15125 (N_15125,N_14904,N_14877);
nor U15126 (N_15126,N_14657,N_14902);
and U15127 (N_15127,N_14990,N_14849);
nand U15128 (N_15128,N_14586,N_14950);
xor U15129 (N_15129,N_14450,N_14548);
nor U15130 (N_15130,N_14680,N_14977);
or U15131 (N_15131,N_14926,N_14550);
nand U15132 (N_15132,N_14985,N_14488);
nand U15133 (N_15133,N_14888,N_14776);
or U15134 (N_15134,N_14919,N_14588);
nor U15135 (N_15135,N_14915,N_14821);
or U15136 (N_15136,N_14859,N_14941);
xnor U15137 (N_15137,N_14647,N_14415);
nand U15138 (N_15138,N_14682,N_14665);
or U15139 (N_15139,N_14544,N_14422);
nand U15140 (N_15140,N_14679,N_14574);
or U15141 (N_15141,N_14475,N_14506);
nand U15142 (N_15142,N_14604,N_14829);
nor U15143 (N_15143,N_14429,N_14835);
xor U15144 (N_15144,N_14786,N_14970);
nor U15145 (N_15145,N_14787,N_14481);
nand U15146 (N_15146,N_14498,N_14452);
or U15147 (N_15147,N_14954,N_14560);
and U15148 (N_15148,N_14535,N_14914);
or U15149 (N_15149,N_14965,N_14596);
nor U15150 (N_15150,N_14583,N_14700);
or U15151 (N_15151,N_14532,N_14881);
nor U15152 (N_15152,N_14593,N_14839);
nor U15153 (N_15153,N_14690,N_14761);
and U15154 (N_15154,N_14767,N_14930);
or U15155 (N_15155,N_14751,N_14779);
nand U15156 (N_15156,N_14513,N_14515);
nor U15157 (N_15157,N_14558,N_14688);
nor U15158 (N_15158,N_14576,N_14719);
xnor U15159 (N_15159,N_14597,N_14696);
or U15160 (N_15160,N_14663,N_14782);
nor U15161 (N_15161,N_14531,N_14742);
nor U15162 (N_15162,N_14505,N_14697);
nor U15163 (N_15163,N_14619,N_14975);
nor U15164 (N_15164,N_14971,N_14503);
nor U15165 (N_15165,N_14942,N_14482);
xnor U15166 (N_15166,N_14578,N_14463);
xnor U15167 (N_15167,N_14741,N_14487);
or U15168 (N_15168,N_14721,N_14561);
nor U15169 (N_15169,N_14436,N_14684);
or U15170 (N_15170,N_14922,N_14830);
nor U15171 (N_15171,N_14760,N_14885);
and U15172 (N_15172,N_14805,N_14617);
and U15173 (N_15173,N_14935,N_14860);
and U15174 (N_15174,N_14410,N_14494);
xnor U15175 (N_15175,N_14804,N_14791);
xnor U15176 (N_15176,N_14528,N_14763);
nand U15177 (N_15177,N_14573,N_14409);
nand U15178 (N_15178,N_14803,N_14903);
or U15179 (N_15179,N_14526,N_14880);
and U15180 (N_15180,N_14406,N_14927);
and U15181 (N_15181,N_14603,N_14861);
nand U15182 (N_15182,N_14772,N_14718);
xnor U15183 (N_15183,N_14704,N_14418);
xnor U15184 (N_15184,N_14886,N_14709);
xor U15185 (N_15185,N_14648,N_14567);
nand U15186 (N_15186,N_14853,N_14571);
and U15187 (N_15187,N_14633,N_14642);
nor U15188 (N_15188,N_14411,N_14400);
and U15189 (N_15189,N_14537,N_14857);
nand U15190 (N_15190,N_14615,N_14909);
xor U15191 (N_15191,N_14991,N_14431);
xor U15192 (N_15192,N_14995,N_14511);
xor U15193 (N_15193,N_14945,N_14557);
nand U15194 (N_15194,N_14899,N_14848);
and U15195 (N_15195,N_14756,N_14445);
nor U15196 (N_15196,N_14480,N_14789);
nor U15197 (N_15197,N_14923,N_14916);
and U15198 (N_15198,N_14458,N_14948);
xnor U15199 (N_15199,N_14538,N_14834);
nand U15200 (N_15200,N_14800,N_14823);
and U15201 (N_15201,N_14447,N_14656);
xnor U15202 (N_15202,N_14833,N_14518);
nand U15203 (N_15203,N_14778,N_14643);
nand U15204 (N_15204,N_14933,N_14632);
and U15205 (N_15205,N_14668,N_14683);
xnor U15206 (N_15206,N_14921,N_14471);
nor U15207 (N_15207,N_14745,N_14527);
nor U15208 (N_15208,N_14871,N_14545);
or U15209 (N_15209,N_14972,N_14652);
nand U15210 (N_15210,N_14951,N_14928);
or U15211 (N_15211,N_14435,N_14764);
nor U15212 (N_15212,N_14473,N_14743);
xnor U15213 (N_15213,N_14525,N_14637);
or U15214 (N_15214,N_14911,N_14467);
nand U15215 (N_15215,N_14602,N_14523);
xnor U15216 (N_15216,N_14694,N_14832);
or U15217 (N_15217,N_14842,N_14980);
nor U15218 (N_15218,N_14932,N_14685);
nand U15219 (N_15219,N_14556,N_14490);
and U15220 (N_15220,N_14651,N_14613);
xnor U15221 (N_15221,N_14964,N_14966);
and U15222 (N_15222,N_14755,N_14662);
nand U15223 (N_15223,N_14953,N_14729);
xnor U15224 (N_15224,N_14645,N_14769);
nand U15225 (N_15225,N_14865,N_14748);
and U15226 (N_15226,N_14715,N_14417);
xnor U15227 (N_15227,N_14734,N_14758);
nand U15228 (N_15228,N_14522,N_14521);
nor U15229 (N_15229,N_14714,N_14937);
and U15230 (N_15230,N_14626,N_14448);
nand U15231 (N_15231,N_14771,N_14504);
xor U15232 (N_15232,N_14698,N_14681);
or U15233 (N_15233,N_14824,N_14677);
and U15234 (N_15234,N_14817,N_14717);
nor U15235 (N_15235,N_14461,N_14777);
and U15236 (N_15236,N_14570,N_14614);
nor U15237 (N_15237,N_14802,N_14479);
nand U15238 (N_15238,N_14864,N_14850);
or U15239 (N_15239,N_14720,N_14628);
nor U15240 (N_15240,N_14577,N_14731);
and U15241 (N_15241,N_14841,N_14559);
xor U15242 (N_15242,N_14575,N_14491);
xor U15243 (N_15243,N_14451,N_14529);
nor U15244 (N_15244,N_14867,N_14775);
nand U15245 (N_15245,N_14660,N_14810);
or U15246 (N_15246,N_14998,N_14671);
nor U15247 (N_15247,N_14992,N_14454);
or U15248 (N_15248,N_14661,N_14913);
nor U15249 (N_15249,N_14509,N_14746);
nand U15250 (N_15250,N_14931,N_14836);
or U15251 (N_15251,N_14894,N_14483);
nand U15252 (N_15252,N_14749,N_14873);
nand U15253 (N_15253,N_14783,N_14713);
nor U15254 (N_15254,N_14825,N_14565);
xor U15255 (N_15255,N_14872,N_14944);
and U15256 (N_15256,N_14582,N_14845);
or U15257 (N_15257,N_14724,N_14649);
and U15258 (N_15258,N_14785,N_14474);
and U15259 (N_15259,N_14627,N_14424);
nor U15260 (N_15260,N_14441,N_14591);
xor U15261 (N_15261,N_14958,N_14925);
nor U15262 (N_15262,N_14882,N_14540);
nand U15263 (N_15263,N_14989,N_14404);
xnor U15264 (N_15264,N_14726,N_14423);
nor U15265 (N_15265,N_14826,N_14946);
and U15266 (N_15266,N_14982,N_14428);
or U15267 (N_15267,N_14555,N_14601);
and U15268 (N_15268,N_14905,N_14439);
nand U15269 (N_15269,N_14499,N_14854);
nor U15270 (N_15270,N_14623,N_14403);
xor U15271 (N_15271,N_14641,N_14788);
and U15272 (N_15272,N_14686,N_14666);
xor U15273 (N_15273,N_14879,N_14493);
or U15274 (N_15274,N_14547,N_14725);
xnor U15275 (N_15275,N_14462,N_14553);
and U15276 (N_15276,N_14955,N_14630);
xor U15277 (N_15277,N_14667,N_14907);
xor U15278 (N_15278,N_14412,N_14939);
and U15279 (N_15279,N_14620,N_14512);
nand U15280 (N_15280,N_14670,N_14807);
xnor U15281 (N_15281,N_14874,N_14693);
nor U15282 (N_15282,N_14740,N_14924);
nand U15283 (N_15283,N_14976,N_14878);
nor U15284 (N_15284,N_14413,N_14855);
xor U15285 (N_15285,N_14672,N_14895);
or U15286 (N_15286,N_14520,N_14828);
or U15287 (N_15287,N_14533,N_14809);
nor U15288 (N_15288,N_14798,N_14610);
and U15289 (N_15289,N_14598,N_14456);
and U15290 (N_15290,N_14814,N_14875);
and U15291 (N_15291,N_14566,N_14438);
nand U15292 (N_15292,N_14739,N_14969);
nand U15293 (N_15293,N_14590,N_14773);
xor U15294 (N_15294,N_14624,N_14489);
nor U15295 (N_15295,N_14653,N_14440);
and U15296 (N_15296,N_14780,N_14460);
nand U15297 (N_15297,N_14562,N_14446);
and U15298 (N_15298,N_14768,N_14705);
and U15299 (N_15299,N_14618,N_14635);
or U15300 (N_15300,N_14867,N_14832);
or U15301 (N_15301,N_14878,N_14483);
nor U15302 (N_15302,N_14951,N_14644);
nand U15303 (N_15303,N_14824,N_14561);
and U15304 (N_15304,N_14623,N_14959);
or U15305 (N_15305,N_14897,N_14416);
xor U15306 (N_15306,N_14456,N_14707);
nor U15307 (N_15307,N_14911,N_14713);
or U15308 (N_15308,N_14571,N_14968);
or U15309 (N_15309,N_14891,N_14808);
nand U15310 (N_15310,N_14921,N_14941);
xor U15311 (N_15311,N_14426,N_14909);
and U15312 (N_15312,N_14678,N_14614);
nor U15313 (N_15313,N_14699,N_14822);
nand U15314 (N_15314,N_14477,N_14859);
nor U15315 (N_15315,N_14999,N_14956);
xor U15316 (N_15316,N_14440,N_14473);
nor U15317 (N_15317,N_14787,N_14946);
and U15318 (N_15318,N_14692,N_14650);
and U15319 (N_15319,N_14612,N_14562);
and U15320 (N_15320,N_14860,N_14532);
nor U15321 (N_15321,N_14636,N_14953);
or U15322 (N_15322,N_14831,N_14493);
nand U15323 (N_15323,N_14597,N_14668);
and U15324 (N_15324,N_14774,N_14420);
nor U15325 (N_15325,N_14569,N_14809);
xnor U15326 (N_15326,N_14839,N_14568);
and U15327 (N_15327,N_14947,N_14415);
nor U15328 (N_15328,N_14431,N_14447);
and U15329 (N_15329,N_14606,N_14939);
and U15330 (N_15330,N_14631,N_14409);
nand U15331 (N_15331,N_14685,N_14989);
or U15332 (N_15332,N_14656,N_14750);
nand U15333 (N_15333,N_14533,N_14777);
nand U15334 (N_15334,N_14786,N_14711);
nor U15335 (N_15335,N_14677,N_14704);
or U15336 (N_15336,N_14825,N_14441);
nor U15337 (N_15337,N_14466,N_14597);
nand U15338 (N_15338,N_14717,N_14487);
nor U15339 (N_15339,N_14872,N_14996);
and U15340 (N_15340,N_14434,N_14962);
nand U15341 (N_15341,N_14773,N_14869);
xor U15342 (N_15342,N_14985,N_14942);
xor U15343 (N_15343,N_14414,N_14910);
xnor U15344 (N_15344,N_14477,N_14724);
and U15345 (N_15345,N_14627,N_14959);
and U15346 (N_15346,N_14883,N_14562);
xor U15347 (N_15347,N_14971,N_14870);
nor U15348 (N_15348,N_14661,N_14986);
and U15349 (N_15349,N_14746,N_14912);
nor U15350 (N_15350,N_14934,N_14765);
or U15351 (N_15351,N_14983,N_14949);
xnor U15352 (N_15352,N_14896,N_14591);
xnor U15353 (N_15353,N_14460,N_14708);
and U15354 (N_15354,N_14928,N_14835);
nand U15355 (N_15355,N_14776,N_14690);
xor U15356 (N_15356,N_14989,N_14412);
and U15357 (N_15357,N_14840,N_14486);
nand U15358 (N_15358,N_14730,N_14683);
xnor U15359 (N_15359,N_14473,N_14483);
or U15360 (N_15360,N_14453,N_14472);
nand U15361 (N_15361,N_14589,N_14913);
and U15362 (N_15362,N_14598,N_14681);
or U15363 (N_15363,N_14425,N_14853);
or U15364 (N_15364,N_14541,N_14554);
nand U15365 (N_15365,N_14909,N_14686);
or U15366 (N_15366,N_14855,N_14627);
nand U15367 (N_15367,N_14480,N_14910);
or U15368 (N_15368,N_14539,N_14861);
nor U15369 (N_15369,N_14749,N_14637);
nor U15370 (N_15370,N_14648,N_14630);
nor U15371 (N_15371,N_14543,N_14581);
and U15372 (N_15372,N_14595,N_14944);
and U15373 (N_15373,N_14614,N_14855);
nor U15374 (N_15374,N_14584,N_14495);
or U15375 (N_15375,N_14979,N_14461);
xnor U15376 (N_15376,N_14931,N_14473);
and U15377 (N_15377,N_14614,N_14511);
nand U15378 (N_15378,N_14915,N_14690);
xnor U15379 (N_15379,N_14494,N_14717);
xor U15380 (N_15380,N_14456,N_14471);
nor U15381 (N_15381,N_14885,N_14731);
xnor U15382 (N_15382,N_14742,N_14759);
nand U15383 (N_15383,N_14415,N_14659);
nand U15384 (N_15384,N_14509,N_14517);
xnor U15385 (N_15385,N_14989,N_14575);
nand U15386 (N_15386,N_14844,N_14939);
xnor U15387 (N_15387,N_14515,N_14995);
xnor U15388 (N_15388,N_14800,N_14428);
or U15389 (N_15389,N_14598,N_14980);
nor U15390 (N_15390,N_14881,N_14417);
and U15391 (N_15391,N_14412,N_14680);
xnor U15392 (N_15392,N_14635,N_14568);
and U15393 (N_15393,N_14986,N_14651);
nand U15394 (N_15394,N_14635,N_14538);
xor U15395 (N_15395,N_14894,N_14721);
xor U15396 (N_15396,N_14463,N_14656);
xor U15397 (N_15397,N_14443,N_14935);
nor U15398 (N_15398,N_14621,N_14854);
nor U15399 (N_15399,N_14628,N_14455);
and U15400 (N_15400,N_14722,N_14830);
and U15401 (N_15401,N_14817,N_14928);
nor U15402 (N_15402,N_14400,N_14923);
or U15403 (N_15403,N_14955,N_14668);
nor U15404 (N_15404,N_14608,N_14751);
xnor U15405 (N_15405,N_14724,N_14542);
xnor U15406 (N_15406,N_14455,N_14450);
and U15407 (N_15407,N_14475,N_14788);
or U15408 (N_15408,N_14726,N_14422);
xnor U15409 (N_15409,N_14438,N_14546);
nor U15410 (N_15410,N_14439,N_14407);
nor U15411 (N_15411,N_14558,N_14481);
nor U15412 (N_15412,N_14981,N_14680);
nor U15413 (N_15413,N_14562,N_14656);
nor U15414 (N_15414,N_14814,N_14927);
xor U15415 (N_15415,N_14947,N_14434);
nor U15416 (N_15416,N_14507,N_14745);
nand U15417 (N_15417,N_14889,N_14812);
nand U15418 (N_15418,N_14469,N_14512);
nor U15419 (N_15419,N_14884,N_14771);
nor U15420 (N_15420,N_14614,N_14813);
xor U15421 (N_15421,N_14421,N_14668);
xor U15422 (N_15422,N_14679,N_14584);
nand U15423 (N_15423,N_14664,N_14758);
nand U15424 (N_15424,N_14780,N_14732);
nor U15425 (N_15425,N_14889,N_14976);
nor U15426 (N_15426,N_14943,N_14957);
or U15427 (N_15427,N_14696,N_14606);
nand U15428 (N_15428,N_14577,N_14542);
or U15429 (N_15429,N_14730,N_14702);
nor U15430 (N_15430,N_14865,N_14945);
xor U15431 (N_15431,N_14872,N_14867);
or U15432 (N_15432,N_14912,N_14842);
xnor U15433 (N_15433,N_14428,N_14828);
nand U15434 (N_15434,N_14738,N_14631);
and U15435 (N_15435,N_14716,N_14686);
xnor U15436 (N_15436,N_14475,N_14460);
or U15437 (N_15437,N_14819,N_14553);
nand U15438 (N_15438,N_14762,N_14981);
xor U15439 (N_15439,N_14914,N_14697);
or U15440 (N_15440,N_14598,N_14793);
nand U15441 (N_15441,N_14774,N_14573);
nor U15442 (N_15442,N_14883,N_14593);
nor U15443 (N_15443,N_14501,N_14627);
nand U15444 (N_15444,N_14430,N_14511);
and U15445 (N_15445,N_14738,N_14951);
and U15446 (N_15446,N_14767,N_14939);
or U15447 (N_15447,N_14762,N_14989);
nand U15448 (N_15448,N_14716,N_14778);
and U15449 (N_15449,N_14889,N_14826);
nor U15450 (N_15450,N_14466,N_14810);
xor U15451 (N_15451,N_14623,N_14918);
nand U15452 (N_15452,N_14452,N_14935);
nand U15453 (N_15453,N_14727,N_14634);
xnor U15454 (N_15454,N_14841,N_14953);
xor U15455 (N_15455,N_14661,N_14614);
or U15456 (N_15456,N_14924,N_14693);
or U15457 (N_15457,N_14778,N_14970);
and U15458 (N_15458,N_14551,N_14656);
nor U15459 (N_15459,N_14683,N_14948);
and U15460 (N_15460,N_14854,N_14984);
or U15461 (N_15461,N_14597,N_14501);
and U15462 (N_15462,N_14947,N_14912);
or U15463 (N_15463,N_14671,N_14873);
nor U15464 (N_15464,N_14566,N_14808);
or U15465 (N_15465,N_14979,N_14774);
nor U15466 (N_15466,N_14834,N_14982);
nand U15467 (N_15467,N_14706,N_14635);
xor U15468 (N_15468,N_14620,N_14934);
nand U15469 (N_15469,N_14966,N_14550);
and U15470 (N_15470,N_14572,N_14817);
nor U15471 (N_15471,N_14447,N_14516);
xor U15472 (N_15472,N_14472,N_14676);
nand U15473 (N_15473,N_14678,N_14915);
nand U15474 (N_15474,N_14908,N_14918);
xnor U15475 (N_15475,N_14411,N_14998);
nor U15476 (N_15476,N_14739,N_14492);
nand U15477 (N_15477,N_14886,N_14968);
xor U15478 (N_15478,N_14505,N_14422);
or U15479 (N_15479,N_14838,N_14955);
and U15480 (N_15480,N_14583,N_14855);
or U15481 (N_15481,N_14776,N_14902);
and U15482 (N_15482,N_14517,N_14989);
or U15483 (N_15483,N_14692,N_14697);
nor U15484 (N_15484,N_14429,N_14915);
nand U15485 (N_15485,N_14757,N_14833);
nand U15486 (N_15486,N_14459,N_14947);
and U15487 (N_15487,N_14704,N_14528);
or U15488 (N_15488,N_14563,N_14574);
xnor U15489 (N_15489,N_14461,N_14651);
nor U15490 (N_15490,N_14456,N_14624);
or U15491 (N_15491,N_14679,N_14680);
nand U15492 (N_15492,N_14409,N_14437);
nor U15493 (N_15493,N_14486,N_14561);
xor U15494 (N_15494,N_14634,N_14766);
nor U15495 (N_15495,N_14418,N_14587);
xnor U15496 (N_15496,N_14905,N_14433);
nor U15497 (N_15497,N_14710,N_14476);
xnor U15498 (N_15498,N_14994,N_14837);
and U15499 (N_15499,N_14681,N_14417);
nor U15500 (N_15500,N_14773,N_14708);
nor U15501 (N_15501,N_14426,N_14696);
xnor U15502 (N_15502,N_14556,N_14515);
and U15503 (N_15503,N_14833,N_14513);
or U15504 (N_15504,N_14442,N_14800);
or U15505 (N_15505,N_14872,N_14803);
nand U15506 (N_15506,N_14836,N_14871);
xnor U15507 (N_15507,N_14968,N_14572);
xor U15508 (N_15508,N_14959,N_14919);
or U15509 (N_15509,N_14819,N_14934);
xnor U15510 (N_15510,N_14694,N_14760);
or U15511 (N_15511,N_14766,N_14841);
or U15512 (N_15512,N_14462,N_14862);
nand U15513 (N_15513,N_14741,N_14443);
xor U15514 (N_15514,N_14667,N_14436);
nand U15515 (N_15515,N_14710,N_14594);
or U15516 (N_15516,N_14580,N_14869);
nor U15517 (N_15517,N_14475,N_14581);
nand U15518 (N_15518,N_14699,N_14666);
nand U15519 (N_15519,N_14801,N_14505);
nand U15520 (N_15520,N_14849,N_14418);
nand U15521 (N_15521,N_14654,N_14878);
or U15522 (N_15522,N_14910,N_14601);
nand U15523 (N_15523,N_14649,N_14599);
nand U15524 (N_15524,N_14759,N_14547);
xnor U15525 (N_15525,N_14579,N_14926);
nand U15526 (N_15526,N_14600,N_14692);
xnor U15527 (N_15527,N_14722,N_14772);
xor U15528 (N_15528,N_14882,N_14730);
nand U15529 (N_15529,N_14604,N_14765);
and U15530 (N_15530,N_14563,N_14687);
nand U15531 (N_15531,N_14450,N_14640);
nand U15532 (N_15532,N_14920,N_14494);
nand U15533 (N_15533,N_14579,N_14558);
and U15534 (N_15534,N_14601,N_14436);
nor U15535 (N_15535,N_14982,N_14484);
nand U15536 (N_15536,N_14761,N_14979);
and U15537 (N_15537,N_14652,N_14718);
or U15538 (N_15538,N_14670,N_14531);
and U15539 (N_15539,N_14727,N_14599);
nand U15540 (N_15540,N_14493,N_14670);
nor U15541 (N_15541,N_14934,N_14951);
xor U15542 (N_15542,N_14529,N_14831);
or U15543 (N_15543,N_14900,N_14776);
or U15544 (N_15544,N_14662,N_14968);
or U15545 (N_15545,N_14779,N_14704);
xnor U15546 (N_15546,N_14561,N_14838);
or U15547 (N_15547,N_14580,N_14609);
xor U15548 (N_15548,N_14826,N_14908);
nand U15549 (N_15549,N_14892,N_14490);
nand U15550 (N_15550,N_14571,N_14693);
and U15551 (N_15551,N_14737,N_14731);
nand U15552 (N_15552,N_14500,N_14960);
nor U15553 (N_15553,N_14535,N_14947);
nand U15554 (N_15554,N_14538,N_14702);
xnor U15555 (N_15555,N_14414,N_14865);
and U15556 (N_15556,N_14851,N_14508);
nand U15557 (N_15557,N_14657,N_14589);
nor U15558 (N_15558,N_14460,N_14495);
and U15559 (N_15559,N_14620,N_14553);
nand U15560 (N_15560,N_14460,N_14627);
nor U15561 (N_15561,N_14874,N_14724);
and U15562 (N_15562,N_14511,N_14553);
and U15563 (N_15563,N_14496,N_14552);
and U15564 (N_15564,N_14911,N_14712);
or U15565 (N_15565,N_14720,N_14565);
and U15566 (N_15566,N_14625,N_14859);
and U15567 (N_15567,N_14454,N_14866);
xnor U15568 (N_15568,N_14510,N_14639);
nand U15569 (N_15569,N_14518,N_14687);
nand U15570 (N_15570,N_14421,N_14707);
xor U15571 (N_15571,N_14791,N_14858);
nand U15572 (N_15572,N_14705,N_14477);
xor U15573 (N_15573,N_14515,N_14735);
xnor U15574 (N_15574,N_14446,N_14453);
nor U15575 (N_15575,N_14409,N_14716);
nand U15576 (N_15576,N_14816,N_14921);
nor U15577 (N_15577,N_14405,N_14609);
xor U15578 (N_15578,N_14742,N_14566);
or U15579 (N_15579,N_14550,N_14916);
nand U15580 (N_15580,N_14653,N_14775);
or U15581 (N_15581,N_14798,N_14777);
nand U15582 (N_15582,N_14481,N_14648);
nand U15583 (N_15583,N_14427,N_14846);
nor U15584 (N_15584,N_14497,N_14562);
xor U15585 (N_15585,N_14953,N_14538);
xnor U15586 (N_15586,N_14769,N_14539);
or U15587 (N_15587,N_14940,N_14495);
and U15588 (N_15588,N_14692,N_14533);
and U15589 (N_15589,N_14768,N_14741);
xnor U15590 (N_15590,N_14837,N_14534);
or U15591 (N_15591,N_14416,N_14613);
xor U15592 (N_15592,N_14968,N_14659);
nor U15593 (N_15593,N_14856,N_14803);
or U15594 (N_15594,N_14510,N_14505);
and U15595 (N_15595,N_14481,N_14602);
nor U15596 (N_15596,N_14560,N_14914);
and U15597 (N_15597,N_14416,N_14560);
and U15598 (N_15598,N_14641,N_14691);
nor U15599 (N_15599,N_14691,N_14501);
xor U15600 (N_15600,N_15373,N_15245);
or U15601 (N_15601,N_15504,N_15114);
or U15602 (N_15602,N_15186,N_15367);
nor U15603 (N_15603,N_15382,N_15041);
and U15604 (N_15604,N_15117,N_15001);
xor U15605 (N_15605,N_15031,N_15210);
nand U15606 (N_15606,N_15073,N_15309);
or U15607 (N_15607,N_15107,N_15527);
and U15608 (N_15608,N_15583,N_15328);
nand U15609 (N_15609,N_15493,N_15028);
nand U15610 (N_15610,N_15501,N_15012);
and U15611 (N_15611,N_15195,N_15505);
nor U15612 (N_15612,N_15259,N_15495);
xor U15613 (N_15613,N_15329,N_15469);
xnor U15614 (N_15614,N_15580,N_15099);
or U15615 (N_15615,N_15377,N_15154);
xor U15616 (N_15616,N_15130,N_15502);
and U15617 (N_15617,N_15353,N_15238);
and U15618 (N_15618,N_15576,N_15018);
or U15619 (N_15619,N_15349,N_15554);
or U15620 (N_15620,N_15277,N_15463);
nor U15621 (N_15621,N_15410,N_15038);
or U15622 (N_15622,N_15011,N_15293);
xor U15623 (N_15623,N_15287,N_15026);
nor U15624 (N_15624,N_15413,N_15345);
nand U15625 (N_15625,N_15000,N_15218);
nand U15626 (N_15626,N_15100,N_15437);
nor U15627 (N_15627,N_15153,N_15521);
or U15628 (N_15628,N_15076,N_15584);
or U15629 (N_15629,N_15161,N_15404);
xnor U15630 (N_15630,N_15301,N_15569);
nor U15631 (N_15631,N_15457,N_15202);
nor U15632 (N_15632,N_15201,N_15477);
nor U15633 (N_15633,N_15407,N_15281);
nand U15634 (N_15634,N_15533,N_15282);
nand U15635 (N_15635,N_15178,N_15222);
or U15636 (N_15636,N_15507,N_15403);
or U15637 (N_15637,N_15299,N_15400);
nand U15638 (N_15638,N_15391,N_15479);
and U15639 (N_15639,N_15070,N_15555);
and U15640 (N_15640,N_15461,N_15175);
nand U15641 (N_15641,N_15360,N_15589);
and U15642 (N_15642,N_15416,N_15185);
nor U15643 (N_15643,N_15080,N_15354);
nor U15644 (N_15644,N_15344,N_15020);
xnor U15645 (N_15645,N_15266,N_15489);
xnor U15646 (N_15646,N_15155,N_15448);
or U15647 (N_15647,N_15386,N_15246);
nor U15648 (N_15648,N_15103,N_15213);
or U15649 (N_15649,N_15503,N_15194);
nand U15650 (N_15650,N_15231,N_15468);
nand U15651 (N_15651,N_15430,N_15578);
nor U15652 (N_15652,N_15491,N_15499);
nor U15653 (N_15653,N_15241,N_15455);
and U15654 (N_15654,N_15279,N_15421);
and U15655 (N_15655,N_15159,N_15376);
and U15656 (N_15656,N_15559,N_15192);
nor U15657 (N_15657,N_15226,N_15497);
nor U15658 (N_15658,N_15478,N_15362);
nor U15659 (N_15659,N_15333,N_15494);
nor U15660 (N_15660,N_15306,N_15253);
xor U15661 (N_15661,N_15136,N_15532);
and U15662 (N_15662,N_15326,N_15229);
and U15663 (N_15663,N_15267,N_15243);
xnor U15664 (N_15664,N_15264,N_15086);
or U15665 (N_15665,N_15581,N_15121);
nor U15666 (N_15666,N_15288,N_15567);
nand U15667 (N_15667,N_15037,N_15445);
or U15668 (N_15668,N_15208,N_15393);
nor U15669 (N_15669,N_15337,N_15044);
xor U15670 (N_15670,N_15340,N_15364);
or U15671 (N_15671,N_15061,N_15321);
nand U15672 (N_15672,N_15387,N_15128);
and U15673 (N_15673,N_15204,N_15090);
or U15674 (N_15674,N_15351,N_15460);
nor U15675 (N_15675,N_15055,N_15392);
xor U15676 (N_15676,N_15420,N_15550);
or U15677 (N_15677,N_15357,N_15372);
and U15678 (N_15678,N_15487,N_15034);
or U15679 (N_15679,N_15177,N_15052);
or U15680 (N_15680,N_15275,N_15546);
xnor U15681 (N_15681,N_15004,N_15169);
xnor U15682 (N_15682,N_15059,N_15582);
nor U15683 (N_15683,N_15015,N_15315);
and U15684 (N_15684,N_15079,N_15203);
or U15685 (N_15685,N_15456,N_15484);
nor U15686 (N_15686,N_15378,N_15474);
and U15687 (N_15687,N_15470,N_15170);
nand U15688 (N_15688,N_15379,N_15027);
nor U15689 (N_15689,N_15295,N_15098);
nor U15690 (N_15690,N_15042,N_15007);
and U15691 (N_15691,N_15311,N_15429);
or U15692 (N_15692,N_15514,N_15389);
or U15693 (N_15693,N_15247,N_15571);
nor U15694 (N_15694,N_15078,N_15054);
or U15695 (N_15695,N_15316,N_15046);
nor U15696 (N_15696,N_15261,N_15257);
or U15697 (N_15697,N_15511,N_15111);
and U15698 (N_15698,N_15248,N_15085);
nor U15699 (N_15699,N_15492,N_15465);
or U15700 (N_15700,N_15473,N_15355);
and U15701 (N_15701,N_15163,N_15347);
and U15702 (N_15702,N_15188,N_15242);
nand U15703 (N_15703,N_15566,N_15062);
nor U15704 (N_15704,N_15588,N_15081);
nand U15705 (N_15705,N_15417,N_15214);
xnor U15706 (N_15706,N_15043,N_15384);
nand U15707 (N_15707,N_15069,N_15152);
nor U15708 (N_15708,N_15124,N_15398);
or U15709 (N_15709,N_15008,N_15356);
or U15710 (N_15710,N_15297,N_15166);
or U15711 (N_15711,N_15298,N_15412);
xor U15712 (N_15712,N_15149,N_15439);
nand U15713 (N_15713,N_15165,N_15358);
nand U15714 (N_15714,N_15370,N_15276);
or U15715 (N_15715,N_15476,N_15325);
and U15716 (N_15716,N_15342,N_15181);
nand U15717 (N_15717,N_15255,N_15262);
and U15718 (N_15718,N_15586,N_15334);
nor U15719 (N_15719,N_15211,N_15449);
nor U15720 (N_15720,N_15048,N_15339);
and U15721 (N_15721,N_15017,N_15096);
nor U15722 (N_15722,N_15313,N_15215);
nor U15723 (N_15723,N_15365,N_15411);
or U15724 (N_15724,N_15074,N_15164);
or U15725 (N_15725,N_15225,N_15535);
nor U15726 (N_15726,N_15462,N_15406);
or U15727 (N_15727,N_15481,N_15453);
and U15728 (N_15728,N_15397,N_15068);
and U15729 (N_15729,N_15140,N_15516);
nor U15730 (N_15730,N_15010,N_15539);
and U15731 (N_15731,N_15158,N_15452);
xnor U15732 (N_15732,N_15088,N_15097);
nand U15733 (N_15733,N_15102,N_15402);
nand U15734 (N_15734,N_15363,N_15033);
and U15735 (N_15735,N_15475,N_15396);
nand U15736 (N_15736,N_15022,N_15019);
nand U15737 (N_15737,N_15120,N_15568);
or U15738 (N_15738,N_15436,N_15331);
or U15739 (N_15739,N_15087,N_15224);
nor U15740 (N_15740,N_15065,N_15597);
or U15741 (N_15741,N_15598,N_15144);
or U15742 (N_15742,N_15595,N_15016);
nand U15743 (N_15743,N_15346,N_15250);
nor U15744 (N_15744,N_15036,N_15390);
nand U15745 (N_15745,N_15109,N_15480);
xnor U15746 (N_15746,N_15302,N_15138);
xnor U15747 (N_15747,N_15083,N_15459);
or U15748 (N_15748,N_15296,N_15156);
nor U15749 (N_15749,N_15260,N_15488);
xnor U15750 (N_15750,N_15536,N_15269);
and U15751 (N_15751,N_15119,N_15335);
xor U15752 (N_15752,N_15599,N_15442);
xnor U15753 (N_15753,N_15112,N_15067);
nand U15754 (N_15754,N_15160,N_15519);
or U15755 (N_15755,N_15548,N_15440);
nor U15756 (N_15756,N_15283,N_15561);
nand U15757 (N_15757,N_15558,N_15374);
nand U15758 (N_15758,N_15221,N_15075);
xnor U15759 (N_15759,N_15513,N_15205);
or U15760 (N_15760,N_15591,N_15458);
nor U15761 (N_15761,N_15104,N_15003);
nor U15762 (N_15762,N_15254,N_15196);
and U15763 (N_15763,N_15219,N_15560);
and U15764 (N_15764,N_15101,N_15147);
or U15765 (N_15765,N_15415,N_15332);
nand U15766 (N_15766,N_15388,N_15143);
nor U15767 (N_15767,N_15471,N_15451);
xor U15768 (N_15768,N_15094,N_15431);
nor U15769 (N_15769,N_15496,N_15021);
nor U15770 (N_15770,N_15320,N_15146);
and U15771 (N_15771,N_15425,N_15577);
or U15772 (N_15772,N_15263,N_15162);
nor U15773 (N_15773,N_15444,N_15438);
or U15774 (N_15774,N_15545,N_15005);
and U15775 (N_15775,N_15184,N_15115);
nand U15776 (N_15776,N_15307,N_15009);
or U15777 (N_15777,N_15542,N_15234);
and U15778 (N_15778,N_15095,N_15148);
nor U15779 (N_15779,N_15056,N_15557);
xnor U15780 (N_15780,N_15082,N_15023);
nor U15781 (N_15781,N_15529,N_15441);
nand U15782 (N_15782,N_15176,N_15314);
xnor U15783 (N_15783,N_15432,N_15030);
or U15784 (N_15784,N_15270,N_15284);
or U15785 (N_15785,N_15552,N_15273);
xor U15786 (N_15786,N_15381,N_15366);
or U15787 (N_15787,N_15024,N_15408);
xnor U15788 (N_15788,N_15330,N_15537);
nand U15789 (N_15789,N_15280,N_15585);
nor U15790 (N_15790,N_15151,N_15050);
nand U15791 (N_15791,N_15522,N_15256);
nor U15792 (N_15792,N_15385,N_15294);
and U15793 (N_15793,N_15077,N_15394);
nor U15794 (N_15794,N_15063,N_15271);
or U15795 (N_15795,N_15350,N_15167);
nand U15796 (N_15796,N_15401,N_15443);
nor U15797 (N_15797,N_15524,N_15498);
nand U15798 (N_15798,N_15187,N_15590);
or U15799 (N_15799,N_15551,N_15324);
xor U15800 (N_15800,N_15127,N_15405);
nor U15801 (N_15801,N_15543,N_15272);
or U15802 (N_15802,N_15232,N_15002);
nor U15803 (N_15803,N_15359,N_15252);
and U15804 (N_15804,N_15399,N_15040);
nor U15805 (N_15805,N_15216,N_15528);
and U15806 (N_15806,N_15422,N_15454);
nor U15807 (N_15807,N_15236,N_15517);
nor U15808 (N_15808,N_15512,N_15191);
nand U15809 (N_15809,N_15508,N_15258);
nand U15810 (N_15810,N_15180,N_15510);
or U15811 (N_15811,N_15369,N_15039);
xor U15812 (N_15812,N_15206,N_15025);
and U15813 (N_15813,N_15239,N_15064);
xnor U15814 (N_15814,N_15538,N_15013);
or U15815 (N_15815,N_15466,N_15172);
nor U15816 (N_15816,N_15228,N_15426);
nor U15817 (N_15817,N_15053,N_15189);
nand U15818 (N_15818,N_15290,N_15500);
xnor U15819 (N_15819,N_15531,N_15193);
nand U15820 (N_15820,N_15348,N_15447);
and U15821 (N_15821,N_15428,N_15251);
xnor U15822 (N_15822,N_15419,N_15534);
nor U15823 (N_15823,N_15223,N_15486);
nor U15824 (N_15824,N_15091,N_15318);
nor U15825 (N_15825,N_15361,N_15207);
nand U15826 (N_15826,N_15515,N_15057);
and U15827 (N_15827,N_15553,N_15574);
nor U15828 (N_15828,N_15066,N_15530);
nor U15829 (N_15829,N_15544,N_15292);
and U15830 (N_15830,N_15141,N_15506);
and U15831 (N_15831,N_15198,N_15485);
xor U15832 (N_15832,N_15424,N_15300);
nand U15833 (N_15833,N_15423,N_15142);
or U15834 (N_15834,N_15520,N_15157);
xor U15835 (N_15835,N_15047,N_15129);
nor U15836 (N_15836,N_15244,N_15118);
nand U15837 (N_15837,N_15304,N_15174);
nand U15838 (N_15838,N_15132,N_15274);
xnor U15839 (N_15839,N_15596,N_15383);
nor U15840 (N_15840,N_15472,N_15490);
nor U15841 (N_15841,N_15072,N_15014);
and U15842 (N_15842,N_15540,N_15467);
nor U15843 (N_15843,N_15035,N_15525);
nand U15844 (N_15844,N_15352,N_15323);
nor U15845 (N_15845,N_15139,N_15123);
nand U15846 (N_15846,N_15171,N_15409);
or U15847 (N_15847,N_15278,N_15368);
xnor U15848 (N_15848,N_15317,N_15071);
nand U15849 (N_15849,N_15575,N_15045);
or U15850 (N_15850,N_15249,N_15547);
or U15851 (N_15851,N_15371,N_15434);
nor U15852 (N_15852,N_15549,N_15464);
nor U15853 (N_15853,N_15594,N_15145);
or U15854 (N_15854,N_15006,N_15116);
nor U15855 (N_15855,N_15110,N_15564);
and U15856 (N_15856,N_15183,N_15433);
nor U15857 (N_15857,N_15197,N_15220);
and U15858 (N_15858,N_15572,N_15322);
and U15859 (N_15859,N_15032,N_15418);
xor U15860 (N_15860,N_15592,N_15212);
nand U15861 (N_15861,N_15049,N_15341);
and U15862 (N_15862,N_15509,N_15150);
nor U15863 (N_15863,N_15084,N_15587);
nor U15864 (N_15864,N_15113,N_15310);
or U15865 (N_15865,N_15200,N_15105);
nand U15866 (N_15866,N_15414,N_15336);
nor U15867 (N_15867,N_15308,N_15237);
xnor U15868 (N_15868,N_15523,N_15126);
xnor U15869 (N_15869,N_15217,N_15285);
nor U15870 (N_15870,N_15092,N_15199);
nor U15871 (N_15871,N_15168,N_15518);
and U15872 (N_15872,N_15179,N_15375);
nor U15873 (N_15873,N_15427,N_15209);
nand U15874 (N_15874,N_15343,N_15122);
and U15875 (N_15875,N_15089,N_15319);
or U15876 (N_15876,N_15380,N_15338);
or U15877 (N_15877,N_15182,N_15579);
or U15878 (N_15878,N_15227,N_15573);
nand U15879 (N_15879,N_15446,N_15305);
or U15880 (N_15880,N_15565,N_15137);
or U15881 (N_15881,N_15286,N_15173);
nor U15882 (N_15882,N_15303,N_15395);
nor U15883 (N_15883,N_15051,N_15265);
and U15884 (N_15884,N_15483,N_15060);
nand U15885 (N_15885,N_15450,N_15106);
and U15886 (N_15886,N_15131,N_15230);
nor U15887 (N_15887,N_15108,N_15327);
xnor U15888 (N_15888,N_15093,N_15268);
and U15889 (N_15889,N_15563,N_15190);
xnor U15890 (N_15890,N_15482,N_15235);
nor U15891 (N_15891,N_15289,N_15058);
nor U15892 (N_15892,N_15240,N_15134);
and U15893 (N_15893,N_15593,N_15435);
xor U15894 (N_15894,N_15135,N_15526);
and U15895 (N_15895,N_15312,N_15233);
or U15896 (N_15896,N_15029,N_15291);
or U15897 (N_15897,N_15570,N_15133);
xnor U15898 (N_15898,N_15541,N_15125);
nand U15899 (N_15899,N_15556,N_15562);
xor U15900 (N_15900,N_15231,N_15376);
nand U15901 (N_15901,N_15507,N_15130);
nand U15902 (N_15902,N_15055,N_15423);
and U15903 (N_15903,N_15214,N_15150);
nor U15904 (N_15904,N_15509,N_15478);
or U15905 (N_15905,N_15373,N_15191);
xnor U15906 (N_15906,N_15507,N_15122);
xor U15907 (N_15907,N_15445,N_15291);
nand U15908 (N_15908,N_15326,N_15268);
and U15909 (N_15909,N_15407,N_15321);
nor U15910 (N_15910,N_15567,N_15211);
and U15911 (N_15911,N_15057,N_15282);
nand U15912 (N_15912,N_15400,N_15518);
nand U15913 (N_15913,N_15219,N_15404);
nand U15914 (N_15914,N_15199,N_15573);
nor U15915 (N_15915,N_15244,N_15025);
and U15916 (N_15916,N_15220,N_15511);
nor U15917 (N_15917,N_15210,N_15118);
nand U15918 (N_15918,N_15272,N_15570);
or U15919 (N_15919,N_15454,N_15212);
or U15920 (N_15920,N_15304,N_15128);
or U15921 (N_15921,N_15225,N_15392);
or U15922 (N_15922,N_15451,N_15412);
xnor U15923 (N_15923,N_15105,N_15318);
nand U15924 (N_15924,N_15247,N_15082);
or U15925 (N_15925,N_15452,N_15583);
nand U15926 (N_15926,N_15130,N_15324);
xnor U15927 (N_15927,N_15055,N_15040);
nor U15928 (N_15928,N_15464,N_15195);
and U15929 (N_15929,N_15567,N_15176);
nor U15930 (N_15930,N_15160,N_15222);
nand U15931 (N_15931,N_15152,N_15416);
xnor U15932 (N_15932,N_15500,N_15598);
xor U15933 (N_15933,N_15531,N_15462);
nor U15934 (N_15934,N_15520,N_15120);
or U15935 (N_15935,N_15461,N_15418);
and U15936 (N_15936,N_15301,N_15208);
nand U15937 (N_15937,N_15274,N_15213);
and U15938 (N_15938,N_15580,N_15593);
xor U15939 (N_15939,N_15010,N_15494);
and U15940 (N_15940,N_15402,N_15412);
and U15941 (N_15941,N_15432,N_15525);
nand U15942 (N_15942,N_15567,N_15144);
nor U15943 (N_15943,N_15428,N_15009);
nand U15944 (N_15944,N_15119,N_15548);
or U15945 (N_15945,N_15200,N_15237);
nand U15946 (N_15946,N_15297,N_15305);
xnor U15947 (N_15947,N_15501,N_15529);
and U15948 (N_15948,N_15374,N_15132);
xor U15949 (N_15949,N_15495,N_15552);
xnor U15950 (N_15950,N_15311,N_15158);
or U15951 (N_15951,N_15381,N_15044);
xor U15952 (N_15952,N_15186,N_15433);
nor U15953 (N_15953,N_15309,N_15335);
nand U15954 (N_15954,N_15100,N_15011);
or U15955 (N_15955,N_15262,N_15399);
or U15956 (N_15956,N_15570,N_15275);
xnor U15957 (N_15957,N_15118,N_15011);
or U15958 (N_15958,N_15283,N_15051);
nor U15959 (N_15959,N_15352,N_15595);
xnor U15960 (N_15960,N_15467,N_15361);
or U15961 (N_15961,N_15093,N_15388);
or U15962 (N_15962,N_15423,N_15013);
nor U15963 (N_15963,N_15129,N_15094);
or U15964 (N_15964,N_15534,N_15167);
and U15965 (N_15965,N_15242,N_15278);
xnor U15966 (N_15966,N_15234,N_15307);
nor U15967 (N_15967,N_15153,N_15598);
and U15968 (N_15968,N_15442,N_15388);
xnor U15969 (N_15969,N_15441,N_15016);
nor U15970 (N_15970,N_15223,N_15405);
nand U15971 (N_15971,N_15014,N_15442);
nand U15972 (N_15972,N_15325,N_15253);
xor U15973 (N_15973,N_15236,N_15417);
and U15974 (N_15974,N_15276,N_15250);
nor U15975 (N_15975,N_15218,N_15508);
xnor U15976 (N_15976,N_15496,N_15549);
or U15977 (N_15977,N_15328,N_15280);
and U15978 (N_15978,N_15583,N_15193);
xnor U15979 (N_15979,N_15592,N_15074);
or U15980 (N_15980,N_15406,N_15582);
nand U15981 (N_15981,N_15307,N_15070);
and U15982 (N_15982,N_15550,N_15412);
or U15983 (N_15983,N_15322,N_15038);
and U15984 (N_15984,N_15326,N_15578);
nor U15985 (N_15985,N_15081,N_15255);
xor U15986 (N_15986,N_15589,N_15524);
nor U15987 (N_15987,N_15386,N_15464);
xnor U15988 (N_15988,N_15109,N_15151);
xor U15989 (N_15989,N_15243,N_15599);
and U15990 (N_15990,N_15594,N_15475);
and U15991 (N_15991,N_15343,N_15210);
nand U15992 (N_15992,N_15135,N_15321);
and U15993 (N_15993,N_15511,N_15035);
nor U15994 (N_15994,N_15365,N_15262);
and U15995 (N_15995,N_15412,N_15256);
nand U15996 (N_15996,N_15468,N_15076);
nor U15997 (N_15997,N_15069,N_15387);
xnor U15998 (N_15998,N_15431,N_15010);
nand U15999 (N_15999,N_15044,N_15248);
and U16000 (N_16000,N_15203,N_15177);
and U16001 (N_16001,N_15138,N_15409);
nand U16002 (N_16002,N_15157,N_15159);
or U16003 (N_16003,N_15313,N_15237);
or U16004 (N_16004,N_15388,N_15001);
nor U16005 (N_16005,N_15050,N_15354);
nand U16006 (N_16006,N_15001,N_15142);
nor U16007 (N_16007,N_15568,N_15301);
nor U16008 (N_16008,N_15529,N_15123);
nand U16009 (N_16009,N_15294,N_15280);
nand U16010 (N_16010,N_15552,N_15047);
and U16011 (N_16011,N_15228,N_15597);
nand U16012 (N_16012,N_15083,N_15105);
nand U16013 (N_16013,N_15494,N_15577);
nand U16014 (N_16014,N_15194,N_15567);
and U16015 (N_16015,N_15102,N_15080);
nor U16016 (N_16016,N_15331,N_15283);
and U16017 (N_16017,N_15281,N_15218);
nand U16018 (N_16018,N_15533,N_15318);
xor U16019 (N_16019,N_15292,N_15526);
and U16020 (N_16020,N_15550,N_15439);
nor U16021 (N_16021,N_15393,N_15437);
or U16022 (N_16022,N_15424,N_15445);
and U16023 (N_16023,N_15266,N_15479);
nor U16024 (N_16024,N_15467,N_15016);
nand U16025 (N_16025,N_15493,N_15387);
xor U16026 (N_16026,N_15494,N_15493);
xor U16027 (N_16027,N_15138,N_15234);
and U16028 (N_16028,N_15341,N_15185);
and U16029 (N_16029,N_15514,N_15003);
or U16030 (N_16030,N_15519,N_15223);
nor U16031 (N_16031,N_15362,N_15003);
and U16032 (N_16032,N_15051,N_15348);
nor U16033 (N_16033,N_15241,N_15227);
and U16034 (N_16034,N_15528,N_15119);
xor U16035 (N_16035,N_15249,N_15011);
nor U16036 (N_16036,N_15207,N_15405);
or U16037 (N_16037,N_15071,N_15440);
nand U16038 (N_16038,N_15289,N_15542);
nor U16039 (N_16039,N_15415,N_15197);
and U16040 (N_16040,N_15328,N_15040);
xnor U16041 (N_16041,N_15480,N_15186);
xor U16042 (N_16042,N_15011,N_15000);
nor U16043 (N_16043,N_15120,N_15084);
nor U16044 (N_16044,N_15259,N_15315);
nor U16045 (N_16045,N_15261,N_15069);
nand U16046 (N_16046,N_15345,N_15414);
xnor U16047 (N_16047,N_15397,N_15526);
or U16048 (N_16048,N_15201,N_15480);
xor U16049 (N_16049,N_15157,N_15582);
or U16050 (N_16050,N_15112,N_15117);
nor U16051 (N_16051,N_15273,N_15152);
xor U16052 (N_16052,N_15191,N_15358);
nor U16053 (N_16053,N_15364,N_15523);
nand U16054 (N_16054,N_15255,N_15235);
nand U16055 (N_16055,N_15015,N_15270);
nand U16056 (N_16056,N_15064,N_15408);
nor U16057 (N_16057,N_15543,N_15148);
nand U16058 (N_16058,N_15549,N_15095);
or U16059 (N_16059,N_15399,N_15278);
xnor U16060 (N_16060,N_15447,N_15021);
nand U16061 (N_16061,N_15087,N_15557);
nor U16062 (N_16062,N_15356,N_15084);
and U16063 (N_16063,N_15301,N_15250);
or U16064 (N_16064,N_15277,N_15514);
nand U16065 (N_16065,N_15038,N_15356);
and U16066 (N_16066,N_15576,N_15313);
nor U16067 (N_16067,N_15065,N_15014);
or U16068 (N_16068,N_15434,N_15486);
or U16069 (N_16069,N_15073,N_15173);
and U16070 (N_16070,N_15320,N_15517);
or U16071 (N_16071,N_15005,N_15580);
or U16072 (N_16072,N_15420,N_15430);
or U16073 (N_16073,N_15472,N_15536);
xor U16074 (N_16074,N_15506,N_15257);
nand U16075 (N_16075,N_15347,N_15517);
nand U16076 (N_16076,N_15464,N_15239);
xnor U16077 (N_16077,N_15323,N_15250);
xnor U16078 (N_16078,N_15352,N_15018);
and U16079 (N_16079,N_15550,N_15311);
nand U16080 (N_16080,N_15414,N_15025);
or U16081 (N_16081,N_15332,N_15038);
xnor U16082 (N_16082,N_15056,N_15143);
nor U16083 (N_16083,N_15096,N_15015);
and U16084 (N_16084,N_15492,N_15366);
nand U16085 (N_16085,N_15096,N_15191);
xor U16086 (N_16086,N_15214,N_15318);
nand U16087 (N_16087,N_15359,N_15429);
nand U16088 (N_16088,N_15523,N_15268);
xnor U16089 (N_16089,N_15141,N_15136);
or U16090 (N_16090,N_15347,N_15390);
xnor U16091 (N_16091,N_15435,N_15348);
xor U16092 (N_16092,N_15023,N_15370);
or U16093 (N_16093,N_15181,N_15320);
or U16094 (N_16094,N_15419,N_15553);
or U16095 (N_16095,N_15567,N_15135);
and U16096 (N_16096,N_15362,N_15309);
xor U16097 (N_16097,N_15208,N_15514);
nor U16098 (N_16098,N_15498,N_15000);
nor U16099 (N_16099,N_15149,N_15197);
nand U16100 (N_16100,N_15583,N_15543);
or U16101 (N_16101,N_15379,N_15139);
xor U16102 (N_16102,N_15374,N_15340);
xnor U16103 (N_16103,N_15079,N_15201);
or U16104 (N_16104,N_15049,N_15303);
and U16105 (N_16105,N_15436,N_15146);
nand U16106 (N_16106,N_15211,N_15053);
nand U16107 (N_16107,N_15232,N_15436);
nor U16108 (N_16108,N_15288,N_15107);
nor U16109 (N_16109,N_15371,N_15455);
nor U16110 (N_16110,N_15417,N_15524);
or U16111 (N_16111,N_15096,N_15120);
and U16112 (N_16112,N_15442,N_15217);
or U16113 (N_16113,N_15506,N_15528);
xor U16114 (N_16114,N_15529,N_15207);
or U16115 (N_16115,N_15221,N_15386);
nor U16116 (N_16116,N_15281,N_15369);
nor U16117 (N_16117,N_15445,N_15113);
nand U16118 (N_16118,N_15029,N_15580);
and U16119 (N_16119,N_15364,N_15013);
xor U16120 (N_16120,N_15437,N_15250);
or U16121 (N_16121,N_15434,N_15088);
xnor U16122 (N_16122,N_15317,N_15307);
and U16123 (N_16123,N_15162,N_15270);
nand U16124 (N_16124,N_15284,N_15400);
and U16125 (N_16125,N_15524,N_15057);
xnor U16126 (N_16126,N_15015,N_15488);
nand U16127 (N_16127,N_15492,N_15183);
nand U16128 (N_16128,N_15259,N_15083);
xor U16129 (N_16129,N_15520,N_15223);
nand U16130 (N_16130,N_15552,N_15453);
and U16131 (N_16131,N_15496,N_15403);
nor U16132 (N_16132,N_15309,N_15325);
xor U16133 (N_16133,N_15474,N_15171);
and U16134 (N_16134,N_15377,N_15599);
nor U16135 (N_16135,N_15492,N_15397);
and U16136 (N_16136,N_15357,N_15522);
nor U16137 (N_16137,N_15356,N_15289);
nor U16138 (N_16138,N_15495,N_15557);
xor U16139 (N_16139,N_15177,N_15190);
nand U16140 (N_16140,N_15295,N_15122);
nor U16141 (N_16141,N_15574,N_15036);
nor U16142 (N_16142,N_15091,N_15378);
xnor U16143 (N_16143,N_15244,N_15357);
nand U16144 (N_16144,N_15339,N_15118);
nor U16145 (N_16145,N_15164,N_15103);
nor U16146 (N_16146,N_15458,N_15445);
or U16147 (N_16147,N_15418,N_15437);
or U16148 (N_16148,N_15209,N_15289);
and U16149 (N_16149,N_15549,N_15120);
nand U16150 (N_16150,N_15439,N_15389);
nor U16151 (N_16151,N_15520,N_15043);
nor U16152 (N_16152,N_15439,N_15507);
xnor U16153 (N_16153,N_15084,N_15377);
nand U16154 (N_16154,N_15231,N_15596);
and U16155 (N_16155,N_15295,N_15512);
or U16156 (N_16156,N_15240,N_15052);
or U16157 (N_16157,N_15409,N_15436);
or U16158 (N_16158,N_15567,N_15438);
nand U16159 (N_16159,N_15230,N_15478);
nand U16160 (N_16160,N_15523,N_15171);
or U16161 (N_16161,N_15446,N_15343);
nand U16162 (N_16162,N_15467,N_15512);
xor U16163 (N_16163,N_15518,N_15399);
xor U16164 (N_16164,N_15222,N_15022);
or U16165 (N_16165,N_15480,N_15494);
nor U16166 (N_16166,N_15013,N_15496);
or U16167 (N_16167,N_15528,N_15369);
nand U16168 (N_16168,N_15503,N_15053);
or U16169 (N_16169,N_15227,N_15372);
xnor U16170 (N_16170,N_15117,N_15553);
nor U16171 (N_16171,N_15519,N_15516);
xnor U16172 (N_16172,N_15016,N_15288);
nand U16173 (N_16173,N_15285,N_15392);
and U16174 (N_16174,N_15529,N_15312);
or U16175 (N_16175,N_15486,N_15290);
or U16176 (N_16176,N_15209,N_15101);
xnor U16177 (N_16177,N_15062,N_15408);
nor U16178 (N_16178,N_15053,N_15102);
xor U16179 (N_16179,N_15252,N_15121);
nand U16180 (N_16180,N_15288,N_15020);
and U16181 (N_16181,N_15502,N_15110);
nor U16182 (N_16182,N_15374,N_15309);
nand U16183 (N_16183,N_15002,N_15268);
or U16184 (N_16184,N_15128,N_15570);
or U16185 (N_16185,N_15333,N_15091);
and U16186 (N_16186,N_15128,N_15544);
xor U16187 (N_16187,N_15380,N_15560);
and U16188 (N_16188,N_15328,N_15005);
nor U16189 (N_16189,N_15261,N_15266);
and U16190 (N_16190,N_15447,N_15155);
and U16191 (N_16191,N_15099,N_15042);
or U16192 (N_16192,N_15204,N_15050);
and U16193 (N_16193,N_15559,N_15441);
nand U16194 (N_16194,N_15232,N_15504);
xnor U16195 (N_16195,N_15210,N_15372);
nor U16196 (N_16196,N_15579,N_15512);
and U16197 (N_16197,N_15324,N_15427);
or U16198 (N_16198,N_15265,N_15303);
nor U16199 (N_16199,N_15516,N_15286);
or U16200 (N_16200,N_16191,N_16155);
or U16201 (N_16201,N_15955,N_16090);
or U16202 (N_16202,N_15893,N_15908);
and U16203 (N_16203,N_15719,N_15660);
or U16204 (N_16204,N_15783,N_15808);
or U16205 (N_16205,N_16022,N_15643);
or U16206 (N_16206,N_15689,N_15737);
xor U16207 (N_16207,N_16016,N_15606);
xor U16208 (N_16208,N_15876,N_16054);
xor U16209 (N_16209,N_15639,N_15611);
xnor U16210 (N_16210,N_16036,N_15802);
xor U16211 (N_16211,N_16183,N_16056);
and U16212 (N_16212,N_16025,N_15868);
xor U16213 (N_16213,N_15984,N_15866);
nand U16214 (N_16214,N_16119,N_15712);
and U16215 (N_16215,N_15964,N_16188);
or U16216 (N_16216,N_16028,N_16070);
nor U16217 (N_16217,N_16175,N_15726);
nor U16218 (N_16218,N_16053,N_15976);
nand U16219 (N_16219,N_15778,N_15618);
and U16220 (N_16220,N_16082,N_15775);
nor U16221 (N_16221,N_15718,N_15785);
or U16222 (N_16222,N_15943,N_15940);
nand U16223 (N_16223,N_16150,N_15627);
nor U16224 (N_16224,N_16174,N_15659);
nand U16225 (N_16225,N_15735,N_15888);
or U16226 (N_16226,N_16026,N_15797);
nor U16227 (N_16227,N_15668,N_15721);
nand U16228 (N_16228,N_15610,N_16140);
nor U16229 (N_16229,N_15637,N_16018);
nor U16230 (N_16230,N_15736,N_15999);
xnor U16231 (N_16231,N_16072,N_15881);
and U16232 (N_16232,N_16037,N_15795);
nor U16233 (N_16233,N_16094,N_15609);
xor U16234 (N_16234,N_16158,N_15832);
xnor U16235 (N_16235,N_15862,N_16114);
xnor U16236 (N_16236,N_15741,N_16074);
xor U16237 (N_16237,N_16079,N_15951);
and U16238 (N_16238,N_15750,N_15905);
xnor U16239 (N_16239,N_16096,N_15898);
or U16240 (N_16240,N_15697,N_15926);
nand U16241 (N_16241,N_16006,N_15789);
nor U16242 (N_16242,N_15946,N_15872);
nor U16243 (N_16243,N_15681,N_16179);
nand U16244 (N_16244,N_15701,N_15693);
nor U16245 (N_16245,N_15944,N_16103);
xnor U16246 (N_16246,N_16180,N_15669);
or U16247 (N_16247,N_16194,N_16192);
or U16248 (N_16248,N_15842,N_15959);
nand U16249 (N_16249,N_16157,N_15685);
and U16250 (N_16250,N_15988,N_15720);
xnor U16251 (N_16251,N_16159,N_16167);
nor U16252 (N_16252,N_15769,N_15772);
nand U16253 (N_16253,N_16134,N_16117);
nand U16254 (N_16254,N_15875,N_16088);
xnor U16255 (N_16255,N_16101,N_15927);
or U16256 (N_16256,N_16173,N_15657);
or U16257 (N_16257,N_16198,N_16132);
nand U16258 (N_16258,N_16065,N_15755);
nor U16259 (N_16259,N_16019,N_15987);
or U16260 (N_16260,N_16017,N_15622);
and U16261 (N_16261,N_15710,N_16197);
xor U16262 (N_16262,N_16143,N_15891);
nor U16263 (N_16263,N_15828,N_15608);
and U16264 (N_16264,N_16177,N_16092);
or U16265 (N_16265,N_15889,N_15945);
nor U16266 (N_16266,N_15801,N_15645);
and U16267 (N_16267,N_16145,N_15728);
or U16268 (N_16268,N_15733,N_15909);
nor U16269 (N_16269,N_15989,N_15732);
nand U16270 (N_16270,N_16156,N_15849);
xnor U16271 (N_16271,N_15653,N_15892);
and U16272 (N_16272,N_16170,N_15825);
nor U16273 (N_16273,N_15759,N_15784);
nand U16274 (N_16274,N_15890,N_16109);
and U16275 (N_16275,N_16038,N_15754);
nor U16276 (N_16276,N_15615,N_16055);
xor U16277 (N_16277,N_16011,N_15666);
nand U16278 (N_16278,N_15855,N_16153);
or U16279 (N_16279,N_15635,N_15974);
xor U16280 (N_16280,N_15641,N_15827);
and U16281 (N_16281,N_15623,N_15993);
nor U16282 (N_16282,N_15931,N_15820);
nand U16283 (N_16283,N_16102,N_16085);
and U16284 (N_16284,N_15724,N_16000);
xor U16285 (N_16285,N_16147,N_16091);
nand U16286 (N_16286,N_16081,N_15804);
nor U16287 (N_16287,N_15674,N_15706);
nor U16288 (N_16288,N_15879,N_16146);
xor U16289 (N_16289,N_15803,N_15771);
and U16290 (N_16290,N_15647,N_16078);
nand U16291 (N_16291,N_16086,N_15970);
or U16292 (N_16292,N_15644,N_15773);
nand U16293 (N_16293,N_16136,N_16139);
or U16294 (N_16294,N_16061,N_15794);
xor U16295 (N_16295,N_16020,N_15781);
and U16296 (N_16296,N_16107,N_16189);
and U16297 (N_16297,N_16035,N_16027);
xor U16298 (N_16298,N_15762,N_15932);
nor U16299 (N_16299,N_15950,N_15824);
or U16300 (N_16300,N_15665,N_15992);
nand U16301 (N_16301,N_16033,N_16181);
nor U16302 (N_16302,N_15949,N_15843);
nand U16303 (N_16303,N_16024,N_16113);
xor U16304 (N_16304,N_15687,N_16098);
nand U16305 (N_16305,N_16112,N_15925);
nor U16306 (N_16306,N_15672,N_16031);
xnor U16307 (N_16307,N_15777,N_15679);
xnor U16308 (N_16308,N_16013,N_15760);
xor U16309 (N_16309,N_15730,N_15851);
xnor U16310 (N_16310,N_16111,N_15699);
nor U16311 (N_16311,N_15723,N_15838);
nand U16312 (N_16312,N_15956,N_15861);
or U16313 (N_16313,N_15815,N_15845);
or U16314 (N_16314,N_15698,N_15640);
nand U16315 (N_16315,N_15776,N_16076);
or U16316 (N_16316,N_15933,N_15822);
xnor U16317 (N_16317,N_15756,N_15997);
xnor U16318 (N_16318,N_15716,N_15968);
xnor U16319 (N_16319,N_15800,N_15700);
xnor U16320 (N_16320,N_15603,N_15912);
nor U16321 (N_16321,N_16195,N_16021);
nand U16322 (N_16322,N_16160,N_15979);
nor U16323 (N_16323,N_16123,N_16040);
xnor U16324 (N_16324,N_16115,N_15840);
and U16325 (N_16325,N_15768,N_16187);
nand U16326 (N_16326,N_15780,N_15821);
nand U16327 (N_16327,N_15885,N_15919);
nor U16328 (N_16328,N_15694,N_15628);
and U16329 (N_16329,N_16127,N_16046);
and U16330 (N_16330,N_15865,N_15920);
or U16331 (N_16331,N_15763,N_15652);
nand U16332 (N_16332,N_15913,N_15998);
xnor U16333 (N_16333,N_15915,N_16172);
and U16334 (N_16334,N_15629,N_16166);
and U16335 (N_16335,N_15717,N_15725);
or U16336 (N_16336,N_15853,N_15939);
nand U16337 (N_16337,N_15633,N_16138);
xor U16338 (N_16338,N_15994,N_15686);
and U16339 (N_16339,N_15811,N_15911);
xor U16340 (N_16340,N_15695,N_15727);
or U16341 (N_16341,N_15764,N_16105);
and U16342 (N_16342,N_15704,N_15617);
and U16343 (N_16343,N_16051,N_15907);
nand U16344 (N_16344,N_16135,N_15807);
and U16345 (N_16345,N_15880,N_16193);
xor U16346 (N_16346,N_15924,N_15658);
or U16347 (N_16347,N_15973,N_16168);
xor U16348 (N_16348,N_16142,N_15839);
or U16349 (N_16349,N_15857,N_15856);
or U16350 (N_16350,N_16100,N_15678);
nor U16351 (N_16351,N_15859,N_15810);
nand U16352 (N_16352,N_16152,N_15995);
xor U16353 (N_16353,N_15675,N_15982);
xor U16354 (N_16354,N_15655,N_15850);
nand U16355 (N_16355,N_15671,N_15702);
and U16356 (N_16356,N_16199,N_16064);
nand U16357 (N_16357,N_15921,N_16023);
nand U16358 (N_16358,N_15829,N_16069);
or U16359 (N_16359,N_16002,N_15864);
nor U16360 (N_16360,N_15711,N_15682);
or U16361 (N_16361,N_15767,N_15731);
and U16362 (N_16362,N_15753,N_16066);
nor U16363 (N_16363,N_15744,N_15656);
nand U16364 (N_16364,N_16151,N_15749);
or U16365 (N_16365,N_16048,N_16008);
xor U16366 (N_16366,N_16049,N_15830);
and U16367 (N_16367,N_15928,N_15673);
and U16368 (N_16368,N_15638,N_15996);
and U16369 (N_16369,N_15648,N_15743);
nand U16370 (N_16370,N_16003,N_15747);
nand U16371 (N_16371,N_15680,N_16001);
and U16372 (N_16372,N_16099,N_15796);
nor U16373 (N_16373,N_15662,N_15651);
and U16374 (N_16374,N_15751,N_15961);
nand U16375 (N_16375,N_15903,N_15869);
xnor U16376 (N_16376,N_16043,N_16154);
or U16377 (N_16377,N_16122,N_15841);
xor U16378 (N_16378,N_15978,N_15624);
xor U16379 (N_16379,N_16014,N_15863);
and U16380 (N_16380,N_16050,N_15823);
nor U16381 (N_16381,N_15936,N_15782);
and U16382 (N_16382,N_16128,N_15910);
nor U16383 (N_16383,N_15806,N_16083);
xnor U16384 (N_16384,N_15742,N_15620);
and U16385 (N_16385,N_15977,N_15844);
nand U16386 (N_16386,N_15696,N_15901);
and U16387 (N_16387,N_16149,N_16110);
or U16388 (N_16388,N_16059,N_15600);
nor U16389 (N_16389,N_15670,N_16058);
or U16390 (N_16390,N_16196,N_15900);
nor U16391 (N_16391,N_15873,N_16125);
or U16392 (N_16392,N_15605,N_15835);
and U16393 (N_16393,N_15991,N_16178);
xnor U16394 (N_16394,N_16176,N_16030);
and U16395 (N_16395,N_15965,N_15602);
or U16396 (N_16396,N_15871,N_15746);
or U16397 (N_16397,N_15621,N_15896);
nor U16398 (N_16398,N_16186,N_15981);
and U16399 (N_16399,N_15734,N_15713);
nor U16400 (N_16400,N_15636,N_15948);
nor U16401 (N_16401,N_16097,N_16068);
nor U16402 (N_16402,N_16032,N_16118);
and U16403 (N_16403,N_15817,N_15774);
nand U16404 (N_16404,N_15690,N_15707);
nor U16405 (N_16405,N_15957,N_15899);
and U16406 (N_16406,N_15798,N_15630);
or U16407 (N_16407,N_15960,N_15616);
nand U16408 (N_16408,N_16067,N_15834);
and U16409 (N_16409,N_16108,N_15715);
and U16410 (N_16410,N_15934,N_15874);
or U16411 (N_16411,N_15941,N_16087);
nand U16412 (N_16412,N_16073,N_15971);
or U16413 (N_16413,N_15870,N_15895);
nor U16414 (N_16414,N_15809,N_15626);
xor U16415 (N_16415,N_15676,N_15661);
nor U16416 (N_16416,N_16077,N_15860);
xnor U16417 (N_16417,N_15990,N_15958);
and U16418 (N_16418,N_15705,N_15632);
or U16419 (N_16419,N_15967,N_16130);
nand U16420 (N_16420,N_15917,N_15779);
nor U16421 (N_16421,N_16171,N_16137);
nor U16422 (N_16422,N_15894,N_15813);
or U16423 (N_16423,N_15877,N_16007);
nand U16424 (N_16424,N_15684,N_15601);
xnor U16425 (N_16425,N_15683,N_15692);
and U16426 (N_16426,N_15765,N_16071);
or U16427 (N_16427,N_15858,N_15848);
and U16428 (N_16428,N_15677,N_16044);
or U16429 (N_16429,N_16004,N_15837);
xnor U16430 (N_16430,N_15739,N_15897);
nor U16431 (N_16431,N_15963,N_16104);
or U16432 (N_16432,N_15852,N_16141);
or U16433 (N_16433,N_15902,N_15942);
nand U16434 (N_16434,N_15929,N_15703);
nand U16435 (N_16435,N_15788,N_15818);
or U16436 (N_16436,N_15882,N_15654);
and U16437 (N_16437,N_15787,N_15625);
nand U16438 (N_16438,N_15953,N_15972);
nor U16439 (N_16439,N_15836,N_16163);
or U16440 (N_16440,N_16165,N_15966);
nor U16441 (N_16441,N_16161,N_15790);
or U16442 (N_16442,N_16126,N_15969);
nand U16443 (N_16443,N_15793,N_15914);
nand U16444 (N_16444,N_16060,N_15833);
or U16445 (N_16445,N_16182,N_16012);
or U16446 (N_16446,N_16039,N_15740);
nand U16447 (N_16447,N_16063,N_15938);
nand U16448 (N_16448,N_16133,N_15766);
or U16449 (N_16449,N_15791,N_16129);
and U16450 (N_16450,N_15757,N_15738);
nor U16451 (N_16451,N_16089,N_15937);
nor U16452 (N_16452,N_15805,N_16075);
nor U16453 (N_16453,N_16144,N_16010);
xnor U16454 (N_16454,N_15980,N_15812);
nor U16455 (N_16455,N_15761,N_15786);
or U16456 (N_16456,N_15709,N_16190);
xnor U16457 (N_16457,N_15752,N_15814);
xnor U16458 (N_16458,N_16120,N_15799);
nand U16459 (N_16459,N_16093,N_15826);
xor U16460 (N_16460,N_15607,N_16095);
xor U16461 (N_16461,N_15819,N_16062);
or U16462 (N_16462,N_16047,N_15904);
nand U16463 (N_16463,N_16042,N_15748);
xor U16464 (N_16464,N_16080,N_15650);
or U16465 (N_16465,N_15758,N_16009);
nor U16466 (N_16466,N_15691,N_15714);
or U16467 (N_16467,N_16106,N_15985);
and U16468 (N_16468,N_15930,N_16185);
xor U16469 (N_16469,N_15884,N_16121);
and U16470 (N_16470,N_15667,N_15923);
nand U16471 (N_16471,N_15729,N_15612);
xnor U16472 (N_16472,N_16015,N_16034);
and U16473 (N_16473,N_15663,N_16057);
nor U16474 (N_16474,N_15619,N_15954);
nand U16475 (N_16475,N_16005,N_15846);
and U16476 (N_16476,N_15613,N_15631);
nor U16477 (N_16477,N_15722,N_15935);
nor U16478 (N_16478,N_15886,N_16116);
and U16479 (N_16479,N_15952,N_16184);
or U16480 (N_16480,N_15962,N_15816);
nor U16481 (N_16481,N_15878,N_15986);
or U16482 (N_16482,N_15918,N_15831);
nor U16483 (N_16483,N_16162,N_16029);
xor U16484 (N_16484,N_15745,N_15906);
or U16485 (N_16485,N_15708,N_15847);
nor U16486 (N_16486,N_15614,N_16052);
nand U16487 (N_16487,N_15916,N_16169);
nand U16488 (N_16488,N_16084,N_16045);
or U16489 (N_16489,N_15688,N_16148);
or U16490 (N_16490,N_15922,N_15883);
xor U16491 (N_16491,N_16164,N_15634);
nand U16492 (N_16492,N_16124,N_15646);
and U16493 (N_16493,N_15975,N_15887);
and U16494 (N_16494,N_15983,N_15604);
nand U16495 (N_16495,N_15770,N_15947);
or U16496 (N_16496,N_15792,N_15642);
nand U16497 (N_16497,N_15649,N_16041);
or U16498 (N_16498,N_15664,N_15867);
nand U16499 (N_16499,N_16131,N_15854);
nand U16500 (N_16500,N_15663,N_15926);
nand U16501 (N_16501,N_16110,N_16091);
nor U16502 (N_16502,N_16176,N_15995);
nand U16503 (N_16503,N_15913,N_15821);
and U16504 (N_16504,N_16160,N_16104);
nand U16505 (N_16505,N_15922,N_15988);
or U16506 (N_16506,N_15996,N_15953);
and U16507 (N_16507,N_15651,N_15910);
and U16508 (N_16508,N_15679,N_16075);
and U16509 (N_16509,N_15962,N_16057);
or U16510 (N_16510,N_15815,N_15900);
nor U16511 (N_16511,N_15625,N_15992);
xnor U16512 (N_16512,N_16011,N_16078);
xor U16513 (N_16513,N_15817,N_15989);
xor U16514 (N_16514,N_15963,N_16176);
and U16515 (N_16515,N_16073,N_15966);
nor U16516 (N_16516,N_15667,N_15848);
or U16517 (N_16517,N_16046,N_16171);
or U16518 (N_16518,N_15943,N_15776);
xor U16519 (N_16519,N_16073,N_15645);
or U16520 (N_16520,N_16154,N_16047);
nand U16521 (N_16521,N_15727,N_15701);
and U16522 (N_16522,N_15945,N_16027);
and U16523 (N_16523,N_15716,N_15988);
nor U16524 (N_16524,N_15938,N_15779);
xnor U16525 (N_16525,N_15969,N_15873);
nor U16526 (N_16526,N_15861,N_15931);
nand U16527 (N_16527,N_15686,N_16049);
or U16528 (N_16528,N_15940,N_16197);
xor U16529 (N_16529,N_15922,N_16025);
nand U16530 (N_16530,N_16066,N_15745);
or U16531 (N_16531,N_16025,N_15826);
and U16532 (N_16532,N_16130,N_15713);
nor U16533 (N_16533,N_15658,N_15715);
and U16534 (N_16534,N_16148,N_16028);
nand U16535 (N_16535,N_15720,N_16029);
nand U16536 (N_16536,N_15726,N_16150);
nand U16537 (N_16537,N_15610,N_15795);
and U16538 (N_16538,N_15923,N_15756);
and U16539 (N_16539,N_15640,N_15606);
and U16540 (N_16540,N_15736,N_16191);
nor U16541 (N_16541,N_15839,N_15603);
nor U16542 (N_16542,N_15742,N_15720);
and U16543 (N_16543,N_16064,N_15996);
nor U16544 (N_16544,N_16044,N_15791);
nand U16545 (N_16545,N_16017,N_15818);
nor U16546 (N_16546,N_15773,N_15981);
or U16547 (N_16547,N_15866,N_15601);
xnor U16548 (N_16548,N_15730,N_15841);
and U16549 (N_16549,N_16181,N_16169);
or U16550 (N_16550,N_16002,N_15718);
nand U16551 (N_16551,N_16199,N_15977);
nor U16552 (N_16552,N_15724,N_15628);
or U16553 (N_16553,N_15711,N_16101);
xor U16554 (N_16554,N_16115,N_15653);
xor U16555 (N_16555,N_16084,N_15947);
or U16556 (N_16556,N_15823,N_16170);
nor U16557 (N_16557,N_15788,N_16012);
or U16558 (N_16558,N_15890,N_16175);
or U16559 (N_16559,N_16098,N_15650);
xor U16560 (N_16560,N_16089,N_15719);
nor U16561 (N_16561,N_15636,N_15791);
and U16562 (N_16562,N_15902,N_16056);
and U16563 (N_16563,N_15607,N_15966);
xor U16564 (N_16564,N_15744,N_15737);
and U16565 (N_16565,N_15897,N_15864);
or U16566 (N_16566,N_15818,N_15704);
xor U16567 (N_16567,N_15742,N_15942);
or U16568 (N_16568,N_15732,N_15931);
xor U16569 (N_16569,N_15828,N_15735);
and U16570 (N_16570,N_15941,N_16044);
nand U16571 (N_16571,N_15761,N_15982);
nor U16572 (N_16572,N_16152,N_15666);
and U16573 (N_16573,N_16140,N_16034);
xor U16574 (N_16574,N_15855,N_15858);
nand U16575 (N_16575,N_15824,N_15851);
nand U16576 (N_16576,N_16126,N_16116);
and U16577 (N_16577,N_15605,N_15911);
or U16578 (N_16578,N_16097,N_15759);
and U16579 (N_16579,N_16125,N_15652);
or U16580 (N_16580,N_15732,N_15816);
xnor U16581 (N_16581,N_15754,N_15892);
and U16582 (N_16582,N_15909,N_16085);
xor U16583 (N_16583,N_15609,N_16122);
nor U16584 (N_16584,N_15784,N_15719);
xnor U16585 (N_16585,N_15753,N_15941);
nor U16586 (N_16586,N_15755,N_15964);
or U16587 (N_16587,N_15657,N_15802);
or U16588 (N_16588,N_15766,N_15917);
and U16589 (N_16589,N_16026,N_16096);
and U16590 (N_16590,N_16046,N_15667);
nor U16591 (N_16591,N_16128,N_15844);
nor U16592 (N_16592,N_15865,N_15862);
nor U16593 (N_16593,N_15796,N_16129);
nand U16594 (N_16594,N_15865,N_15691);
or U16595 (N_16595,N_15639,N_15720);
nand U16596 (N_16596,N_15669,N_16087);
xor U16597 (N_16597,N_15681,N_16142);
and U16598 (N_16598,N_15603,N_15919);
nor U16599 (N_16599,N_15941,N_16032);
xnor U16600 (N_16600,N_15983,N_15860);
nor U16601 (N_16601,N_15978,N_15816);
and U16602 (N_16602,N_16045,N_16100);
and U16603 (N_16603,N_15678,N_15636);
or U16604 (N_16604,N_15702,N_16055);
nor U16605 (N_16605,N_16164,N_15841);
nand U16606 (N_16606,N_15669,N_16131);
xor U16607 (N_16607,N_15935,N_15952);
nand U16608 (N_16608,N_15605,N_16057);
nand U16609 (N_16609,N_15648,N_15629);
nand U16610 (N_16610,N_15991,N_15954);
xor U16611 (N_16611,N_15970,N_15918);
or U16612 (N_16612,N_15913,N_15833);
xnor U16613 (N_16613,N_15606,N_15805);
nor U16614 (N_16614,N_16116,N_15939);
xnor U16615 (N_16615,N_16133,N_15989);
nand U16616 (N_16616,N_16080,N_15749);
nand U16617 (N_16617,N_15786,N_16157);
nand U16618 (N_16618,N_15780,N_16037);
xor U16619 (N_16619,N_15975,N_15708);
xor U16620 (N_16620,N_15768,N_16081);
xnor U16621 (N_16621,N_15780,N_15678);
and U16622 (N_16622,N_16076,N_15999);
xor U16623 (N_16623,N_16182,N_15696);
or U16624 (N_16624,N_16065,N_15720);
xor U16625 (N_16625,N_15983,N_16055);
nor U16626 (N_16626,N_16020,N_16019);
nand U16627 (N_16627,N_16060,N_15623);
xnor U16628 (N_16628,N_15681,N_15733);
or U16629 (N_16629,N_15846,N_16165);
xor U16630 (N_16630,N_16139,N_16107);
nor U16631 (N_16631,N_15712,N_15971);
or U16632 (N_16632,N_15973,N_15919);
and U16633 (N_16633,N_15892,N_16170);
nand U16634 (N_16634,N_15796,N_16177);
nor U16635 (N_16635,N_15994,N_15649);
nand U16636 (N_16636,N_15934,N_15780);
or U16637 (N_16637,N_16189,N_16190);
and U16638 (N_16638,N_15950,N_16046);
or U16639 (N_16639,N_15694,N_15836);
or U16640 (N_16640,N_15723,N_16017);
and U16641 (N_16641,N_15900,N_16118);
xnor U16642 (N_16642,N_16062,N_16021);
xor U16643 (N_16643,N_15638,N_16130);
and U16644 (N_16644,N_16019,N_15817);
nand U16645 (N_16645,N_16196,N_15695);
xnor U16646 (N_16646,N_15640,N_16103);
xnor U16647 (N_16647,N_16186,N_16096);
xnor U16648 (N_16648,N_15839,N_15694);
nand U16649 (N_16649,N_16134,N_15870);
and U16650 (N_16650,N_16118,N_16020);
or U16651 (N_16651,N_15917,N_15895);
nand U16652 (N_16652,N_15910,N_16129);
nor U16653 (N_16653,N_15784,N_15604);
or U16654 (N_16654,N_16120,N_15944);
and U16655 (N_16655,N_15784,N_15829);
xnor U16656 (N_16656,N_15839,N_16158);
or U16657 (N_16657,N_16019,N_15981);
nand U16658 (N_16658,N_15671,N_15875);
or U16659 (N_16659,N_15946,N_16007);
nor U16660 (N_16660,N_15883,N_15784);
nor U16661 (N_16661,N_15918,N_15798);
nand U16662 (N_16662,N_16068,N_15959);
xnor U16663 (N_16663,N_15992,N_16002);
or U16664 (N_16664,N_15814,N_15914);
or U16665 (N_16665,N_15984,N_15614);
or U16666 (N_16666,N_16159,N_15659);
xnor U16667 (N_16667,N_15743,N_16020);
nor U16668 (N_16668,N_16179,N_15750);
nor U16669 (N_16669,N_15784,N_16081);
xnor U16670 (N_16670,N_16095,N_15691);
nand U16671 (N_16671,N_15628,N_15830);
or U16672 (N_16672,N_15994,N_15856);
nor U16673 (N_16673,N_15712,N_15855);
nor U16674 (N_16674,N_15817,N_15745);
and U16675 (N_16675,N_15928,N_15700);
nor U16676 (N_16676,N_15702,N_15630);
nand U16677 (N_16677,N_15607,N_15680);
nand U16678 (N_16678,N_16084,N_15841);
and U16679 (N_16679,N_15926,N_16053);
nor U16680 (N_16680,N_15969,N_16197);
nand U16681 (N_16681,N_16179,N_15602);
nor U16682 (N_16682,N_15855,N_15935);
nor U16683 (N_16683,N_15750,N_15883);
nor U16684 (N_16684,N_15729,N_16181);
nor U16685 (N_16685,N_15799,N_16099);
and U16686 (N_16686,N_15865,N_15645);
nand U16687 (N_16687,N_16057,N_16130);
nand U16688 (N_16688,N_15990,N_16175);
or U16689 (N_16689,N_15761,N_15915);
and U16690 (N_16690,N_15712,N_15801);
and U16691 (N_16691,N_15827,N_15903);
nand U16692 (N_16692,N_15672,N_15855);
and U16693 (N_16693,N_15725,N_15864);
nor U16694 (N_16694,N_15693,N_16136);
or U16695 (N_16695,N_15665,N_16149);
xnor U16696 (N_16696,N_15998,N_15735);
or U16697 (N_16697,N_15899,N_15614);
or U16698 (N_16698,N_15817,N_15881);
nor U16699 (N_16699,N_16042,N_15968);
and U16700 (N_16700,N_15933,N_15816);
nor U16701 (N_16701,N_15752,N_15899);
xor U16702 (N_16702,N_16120,N_16099);
xnor U16703 (N_16703,N_15910,N_16045);
or U16704 (N_16704,N_15939,N_16110);
xnor U16705 (N_16705,N_16070,N_15806);
and U16706 (N_16706,N_16100,N_15858);
or U16707 (N_16707,N_15803,N_15631);
or U16708 (N_16708,N_16194,N_15958);
nand U16709 (N_16709,N_15780,N_15625);
nand U16710 (N_16710,N_15778,N_15652);
or U16711 (N_16711,N_15919,N_15793);
nor U16712 (N_16712,N_16137,N_15731);
and U16713 (N_16713,N_16111,N_15898);
nor U16714 (N_16714,N_15614,N_16015);
nand U16715 (N_16715,N_15869,N_15794);
and U16716 (N_16716,N_16093,N_15756);
nor U16717 (N_16717,N_16114,N_15640);
or U16718 (N_16718,N_15815,N_15917);
or U16719 (N_16719,N_16183,N_15695);
nand U16720 (N_16720,N_15808,N_16176);
xnor U16721 (N_16721,N_15774,N_15765);
or U16722 (N_16722,N_15678,N_15666);
or U16723 (N_16723,N_15617,N_15730);
nand U16724 (N_16724,N_15827,N_15807);
xor U16725 (N_16725,N_15736,N_15879);
and U16726 (N_16726,N_15944,N_15877);
and U16727 (N_16727,N_15934,N_16180);
nand U16728 (N_16728,N_15682,N_15847);
xor U16729 (N_16729,N_15896,N_16181);
nand U16730 (N_16730,N_15864,N_15609);
nand U16731 (N_16731,N_15939,N_16192);
or U16732 (N_16732,N_15643,N_16025);
or U16733 (N_16733,N_16080,N_15958);
or U16734 (N_16734,N_15657,N_15960);
and U16735 (N_16735,N_15977,N_15712);
xor U16736 (N_16736,N_15681,N_15919);
and U16737 (N_16737,N_15767,N_15736);
or U16738 (N_16738,N_15913,N_15819);
xnor U16739 (N_16739,N_15856,N_15999);
nor U16740 (N_16740,N_16142,N_15735);
or U16741 (N_16741,N_15879,N_16069);
or U16742 (N_16742,N_15959,N_15851);
xnor U16743 (N_16743,N_15647,N_16129);
and U16744 (N_16744,N_15915,N_16065);
xnor U16745 (N_16745,N_16080,N_15881);
xnor U16746 (N_16746,N_15865,N_15963);
and U16747 (N_16747,N_15911,N_15725);
and U16748 (N_16748,N_15996,N_16182);
nand U16749 (N_16749,N_15989,N_15993);
xor U16750 (N_16750,N_15963,N_15910);
nor U16751 (N_16751,N_15832,N_15639);
nor U16752 (N_16752,N_16192,N_15662);
nor U16753 (N_16753,N_15874,N_16174);
or U16754 (N_16754,N_15791,N_15908);
or U16755 (N_16755,N_16181,N_15851);
or U16756 (N_16756,N_15648,N_15841);
or U16757 (N_16757,N_15802,N_16091);
and U16758 (N_16758,N_15714,N_16085);
and U16759 (N_16759,N_15652,N_15741);
nor U16760 (N_16760,N_15921,N_15808);
or U16761 (N_16761,N_15781,N_15861);
and U16762 (N_16762,N_15725,N_15782);
and U16763 (N_16763,N_15637,N_15780);
and U16764 (N_16764,N_16170,N_16109);
or U16765 (N_16765,N_15659,N_15661);
and U16766 (N_16766,N_15601,N_15906);
nand U16767 (N_16767,N_15690,N_16162);
and U16768 (N_16768,N_15981,N_15733);
and U16769 (N_16769,N_16176,N_16048);
nand U16770 (N_16770,N_15994,N_16160);
xor U16771 (N_16771,N_15904,N_15886);
nand U16772 (N_16772,N_15952,N_16071);
and U16773 (N_16773,N_15944,N_15656);
or U16774 (N_16774,N_16069,N_15685);
nand U16775 (N_16775,N_16169,N_16054);
nor U16776 (N_16776,N_16096,N_15954);
and U16777 (N_16777,N_15607,N_16182);
xor U16778 (N_16778,N_15624,N_15710);
nor U16779 (N_16779,N_15869,N_15783);
or U16780 (N_16780,N_15854,N_16005);
or U16781 (N_16781,N_15668,N_16053);
nand U16782 (N_16782,N_15769,N_15951);
or U16783 (N_16783,N_15813,N_15761);
nor U16784 (N_16784,N_16071,N_16156);
and U16785 (N_16785,N_16093,N_15607);
nor U16786 (N_16786,N_16172,N_15681);
nor U16787 (N_16787,N_15891,N_15905);
nand U16788 (N_16788,N_15693,N_16027);
and U16789 (N_16789,N_15637,N_15815);
and U16790 (N_16790,N_15733,N_15755);
xor U16791 (N_16791,N_15821,N_15921);
nor U16792 (N_16792,N_15998,N_15785);
xnor U16793 (N_16793,N_15759,N_15688);
and U16794 (N_16794,N_15663,N_16078);
nand U16795 (N_16795,N_15742,N_15929);
xnor U16796 (N_16796,N_16124,N_16098);
and U16797 (N_16797,N_15885,N_15714);
nor U16798 (N_16798,N_15882,N_15856);
or U16799 (N_16799,N_15641,N_15646);
xnor U16800 (N_16800,N_16722,N_16254);
xor U16801 (N_16801,N_16530,N_16293);
and U16802 (N_16802,N_16288,N_16601);
nor U16803 (N_16803,N_16501,N_16684);
nand U16804 (N_16804,N_16215,N_16306);
or U16805 (N_16805,N_16205,N_16756);
nor U16806 (N_16806,N_16707,N_16490);
xnor U16807 (N_16807,N_16551,N_16588);
nand U16808 (N_16808,N_16364,N_16558);
xor U16809 (N_16809,N_16370,N_16791);
nor U16810 (N_16810,N_16731,N_16708);
nand U16811 (N_16811,N_16214,N_16474);
xor U16812 (N_16812,N_16275,N_16500);
nor U16813 (N_16813,N_16415,N_16308);
or U16814 (N_16814,N_16630,N_16298);
xnor U16815 (N_16815,N_16483,N_16590);
xnor U16816 (N_16816,N_16413,N_16251);
nor U16817 (N_16817,N_16672,N_16663);
or U16818 (N_16818,N_16318,N_16753);
and U16819 (N_16819,N_16286,N_16462);
and U16820 (N_16820,N_16538,N_16648);
or U16821 (N_16821,N_16466,N_16238);
nand U16822 (N_16822,N_16494,N_16556);
and U16823 (N_16823,N_16662,N_16699);
nand U16824 (N_16824,N_16673,N_16777);
or U16825 (N_16825,N_16299,N_16626);
nor U16826 (N_16826,N_16326,N_16635);
nand U16827 (N_16827,N_16495,N_16263);
and U16828 (N_16828,N_16455,N_16411);
or U16829 (N_16829,N_16587,N_16305);
nor U16830 (N_16830,N_16464,N_16217);
xnor U16831 (N_16831,N_16624,N_16422);
xnor U16832 (N_16832,N_16330,N_16343);
and U16833 (N_16833,N_16646,N_16654);
nor U16834 (N_16834,N_16287,N_16712);
and U16835 (N_16835,N_16666,N_16231);
and U16836 (N_16836,N_16525,N_16241);
and U16837 (N_16837,N_16581,N_16645);
xor U16838 (N_16838,N_16797,N_16509);
nor U16839 (N_16839,N_16738,N_16599);
or U16840 (N_16840,N_16657,N_16341);
or U16841 (N_16841,N_16697,N_16467);
xor U16842 (N_16842,N_16638,N_16211);
xnor U16843 (N_16843,N_16683,N_16499);
nor U16844 (N_16844,N_16468,N_16732);
or U16845 (N_16845,N_16799,N_16236);
nand U16846 (N_16846,N_16545,N_16507);
nor U16847 (N_16847,N_16677,N_16442);
nor U16848 (N_16848,N_16356,N_16210);
nor U16849 (N_16849,N_16678,N_16562);
or U16850 (N_16850,N_16594,N_16786);
nand U16851 (N_16851,N_16432,N_16389);
nor U16852 (N_16852,N_16418,N_16276);
nand U16853 (N_16853,N_16283,N_16284);
nor U16854 (N_16854,N_16395,N_16227);
xor U16855 (N_16855,N_16434,N_16213);
or U16856 (N_16856,N_16269,N_16260);
xor U16857 (N_16857,N_16273,N_16573);
nand U16858 (N_16858,N_16569,N_16685);
and U16859 (N_16859,N_16655,N_16519);
and U16860 (N_16860,N_16475,N_16783);
xor U16861 (N_16861,N_16393,N_16259);
or U16862 (N_16862,N_16378,N_16570);
nand U16863 (N_16863,N_16669,N_16255);
nor U16864 (N_16864,N_16261,N_16681);
nand U16865 (N_16865,N_16610,N_16472);
xor U16866 (N_16866,N_16679,N_16511);
and U16867 (N_16867,N_16279,N_16565);
or U16868 (N_16868,N_16307,N_16752);
and U16869 (N_16869,N_16243,N_16785);
nor U16870 (N_16870,N_16513,N_16720);
nor U16871 (N_16871,N_16516,N_16354);
and U16872 (N_16872,N_16268,N_16692);
or U16873 (N_16873,N_16376,N_16314);
nor U16874 (N_16874,N_16717,N_16220);
nand U16875 (N_16875,N_16244,N_16249);
or U16876 (N_16876,N_16576,N_16652);
and U16877 (N_16877,N_16580,N_16774);
or U16878 (N_16878,N_16438,N_16715);
nand U16879 (N_16879,N_16399,N_16333);
xor U16880 (N_16880,N_16613,N_16367);
and U16881 (N_16881,N_16484,N_16651);
nor U16882 (N_16882,N_16765,N_16424);
and U16883 (N_16883,N_16201,N_16271);
and U16884 (N_16884,N_16589,N_16609);
or U16885 (N_16885,N_16470,N_16757);
xor U16886 (N_16886,N_16480,N_16769);
nor U16887 (N_16887,N_16760,N_16705);
or U16888 (N_16888,N_16704,N_16502);
xnor U16889 (N_16889,N_16749,N_16414);
nand U16890 (N_16890,N_16452,N_16232);
and U16891 (N_16891,N_16706,N_16703);
and U16892 (N_16892,N_16459,N_16346);
xnor U16893 (N_16893,N_16543,N_16405);
nor U16894 (N_16894,N_16762,N_16686);
or U16895 (N_16895,N_16453,N_16487);
nor U16896 (N_16896,N_16351,N_16374);
or U16897 (N_16897,N_16301,N_16793);
and U16898 (N_16898,N_16278,N_16242);
nor U16899 (N_16899,N_16397,N_16714);
nor U16900 (N_16900,N_16695,N_16781);
and U16901 (N_16901,N_16579,N_16441);
or U16902 (N_16902,N_16449,N_16221);
and U16903 (N_16903,N_16444,N_16317);
xnor U16904 (N_16904,N_16404,N_16529);
nor U16905 (N_16905,N_16764,N_16741);
and U16906 (N_16906,N_16637,N_16302);
xor U16907 (N_16907,N_16602,N_16312);
or U16908 (N_16908,N_16366,N_16548);
nand U16909 (N_16909,N_16325,N_16554);
xor U16910 (N_16910,N_16571,N_16375);
nor U16911 (N_16911,N_16734,N_16440);
xnor U16912 (N_16912,N_16230,N_16552);
or U16913 (N_16913,N_16748,N_16761);
and U16914 (N_16914,N_16246,N_16329);
xor U16915 (N_16915,N_16469,N_16369);
and U16916 (N_16916,N_16674,N_16607);
nor U16917 (N_16917,N_16402,N_16650);
xor U16918 (N_16918,N_16234,N_16694);
and U16919 (N_16919,N_16612,N_16512);
xnor U16920 (N_16920,N_16533,N_16479);
and U16921 (N_16921,N_16770,N_16547);
nor U16922 (N_16922,N_16553,N_16206);
xnor U16923 (N_16923,N_16471,N_16292);
xnor U16924 (N_16924,N_16486,N_16659);
nand U16925 (N_16925,N_16448,N_16642);
nor U16926 (N_16926,N_16398,N_16661);
nor U16927 (N_16927,N_16429,N_16544);
and U16928 (N_16928,N_16270,N_16372);
nor U16929 (N_16929,N_16400,N_16563);
xnor U16930 (N_16930,N_16394,N_16716);
or U16931 (N_16931,N_16328,N_16361);
and U16932 (N_16932,N_16258,N_16435);
nor U16933 (N_16933,N_16682,N_16639);
or U16934 (N_16934,N_16381,N_16640);
nand U16935 (N_16935,N_16297,N_16225);
xor U16936 (N_16936,N_16758,N_16339);
xor U16937 (N_16937,N_16634,N_16212);
and U16938 (N_16938,N_16790,N_16342);
nor U16939 (N_16939,N_16280,N_16632);
and U16940 (N_16940,N_16537,N_16368);
nor U16941 (N_16941,N_16332,N_16463);
and U16942 (N_16942,N_16226,N_16660);
nor U16943 (N_16943,N_16403,N_16496);
xnor U16944 (N_16944,N_16416,N_16702);
nor U16945 (N_16945,N_16555,N_16606);
xor U16946 (N_16946,N_16627,N_16478);
nand U16947 (N_16947,N_16281,N_16725);
nor U16948 (N_16948,N_16262,N_16207);
and U16949 (N_16949,N_16713,N_16629);
nand U16950 (N_16950,N_16535,N_16505);
and U16951 (N_16951,N_16798,N_16492);
xnor U16952 (N_16952,N_16766,N_16481);
and U16953 (N_16953,N_16727,N_16526);
and U16954 (N_16954,N_16473,N_16387);
and U16955 (N_16955,N_16605,N_16245);
nand U16956 (N_16956,N_16296,N_16322);
xor U16957 (N_16957,N_16506,N_16524);
and U16958 (N_16958,N_16755,N_16460);
or U16959 (N_16959,N_16614,N_16742);
or U16960 (N_16960,N_16250,N_16477);
nand U16961 (N_16961,N_16508,N_16335);
xor U16962 (N_16962,N_16362,N_16643);
and U16963 (N_16963,N_16313,N_16566);
or U16964 (N_16964,N_16355,N_16726);
nand U16965 (N_16965,N_16751,N_16754);
and U16966 (N_16966,N_16349,N_16779);
or U16967 (N_16967,N_16656,N_16363);
xnor U16968 (N_16968,N_16358,N_16598);
or U16969 (N_16969,N_16584,N_16687);
and U16970 (N_16970,N_16745,N_16597);
nand U16971 (N_16971,N_16653,N_16482);
nand U16972 (N_16972,N_16359,N_16750);
or U16973 (N_16973,N_16377,N_16578);
nor U16974 (N_16974,N_16202,N_16736);
or U16975 (N_16975,N_16222,N_16433);
or U16976 (N_16976,N_16491,N_16218);
xor U16977 (N_16977,N_16203,N_16316);
nor U16978 (N_16978,N_16711,N_16267);
nor U16979 (N_16979,N_16353,N_16383);
or U16980 (N_16980,N_16497,N_16796);
xor U16981 (N_16981,N_16721,N_16309);
and U16982 (N_16982,N_16461,N_16304);
nand U16983 (N_16983,N_16410,N_16572);
nor U16984 (N_16984,N_16382,N_16425);
and U16985 (N_16985,N_16303,N_16616);
nor U16986 (N_16986,N_16621,N_16550);
nand U16987 (N_16987,N_16780,N_16690);
xor U16988 (N_16988,N_16515,N_16771);
xnor U16989 (N_16989,N_16772,N_16619);
xor U16990 (N_16990,N_16265,N_16423);
nor U16991 (N_16991,N_16503,N_16560);
or U16992 (N_16992,N_16380,N_16357);
and U16993 (N_16993,N_16264,N_16345);
xor U16994 (N_16994,N_16608,N_16523);
and U16995 (N_16995,N_16493,N_16586);
or U16996 (N_16996,N_16676,N_16379);
xnor U16997 (N_16997,N_16730,N_16527);
and U16998 (N_16998,N_16208,N_16583);
or U16999 (N_16999,N_16295,N_16457);
nand U17000 (N_17000,N_16604,N_16622);
nand U17001 (N_17001,N_16744,N_16360);
xor U17002 (N_17002,N_16253,N_16409);
nor U17003 (N_17003,N_16549,N_16696);
or U17004 (N_17004,N_16784,N_16320);
or U17005 (N_17005,N_16740,N_16216);
nand U17006 (N_17006,N_16788,N_16248);
and U17007 (N_17007,N_16392,N_16504);
xor U17008 (N_17008,N_16311,N_16488);
xnor U17009 (N_17009,N_16794,N_16577);
xnor U17010 (N_17010,N_16615,N_16778);
and U17011 (N_17011,N_16521,N_16561);
nor U17012 (N_17012,N_16291,N_16710);
nor U17013 (N_17013,N_16665,N_16520);
and U17014 (N_17014,N_16200,N_16729);
xnor U17015 (N_17015,N_16628,N_16776);
nand U17016 (N_17016,N_16600,N_16219);
nor U17017 (N_17017,N_16485,N_16795);
and U17018 (N_17018,N_16443,N_16617);
xor U17019 (N_17019,N_16542,N_16417);
nor U17020 (N_17020,N_16340,N_16735);
xnor U17021 (N_17021,N_16228,N_16540);
nand U17022 (N_17022,N_16718,N_16446);
and U17023 (N_17023,N_16739,N_16454);
xor U17024 (N_17024,N_16396,N_16644);
and U17025 (N_17025,N_16240,N_16428);
nand U17026 (N_17026,N_16724,N_16390);
and U17027 (N_17027,N_16277,N_16719);
nand U17028 (N_17028,N_16224,N_16532);
or U17029 (N_17029,N_16746,N_16768);
nand U17030 (N_17030,N_16310,N_16290);
or U17031 (N_17031,N_16235,N_16782);
nor U17032 (N_17032,N_16327,N_16633);
nor U17033 (N_17033,N_16406,N_16625);
and U17034 (N_17034,N_16664,N_16620);
xor U17035 (N_17035,N_16728,N_16559);
nand U17036 (N_17036,N_16531,N_16282);
nand U17037 (N_17037,N_16763,N_16723);
and U17038 (N_17038,N_16266,N_16347);
or U17039 (N_17039,N_16334,N_16239);
xor U17040 (N_17040,N_16568,N_16237);
nor U17041 (N_17041,N_16274,N_16675);
nand U17042 (N_17042,N_16350,N_16336);
nor U17043 (N_17043,N_16591,N_16671);
or U17044 (N_17044,N_16668,N_16450);
and U17045 (N_17045,N_16534,N_16517);
xor U17046 (N_17046,N_16385,N_16384);
xor U17047 (N_17047,N_16585,N_16733);
nor U17048 (N_17048,N_16344,N_16458);
nor U17049 (N_17049,N_16408,N_16518);
nand U17050 (N_17050,N_16421,N_16223);
and U17051 (N_17051,N_16700,N_16787);
xor U17052 (N_17052,N_16430,N_16257);
nand U17053 (N_17053,N_16419,N_16365);
xnor U17054 (N_17054,N_16431,N_16510);
nand U17055 (N_17055,N_16256,N_16593);
or U17056 (N_17056,N_16420,N_16689);
nand U17057 (N_17057,N_16331,N_16658);
nor U17058 (N_17058,N_16747,N_16595);
and U17059 (N_17059,N_16536,N_16528);
nor U17060 (N_17060,N_16759,N_16557);
nor U17061 (N_17061,N_16636,N_16680);
nor U17062 (N_17062,N_16285,N_16348);
nand U17063 (N_17063,N_16436,N_16323);
and U17064 (N_17064,N_16564,N_16514);
and U17065 (N_17065,N_16294,N_16371);
or U17066 (N_17066,N_16670,N_16391);
xnor U17067 (N_17067,N_16596,N_16289);
or U17068 (N_17068,N_16412,N_16247);
or U17069 (N_17069,N_16447,N_16300);
and U17070 (N_17070,N_16603,N_16324);
nor U17071 (N_17071,N_16352,N_16321);
xor U17072 (N_17072,N_16539,N_16465);
or U17073 (N_17073,N_16233,N_16641);
nor U17074 (N_17074,N_16743,N_16337);
xnor U17075 (N_17075,N_16574,N_16775);
nor U17076 (N_17076,N_16618,N_16792);
xnor U17077 (N_17077,N_16407,N_16623);
or U17078 (N_17078,N_16427,N_16575);
and U17079 (N_17079,N_16582,N_16209);
nor U17080 (N_17080,N_16767,N_16698);
xnor U17081 (N_17081,N_16426,N_16204);
and U17082 (N_17082,N_16737,N_16476);
nand U17083 (N_17083,N_16338,N_16691);
xor U17084 (N_17084,N_16647,N_16445);
or U17085 (N_17085,N_16649,N_16451);
nand U17086 (N_17086,N_16546,N_16688);
nand U17087 (N_17087,N_16439,N_16319);
xor U17088 (N_17088,N_16437,N_16386);
or U17089 (N_17089,N_16229,N_16489);
xnor U17090 (N_17090,N_16701,N_16522);
nand U17091 (N_17091,N_16693,N_16631);
nand U17092 (N_17092,N_16709,N_16773);
or U17093 (N_17093,N_16315,N_16272);
nor U17094 (N_17094,N_16498,N_16567);
or U17095 (N_17095,N_16789,N_16401);
nand U17096 (N_17096,N_16456,N_16592);
and U17097 (N_17097,N_16541,N_16373);
xnor U17098 (N_17098,N_16388,N_16252);
and U17099 (N_17099,N_16611,N_16667);
or U17100 (N_17100,N_16640,N_16277);
or U17101 (N_17101,N_16736,N_16200);
nand U17102 (N_17102,N_16623,N_16784);
or U17103 (N_17103,N_16542,N_16372);
xnor U17104 (N_17104,N_16667,N_16464);
xnor U17105 (N_17105,N_16466,N_16641);
nor U17106 (N_17106,N_16722,N_16327);
xor U17107 (N_17107,N_16642,N_16340);
and U17108 (N_17108,N_16309,N_16799);
nand U17109 (N_17109,N_16748,N_16564);
nor U17110 (N_17110,N_16646,N_16360);
or U17111 (N_17111,N_16455,N_16275);
or U17112 (N_17112,N_16386,N_16740);
xnor U17113 (N_17113,N_16250,N_16307);
nor U17114 (N_17114,N_16369,N_16397);
nand U17115 (N_17115,N_16757,N_16722);
xor U17116 (N_17116,N_16668,N_16719);
and U17117 (N_17117,N_16470,N_16519);
xor U17118 (N_17118,N_16686,N_16400);
xnor U17119 (N_17119,N_16747,N_16214);
nor U17120 (N_17120,N_16205,N_16310);
xnor U17121 (N_17121,N_16687,N_16768);
nor U17122 (N_17122,N_16464,N_16385);
xor U17123 (N_17123,N_16232,N_16734);
nand U17124 (N_17124,N_16277,N_16556);
or U17125 (N_17125,N_16524,N_16392);
or U17126 (N_17126,N_16207,N_16629);
nand U17127 (N_17127,N_16682,N_16631);
nor U17128 (N_17128,N_16594,N_16414);
nor U17129 (N_17129,N_16212,N_16216);
or U17130 (N_17130,N_16304,N_16376);
and U17131 (N_17131,N_16269,N_16291);
nor U17132 (N_17132,N_16677,N_16774);
xnor U17133 (N_17133,N_16251,N_16331);
nand U17134 (N_17134,N_16533,N_16308);
nor U17135 (N_17135,N_16561,N_16494);
and U17136 (N_17136,N_16573,N_16422);
nand U17137 (N_17137,N_16789,N_16343);
xor U17138 (N_17138,N_16348,N_16625);
xnor U17139 (N_17139,N_16562,N_16564);
nor U17140 (N_17140,N_16303,N_16217);
xnor U17141 (N_17141,N_16630,N_16643);
nand U17142 (N_17142,N_16719,N_16772);
nor U17143 (N_17143,N_16324,N_16411);
nor U17144 (N_17144,N_16218,N_16247);
nor U17145 (N_17145,N_16601,N_16511);
and U17146 (N_17146,N_16742,N_16344);
and U17147 (N_17147,N_16447,N_16358);
nor U17148 (N_17148,N_16576,N_16439);
xor U17149 (N_17149,N_16733,N_16518);
nor U17150 (N_17150,N_16544,N_16411);
xor U17151 (N_17151,N_16380,N_16315);
and U17152 (N_17152,N_16724,N_16221);
and U17153 (N_17153,N_16663,N_16252);
nor U17154 (N_17154,N_16231,N_16354);
nand U17155 (N_17155,N_16551,N_16410);
and U17156 (N_17156,N_16794,N_16671);
nand U17157 (N_17157,N_16535,N_16293);
and U17158 (N_17158,N_16726,N_16576);
nand U17159 (N_17159,N_16470,N_16636);
nand U17160 (N_17160,N_16577,N_16409);
nand U17161 (N_17161,N_16590,N_16751);
and U17162 (N_17162,N_16703,N_16414);
or U17163 (N_17163,N_16669,N_16643);
and U17164 (N_17164,N_16527,N_16708);
xnor U17165 (N_17165,N_16466,N_16355);
nand U17166 (N_17166,N_16271,N_16463);
and U17167 (N_17167,N_16421,N_16626);
nor U17168 (N_17168,N_16418,N_16402);
or U17169 (N_17169,N_16570,N_16531);
or U17170 (N_17170,N_16680,N_16758);
nor U17171 (N_17171,N_16390,N_16437);
and U17172 (N_17172,N_16272,N_16257);
xnor U17173 (N_17173,N_16557,N_16334);
nor U17174 (N_17174,N_16388,N_16405);
xor U17175 (N_17175,N_16629,N_16436);
xnor U17176 (N_17176,N_16436,N_16406);
nand U17177 (N_17177,N_16521,N_16243);
and U17178 (N_17178,N_16290,N_16794);
and U17179 (N_17179,N_16786,N_16497);
nand U17180 (N_17180,N_16568,N_16646);
nor U17181 (N_17181,N_16657,N_16437);
nor U17182 (N_17182,N_16351,N_16369);
nor U17183 (N_17183,N_16494,N_16461);
xor U17184 (N_17184,N_16389,N_16459);
nor U17185 (N_17185,N_16356,N_16259);
nand U17186 (N_17186,N_16222,N_16545);
nor U17187 (N_17187,N_16763,N_16598);
xor U17188 (N_17188,N_16687,N_16210);
nand U17189 (N_17189,N_16789,N_16271);
nor U17190 (N_17190,N_16497,N_16385);
and U17191 (N_17191,N_16612,N_16589);
or U17192 (N_17192,N_16468,N_16724);
xor U17193 (N_17193,N_16571,N_16308);
xnor U17194 (N_17194,N_16602,N_16464);
nand U17195 (N_17195,N_16246,N_16400);
xnor U17196 (N_17196,N_16564,N_16344);
nor U17197 (N_17197,N_16526,N_16510);
xnor U17198 (N_17198,N_16767,N_16776);
and U17199 (N_17199,N_16426,N_16768);
and U17200 (N_17200,N_16291,N_16369);
xnor U17201 (N_17201,N_16622,N_16415);
xor U17202 (N_17202,N_16354,N_16743);
xnor U17203 (N_17203,N_16644,N_16719);
xnor U17204 (N_17204,N_16700,N_16293);
nand U17205 (N_17205,N_16567,N_16210);
xnor U17206 (N_17206,N_16532,N_16770);
and U17207 (N_17207,N_16502,N_16707);
nor U17208 (N_17208,N_16340,N_16281);
nand U17209 (N_17209,N_16336,N_16522);
and U17210 (N_17210,N_16718,N_16799);
xor U17211 (N_17211,N_16307,N_16600);
nand U17212 (N_17212,N_16548,N_16293);
or U17213 (N_17213,N_16540,N_16641);
nand U17214 (N_17214,N_16243,N_16691);
or U17215 (N_17215,N_16212,N_16229);
or U17216 (N_17216,N_16226,N_16285);
xnor U17217 (N_17217,N_16743,N_16227);
nor U17218 (N_17218,N_16218,N_16203);
or U17219 (N_17219,N_16321,N_16219);
xnor U17220 (N_17220,N_16528,N_16232);
nand U17221 (N_17221,N_16333,N_16352);
nand U17222 (N_17222,N_16585,N_16328);
nand U17223 (N_17223,N_16675,N_16439);
or U17224 (N_17224,N_16383,N_16598);
and U17225 (N_17225,N_16681,N_16554);
xnor U17226 (N_17226,N_16547,N_16386);
nand U17227 (N_17227,N_16362,N_16535);
nand U17228 (N_17228,N_16314,N_16542);
nor U17229 (N_17229,N_16484,N_16629);
and U17230 (N_17230,N_16461,N_16305);
nand U17231 (N_17231,N_16792,N_16298);
and U17232 (N_17232,N_16409,N_16336);
xor U17233 (N_17233,N_16359,N_16284);
nand U17234 (N_17234,N_16772,N_16303);
and U17235 (N_17235,N_16469,N_16224);
and U17236 (N_17236,N_16241,N_16709);
nand U17237 (N_17237,N_16477,N_16531);
and U17238 (N_17238,N_16676,N_16310);
nor U17239 (N_17239,N_16236,N_16486);
xor U17240 (N_17240,N_16538,N_16475);
xnor U17241 (N_17241,N_16369,N_16519);
xnor U17242 (N_17242,N_16304,N_16357);
nand U17243 (N_17243,N_16494,N_16592);
nand U17244 (N_17244,N_16269,N_16721);
nand U17245 (N_17245,N_16446,N_16339);
nand U17246 (N_17246,N_16392,N_16630);
or U17247 (N_17247,N_16421,N_16505);
nor U17248 (N_17248,N_16597,N_16443);
xnor U17249 (N_17249,N_16469,N_16495);
nand U17250 (N_17250,N_16328,N_16565);
or U17251 (N_17251,N_16334,N_16287);
xnor U17252 (N_17252,N_16749,N_16654);
or U17253 (N_17253,N_16515,N_16587);
nand U17254 (N_17254,N_16237,N_16604);
or U17255 (N_17255,N_16287,N_16691);
or U17256 (N_17256,N_16727,N_16304);
nand U17257 (N_17257,N_16367,N_16582);
and U17258 (N_17258,N_16515,N_16362);
and U17259 (N_17259,N_16259,N_16737);
xnor U17260 (N_17260,N_16732,N_16213);
nor U17261 (N_17261,N_16767,N_16341);
xor U17262 (N_17262,N_16351,N_16242);
nor U17263 (N_17263,N_16618,N_16585);
nand U17264 (N_17264,N_16761,N_16459);
nor U17265 (N_17265,N_16792,N_16527);
xnor U17266 (N_17266,N_16791,N_16730);
and U17267 (N_17267,N_16649,N_16434);
nor U17268 (N_17268,N_16407,N_16489);
or U17269 (N_17269,N_16606,N_16435);
or U17270 (N_17270,N_16216,N_16626);
nand U17271 (N_17271,N_16569,N_16485);
nor U17272 (N_17272,N_16415,N_16729);
nand U17273 (N_17273,N_16402,N_16611);
nand U17274 (N_17274,N_16264,N_16292);
or U17275 (N_17275,N_16304,N_16622);
xor U17276 (N_17276,N_16662,N_16354);
or U17277 (N_17277,N_16543,N_16402);
and U17278 (N_17278,N_16518,N_16308);
xnor U17279 (N_17279,N_16684,N_16458);
and U17280 (N_17280,N_16224,N_16610);
nor U17281 (N_17281,N_16335,N_16235);
nor U17282 (N_17282,N_16454,N_16752);
or U17283 (N_17283,N_16396,N_16245);
and U17284 (N_17284,N_16346,N_16692);
nor U17285 (N_17285,N_16388,N_16205);
nor U17286 (N_17286,N_16631,N_16700);
and U17287 (N_17287,N_16426,N_16496);
and U17288 (N_17288,N_16530,N_16220);
nor U17289 (N_17289,N_16796,N_16509);
and U17290 (N_17290,N_16788,N_16221);
nor U17291 (N_17291,N_16710,N_16256);
or U17292 (N_17292,N_16797,N_16439);
nand U17293 (N_17293,N_16489,N_16266);
nor U17294 (N_17294,N_16424,N_16255);
and U17295 (N_17295,N_16382,N_16583);
and U17296 (N_17296,N_16582,N_16781);
xnor U17297 (N_17297,N_16391,N_16300);
nand U17298 (N_17298,N_16491,N_16622);
and U17299 (N_17299,N_16320,N_16615);
xnor U17300 (N_17300,N_16397,N_16297);
nand U17301 (N_17301,N_16328,N_16243);
nand U17302 (N_17302,N_16636,N_16737);
xnor U17303 (N_17303,N_16208,N_16243);
xor U17304 (N_17304,N_16796,N_16751);
xor U17305 (N_17305,N_16768,N_16273);
nand U17306 (N_17306,N_16538,N_16602);
nand U17307 (N_17307,N_16726,N_16676);
xor U17308 (N_17308,N_16603,N_16378);
nand U17309 (N_17309,N_16500,N_16798);
xnor U17310 (N_17310,N_16529,N_16764);
xnor U17311 (N_17311,N_16612,N_16650);
nor U17312 (N_17312,N_16492,N_16446);
and U17313 (N_17313,N_16744,N_16447);
or U17314 (N_17314,N_16338,N_16595);
or U17315 (N_17315,N_16412,N_16512);
or U17316 (N_17316,N_16344,N_16616);
nor U17317 (N_17317,N_16363,N_16406);
nor U17318 (N_17318,N_16393,N_16610);
nor U17319 (N_17319,N_16291,N_16288);
nand U17320 (N_17320,N_16752,N_16510);
or U17321 (N_17321,N_16489,N_16393);
or U17322 (N_17322,N_16461,N_16302);
nor U17323 (N_17323,N_16700,N_16614);
nand U17324 (N_17324,N_16639,N_16537);
nor U17325 (N_17325,N_16386,N_16293);
nor U17326 (N_17326,N_16664,N_16440);
or U17327 (N_17327,N_16640,N_16308);
or U17328 (N_17328,N_16718,N_16290);
nand U17329 (N_17329,N_16614,N_16702);
and U17330 (N_17330,N_16516,N_16723);
and U17331 (N_17331,N_16545,N_16678);
and U17332 (N_17332,N_16227,N_16645);
or U17333 (N_17333,N_16685,N_16465);
or U17334 (N_17334,N_16603,N_16620);
nand U17335 (N_17335,N_16498,N_16488);
xnor U17336 (N_17336,N_16563,N_16454);
xor U17337 (N_17337,N_16487,N_16298);
nand U17338 (N_17338,N_16667,N_16331);
and U17339 (N_17339,N_16218,N_16586);
nor U17340 (N_17340,N_16302,N_16517);
or U17341 (N_17341,N_16550,N_16340);
nor U17342 (N_17342,N_16562,N_16236);
nor U17343 (N_17343,N_16549,N_16497);
or U17344 (N_17344,N_16248,N_16369);
or U17345 (N_17345,N_16395,N_16388);
nand U17346 (N_17346,N_16567,N_16282);
nor U17347 (N_17347,N_16792,N_16682);
nor U17348 (N_17348,N_16549,N_16396);
or U17349 (N_17349,N_16706,N_16435);
or U17350 (N_17350,N_16240,N_16475);
nand U17351 (N_17351,N_16778,N_16570);
nand U17352 (N_17352,N_16438,N_16244);
nor U17353 (N_17353,N_16697,N_16781);
nor U17354 (N_17354,N_16789,N_16565);
nand U17355 (N_17355,N_16214,N_16530);
nand U17356 (N_17356,N_16388,N_16456);
xor U17357 (N_17357,N_16487,N_16576);
nand U17358 (N_17358,N_16452,N_16619);
and U17359 (N_17359,N_16312,N_16440);
nand U17360 (N_17360,N_16370,N_16610);
and U17361 (N_17361,N_16520,N_16401);
nand U17362 (N_17362,N_16324,N_16547);
or U17363 (N_17363,N_16477,N_16262);
nand U17364 (N_17364,N_16528,N_16357);
nor U17365 (N_17365,N_16327,N_16366);
xor U17366 (N_17366,N_16751,N_16388);
and U17367 (N_17367,N_16603,N_16479);
or U17368 (N_17368,N_16377,N_16338);
xnor U17369 (N_17369,N_16212,N_16641);
or U17370 (N_17370,N_16458,N_16503);
or U17371 (N_17371,N_16306,N_16259);
or U17372 (N_17372,N_16784,N_16354);
or U17373 (N_17373,N_16640,N_16551);
xnor U17374 (N_17374,N_16257,N_16281);
or U17375 (N_17375,N_16791,N_16610);
xnor U17376 (N_17376,N_16603,N_16396);
xor U17377 (N_17377,N_16572,N_16641);
nand U17378 (N_17378,N_16785,N_16588);
xnor U17379 (N_17379,N_16295,N_16385);
nor U17380 (N_17380,N_16585,N_16529);
or U17381 (N_17381,N_16209,N_16342);
xor U17382 (N_17382,N_16459,N_16297);
or U17383 (N_17383,N_16395,N_16243);
xor U17384 (N_17384,N_16609,N_16345);
nor U17385 (N_17385,N_16678,N_16286);
and U17386 (N_17386,N_16225,N_16592);
nand U17387 (N_17387,N_16226,N_16690);
nand U17388 (N_17388,N_16302,N_16733);
or U17389 (N_17389,N_16420,N_16409);
nor U17390 (N_17390,N_16366,N_16256);
and U17391 (N_17391,N_16562,N_16314);
nor U17392 (N_17392,N_16411,N_16686);
or U17393 (N_17393,N_16227,N_16587);
or U17394 (N_17394,N_16725,N_16319);
or U17395 (N_17395,N_16623,N_16238);
and U17396 (N_17396,N_16378,N_16344);
nand U17397 (N_17397,N_16433,N_16466);
nor U17398 (N_17398,N_16725,N_16458);
xor U17399 (N_17399,N_16704,N_16765);
or U17400 (N_17400,N_17183,N_16986);
xor U17401 (N_17401,N_16964,N_17107);
nor U17402 (N_17402,N_16934,N_17348);
nor U17403 (N_17403,N_17039,N_17105);
nand U17404 (N_17404,N_16872,N_17067);
or U17405 (N_17405,N_16941,N_16914);
and U17406 (N_17406,N_17365,N_17174);
nand U17407 (N_17407,N_16957,N_16866);
nand U17408 (N_17408,N_17066,N_17180);
nand U17409 (N_17409,N_17239,N_17234);
and U17410 (N_17410,N_16898,N_16968);
xnor U17411 (N_17411,N_17188,N_17237);
and U17412 (N_17412,N_16810,N_17097);
or U17413 (N_17413,N_16924,N_16862);
and U17414 (N_17414,N_17335,N_17372);
or U17415 (N_17415,N_17203,N_17080);
or U17416 (N_17416,N_17255,N_17218);
nor U17417 (N_17417,N_17209,N_16827);
nor U17418 (N_17418,N_17143,N_16920);
nand U17419 (N_17419,N_17046,N_17160);
nand U17420 (N_17420,N_17198,N_17077);
nand U17421 (N_17421,N_17045,N_17224);
or U17422 (N_17422,N_17001,N_17199);
and U17423 (N_17423,N_16988,N_16992);
and U17424 (N_17424,N_17023,N_16916);
nand U17425 (N_17425,N_17125,N_17299);
xor U17426 (N_17426,N_17282,N_17060);
and U17427 (N_17427,N_16907,N_17185);
and U17428 (N_17428,N_16834,N_17337);
nand U17429 (N_17429,N_17018,N_17150);
nand U17430 (N_17430,N_17339,N_17298);
and U17431 (N_17431,N_16856,N_17296);
nor U17432 (N_17432,N_17050,N_16857);
and U17433 (N_17433,N_17280,N_16854);
xnor U17434 (N_17434,N_16825,N_17380);
nand U17435 (N_17435,N_17259,N_17379);
or U17436 (N_17436,N_17386,N_17243);
xnor U17437 (N_17437,N_17257,N_17394);
and U17438 (N_17438,N_17109,N_17363);
or U17439 (N_17439,N_17005,N_17164);
xor U17440 (N_17440,N_16822,N_17307);
and U17441 (N_17441,N_17300,N_17130);
xnor U17442 (N_17442,N_16967,N_17123);
and U17443 (N_17443,N_16930,N_17129);
and U17444 (N_17444,N_17207,N_16838);
nand U17445 (N_17445,N_17321,N_17085);
xor U17446 (N_17446,N_17070,N_17204);
and U17447 (N_17447,N_16929,N_16836);
or U17448 (N_17448,N_17373,N_17026);
nand U17449 (N_17449,N_17213,N_17202);
nor U17450 (N_17450,N_17187,N_17137);
or U17451 (N_17451,N_17162,N_17356);
or U17452 (N_17452,N_17270,N_17121);
nand U17453 (N_17453,N_16998,N_17163);
or U17454 (N_17454,N_16829,N_17169);
nand U17455 (N_17455,N_16855,N_17044);
and U17456 (N_17456,N_17059,N_17319);
or U17457 (N_17457,N_17101,N_17133);
nand U17458 (N_17458,N_16816,N_16864);
or U17459 (N_17459,N_16861,N_17397);
or U17460 (N_17460,N_16993,N_17306);
xnor U17461 (N_17461,N_16927,N_17167);
and U17462 (N_17462,N_17261,N_17030);
and U17463 (N_17463,N_17344,N_17057);
or U17464 (N_17464,N_17193,N_17399);
or U17465 (N_17465,N_16937,N_17336);
and U17466 (N_17466,N_16983,N_17275);
nor U17467 (N_17467,N_17233,N_17368);
or U17468 (N_17468,N_16972,N_17178);
xnor U17469 (N_17469,N_17036,N_16889);
nor U17470 (N_17470,N_17112,N_17278);
nor U17471 (N_17471,N_17008,N_17272);
and U17472 (N_17472,N_16812,N_17245);
and U17473 (N_17473,N_16936,N_17349);
nor U17474 (N_17474,N_17314,N_17113);
nor U17475 (N_17475,N_17342,N_16865);
xnor U17476 (N_17476,N_17316,N_17049);
xnor U17477 (N_17477,N_16935,N_16890);
nand U17478 (N_17478,N_16903,N_17020);
xnor U17479 (N_17479,N_17111,N_17327);
or U17480 (N_17480,N_16915,N_16805);
nor U17481 (N_17481,N_16840,N_17241);
and U17482 (N_17482,N_17040,N_17326);
and U17483 (N_17483,N_17374,N_17117);
and U17484 (N_17484,N_17144,N_17361);
nor U17485 (N_17485,N_17103,N_17012);
nand U17486 (N_17486,N_16945,N_17251);
and U17487 (N_17487,N_17106,N_16837);
xnor U17488 (N_17488,N_16876,N_16895);
xnor U17489 (N_17489,N_17014,N_16875);
nand U17490 (N_17490,N_16842,N_16873);
nand U17491 (N_17491,N_16852,N_16801);
xor U17492 (N_17492,N_16922,N_16959);
nand U17493 (N_17493,N_16991,N_16910);
nand U17494 (N_17494,N_16891,N_17093);
xor U17495 (N_17495,N_16996,N_17279);
xnor U17496 (N_17496,N_16943,N_17376);
xnor U17497 (N_17497,N_16860,N_17396);
and U17498 (N_17498,N_17242,N_16870);
and U17499 (N_17499,N_17208,N_16877);
nor U17500 (N_17500,N_17249,N_17304);
and U17501 (N_17501,N_17051,N_17263);
nor U17502 (N_17502,N_16949,N_17171);
and U17503 (N_17503,N_17041,N_17016);
and U17504 (N_17504,N_17353,N_17090);
nor U17505 (N_17505,N_17095,N_17240);
nand U17506 (N_17506,N_16974,N_17392);
nor U17507 (N_17507,N_16868,N_17317);
nor U17508 (N_17508,N_16995,N_17177);
nor U17509 (N_17509,N_16806,N_16802);
or U17510 (N_17510,N_16883,N_17158);
and U17511 (N_17511,N_17191,N_17276);
nand U17512 (N_17512,N_17220,N_16928);
nor U17513 (N_17513,N_16853,N_16939);
xor U17514 (N_17514,N_16884,N_17384);
or U17515 (N_17515,N_17146,N_17345);
and U17516 (N_17516,N_17000,N_17291);
and U17517 (N_17517,N_16824,N_17247);
nand U17518 (N_17518,N_16811,N_17389);
or U17519 (N_17519,N_17084,N_17205);
xor U17520 (N_17520,N_17217,N_16878);
xor U17521 (N_17521,N_17024,N_17056);
nor U17522 (N_17522,N_17294,N_16859);
xnor U17523 (N_17523,N_17229,N_17352);
nand U17524 (N_17524,N_17082,N_16841);
nand U17525 (N_17525,N_17140,N_17295);
nor U17526 (N_17526,N_17212,N_16953);
nand U17527 (N_17527,N_17385,N_16833);
or U17528 (N_17528,N_17227,N_17287);
or U17529 (N_17529,N_17366,N_16893);
and U17530 (N_17530,N_16908,N_17281);
and U17531 (N_17531,N_17273,N_16963);
xor U17532 (N_17532,N_17153,N_16880);
nor U17533 (N_17533,N_16932,N_17215);
or U17534 (N_17534,N_16913,N_17290);
or U17535 (N_17535,N_17110,N_17078);
xor U17536 (N_17536,N_17010,N_17232);
and U17537 (N_17537,N_17266,N_17250);
xor U17538 (N_17538,N_17214,N_17268);
or U17539 (N_17539,N_16980,N_16948);
nand U17540 (N_17540,N_17230,N_17099);
or U17541 (N_17541,N_16828,N_17116);
or U17542 (N_17542,N_17347,N_17136);
xnor U17543 (N_17543,N_17079,N_16808);
and U17544 (N_17544,N_16897,N_17120);
and U17545 (N_17545,N_17343,N_17302);
or U17546 (N_17546,N_16831,N_16814);
or U17547 (N_17547,N_17122,N_16809);
xor U17548 (N_17548,N_16848,N_17108);
or U17549 (N_17549,N_17391,N_17388);
or U17550 (N_17550,N_17246,N_17331);
nand U17551 (N_17551,N_17308,N_16997);
nand U17552 (N_17552,N_17312,N_17038);
nand U17553 (N_17553,N_17225,N_17328);
nand U17554 (N_17554,N_17069,N_17100);
nand U17555 (N_17555,N_16871,N_17081);
nor U17556 (N_17556,N_17252,N_16950);
and U17557 (N_17557,N_16961,N_16926);
and U17558 (N_17558,N_17064,N_17371);
or U17559 (N_17559,N_17118,N_17194);
xor U17560 (N_17560,N_17340,N_16817);
nand U17561 (N_17561,N_16919,N_16851);
nand U17562 (N_17562,N_16955,N_16905);
nand U17563 (N_17563,N_16844,N_17219);
xnor U17564 (N_17564,N_17184,N_17350);
or U17565 (N_17565,N_16940,N_17115);
nand U17566 (N_17566,N_16847,N_16909);
and U17567 (N_17567,N_16902,N_16921);
nand U17568 (N_17568,N_17310,N_17236);
or U17569 (N_17569,N_17285,N_16896);
or U17570 (N_17570,N_17009,N_16882);
or U17571 (N_17571,N_17062,N_17021);
xor U17572 (N_17572,N_17152,N_17139);
or U17573 (N_17573,N_17293,N_17387);
nor U17574 (N_17574,N_17223,N_16911);
and U17575 (N_17575,N_17311,N_17284);
and U17576 (N_17576,N_17025,N_16942);
nand U17577 (N_17577,N_16982,N_17119);
nor U17578 (N_17578,N_17052,N_17309);
nand U17579 (N_17579,N_16839,N_17149);
xor U17580 (N_17580,N_17341,N_16973);
nor U17581 (N_17581,N_17019,N_17135);
nor U17582 (N_17582,N_17271,N_17359);
xor U17583 (N_17583,N_17151,N_17034);
nor U17584 (N_17584,N_17269,N_17189);
and U17585 (N_17585,N_17313,N_16830);
or U17586 (N_17586,N_16999,N_17221);
nor U17587 (N_17587,N_16892,N_17186);
or U17588 (N_17588,N_17211,N_17173);
xnor U17589 (N_17589,N_17017,N_17053);
nor U17590 (N_17590,N_16804,N_17395);
nand U17591 (N_17591,N_16989,N_17170);
xnor U17592 (N_17592,N_17011,N_16901);
or U17593 (N_17593,N_17102,N_17007);
and U17594 (N_17594,N_17002,N_17004);
nand U17595 (N_17595,N_17088,N_16843);
and U17596 (N_17596,N_16969,N_17141);
nor U17597 (N_17597,N_17244,N_16931);
and U17598 (N_17598,N_17238,N_17231);
and U17599 (N_17599,N_16918,N_16849);
nor U17600 (N_17600,N_17006,N_16858);
and U17601 (N_17601,N_17159,N_16881);
or U17602 (N_17602,N_17092,N_17022);
xor U17603 (N_17603,N_16966,N_17325);
xnor U17604 (N_17604,N_16886,N_17003);
xnor U17605 (N_17605,N_17318,N_16826);
xor U17606 (N_17606,N_17351,N_16800);
nor U17607 (N_17607,N_17127,N_17334);
xor U17608 (N_17608,N_17201,N_16985);
or U17609 (N_17609,N_17283,N_17124);
and U17610 (N_17610,N_17148,N_17083);
and U17611 (N_17611,N_17155,N_17068);
nand U17612 (N_17612,N_16813,N_17200);
nand U17613 (N_17613,N_17377,N_16965);
and U17614 (N_17614,N_17333,N_17197);
and U17615 (N_17615,N_16832,N_16904);
nor U17616 (N_17616,N_17381,N_16888);
xor U17617 (N_17617,N_17383,N_16951);
xor U17618 (N_17618,N_17032,N_17104);
and U17619 (N_17619,N_16933,N_16899);
and U17620 (N_17620,N_16879,N_17364);
and U17621 (N_17621,N_16984,N_16962);
nand U17622 (N_17622,N_16917,N_17128);
xor U17623 (N_17623,N_17301,N_17226);
or U17624 (N_17624,N_17072,N_17027);
and U17625 (N_17625,N_17390,N_17013);
nand U17626 (N_17626,N_17235,N_16954);
nor U17627 (N_17627,N_17035,N_17055);
xor U17628 (N_17628,N_17132,N_17075);
and U17629 (N_17629,N_16887,N_17254);
nand U17630 (N_17630,N_16970,N_17156);
or U17631 (N_17631,N_17248,N_17031);
or U17632 (N_17632,N_17190,N_17286);
or U17633 (N_17633,N_17360,N_16947);
nor U17634 (N_17634,N_17096,N_16923);
and U17635 (N_17635,N_17074,N_17161);
xor U17636 (N_17636,N_17338,N_17357);
nor U17637 (N_17637,N_17288,N_17033);
nand U17638 (N_17638,N_17076,N_17058);
or U17639 (N_17639,N_17274,N_17166);
and U17640 (N_17640,N_17398,N_17047);
nand U17641 (N_17641,N_17165,N_16863);
or U17642 (N_17642,N_16867,N_17182);
nor U17643 (N_17643,N_17222,N_17126);
xnor U17644 (N_17644,N_17089,N_17065);
or U17645 (N_17645,N_17114,N_16981);
nand U17646 (N_17646,N_17332,N_16874);
nor U17647 (N_17647,N_16946,N_17196);
and U17648 (N_17648,N_16869,N_17206);
nor U17649 (N_17649,N_17098,N_17358);
nand U17650 (N_17650,N_17329,N_16885);
nor U17651 (N_17651,N_16820,N_16987);
nor U17652 (N_17652,N_16958,N_17265);
xor U17653 (N_17653,N_16906,N_16979);
xor U17654 (N_17654,N_17063,N_16971);
and U17655 (N_17655,N_17320,N_17362);
or U17656 (N_17656,N_16807,N_17382);
nor U17657 (N_17657,N_17073,N_17176);
xnor U17658 (N_17658,N_17131,N_17134);
and U17659 (N_17659,N_16925,N_17393);
or U17660 (N_17660,N_17256,N_16977);
or U17661 (N_17661,N_17355,N_17322);
or U17662 (N_17662,N_17289,N_17267);
or U17663 (N_17663,N_17142,N_17210);
or U17664 (N_17664,N_16821,N_17375);
nand U17665 (N_17665,N_17367,N_16900);
nor U17666 (N_17666,N_17369,N_17091);
or U17667 (N_17667,N_16819,N_16835);
and U17668 (N_17668,N_17253,N_17037);
nand U17669 (N_17669,N_17297,N_16990);
or U17670 (N_17670,N_17043,N_16846);
nor U17671 (N_17671,N_17029,N_17264);
nand U17672 (N_17672,N_17048,N_17094);
nand U17673 (N_17673,N_17216,N_17330);
xor U17674 (N_17674,N_17071,N_17172);
nor U17675 (N_17675,N_16994,N_17228);
nor U17676 (N_17676,N_16894,N_17147);
or U17677 (N_17677,N_17015,N_16960);
nor U17678 (N_17678,N_17138,N_17195);
or U17679 (N_17679,N_16956,N_16823);
and U17680 (N_17680,N_17324,N_17303);
nor U17681 (N_17681,N_17258,N_16850);
nor U17682 (N_17682,N_17378,N_17157);
nand U17683 (N_17683,N_17154,N_17315);
nand U17684 (N_17684,N_17087,N_17042);
nor U17685 (N_17685,N_16815,N_17323);
nor U17686 (N_17686,N_17181,N_16845);
nand U17687 (N_17687,N_17179,N_16818);
or U17688 (N_17688,N_17277,N_17054);
or U17689 (N_17689,N_17175,N_17061);
nor U17690 (N_17690,N_16975,N_17354);
or U17691 (N_17691,N_17292,N_16803);
or U17692 (N_17692,N_17145,N_17346);
nand U17693 (N_17693,N_16944,N_17086);
and U17694 (N_17694,N_16952,N_17168);
and U17695 (N_17695,N_17262,N_16978);
nand U17696 (N_17696,N_17192,N_17305);
xnor U17697 (N_17697,N_17370,N_16912);
nor U17698 (N_17698,N_16976,N_17260);
xor U17699 (N_17699,N_17028,N_16938);
xor U17700 (N_17700,N_16854,N_16837);
xor U17701 (N_17701,N_17144,N_17220);
xnor U17702 (N_17702,N_17262,N_17156);
or U17703 (N_17703,N_17184,N_17109);
nor U17704 (N_17704,N_17205,N_17012);
xor U17705 (N_17705,N_17124,N_16865);
nand U17706 (N_17706,N_17225,N_17363);
nand U17707 (N_17707,N_16801,N_17021);
and U17708 (N_17708,N_16804,N_17139);
or U17709 (N_17709,N_17261,N_16803);
nand U17710 (N_17710,N_16865,N_16802);
and U17711 (N_17711,N_17224,N_17167);
and U17712 (N_17712,N_17198,N_17060);
xor U17713 (N_17713,N_17195,N_17051);
and U17714 (N_17714,N_16805,N_16948);
nand U17715 (N_17715,N_17193,N_17342);
or U17716 (N_17716,N_17329,N_17248);
nor U17717 (N_17717,N_16991,N_17005);
and U17718 (N_17718,N_17108,N_17201);
nand U17719 (N_17719,N_16911,N_16822);
nor U17720 (N_17720,N_17316,N_16862);
nand U17721 (N_17721,N_17036,N_17015);
and U17722 (N_17722,N_16890,N_16888);
or U17723 (N_17723,N_16963,N_16948);
and U17724 (N_17724,N_17373,N_17374);
nor U17725 (N_17725,N_17235,N_16848);
and U17726 (N_17726,N_16906,N_16973);
or U17727 (N_17727,N_17317,N_16952);
or U17728 (N_17728,N_16969,N_16952);
xnor U17729 (N_17729,N_16807,N_17243);
nand U17730 (N_17730,N_16993,N_17036);
xor U17731 (N_17731,N_17365,N_16844);
xor U17732 (N_17732,N_17308,N_16977);
and U17733 (N_17733,N_16953,N_17287);
nand U17734 (N_17734,N_17251,N_17248);
or U17735 (N_17735,N_17123,N_17023);
nor U17736 (N_17736,N_17162,N_16876);
nor U17737 (N_17737,N_16936,N_16917);
xnor U17738 (N_17738,N_16847,N_17170);
nor U17739 (N_17739,N_17320,N_16980);
nor U17740 (N_17740,N_17102,N_17049);
nand U17741 (N_17741,N_17377,N_17261);
nand U17742 (N_17742,N_17049,N_16854);
or U17743 (N_17743,N_17304,N_17137);
nor U17744 (N_17744,N_17054,N_17306);
and U17745 (N_17745,N_17398,N_16875);
nand U17746 (N_17746,N_17308,N_17296);
nand U17747 (N_17747,N_17285,N_17366);
or U17748 (N_17748,N_17158,N_17310);
nand U17749 (N_17749,N_16890,N_16859);
xnor U17750 (N_17750,N_17103,N_16840);
xor U17751 (N_17751,N_16811,N_17058);
or U17752 (N_17752,N_17342,N_17235);
or U17753 (N_17753,N_17239,N_16877);
and U17754 (N_17754,N_16931,N_17347);
xor U17755 (N_17755,N_16869,N_16802);
nor U17756 (N_17756,N_16876,N_17278);
and U17757 (N_17757,N_16926,N_17184);
nand U17758 (N_17758,N_17048,N_17068);
xnor U17759 (N_17759,N_16929,N_16893);
xnor U17760 (N_17760,N_16871,N_17382);
and U17761 (N_17761,N_17024,N_17325);
or U17762 (N_17762,N_17086,N_17247);
xnor U17763 (N_17763,N_17268,N_16879);
and U17764 (N_17764,N_16889,N_16930);
xor U17765 (N_17765,N_16938,N_17294);
xor U17766 (N_17766,N_17267,N_17333);
nor U17767 (N_17767,N_16823,N_17094);
and U17768 (N_17768,N_17108,N_16832);
or U17769 (N_17769,N_16919,N_17208);
nand U17770 (N_17770,N_17269,N_17320);
xnor U17771 (N_17771,N_17061,N_17382);
or U17772 (N_17772,N_17014,N_16902);
or U17773 (N_17773,N_17102,N_17081);
nand U17774 (N_17774,N_17213,N_16940);
nand U17775 (N_17775,N_16997,N_17023);
nor U17776 (N_17776,N_17073,N_17145);
or U17777 (N_17777,N_17010,N_17134);
nor U17778 (N_17778,N_17370,N_16832);
nor U17779 (N_17779,N_16921,N_17387);
nand U17780 (N_17780,N_17306,N_17007);
and U17781 (N_17781,N_17200,N_17095);
xnor U17782 (N_17782,N_16885,N_16811);
or U17783 (N_17783,N_17087,N_16970);
xnor U17784 (N_17784,N_16975,N_17089);
nor U17785 (N_17785,N_16937,N_17202);
and U17786 (N_17786,N_17028,N_17081);
and U17787 (N_17787,N_16803,N_17204);
nor U17788 (N_17788,N_16803,N_17233);
or U17789 (N_17789,N_16864,N_16930);
xnor U17790 (N_17790,N_16830,N_17084);
nor U17791 (N_17791,N_16910,N_17147);
nand U17792 (N_17792,N_17081,N_17334);
or U17793 (N_17793,N_17207,N_16977);
or U17794 (N_17794,N_17156,N_17067);
and U17795 (N_17795,N_17087,N_16804);
nor U17796 (N_17796,N_16894,N_16846);
xnor U17797 (N_17797,N_17153,N_16859);
xnor U17798 (N_17798,N_17112,N_16973);
nand U17799 (N_17799,N_16839,N_16876);
nor U17800 (N_17800,N_17028,N_17002);
xor U17801 (N_17801,N_16933,N_16833);
xor U17802 (N_17802,N_17080,N_17344);
nor U17803 (N_17803,N_16860,N_16894);
nand U17804 (N_17804,N_17028,N_17183);
or U17805 (N_17805,N_16910,N_16848);
xnor U17806 (N_17806,N_17370,N_17187);
xnor U17807 (N_17807,N_17289,N_17183);
and U17808 (N_17808,N_17276,N_17090);
nand U17809 (N_17809,N_17064,N_17164);
xor U17810 (N_17810,N_17100,N_16998);
or U17811 (N_17811,N_16877,N_16921);
nor U17812 (N_17812,N_17351,N_17146);
nor U17813 (N_17813,N_17352,N_17118);
nand U17814 (N_17814,N_17110,N_17096);
and U17815 (N_17815,N_17229,N_16843);
and U17816 (N_17816,N_16833,N_16944);
or U17817 (N_17817,N_17289,N_17016);
xnor U17818 (N_17818,N_17042,N_16928);
xor U17819 (N_17819,N_17292,N_16860);
or U17820 (N_17820,N_17226,N_17387);
nor U17821 (N_17821,N_16841,N_17360);
nor U17822 (N_17822,N_17116,N_17148);
nor U17823 (N_17823,N_16836,N_17333);
or U17824 (N_17824,N_17351,N_17167);
nand U17825 (N_17825,N_16951,N_16914);
nor U17826 (N_17826,N_16956,N_17012);
and U17827 (N_17827,N_16915,N_16955);
xor U17828 (N_17828,N_16804,N_17227);
xor U17829 (N_17829,N_17371,N_16956);
nand U17830 (N_17830,N_17306,N_17195);
and U17831 (N_17831,N_17095,N_16812);
nor U17832 (N_17832,N_17297,N_17164);
nand U17833 (N_17833,N_16966,N_17248);
nor U17834 (N_17834,N_17054,N_16969);
or U17835 (N_17835,N_17278,N_17170);
or U17836 (N_17836,N_17201,N_16952);
nand U17837 (N_17837,N_16906,N_16881);
nor U17838 (N_17838,N_17218,N_17393);
xor U17839 (N_17839,N_17150,N_17324);
and U17840 (N_17840,N_16868,N_16907);
xnor U17841 (N_17841,N_17175,N_17378);
nor U17842 (N_17842,N_17156,N_17010);
nand U17843 (N_17843,N_17358,N_16926);
nor U17844 (N_17844,N_16852,N_17022);
nand U17845 (N_17845,N_17038,N_17012);
and U17846 (N_17846,N_17397,N_17126);
xnor U17847 (N_17847,N_17194,N_17276);
or U17848 (N_17848,N_16850,N_17180);
and U17849 (N_17849,N_17213,N_16837);
and U17850 (N_17850,N_16993,N_17366);
or U17851 (N_17851,N_16991,N_17050);
nand U17852 (N_17852,N_17312,N_17274);
nand U17853 (N_17853,N_17306,N_17290);
and U17854 (N_17854,N_17342,N_17256);
and U17855 (N_17855,N_16839,N_17307);
nand U17856 (N_17856,N_17024,N_17187);
nor U17857 (N_17857,N_17226,N_17347);
xor U17858 (N_17858,N_16960,N_17053);
xnor U17859 (N_17859,N_17011,N_17100);
nand U17860 (N_17860,N_17278,N_16974);
or U17861 (N_17861,N_16891,N_17096);
nor U17862 (N_17862,N_17336,N_17014);
or U17863 (N_17863,N_17215,N_16948);
xor U17864 (N_17864,N_17166,N_17029);
nand U17865 (N_17865,N_17128,N_17016);
or U17866 (N_17866,N_17166,N_17125);
or U17867 (N_17867,N_17083,N_17318);
nor U17868 (N_17868,N_17010,N_17072);
xnor U17869 (N_17869,N_16874,N_16870);
nor U17870 (N_17870,N_17392,N_17255);
nor U17871 (N_17871,N_17026,N_17179);
xnor U17872 (N_17872,N_17349,N_16970);
and U17873 (N_17873,N_16986,N_16918);
or U17874 (N_17874,N_17241,N_17275);
xor U17875 (N_17875,N_16824,N_17025);
xor U17876 (N_17876,N_17378,N_16932);
xnor U17877 (N_17877,N_17360,N_17209);
and U17878 (N_17878,N_17279,N_17182);
and U17879 (N_17879,N_17034,N_17232);
xor U17880 (N_17880,N_17261,N_17382);
and U17881 (N_17881,N_16882,N_17013);
and U17882 (N_17882,N_17330,N_16844);
or U17883 (N_17883,N_17143,N_17293);
xnor U17884 (N_17884,N_16990,N_16828);
xor U17885 (N_17885,N_17150,N_17291);
or U17886 (N_17886,N_17053,N_17165);
nor U17887 (N_17887,N_17382,N_17011);
xnor U17888 (N_17888,N_17341,N_16956);
or U17889 (N_17889,N_17031,N_17168);
and U17890 (N_17890,N_16870,N_16806);
nor U17891 (N_17891,N_16920,N_16914);
nand U17892 (N_17892,N_16826,N_17058);
xor U17893 (N_17893,N_17349,N_16824);
nor U17894 (N_17894,N_17111,N_16857);
nor U17895 (N_17895,N_17255,N_16975);
xor U17896 (N_17896,N_16824,N_17052);
xnor U17897 (N_17897,N_17106,N_16804);
nand U17898 (N_17898,N_16913,N_16876);
xor U17899 (N_17899,N_17189,N_17253);
nand U17900 (N_17900,N_16904,N_17188);
and U17901 (N_17901,N_17120,N_17046);
nand U17902 (N_17902,N_17016,N_17091);
or U17903 (N_17903,N_16820,N_16902);
nor U17904 (N_17904,N_16973,N_16904);
nand U17905 (N_17905,N_16863,N_17041);
nand U17906 (N_17906,N_16974,N_16880);
and U17907 (N_17907,N_16977,N_17036);
and U17908 (N_17908,N_16914,N_17243);
and U17909 (N_17909,N_16973,N_16901);
nor U17910 (N_17910,N_17007,N_17292);
and U17911 (N_17911,N_17144,N_17213);
nor U17912 (N_17912,N_16921,N_17344);
and U17913 (N_17913,N_17110,N_17060);
xnor U17914 (N_17914,N_17127,N_17025);
and U17915 (N_17915,N_17042,N_17222);
nor U17916 (N_17916,N_17333,N_17004);
nor U17917 (N_17917,N_17318,N_17030);
and U17918 (N_17918,N_17045,N_17218);
xnor U17919 (N_17919,N_17036,N_17017);
and U17920 (N_17920,N_17305,N_16991);
xor U17921 (N_17921,N_17233,N_17039);
nor U17922 (N_17922,N_17137,N_16813);
nor U17923 (N_17923,N_17130,N_17123);
xor U17924 (N_17924,N_17312,N_16817);
xnor U17925 (N_17925,N_17301,N_17361);
xor U17926 (N_17926,N_17170,N_17046);
or U17927 (N_17927,N_16884,N_17080);
and U17928 (N_17928,N_17313,N_16899);
nand U17929 (N_17929,N_17319,N_16804);
nor U17930 (N_17930,N_16860,N_17260);
xor U17931 (N_17931,N_17181,N_16901);
or U17932 (N_17932,N_17013,N_17360);
or U17933 (N_17933,N_16976,N_16971);
xor U17934 (N_17934,N_17178,N_17187);
xor U17935 (N_17935,N_16933,N_17229);
xor U17936 (N_17936,N_17264,N_17173);
xnor U17937 (N_17937,N_17237,N_17380);
and U17938 (N_17938,N_17022,N_17345);
nand U17939 (N_17939,N_16823,N_17326);
nor U17940 (N_17940,N_17049,N_17084);
or U17941 (N_17941,N_17266,N_16812);
and U17942 (N_17942,N_17026,N_17068);
nor U17943 (N_17943,N_17284,N_17032);
or U17944 (N_17944,N_17243,N_16814);
nor U17945 (N_17945,N_16827,N_17326);
and U17946 (N_17946,N_17303,N_16892);
xor U17947 (N_17947,N_17073,N_17173);
nor U17948 (N_17948,N_17060,N_16847);
or U17949 (N_17949,N_17328,N_17058);
and U17950 (N_17950,N_17188,N_16960);
nor U17951 (N_17951,N_17370,N_17295);
nand U17952 (N_17952,N_17041,N_16952);
nor U17953 (N_17953,N_16947,N_17375);
xnor U17954 (N_17954,N_16984,N_16832);
or U17955 (N_17955,N_16898,N_17056);
or U17956 (N_17956,N_17066,N_16991);
xnor U17957 (N_17957,N_17215,N_16830);
nor U17958 (N_17958,N_16826,N_16917);
nand U17959 (N_17959,N_16912,N_17237);
xnor U17960 (N_17960,N_17399,N_17395);
and U17961 (N_17961,N_17072,N_16865);
or U17962 (N_17962,N_17353,N_17397);
nor U17963 (N_17963,N_17159,N_17183);
and U17964 (N_17964,N_17374,N_17343);
nor U17965 (N_17965,N_17228,N_17363);
nor U17966 (N_17966,N_17075,N_17129);
and U17967 (N_17967,N_17116,N_16913);
and U17968 (N_17968,N_17118,N_17181);
and U17969 (N_17969,N_16826,N_17082);
xnor U17970 (N_17970,N_17079,N_17083);
or U17971 (N_17971,N_16842,N_16805);
nand U17972 (N_17972,N_17103,N_17388);
nor U17973 (N_17973,N_17266,N_17278);
xor U17974 (N_17974,N_17138,N_16990);
and U17975 (N_17975,N_17058,N_16869);
xor U17976 (N_17976,N_16889,N_17067);
nor U17977 (N_17977,N_17292,N_17085);
nor U17978 (N_17978,N_16904,N_17241);
or U17979 (N_17979,N_17009,N_17149);
or U17980 (N_17980,N_16903,N_17270);
and U17981 (N_17981,N_17241,N_16934);
nor U17982 (N_17982,N_17302,N_16900);
nand U17983 (N_17983,N_16813,N_17373);
or U17984 (N_17984,N_17062,N_17084);
nor U17985 (N_17985,N_17247,N_17191);
and U17986 (N_17986,N_17038,N_17067);
and U17987 (N_17987,N_17389,N_16880);
xor U17988 (N_17988,N_16880,N_17112);
nand U17989 (N_17989,N_17200,N_17069);
nand U17990 (N_17990,N_16916,N_16954);
xnor U17991 (N_17991,N_16968,N_17117);
or U17992 (N_17992,N_17182,N_17025);
xnor U17993 (N_17993,N_16874,N_17011);
nand U17994 (N_17994,N_16861,N_16978);
xor U17995 (N_17995,N_17362,N_16908);
nor U17996 (N_17996,N_17205,N_16953);
nor U17997 (N_17997,N_16983,N_16900);
and U17998 (N_17998,N_17307,N_17235);
nand U17999 (N_17999,N_16856,N_17207);
or U18000 (N_18000,N_17850,N_17459);
and U18001 (N_18001,N_17609,N_17889);
and U18002 (N_18002,N_17864,N_17467);
xor U18003 (N_18003,N_17684,N_17464);
nor U18004 (N_18004,N_17800,N_17765);
nor U18005 (N_18005,N_17652,N_17469);
and U18006 (N_18006,N_17404,N_17967);
nor U18007 (N_18007,N_17568,N_17754);
nor U18008 (N_18008,N_17851,N_17852);
and U18009 (N_18009,N_17751,N_17854);
nand U18010 (N_18010,N_17816,N_17458);
xnor U18011 (N_18011,N_17735,N_17588);
nand U18012 (N_18012,N_17874,N_17471);
or U18013 (N_18013,N_17927,N_17463);
xor U18014 (N_18014,N_17779,N_17837);
nand U18015 (N_18015,N_17466,N_17758);
nor U18016 (N_18016,N_17631,N_17776);
nor U18017 (N_18017,N_17741,N_17576);
xnor U18018 (N_18018,N_17481,N_17785);
nor U18019 (N_18019,N_17830,N_17728);
or U18020 (N_18020,N_17766,N_17817);
xnor U18021 (N_18021,N_17629,N_17422);
xnor U18022 (N_18022,N_17493,N_17418);
nor U18023 (N_18023,N_17675,N_17944);
xnor U18024 (N_18024,N_17999,N_17801);
xnor U18025 (N_18025,N_17718,N_17863);
nor U18026 (N_18026,N_17616,N_17527);
xor U18027 (N_18027,N_17604,N_17945);
xor U18028 (N_18028,N_17487,N_17884);
xor U18029 (N_18029,N_17804,N_17678);
or U18030 (N_18030,N_17737,N_17662);
nand U18031 (N_18031,N_17748,N_17460);
xor U18032 (N_18032,N_17904,N_17794);
or U18033 (N_18033,N_17842,N_17554);
xnor U18034 (N_18034,N_17465,N_17462);
and U18035 (N_18035,N_17613,N_17950);
or U18036 (N_18036,N_17755,N_17611);
and U18037 (N_18037,N_17571,N_17709);
nor U18038 (N_18038,N_17557,N_17690);
nand U18039 (N_18039,N_17507,N_17476);
nand U18040 (N_18040,N_17529,N_17639);
xnor U18041 (N_18041,N_17905,N_17743);
nor U18042 (N_18042,N_17907,N_17440);
nor U18043 (N_18043,N_17583,N_17562);
xor U18044 (N_18044,N_17663,N_17723);
or U18045 (N_18045,N_17667,N_17856);
nor U18046 (N_18046,N_17516,N_17964);
nor U18047 (N_18047,N_17757,N_17977);
xor U18048 (N_18048,N_17888,N_17902);
nor U18049 (N_18049,N_17602,N_17485);
nand U18050 (N_18050,N_17506,N_17897);
xor U18051 (N_18051,N_17406,N_17607);
xor U18052 (N_18052,N_17490,N_17798);
xnor U18053 (N_18053,N_17915,N_17929);
or U18054 (N_18054,N_17879,N_17574);
nand U18055 (N_18055,N_17722,N_17784);
or U18056 (N_18056,N_17677,N_17447);
nand U18057 (N_18057,N_17858,N_17657);
or U18058 (N_18058,N_17505,N_17708);
nor U18059 (N_18059,N_17513,N_17720);
and U18060 (N_18060,N_17514,N_17425);
or U18061 (N_18061,N_17787,N_17530);
and U18062 (N_18062,N_17873,N_17986);
nand U18063 (N_18063,N_17764,N_17700);
xnor U18064 (N_18064,N_17955,N_17760);
or U18065 (N_18065,N_17893,N_17815);
nand U18066 (N_18066,N_17685,N_17540);
nand U18067 (N_18067,N_17747,N_17970);
xnor U18068 (N_18068,N_17402,N_17991);
nor U18069 (N_18069,N_17846,N_17622);
and U18070 (N_18070,N_17995,N_17957);
nand U18071 (N_18071,N_17564,N_17729);
xnor U18072 (N_18072,N_17865,N_17563);
or U18073 (N_18073,N_17809,N_17962);
xnor U18074 (N_18074,N_17472,N_17810);
or U18075 (N_18075,N_17828,N_17732);
xor U18076 (N_18076,N_17625,N_17772);
nand U18077 (N_18077,N_17570,N_17695);
or U18078 (N_18078,N_17844,N_17792);
or U18079 (N_18079,N_17827,N_17612);
and U18080 (N_18080,N_17831,N_17648);
xnor U18081 (N_18081,N_17468,N_17618);
and U18082 (N_18082,N_17849,N_17566);
xnor U18083 (N_18083,N_17871,N_17585);
nor U18084 (N_18084,N_17681,N_17870);
and U18085 (N_18085,N_17666,N_17532);
nand U18086 (N_18086,N_17705,N_17594);
xor U18087 (N_18087,N_17496,N_17998);
nand U18088 (N_18088,N_17932,N_17595);
and U18089 (N_18089,N_17716,N_17813);
nand U18090 (N_18090,N_17994,N_17836);
and U18091 (N_18091,N_17670,N_17692);
xnor U18092 (N_18092,N_17452,N_17433);
and U18093 (N_18093,N_17548,N_17510);
nand U18094 (N_18094,N_17908,N_17711);
or U18095 (N_18095,N_17996,N_17664);
and U18096 (N_18096,N_17619,N_17937);
nor U18097 (N_18097,N_17742,N_17446);
xnor U18098 (N_18098,N_17824,N_17508);
nor U18099 (N_18099,N_17650,N_17974);
or U18100 (N_18100,N_17579,N_17761);
xor U18101 (N_18101,N_17546,N_17895);
nor U18102 (N_18102,N_17428,N_17598);
xnor U18103 (N_18103,N_17948,N_17811);
or U18104 (N_18104,N_17614,N_17959);
and U18105 (N_18105,N_17917,N_17878);
nor U18106 (N_18106,N_17597,N_17832);
or U18107 (N_18107,N_17649,N_17615);
and U18108 (N_18108,N_17968,N_17414);
nor U18109 (N_18109,N_17825,N_17829);
xor U18110 (N_18110,N_17504,N_17424);
and U18111 (N_18111,N_17682,N_17925);
nor U18112 (N_18112,N_17478,N_17980);
nand U18113 (N_18113,N_17972,N_17483);
nand U18114 (N_18114,N_17599,N_17545);
and U18115 (N_18115,N_17627,N_17531);
and U18116 (N_18116,N_17580,N_17866);
nor U18117 (N_18117,N_17543,N_17555);
xnor U18118 (N_18118,N_17450,N_17638);
nand U18119 (N_18119,N_17790,N_17489);
nor U18120 (N_18120,N_17587,N_17525);
nor U18121 (N_18121,N_17926,N_17763);
nand U18122 (N_18122,N_17988,N_17606);
xnor U18123 (N_18123,N_17634,N_17872);
nor U18124 (N_18124,N_17412,N_17973);
and U18125 (N_18125,N_17600,N_17444);
nor U18126 (N_18126,N_17492,N_17821);
nand U18127 (N_18127,N_17845,N_17714);
nand U18128 (N_18128,N_17470,N_17788);
or U18129 (N_18129,N_17647,N_17807);
nor U18130 (N_18130,N_17891,N_17669);
nor U18131 (N_18131,N_17573,N_17408);
xnor U18132 (N_18132,N_17538,N_17738);
nor U18133 (N_18133,N_17498,N_17750);
and U18134 (N_18134,N_17910,N_17411);
nand U18135 (N_18135,N_17936,N_17969);
nor U18136 (N_18136,N_17985,N_17620);
and U18137 (N_18137,N_17861,N_17782);
and U18138 (N_18138,N_17847,N_17783);
or U18139 (N_18139,N_17710,N_17997);
or U18140 (N_18140,N_17819,N_17803);
xnor U18141 (N_18141,N_17731,N_17486);
nand U18142 (N_18142,N_17642,N_17961);
xor U18143 (N_18143,N_17644,N_17943);
or U18144 (N_18144,N_17952,N_17423);
xor U18145 (N_18145,N_17537,N_17437);
or U18146 (N_18146,N_17439,N_17436);
nand U18147 (N_18147,N_17777,N_17448);
nand U18148 (N_18148,N_17651,N_17975);
and U18149 (N_18149,N_17558,N_17536);
nand U18150 (N_18150,N_17886,N_17859);
nor U18151 (N_18151,N_17429,N_17517);
or U18152 (N_18152,N_17660,N_17591);
xnor U18153 (N_18153,N_17706,N_17963);
and U18154 (N_18154,N_17880,N_17500);
nand U18155 (N_18155,N_17628,N_17415);
xnor U18156 (N_18156,N_17430,N_17590);
or U18157 (N_18157,N_17656,N_17432);
nand U18158 (N_18158,N_17547,N_17928);
or U18159 (N_18159,N_17935,N_17778);
xnor U18160 (N_18160,N_17417,N_17984);
nor U18161 (N_18161,N_17694,N_17713);
and U18162 (N_18162,N_17551,N_17549);
xor U18163 (N_18163,N_17409,N_17671);
nand U18164 (N_18164,N_17686,N_17981);
or U18165 (N_18165,N_17443,N_17427);
nor U18166 (N_18166,N_17894,N_17941);
xnor U18167 (N_18167,N_17877,N_17900);
and U18168 (N_18168,N_17702,N_17982);
xor U18169 (N_18169,N_17835,N_17746);
or U18170 (N_18170,N_17903,N_17942);
nor U18171 (N_18171,N_17535,N_17561);
and U18172 (N_18172,N_17449,N_17689);
or U18173 (N_18173,N_17916,N_17626);
or U18174 (N_18174,N_17518,N_17703);
nor U18175 (N_18175,N_17501,N_17774);
nor U18176 (N_18176,N_17410,N_17477);
and U18177 (N_18177,N_17473,N_17655);
nor U18178 (N_18178,N_17539,N_17826);
nand U18179 (N_18179,N_17739,N_17976);
or U18180 (N_18180,N_17645,N_17938);
and U18181 (N_18181,N_17721,N_17608);
nor U18182 (N_18182,N_17680,N_17767);
xnor U18183 (N_18183,N_17914,N_17913);
xor U18184 (N_18184,N_17693,N_17931);
or U18185 (N_18185,N_17793,N_17623);
and U18186 (N_18186,N_17876,N_17899);
and U18187 (N_18187,N_17795,N_17491);
xor U18188 (N_18188,N_17733,N_17726);
or U18189 (N_18189,N_17812,N_17841);
nor U18190 (N_18190,N_17853,N_17636);
or U18191 (N_18191,N_17808,N_17673);
or U18192 (N_18192,N_17701,N_17992);
xnor U18193 (N_18193,N_17930,N_17533);
or U18194 (N_18194,N_17920,N_17960);
and U18195 (N_18195,N_17691,N_17883);
xnor U18196 (N_18196,N_17567,N_17781);
xor U18197 (N_18197,N_17715,N_17947);
nor U18198 (N_18198,N_17400,N_17584);
nor U18199 (N_18199,N_17727,N_17730);
nand U18200 (N_18200,N_17896,N_17416);
nor U18201 (N_18201,N_17882,N_17683);
or U18202 (N_18202,N_17451,N_17640);
nand U18203 (N_18203,N_17993,N_17820);
nor U18204 (N_18204,N_17654,N_17637);
nor U18205 (N_18205,N_17407,N_17577);
and U18206 (N_18206,N_17823,N_17770);
nor U18207 (N_18207,N_17524,N_17522);
or U18208 (N_18208,N_17867,N_17441);
xor U18209 (N_18209,N_17707,N_17834);
or U18210 (N_18210,N_17887,N_17966);
nand U18211 (N_18211,N_17635,N_17454);
nor U18212 (N_18212,N_17668,N_17419);
nand U18213 (N_18213,N_17565,N_17946);
or U18214 (N_18214,N_17717,N_17617);
xnor U18215 (N_18215,N_17814,N_17901);
xor U18216 (N_18216,N_17661,N_17934);
nor U18217 (N_18217,N_17818,N_17641);
xnor U18218 (N_18218,N_17923,N_17484);
and U18219 (N_18219,N_17768,N_17749);
nand U18220 (N_18220,N_17744,N_17575);
and U18221 (N_18221,N_17633,N_17475);
or U18222 (N_18222,N_17875,N_17541);
or U18223 (N_18223,N_17939,N_17653);
nand U18224 (N_18224,N_17796,N_17840);
and U18225 (N_18225,N_17621,N_17499);
nor U18226 (N_18226,N_17593,N_17456);
nand U18227 (N_18227,N_17919,N_17520);
and U18228 (N_18228,N_17990,N_17698);
or U18229 (N_18229,N_17552,N_17885);
nor U18230 (N_18230,N_17578,N_17658);
and U18231 (N_18231,N_17519,N_17509);
nor U18232 (N_18232,N_17855,N_17924);
or U18233 (N_18233,N_17949,N_17860);
nand U18234 (N_18234,N_17989,N_17665);
or U18235 (N_18235,N_17775,N_17933);
xor U18236 (N_18236,N_17951,N_17838);
or U18237 (N_18237,N_17773,N_17646);
nor U18238 (N_18238,N_17488,N_17403);
or U18239 (N_18239,N_17906,N_17769);
or U18240 (N_18240,N_17956,N_17632);
xor U18241 (N_18241,N_17474,N_17921);
and U18242 (N_18242,N_17759,N_17445);
or U18243 (N_18243,N_17753,N_17797);
or U18244 (N_18244,N_17869,N_17589);
nand U18245 (N_18245,N_17553,N_17405);
and U18246 (N_18246,N_17596,N_17572);
xnor U18247 (N_18247,N_17434,N_17442);
xnor U18248 (N_18248,N_17605,N_17712);
and U18249 (N_18249,N_17401,N_17786);
nand U18250 (N_18250,N_17457,N_17953);
or U18251 (N_18251,N_17780,N_17542);
and U18252 (N_18252,N_17526,N_17512);
or U18253 (N_18253,N_17892,N_17862);
nand U18254 (N_18254,N_17745,N_17581);
or U18255 (N_18255,N_17719,N_17610);
nor U18256 (N_18256,N_17724,N_17630);
and U18257 (N_18257,N_17979,N_17586);
nor U18258 (N_18258,N_17453,N_17643);
and U18259 (N_18259,N_17503,N_17762);
nand U18260 (N_18260,N_17592,N_17550);
or U18261 (N_18261,N_17971,N_17676);
or U18262 (N_18262,N_17965,N_17479);
or U18263 (N_18263,N_17688,N_17461);
xor U18264 (N_18264,N_17697,N_17833);
nand U18265 (N_18265,N_17523,N_17848);
nand U18266 (N_18266,N_17560,N_17699);
and U18267 (N_18267,N_17413,N_17898);
or U18268 (N_18268,N_17674,N_17421);
nor U18269 (N_18269,N_17431,N_17881);
nor U18270 (N_18270,N_17511,N_17789);
xnor U18271 (N_18271,N_17958,N_17799);
and U18272 (N_18272,N_17559,N_17704);
or U18273 (N_18273,N_17791,N_17515);
or U18274 (N_18274,N_17696,N_17556);
and U18275 (N_18275,N_17497,N_17494);
nand U18276 (N_18276,N_17659,N_17435);
xnor U18277 (N_18277,N_17909,N_17868);
or U18278 (N_18278,N_17534,N_17569);
and U18279 (N_18279,N_17954,N_17756);
or U18280 (N_18280,N_17912,N_17805);
and U18281 (N_18281,N_17802,N_17740);
nor U18282 (N_18282,N_17734,N_17480);
and U18283 (N_18283,N_17420,N_17987);
and U18284 (N_18284,N_17672,N_17839);
xnor U18285 (N_18285,N_17822,N_17482);
nand U18286 (N_18286,N_17426,N_17725);
nand U18287 (N_18287,N_17983,N_17978);
nand U18288 (N_18288,N_17806,N_17918);
nor U18289 (N_18289,N_17857,N_17528);
xnor U18290 (N_18290,N_17544,N_17679);
nand U18291 (N_18291,N_17502,N_17603);
xnor U18292 (N_18292,N_17455,N_17911);
nor U18293 (N_18293,N_17922,N_17752);
nor U18294 (N_18294,N_17601,N_17624);
xnor U18295 (N_18295,N_17521,N_17495);
nand U18296 (N_18296,N_17843,N_17771);
and U18297 (N_18297,N_17890,N_17940);
nor U18298 (N_18298,N_17438,N_17582);
and U18299 (N_18299,N_17687,N_17736);
and U18300 (N_18300,N_17618,N_17421);
xnor U18301 (N_18301,N_17595,N_17706);
xnor U18302 (N_18302,N_17861,N_17499);
and U18303 (N_18303,N_17949,N_17812);
nor U18304 (N_18304,N_17976,N_17541);
and U18305 (N_18305,N_17445,N_17904);
nor U18306 (N_18306,N_17466,N_17707);
or U18307 (N_18307,N_17797,N_17675);
xor U18308 (N_18308,N_17496,N_17640);
and U18309 (N_18309,N_17959,N_17764);
nand U18310 (N_18310,N_17443,N_17852);
and U18311 (N_18311,N_17509,N_17932);
nor U18312 (N_18312,N_17610,N_17536);
nand U18313 (N_18313,N_17491,N_17600);
and U18314 (N_18314,N_17672,N_17675);
nand U18315 (N_18315,N_17761,N_17966);
or U18316 (N_18316,N_17422,N_17679);
xnor U18317 (N_18317,N_17980,N_17809);
or U18318 (N_18318,N_17798,N_17433);
and U18319 (N_18319,N_17437,N_17979);
nand U18320 (N_18320,N_17688,N_17774);
nand U18321 (N_18321,N_17996,N_17489);
nand U18322 (N_18322,N_17604,N_17876);
nand U18323 (N_18323,N_17831,N_17590);
xnor U18324 (N_18324,N_17632,N_17581);
xor U18325 (N_18325,N_17554,N_17980);
nor U18326 (N_18326,N_17422,N_17491);
xor U18327 (N_18327,N_17473,N_17591);
and U18328 (N_18328,N_17565,N_17438);
or U18329 (N_18329,N_17430,N_17906);
nand U18330 (N_18330,N_17541,N_17750);
and U18331 (N_18331,N_17419,N_17664);
and U18332 (N_18332,N_17584,N_17522);
or U18333 (N_18333,N_17499,N_17752);
and U18334 (N_18334,N_17522,N_17844);
or U18335 (N_18335,N_17669,N_17525);
nand U18336 (N_18336,N_17791,N_17621);
and U18337 (N_18337,N_17860,N_17962);
and U18338 (N_18338,N_17862,N_17660);
or U18339 (N_18339,N_17931,N_17541);
nand U18340 (N_18340,N_17559,N_17432);
or U18341 (N_18341,N_17955,N_17608);
and U18342 (N_18342,N_17650,N_17899);
or U18343 (N_18343,N_17741,N_17525);
xor U18344 (N_18344,N_17515,N_17672);
or U18345 (N_18345,N_17644,N_17510);
xor U18346 (N_18346,N_17428,N_17972);
and U18347 (N_18347,N_17473,N_17775);
and U18348 (N_18348,N_17669,N_17455);
and U18349 (N_18349,N_17442,N_17710);
or U18350 (N_18350,N_17696,N_17478);
nand U18351 (N_18351,N_17945,N_17990);
xnor U18352 (N_18352,N_17892,N_17846);
xnor U18353 (N_18353,N_17921,N_17868);
xor U18354 (N_18354,N_17605,N_17419);
nor U18355 (N_18355,N_17880,N_17570);
xor U18356 (N_18356,N_17578,N_17974);
or U18357 (N_18357,N_17943,N_17872);
nor U18358 (N_18358,N_17681,N_17714);
and U18359 (N_18359,N_17857,N_17570);
and U18360 (N_18360,N_17884,N_17430);
and U18361 (N_18361,N_17413,N_17621);
or U18362 (N_18362,N_17972,N_17870);
and U18363 (N_18363,N_17939,N_17484);
xor U18364 (N_18364,N_17403,N_17505);
nor U18365 (N_18365,N_17461,N_17925);
or U18366 (N_18366,N_17684,N_17500);
nand U18367 (N_18367,N_17860,N_17757);
xnor U18368 (N_18368,N_17471,N_17485);
and U18369 (N_18369,N_17809,N_17409);
xnor U18370 (N_18370,N_17757,N_17819);
nand U18371 (N_18371,N_17912,N_17436);
nor U18372 (N_18372,N_17909,N_17864);
xnor U18373 (N_18373,N_17586,N_17787);
nor U18374 (N_18374,N_17887,N_17572);
nor U18375 (N_18375,N_17514,N_17449);
xor U18376 (N_18376,N_17698,N_17473);
nand U18377 (N_18377,N_17897,N_17965);
or U18378 (N_18378,N_17927,N_17583);
xor U18379 (N_18379,N_17571,N_17969);
nor U18380 (N_18380,N_17989,N_17445);
nand U18381 (N_18381,N_17995,N_17837);
nand U18382 (N_18382,N_17801,N_17855);
nor U18383 (N_18383,N_17753,N_17749);
xnor U18384 (N_18384,N_17496,N_17555);
xnor U18385 (N_18385,N_17985,N_17948);
nor U18386 (N_18386,N_17948,N_17978);
xnor U18387 (N_18387,N_17425,N_17817);
or U18388 (N_18388,N_17866,N_17807);
and U18389 (N_18389,N_17486,N_17500);
and U18390 (N_18390,N_17639,N_17550);
or U18391 (N_18391,N_17641,N_17539);
and U18392 (N_18392,N_17411,N_17506);
nor U18393 (N_18393,N_17821,N_17668);
nand U18394 (N_18394,N_17516,N_17880);
xnor U18395 (N_18395,N_17506,N_17652);
nor U18396 (N_18396,N_17413,N_17436);
xnor U18397 (N_18397,N_17752,N_17637);
xnor U18398 (N_18398,N_17906,N_17607);
and U18399 (N_18399,N_17616,N_17656);
nor U18400 (N_18400,N_17520,N_17689);
or U18401 (N_18401,N_17490,N_17811);
or U18402 (N_18402,N_17563,N_17836);
xor U18403 (N_18403,N_17633,N_17680);
nand U18404 (N_18404,N_17919,N_17414);
or U18405 (N_18405,N_17954,N_17799);
nor U18406 (N_18406,N_17484,N_17410);
nand U18407 (N_18407,N_17633,N_17411);
nor U18408 (N_18408,N_17461,N_17901);
xnor U18409 (N_18409,N_17744,N_17976);
nor U18410 (N_18410,N_17819,N_17858);
nor U18411 (N_18411,N_17520,N_17882);
or U18412 (N_18412,N_17543,N_17826);
and U18413 (N_18413,N_17829,N_17465);
and U18414 (N_18414,N_17815,N_17983);
and U18415 (N_18415,N_17557,N_17742);
and U18416 (N_18416,N_17914,N_17569);
xor U18417 (N_18417,N_17492,N_17878);
nand U18418 (N_18418,N_17666,N_17744);
nand U18419 (N_18419,N_17551,N_17948);
nor U18420 (N_18420,N_17784,N_17918);
xor U18421 (N_18421,N_17807,N_17843);
and U18422 (N_18422,N_17675,N_17464);
nand U18423 (N_18423,N_17939,N_17935);
or U18424 (N_18424,N_17668,N_17509);
xor U18425 (N_18425,N_17558,N_17635);
nand U18426 (N_18426,N_17748,N_17688);
or U18427 (N_18427,N_17815,N_17615);
nor U18428 (N_18428,N_17810,N_17493);
or U18429 (N_18429,N_17833,N_17765);
xnor U18430 (N_18430,N_17458,N_17763);
and U18431 (N_18431,N_17880,N_17970);
or U18432 (N_18432,N_17422,N_17849);
and U18433 (N_18433,N_17619,N_17857);
nor U18434 (N_18434,N_17992,N_17849);
and U18435 (N_18435,N_17993,N_17551);
or U18436 (N_18436,N_17845,N_17479);
and U18437 (N_18437,N_17476,N_17448);
xor U18438 (N_18438,N_17428,N_17582);
nor U18439 (N_18439,N_17813,N_17911);
xnor U18440 (N_18440,N_17544,N_17825);
and U18441 (N_18441,N_17719,N_17718);
and U18442 (N_18442,N_17955,N_17898);
or U18443 (N_18443,N_17442,N_17745);
nor U18444 (N_18444,N_17752,N_17712);
and U18445 (N_18445,N_17822,N_17875);
nand U18446 (N_18446,N_17891,N_17687);
nor U18447 (N_18447,N_17433,N_17686);
and U18448 (N_18448,N_17757,N_17856);
nor U18449 (N_18449,N_17988,N_17738);
xor U18450 (N_18450,N_17912,N_17838);
or U18451 (N_18451,N_17788,N_17924);
or U18452 (N_18452,N_17740,N_17879);
or U18453 (N_18453,N_17465,N_17550);
xor U18454 (N_18454,N_17409,N_17829);
nor U18455 (N_18455,N_17979,N_17537);
or U18456 (N_18456,N_17542,N_17550);
nand U18457 (N_18457,N_17715,N_17732);
nor U18458 (N_18458,N_17468,N_17693);
xor U18459 (N_18459,N_17555,N_17663);
nor U18460 (N_18460,N_17720,N_17707);
nand U18461 (N_18461,N_17565,N_17623);
xor U18462 (N_18462,N_17997,N_17555);
and U18463 (N_18463,N_17494,N_17401);
nand U18464 (N_18464,N_17839,N_17854);
or U18465 (N_18465,N_17549,N_17521);
and U18466 (N_18466,N_17937,N_17492);
or U18467 (N_18467,N_17551,N_17758);
or U18468 (N_18468,N_17741,N_17809);
or U18469 (N_18469,N_17828,N_17986);
nor U18470 (N_18470,N_17657,N_17574);
nor U18471 (N_18471,N_17774,N_17837);
and U18472 (N_18472,N_17499,N_17935);
nand U18473 (N_18473,N_17650,N_17564);
or U18474 (N_18474,N_17814,N_17995);
or U18475 (N_18475,N_17674,N_17752);
xnor U18476 (N_18476,N_17607,N_17663);
xor U18477 (N_18477,N_17477,N_17409);
or U18478 (N_18478,N_17800,N_17640);
and U18479 (N_18479,N_17893,N_17684);
nand U18480 (N_18480,N_17459,N_17407);
nor U18481 (N_18481,N_17461,N_17672);
and U18482 (N_18482,N_17512,N_17590);
nand U18483 (N_18483,N_17589,N_17855);
and U18484 (N_18484,N_17875,N_17642);
nand U18485 (N_18485,N_17962,N_17628);
or U18486 (N_18486,N_17556,N_17825);
xor U18487 (N_18487,N_17819,N_17702);
xor U18488 (N_18488,N_17838,N_17941);
and U18489 (N_18489,N_17462,N_17575);
and U18490 (N_18490,N_17918,N_17809);
and U18491 (N_18491,N_17643,N_17867);
xor U18492 (N_18492,N_17799,N_17649);
nand U18493 (N_18493,N_17969,N_17720);
or U18494 (N_18494,N_17863,N_17503);
nor U18495 (N_18495,N_17487,N_17455);
or U18496 (N_18496,N_17875,N_17508);
xor U18497 (N_18497,N_17786,N_17778);
and U18498 (N_18498,N_17627,N_17602);
nor U18499 (N_18499,N_17722,N_17773);
nand U18500 (N_18500,N_17864,N_17862);
nand U18501 (N_18501,N_17463,N_17499);
xor U18502 (N_18502,N_17859,N_17468);
nor U18503 (N_18503,N_17993,N_17429);
nor U18504 (N_18504,N_17880,N_17837);
and U18505 (N_18505,N_17942,N_17856);
and U18506 (N_18506,N_17871,N_17798);
or U18507 (N_18507,N_17854,N_17679);
nand U18508 (N_18508,N_17516,N_17860);
or U18509 (N_18509,N_17954,N_17901);
and U18510 (N_18510,N_17694,N_17756);
or U18511 (N_18511,N_17431,N_17863);
xor U18512 (N_18512,N_17492,N_17610);
or U18513 (N_18513,N_17947,N_17589);
xor U18514 (N_18514,N_17691,N_17524);
or U18515 (N_18515,N_17558,N_17561);
nor U18516 (N_18516,N_17438,N_17634);
or U18517 (N_18517,N_17810,N_17424);
nand U18518 (N_18518,N_17464,N_17693);
xnor U18519 (N_18519,N_17480,N_17581);
nand U18520 (N_18520,N_17706,N_17797);
or U18521 (N_18521,N_17643,N_17717);
and U18522 (N_18522,N_17495,N_17868);
or U18523 (N_18523,N_17484,N_17472);
nor U18524 (N_18524,N_17487,N_17509);
or U18525 (N_18525,N_17996,N_17488);
and U18526 (N_18526,N_17976,N_17731);
xnor U18527 (N_18527,N_17661,N_17724);
nor U18528 (N_18528,N_17769,N_17833);
and U18529 (N_18529,N_17859,N_17773);
nor U18530 (N_18530,N_17671,N_17738);
or U18531 (N_18531,N_17623,N_17654);
and U18532 (N_18532,N_17664,N_17856);
and U18533 (N_18533,N_17746,N_17491);
nor U18534 (N_18534,N_17971,N_17667);
nor U18535 (N_18535,N_17994,N_17728);
nand U18536 (N_18536,N_17481,N_17531);
nor U18537 (N_18537,N_17848,N_17809);
and U18538 (N_18538,N_17969,N_17876);
or U18539 (N_18539,N_17792,N_17557);
nand U18540 (N_18540,N_17648,N_17649);
nand U18541 (N_18541,N_17401,N_17909);
nand U18542 (N_18542,N_17696,N_17714);
xnor U18543 (N_18543,N_17959,N_17821);
and U18544 (N_18544,N_17474,N_17941);
or U18545 (N_18545,N_17680,N_17759);
xnor U18546 (N_18546,N_17580,N_17718);
nand U18547 (N_18547,N_17889,N_17865);
or U18548 (N_18548,N_17951,N_17803);
nand U18549 (N_18549,N_17402,N_17577);
nand U18550 (N_18550,N_17501,N_17447);
and U18551 (N_18551,N_17720,N_17637);
or U18552 (N_18552,N_17543,N_17781);
and U18553 (N_18553,N_17401,N_17556);
or U18554 (N_18554,N_17816,N_17759);
and U18555 (N_18555,N_17668,N_17619);
xnor U18556 (N_18556,N_17433,N_17931);
nand U18557 (N_18557,N_17652,N_17853);
xor U18558 (N_18558,N_17813,N_17956);
and U18559 (N_18559,N_17468,N_17888);
and U18560 (N_18560,N_17998,N_17613);
nand U18561 (N_18561,N_17901,N_17914);
and U18562 (N_18562,N_17931,N_17777);
nor U18563 (N_18563,N_17708,N_17630);
and U18564 (N_18564,N_17684,N_17415);
and U18565 (N_18565,N_17976,N_17812);
or U18566 (N_18566,N_17491,N_17620);
and U18567 (N_18567,N_17546,N_17754);
nor U18568 (N_18568,N_17910,N_17429);
xnor U18569 (N_18569,N_17736,N_17427);
nand U18570 (N_18570,N_17863,N_17715);
or U18571 (N_18571,N_17432,N_17712);
and U18572 (N_18572,N_17776,N_17432);
and U18573 (N_18573,N_17561,N_17930);
and U18574 (N_18574,N_17481,N_17761);
and U18575 (N_18575,N_17975,N_17473);
and U18576 (N_18576,N_17452,N_17547);
or U18577 (N_18577,N_17730,N_17405);
nand U18578 (N_18578,N_17727,N_17946);
nor U18579 (N_18579,N_17927,N_17799);
nand U18580 (N_18580,N_17816,N_17792);
xor U18581 (N_18581,N_17944,N_17509);
xor U18582 (N_18582,N_17739,N_17929);
xnor U18583 (N_18583,N_17491,N_17538);
nor U18584 (N_18584,N_17640,N_17723);
nand U18585 (N_18585,N_17483,N_17619);
and U18586 (N_18586,N_17898,N_17852);
or U18587 (N_18587,N_17582,N_17947);
xor U18588 (N_18588,N_17793,N_17568);
nand U18589 (N_18589,N_17973,N_17414);
nor U18590 (N_18590,N_17871,N_17665);
nand U18591 (N_18591,N_17736,N_17802);
or U18592 (N_18592,N_17884,N_17410);
and U18593 (N_18593,N_17848,N_17869);
xnor U18594 (N_18594,N_17419,N_17934);
nor U18595 (N_18595,N_17875,N_17625);
or U18596 (N_18596,N_17623,N_17574);
xor U18597 (N_18597,N_17617,N_17983);
or U18598 (N_18598,N_17890,N_17630);
nor U18599 (N_18599,N_17568,N_17634);
and U18600 (N_18600,N_18564,N_18277);
xnor U18601 (N_18601,N_18334,N_18455);
nand U18602 (N_18602,N_18264,N_18388);
xor U18603 (N_18603,N_18020,N_18183);
nand U18604 (N_18604,N_18326,N_18384);
nand U18605 (N_18605,N_18092,N_18132);
or U18606 (N_18606,N_18109,N_18169);
and U18607 (N_18607,N_18454,N_18332);
xor U18608 (N_18608,N_18440,N_18337);
xnor U18609 (N_18609,N_18345,N_18483);
and U18610 (N_18610,N_18000,N_18140);
or U18611 (N_18611,N_18579,N_18193);
and U18612 (N_18612,N_18047,N_18517);
xnor U18613 (N_18613,N_18048,N_18422);
xnor U18614 (N_18614,N_18586,N_18199);
nand U18615 (N_18615,N_18236,N_18429);
and U18616 (N_18616,N_18534,N_18099);
and U18617 (N_18617,N_18465,N_18008);
nor U18618 (N_18618,N_18243,N_18363);
xnor U18619 (N_18619,N_18447,N_18211);
and U18620 (N_18620,N_18280,N_18542);
nand U18621 (N_18621,N_18073,N_18435);
or U18622 (N_18622,N_18516,N_18569);
and U18623 (N_18623,N_18197,N_18335);
xor U18624 (N_18624,N_18500,N_18387);
nand U18625 (N_18625,N_18214,N_18090);
or U18626 (N_18626,N_18595,N_18432);
and U18627 (N_18627,N_18568,N_18421);
nor U18628 (N_18628,N_18049,N_18240);
and U18629 (N_18629,N_18330,N_18368);
xor U18630 (N_18630,N_18472,N_18279);
xor U18631 (N_18631,N_18294,N_18081);
or U18632 (N_18632,N_18200,N_18573);
or U18633 (N_18633,N_18098,N_18307);
nand U18634 (N_18634,N_18269,N_18347);
nor U18635 (N_18635,N_18055,N_18425);
or U18636 (N_18636,N_18017,N_18231);
nor U18637 (N_18637,N_18340,N_18379);
or U18638 (N_18638,N_18273,N_18050);
or U18639 (N_18639,N_18362,N_18574);
and U18640 (N_18640,N_18064,N_18589);
and U18641 (N_18641,N_18030,N_18383);
or U18642 (N_18642,N_18489,N_18145);
xor U18643 (N_18643,N_18572,N_18505);
nor U18644 (N_18644,N_18293,N_18498);
and U18645 (N_18645,N_18309,N_18485);
nor U18646 (N_18646,N_18353,N_18146);
or U18647 (N_18647,N_18381,N_18223);
nand U18648 (N_18648,N_18333,N_18233);
nand U18649 (N_18649,N_18343,N_18592);
or U18650 (N_18650,N_18359,N_18043);
or U18651 (N_18651,N_18533,N_18253);
nor U18652 (N_18652,N_18141,N_18470);
and U18653 (N_18653,N_18229,N_18265);
nand U18654 (N_18654,N_18419,N_18427);
xor U18655 (N_18655,N_18514,N_18522);
and U18656 (N_18656,N_18018,N_18181);
or U18657 (N_18657,N_18248,N_18393);
xor U18658 (N_18658,N_18077,N_18295);
nand U18659 (N_18659,N_18394,N_18210);
xor U18660 (N_18660,N_18420,N_18409);
nor U18661 (N_18661,N_18323,N_18093);
nand U18662 (N_18662,N_18138,N_18084);
nand U18663 (N_18663,N_18545,N_18527);
and U18664 (N_18664,N_18178,N_18342);
xor U18665 (N_18665,N_18357,N_18228);
nor U18666 (N_18666,N_18433,N_18163);
or U18667 (N_18667,N_18320,N_18355);
or U18668 (N_18668,N_18096,N_18150);
or U18669 (N_18669,N_18148,N_18597);
nor U18670 (N_18670,N_18142,N_18196);
xor U18671 (N_18671,N_18222,N_18135);
and U18672 (N_18672,N_18065,N_18496);
and U18673 (N_18673,N_18424,N_18525);
and U18674 (N_18674,N_18202,N_18546);
nor U18675 (N_18675,N_18283,N_18467);
and U18676 (N_18676,N_18459,N_18329);
xnor U18677 (N_18677,N_18053,N_18490);
nand U18678 (N_18678,N_18439,N_18070);
and U18679 (N_18679,N_18028,N_18299);
and U18680 (N_18680,N_18354,N_18451);
nand U18681 (N_18681,N_18182,N_18469);
xnor U18682 (N_18682,N_18205,N_18126);
nand U18683 (N_18683,N_18276,N_18094);
nor U18684 (N_18684,N_18241,N_18207);
and U18685 (N_18685,N_18322,N_18152);
nor U18686 (N_18686,N_18262,N_18587);
or U18687 (N_18687,N_18400,N_18404);
xnor U18688 (N_18688,N_18570,N_18234);
xor U18689 (N_18689,N_18190,N_18539);
and U18690 (N_18690,N_18378,N_18116);
and U18691 (N_18691,N_18104,N_18434);
nand U18692 (N_18692,N_18554,N_18518);
nand U18693 (N_18693,N_18284,N_18230);
xnor U18694 (N_18694,N_18212,N_18097);
nand U18695 (N_18695,N_18054,N_18594);
nor U18696 (N_18696,N_18487,N_18171);
or U18697 (N_18697,N_18367,N_18479);
xor U18698 (N_18698,N_18303,N_18302);
or U18699 (N_18699,N_18315,N_18312);
xor U18700 (N_18700,N_18561,N_18268);
nor U18701 (N_18701,N_18328,N_18375);
xor U18702 (N_18702,N_18201,N_18166);
or U18703 (N_18703,N_18426,N_18188);
xnor U18704 (N_18704,N_18411,N_18003);
xor U18705 (N_18705,N_18177,N_18258);
or U18706 (N_18706,N_18477,N_18399);
nor U18707 (N_18707,N_18390,N_18585);
xor U18708 (N_18708,N_18208,N_18346);
nand U18709 (N_18709,N_18153,N_18305);
and U18710 (N_18710,N_18079,N_18325);
xor U18711 (N_18711,N_18071,N_18010);
or U18712 (N_18712,N_18290,N_18180);
and U18713 (N_18713,N_18121,N_18118);
xor U18714 (N_18714,N_18510,N_18417);
nand U18715 (N_18715,N_18406,N_18137);
nand U18716 (N_18716,N_18068,N_18235);
or U18717 (N_18717,N_18136,N_18578);
nor U18718 (N_18718,N_18058,N_18014);
and U18719 (N_18719,N_18364,N_18519);
xnor U18720 (N_18720,N_18215,N_18474);
nor U18721 (N_18721,N_18504,N_18503);
or U18722 (N_18722,N_18461,N_18051);
nor U18723 (N_18723,N_18168,N_18144);
nor U18724 (N_18724,N_18078,N_18060);
nor U18725 (N_18725,N_18066,N_18398);
or U18726 (N_18726,N_18306,N_18184);
xor U18727 (N_18727,N_18576,N_18195);
or U18728 (N_18728,N_18555,N_18511);
nor U18729 (N_18729,N_18286,N_18529);
xnor U18730 (N_18730,N_18015,N_18012);
and U18731 (N_18731,N_18038,N_18593);
or U18732 (N_18732,N_18556,N_18319);
xnor U18733 (N_18733,N_18256,N_18088);
or U18734 (N_18734,N_18560,N_18558);
nand U18735 (N_18735,N_18219,N_18316);
and U18736 (N_18736,N_18415,N_18270);
or U18737 (N_18737,N_18164,N_18449);
nor U18738 (N_18738,N_18566,N_18386);
nor U18739 (N_18739,N_18494,N_18046);
nand U18740 (N_18740,N_18263,N_18074);
nand U18741 (N_18741,N_18414,N_18083);
nor U18742 (N_18742,N_18350,N_18159);
and U18743 (N_18743,N_18413,N_18584);
xnor U18744 (N_18744,N_18336,N_18172);
or U18745 (N_18745,N_18063,N_18582);
nor U18746 (N_18746,N_18061,N_18022);
or U18747 (N_18747,N_18037,N_18590);
or U18748 (N_18748,N_18103,N_18391);
nand U18749 (N_18749,N_18296,N_18370);
or U18750 (N_18750,N_18250,N_18544);
or U18751 (N_18751,N_18339,N_18385);
xnor U18752 (N_18752,N_18218,N_18105);
or U18753 (N_18753,N_18428,N_18532);
nand U18754 (N_18754,N_18365,N_18547);
or U18755 (N_18755,N_18351,N_18179);
and U18756 (N_18756,N_18127,N_18289);
nor U18757 (N_18757,N_18119,N_18535);
nand U18758 (N_18758,N_18216,N_18338);
nand U18759 (N_18759,N_18024,N_18271);
or U18760 (N_18760,N_18278,N_18112);
nand U18761 (N_18761,N_18310,N_18313);
nor U18762 (N_18762,N_18380,N_18282);
xnor U18763 (N_18763,N_18552,N_18520);
and U18764 (N_18764,N_18013,N_18395);
or U18765 (N_18765,N_18407,N_18194);
or U18766 (N_18766,N_18085,N_18412);
nand U18767 (N_18767,N_18175,N_18358);
and U18768 (N_18768,N_18108,N_18486);
and U18769 (N_18769,N_18291,N_18495);
xor U18770 (N_18770,N_18034,N_18232);
xor U18771 (N_18771,N_18189,N_18087);
and U18772 (N_18772,N_18550,N_18360);
or U18773 (N_18773,N_18032,N_18267);
nor U18774 (N_18774,N_18452,N_18540);
and U18775 (N_18775,N_18275,N_18416);
xnor U18776 (N_18776,N_18086,N_18095);
xnor U18777 (N_18777,N_18245,N_18372);
or U18778 (N_18778,N_18466,N_18117);
and U18779 (N_18779,N_18430,N_18082);
nand U18780 (N_18780,N_18538,N_18553);
nand U18781 (N_18781,N_18115,N_18292);
nor U18782 (N_18782,N_18007,N_18423);
xor U18783 (N_18783,N_18285,N_18528);
or U18784 (N_18784,N_18396,N_18438);
xnor U18785 (N_18785,N_18446,N_18287);
nor U18786 (N_18786,N_18237,N_18565);
xnor U18787 (N_18787,N_18531,N_18512);
nor U18788 (N_18788,N_18297,N_18499);
xnor U18789 (N_18789,N_18151,N_18304);
or U18790 (N_18790,N_18369,N_18041);
xnor U18791 (N_18791,N_18057,N_18562);
and U18792 (N_18792,N_18005,N_18133);
nand U18793 (N_18793,N_18374,N_18403);
nor U18794 (N_18794,N_18596,N_18588);
nor U18795 (N_18795,N_18033,N_18464);
or U18796 (N_18796,N_18541,N_18044);
or U18797 (N_18797,N_18341,N_18448);
and U18798 (N_18798,N_18298,N_18120);
nor U18799 (N_18799,N_18185,N_18158);
and U18800 (N_18800,N_18029,N_18314);
and U18801 (N_18801,N_18526,N_18165);
xnor U18802 (N_18802,N_18176,N_18318);
xor U18803 (N_18803,N_18344,N_18389);
nor U18804 (N_18804,N_18473,N_18156);
and U18805 (N_18805,N_18209,N_18444);
nand U18806 (N_18806,N_18128,N_18255);
nand U18807 (N_18807,N_18274,N_18040);
nand U18808 (N_18808,N_18497,N_18069);
nand U18809 (N_18809,N_18149,N_18371);
nor U18810 (N_18810,N_18481,N_18580);
or U18811 (N_18811,N_18458,N_18080);
nand U18812 (N_18812,N_18300,N_18456);
nor U18813 (N_18813,N_18123,N_18246);
nand U18814 (N_18814,N_18348,N_18509);
and U18815 (N_18815,N_18025,N_18021);
nand U18816 (N_18816,N_18124,N_18484);
and U18817 (N_18817,N_18075,N_18557);
nor U18818 (N_18818,N_18161,N_18571);
xnor U18819 (N_18819,N_18463,N_18220);
xnor U18820 (N_18820,N_18373,N_18402);
nand U18821 (N_18821,N_18392,N_18445);
or U18822 (N_18822,N_18252,N_18599);
xnor U18823 (N_18823,N_18011,N_18100);
nor U18824 (N_18824,N_18143,N_18460);
xor U18825 (N_18825,N_18191,N_18122);
and U18826 (N_18826,N_18382,N_18462);
xnor U18827 (N_18827,N_18059,N_18259);
xnor U18828 (N_18828,N_18501,N_18036);
xnor U18829 (N_18829,N_18515,N_18198);
nand U18830 (N_18830,N_18352,N_18134);
nor U18831 (N_18831,N_18173,N_18548);
and U18832 (N_18832,N_18361,N_18575);
xor U18833 (N_18833,N_18507,N_18027);
nor U18834 (N_18834,N_18131,N_18327);
xnor U18835 (N_18835,N_18468,N_18450);
or U18836 (N_18836,N_18317,N_18247);
xor U18837 (N_18837,N_18225,N_18471);
xor U18838 (N_18838,N_18076,N_18023);
and U18839 (N_18839,N_18110,N_18139);
nor U18840 (N_18840,N_18056,N_18239);
nand U18841 (N_18841,N_18217,N_18376);
nor U18842 (N_18842,N_18244,N_18308);
or U18843 (N_18843,N_18488,N_18559);
xor U18844 (N_18844,N_18537,N_18523);
nand U18845 (N_18845,N_18521,N_18125);
and U18846 (N_18846,N_18106,N_18009);
nor U18847 (N_18847,N_18251,N_18281);
xor U18848 (N_18848,N_18004,N_18549);
or U18849 (N_18849,N_18031,N_18002);
xor U18850 (N_18850,N_18035,N_18260);
nand U18851 (N_18851,N_18453,N_18441);
xor U18852 (N_18852,N_18431,N_18502);
nand U18853 (N_18853,N_18577,N_18349);
and U18854 (N_18854,N_18366,N_18019);
or U18855 (N_18855,N_18042,N_18155);
xor U18856 (N_18856,N_18204,N_18331);
nor U18857 (N_18857,N_18257,N_18111);
xnor U18858 (N_18858,N_18583,N_18067);
xor U18859 (N_18859,N_18405,N_18524);
or U18860 (N_18860,N_18478,N_18492);
nand U18861 (N_18861,N_18591,N_18052);
nand U18862 (N_18862,N_18114,N_18226);
nand U18863 (N_18863,N_18408,N_18272);
and U18864 (N_18864,N_18174,N_18089);
nor U18865 (N_18865,N_18107,N_18213);
or U18866 (N_18866,N_18170,N_18224);
nand U18867 (N_18867,N_18091,N_18377);
and U18868 (N_18868,N_18072,N_18443);
or U18869 (N_18869,N_18476,N_18026);
or U18870 (N_18870,N_18543,N_18480);
and U18871 (N_18871,N_18249,N_18567);
and U18872 (N_18872,N_18016,N_18536);
nor U18873 (N_18873,N_18506,N_18530);
and U18874 (N_18874,N_18513,N_18147);
or U18875 (N_18875,N_18261,N_18266);
or U18876 (N_18876,N_18102,N_18238);
nand U18877 (N_18877,N_18311,N_18493);
xor U18878 (N_18878,N_18598,N_18242);
xnor U18879 (N_18879,N_18006,N_18410);
nand U18880 (N_18880,N_18045,N_18062);
nor U18881 (N_18881,N_18581,N_18508);
and U18882 (N_18882,N_18491,N_18157);
nand U18883 (N_18883,N_18206,N_18113);
xor U18884 (N_18884,N_18563,N_18187);
xnor U18885 (N_18885,N_18288,N_18227);
xor U18886 (N_18886,N_18154,N_18101);
nand U18887 (N_18887,N_18301,N_18160);
and U18888 (N_18888,N_18551,N_18475);
nor U18889 (N_18889,N_18039,N_18162);
nand U18890 (N_18890,N_18001,N_18254);
nor U18891 (N_18891,N_18203,N_18482);
xnor U18892 (N_18892,N_18192,N_18397);
nand U18893 (N_18893,N_18167,N_18324);
nor U18894 (N_18894,N_18401,N_18437);
nor U18895 (N_18895,N_18442,N_18457);
xnor U18896 (N_18896,N_18356,N_18186);
nand U18897 (N_18897,N_18436,N_18321);
nand U18898 (N_18898,N_18129,N_18130);
nand U18899 (N_18899,N_18418,N_18221);
nand U18900 (N_18900,N_18277,N_18492);
nor U18901 (N_18901,N_18031,N_18289);
and U18902 (N_18902,N_18334,N_18369);
nor U18903 (N_18903,N_18541,N_18396);
or U18904 (N_18904,N_18300,N_18443);
or U18905 (N_18905,N_18510,N_18225);
and U18906 (N_18906,N_18245,N_18057);
and U18907 (N_18907,N_18554,N_18210);
nand U18908 (N_18908,N_18348,N_18170);
and U18909 (N_18909,N_18049,N_18331);
xnor U18910 (N_18910,N_18541,N_18172);
or U18911 (N_18911,N_18562,N_18465);
or U18912 (N_18912,N_18164,N_18246);
xor U18913 (N_18913,N_18332,N_18147);
nand U18914 (N_18914,N_18204,N_18446);
or U18915 (N_18915,N_18479,N_18442);
nor U18916 (N_18916,N_18063,N_18156);
or U18917 (N_18917,N_18429,N_18366);
xor U18918 (N_18918,N_18099,N_18385);
nor U18919 (N_18919,N_18054,N_18516);
and U18920 (N_18920,N_18302,N_18406);
or U18921 (N_18921,N_18389,N_18107);
nor U18922 (N_18922,N_18432,N_18436);
xor U18923 (N_18923,N_18473,N_18426);
nor U18924 (N_18924,N_18516,N_18593);
xnor U18925 (N_18925,N_18526,N_18481);
or U18926 (N_18926,N_18568,N_18248);
and U18927 (N_18927,N_18495,N_18058);
and U18928 (N_18928,N_18499,N_18037);
nor U18929 (N_18929,N_18515,N_18335);
nor U18930 (N_18930,N_18522,N_18075);
or U18931 (N_18931,N_18007,N_18450);
and U18932 (N_18932,N_18335,N_18361);
nand U18933 (N_18933,N_18054,N_18365);
and U18934 (N_18934,N_18129,N_18074);
nand U18935 (N_18935,N_18004,N_18240);
or U18936 (N_18936,N_18384,N_18483);
and U18937 (N_18937,N_18525,N_18096);
and U18938 (N_18938,N_18146,N_18572);
and U18939 (N_18939,N_18074,N_18500);
xor U18940 (N_18940,N_18055,N_18315);
nor U18941 (N_18941,N_18232,N_18217);
and U18942 (N_18942,N_18384,N_18018);
xnor U18943 (N_18943,N_18570,N_18062);
nor U18944 (N_18944,N_18142,N_18100);
or U18945 (N_18945,N_18383,N_18532);
and U18946 (N_18946,N_18491,N_18545);
and U18947 (N_18947,N_18214,N_18436);
xnor U18948 (N_18948,N_18057,N_18173);
and U18949 (N_18949,N_18336,N_18260);
nand U18950 (N_18950,N_18488,N_18449);
nor U18951 (N_18951,N_18352,N_18348);
nor U18952 (N_18952,N_18322,N_18418);
xor U18953 (N_18953,N_18356,N_18316);
nand U18954 (N_18954,N_18103,N_18259);
xor U18955 (N_18955,N_18155,N_18112);
nor U18956 (N_18956,N_18503,N_18582);
and U18957 (N_18957,N_18583,N_18045);
nor U18958 (N_18958,N_18443,N_18089);
and U18959 (N_18959,N_18239,N_18467);
xor U18960 (N_18960,N_18490,N_18114);
nor U18961 (N_18961,N_18237,N_18597);
xnor U18962 (N_18962,N_18505,N_18100);
or U18963 (N_18963,N_18221,N_18484);
and U18964 (N_18964,N_18376,N_18406);
xor U18965 (N_18965,N_18536,N_18049);
nor U18966 (N_18966,N_18062,N_18033);
nor U18967 (N_18967,N_18480,N_18542);
nor U18968 (N_18968,N_18166,N_18070);
and U18969 (N_18969,N_18121,N_18273);
or U18970 (N_18970,N_18202,N_18046);
and U18971 (N_18971,N_18390,N_18538);
or U18972 (N_18972,N_18252,N_18108);
xor U18973 (N_18973,N_18102,N_18553);
xnor U18974 (N_18974,N_18436,N_18196);
and U18975 (N_18975,N_18519,N_18440);
or U18976 (N_18976,N_18110,N_18017);
xor U18977 (N_18977,N_18237,N_18070);
xnor U18978 (N_18978,N_18043,N_18594);
nand U18979 (N_18979,N_18173,N_18539);
and U18980 (N_18980,N_18067,N_18139);
nor U18981 (N_18981,N_18461,N_18079);
nor U18982 (N_18982,N_18009,N_18186);
xnor U18983 (N_18983,N_18144,N_18454);
nor U18984 (N_18984,N_18215,N_18309);
xnor U18985 (N_18985,N_18239,N_18191);
nor U18986 (N_18986,N_18055,N_18142);
and U18987 (N_18987,N_18278,N_18281);
nand U18988 (N_18988,N_18242,N_18583);
and U18989 (N_18989,N_18275,N_18122);
xor U18990 (N_18990,N_18502,N_18011);
nor U18991 (N_18991,N_18440,N_18083);
nand U18992 (N_18992,N_18143,N_18553);
and U18993 (N_18993,N_18530,N_18195);
nor U18994 (N_18994,N_18523,N_18392);
or U18995 (N_18995,N_18073,N_18029);
or U18996 (N_18996,N_18528,N_18513);
or U18997 (N_18997,N_18143,N_18033);
nor U18998 (N_18998,N_18599,N_18405);
nor U18999 (N_18999,N_18357,N_18025);
or U19000 (N_19000,N_18247,N_18197);
and U19001 (N_19001,N_18332,N_18492);
nor U19002 (N_19002,N_18261,N_18439);
and U19003 (N_19003,N_18561,N_18217);
nor U19004 (N_19004,N_18505,N_18442);
xor U19005 (N_19005,N_18202,N_18478);
or U19006 (N_19006,N_18079,N_18045);
xor U19007 (N_19007,N_18280,N_18251);
or U19008 (N_19008,N_18275,N_18182);
nand U19009 (N_19009,N_18529,N_18579);
and U19010 (N_19010,N_18233,N_18444);
and U19011 (N_19011,N_18396,N_18217);
and U19012 (N_19012,N_18495,N_18329);
xnor U19013 (N_19013,N_18464,N_18232);
xor U19014 (N_19014,N_18076,N_18051);
nor U19015 (N_19015,N_18572,N_18516);
nor U19016 (N_19016,N_18211,N_18154);
or U19017 (N_19017,N_18437,N_18525);
or U19018 (N_19018,N_18156,N_18210);
or U19019 (N_19019,N_18400,N_18097);
and U19020 (N_19020,N_18493,N_18437);
or U19021 (N_19021,N_18203,N_18532);
or U19022 (N_19022,N_18331,N_18520);
nand U19023 (N_19023,N_18279,N_18514);
and U19024 (N_19024,N_18413,N_18453);
or U19025 (N_19025,N_18142,N_18484);
nor U19026 (N_19026,N_18369,N_18373);
nand U19027 (N_19027,N_18283,N_18424);
nand U19028 (N_19028,N_18272,N_18430);
and U19029 (N_19029,N_18343,N_18555);
and U19030 (N_19030,N_18092,N_18385);
or U19031 (N_19031,N_18319,N_18468);
or U19032 (N_19032,N_18073,N_18132);
xnor U19033 (N_19033,N_18456,N_18310);
nor U19034 (N_19034,N_18582,N_18071);
and U19035 (N_19035,N_18259,N_18354);
xnor U19036 (N_19036,N_18470,N_18582);
nand U19037 (N_19037,N_18459,N_18226);
nand U19038 (N_19038,N_18286,N_18122);
xor U19039 (N_19039,N_18515,N_18595);
and U19040 (N_19040,N_18511,N_18414);
nor U19041 (N_19041,N_18348,N_18240);
nand U19042 (N_19042,N_18075,N_18431);
nor U19043 (N_19043,N_18563,N_18212);
or U19044 (N_19044,N_18250,N_18419);
or U19045 (N_19045,N_18563,N_18291);
nand U19046 (N_19046,N_18285,N_18475);
xor U19047 (N_19047,N_18194,N_18269);
or U19048 (N_19048,N_18001,N_18317);
nor U19049 (N_19049,N_18345,N_18167);
xor U19050 (N_19050,N_18027,N_18091);
nand U19051 (N_19051,N_18220,N_18285);
and U19052 (N_19052,N_18492,N_18192);
xor U19053 (N_19053,N_18211,N_18281);
nor U19054 (N_19054,N_18327,N_18450);
or U19055 (N_19055,N_18395,N_18230);
and U19056 (N_19056,N_18464,N_18541);
or U19057 (N_19057,N_18541,N_18589);
nor U19058 (N_19058,N_18577,N_18549);
and U19059 (N_19059,N_18034,N_18420);
xnor U19060 (N_19060,N_18198,N_18006);
and U19061 (N_19061,N_18564,N_18289);
xnor U19062 (N_19062,N_18458,N_18182);
nor U19063 (N_19063,N_18233,N_18147);
nor U19064 (N_19064,N_18243,N_18246);
nor U19065 (N_19065,N_18045,N_18342);
or U19066 (N_19066,N_18096,N_18468);
nand U19067 (N_19067,N_18456,N_18421);
xnor U19068 (N_19068,N_18040,N_18516);
and U19069 (N_19069,N_18193,N_18352);
nor U19070 (N_19070,N_18100,N_18324);
nor U19071 (N_19071,N_18442,N_18069);
and U19072 (N_19072,N_18350,N_18534);
nand U19073 (N_19073,N_18093,N_18391);
nand U19074 (N_19074,N_18583,N_18551);
or U19075 (N_19075,N_18032,N_18055);
and U19076 (N_19076,N_18397,N_18467);
nand U19077 (N_19077,N_18453,N_18088);
nor U19078 (N_19078,N_18250,N_18361);
and U19079 (N_19079,N_18415,N_18233);
nor U19080 (N_19080,N_18174,N_18422);
or U19081 (N_19081,N_18234,N_18551);
nor U19082 (N_19082,N_18474,N_18380);
and U19083 (N_19083,N_18154,N_18462);
or U19084 (N_19084,N_18446,N_18061);
and U19085 (N_19085,N_18117,N_18014);
and U19086 (N_19086,N_18405,N_18034);
or U19087 (N_19087,N_18327,N_18175);
and U19088 (N_19088,N_18149,N_18366);
and U19089 (N_19089,N_18116,N_18449);
nand U19090 (N_19090,N_18057,N_18587);
or U19091 (N_19091,N_18043,N_18111);
and U19092 (N_19092,N_18327,N_18578);
nor U19093 (N_19093,N_18335,N_18098);
xor U19094 (N_19094,N_18308,N_18572);
or U19095 (N_19095,N_18496,N_18086);
xnor U19096 (N_19096,N_18418,N_18324);
xor U19097 (N_19097,N_18309,N_18196);
or U19098 (N_19098,N_18134,N_18291);
nor U19099 (N_19099,N_18412,N_18138);
and U19100 (N_19100,N_18006,N_18110);
or U19101 (N_19101,N_18110,N_18140);
nor U19102 (N_19102,N_18551,N_18174);
or U19103 (N_19103,N_18124,N_18572);
and U19104 (N_19104,N_18011,N_18176);
xnor U19105 (N_19105,N_18018,N_18570);
or U19106 (N_19106,N_18270,N_18258);
xor U19107 (N_19107,N_18156,N_18491);
nand U19108 (N_19108,N_18046,N_18309);
nor U19109 (N_19109,N_18247,N_18171);
nand U19110 (N_19110,N_18503,N_18174);
and U19111 (N_19111,N_18270,N_18019);
and U19112 (N_19112,N_18504,N_18095);
or U19113 (N_19113,N_18043,N_18375);
and U19114 (N_19114,N_18001,N_18537);
xnor U19115 (N_19115,N_18567,N_18594);
and U19116 (N_19116,N_18126,N_18035);
nor U19117 (N_19117,N_18438,N_18377);
nor U19118 (N_19118,N_18496,N_18011);
nand U19119 (N_19119,N_18326,N_18231);
or U19120 (N_19120,N_18444,N_18514);
or U19121 (N_19121,N_18578,N_18524);
nor U19122 (N_19122,N_18104,N_18079);
or U19123 (N_19123,N_18548,N_18002);
and U19124 (N_19124,N_18229,N_18215);
and U19125 (N_19125,N_18339,N_18406);
or U19126 (N_19126,N_18160,N_18528);
xnor U19127 (N_19127,N_18476,N_18235);
or U19128 (N_19128,N_18570,N_18552);
or U19129 (N_19129,N_18235,N_18429);
nor U19130 (N_19130,N_18329,N_18152);
or U19131 (N_19131,N_18424,N_18553);
nand U19132 (N_19132,N_18272,N_18253);
nor U19133 (N_19133,N_18345,N_18271);
or U19134 (N_19134,N_18573,N_18291);
nand U19135 (N_19135,N_18254,N_18419);
xnor U19136 (N_19136,N_18112,N_18346);
xor U19137 (N_19137,N_18201,N_18412);
and U19138 (N_19138,N_18535,N_18569);
and U19139 (N_19139,N_18242,N_18205);
xor U19140 (N_19140,N_18190,N_18546);
and U19141 (N_19141,N_18148,N_18573);
nand U19142 (N_19142,N_18322,N_18031);
nor U19143 (N_19143,N_18253,N_18357);
xor U19144 (N_19144,N_18094,N_18294);
or U19145 (N_19145,N_18042,N_18480);
nand U19146 (N_19146,N_18437,N_18396);
xnor U19147 (N_19147,N_18354,N_18371);
nand U19148 (N_19148,N_18300,N_18142);
nand U19149 (N_19149,N_18562,N_18555);
or U19150 (N_19150,N_18419,N_18045);
or U19151 (N_19151,N_18375,N_18167);
or U19152 (N_19152,N_18452,N_18059);
or U19153 (N_19153,N_18271,N_18102);
xnor U19154 (N_19154,N_18456,N_18319);
xor U19155 (N_19155,N_18264,N_18423);
and U19156 (N_19156,N_18162,N_18412);
nor U19157 (N_19157,N_18530,N_18196);
or U19158 (N_19158,N_18464,N_18136);
nor U19159 (N_19159,N_18444,N_18353);
nand U19160 (N_19160,N_18395,N_18051);
xor U19161 (N_19161,N_18118,N_18327);
and U19162 (N_19162,N_18069,N_18448);
and U19163 (N_19163,N_18131,N_18165);
xnor U19164 (N_19164,N_18577,N_18595);
xor U19165 (N_19165,N_18388,N_18235);
or U19166 (N_19166,N_18070,N_18262);
nor U19167 (N_19167,N_18361,N_18198);
nor U19168 (N_19168,N_18173,N_18233);
nor U19169 (N_19169,N_18508,N_18327);
nor U19170 (N_19170,N_18038,N_18582);
or U19171 (N_19171,N_18118,N_18157);
and U19172 (N_19172,N_18131,N_18540);
xnor U19173 (N_19173,N_18151,N_18364);
and U19174 (N_19174,N_18423,N_18087);
or U19175 (N_19175,N_18131,N_18148);
or U19176 (N_19176,N_18597,N_18467);
xnor U19177 (N_19177,N_18109,N_18502);
and U19178 (N_19178,N_18305,N_18464);
nor U19179 (N_19179,N_18097,N_18135);
or U19180 (N_19180,N_18026,N_18073);
and U19181 (N_19181,N_18121,N_18480);
or U19182 (N_19182,N_18362,N_18268);
and U19183 (N_19183,N_18449,N_18282);
xor U19184 (N_19184,N_18532,N_18232);
nand U19185 (N_19185,N_18086,N_18028);
or U19186 (N_19186,N_18266,N_18226);
nor U19187 (N_19187,N_18325,N_18375);
or U19188 (N_19188,N_18454,N_18545);
or U19189 (N_19189,N_18358,N_18133);
or U19190 (N_19190,N_18094,N_18482);
or U19191 (N_19191,N_18246,N_18542);
nor U19192 (N_19192,N_18437,N_18503);
and U19193 (N_19193,N_18264,N_18393);
nand U19194 (N_19194,N_18327,N_18129);
xor U19195 (N_19195,N_18491,N_18216);
and U19196 (N_19196,N_18519,N_18417);
and U19197 (N_19197,N_18369,N_18436);
and U19198 (N_19198,N_18503,N_18335);
xor U19199 (N_19199,N_18222,N_18032);
or U19200 (N_19200,N_19044,N_18667);
nor U19201 (N_19201,N_18974,N_19049);
or U19202 (N_19202,N_18799,N_18782);
and U19203 (N_19203,N_18649,N_18657);
nand U19204 (N_19204,N_18941,N_18745);
and U19205 (N_19205,N_18837,N_18728);
nand U19206 (N_19206,N_18931,N_18961);
nand U19207 (N_19207,N_18988,N_18817);
nand U19208 (N_19208,N_18874,N_18852);
nand U19209 (N_19209,N_18865,N_18828);
nand U19210 (N_19210,N_18990,N_18833);
or U19211 (N_19211,N_18731,N_18840);
nor U19212 (N_19212,N_19133,N_19003);
xnor U19213 (N_19213,N_19170,N_18999);
nand U19214 (N_19214,N_18654,N_18686);
nor U19215 (N_19215,N_18704,N_18643);
nand U19216 (N_19216,N_18979,N_18897);
nor U19217 (N_19217,N_19193,N_19179);
nand U19218 (N_19218,N_19165,N_18744);
nor U19219 (N_19219,N_18775,N_18638);
xor U19220 (N_19220,N_18732,N_18724);
and U19221 (N_19221,N_19141,N_18622);
nand U19222 (N_19222,N_18738,N_18829);
nand U19223 (N_19223,N_19055,N_19145);
or U19224 (N_19224,N_19053,N_18757);
and U19225 (N_19225,N_19092,N_18860);
nor U19226 (N_19226,N_18642,N_18832);
xor U19227 (N_19227,N_18664,N_19050);
nand U19228 (N_19228,N_18838,N_19006);
xnor U19229 (N_19229,N_18971,N_19109);
xor U19230 (N_19230,N_18703,N_18675);
xor U19231 (N_19231,N_19105,N_18623);
and U19232 (N_19232,N_19030,N_19103);
or U19233 (N_19233,N_19144,N_19172);
and U19234 (N_19234,N_19039,N_19000);
nor U19235 (N_19235,N_18945,N_19072);
and U19236 (N_19236,N_18952,N_19199);
nand U19237 (N_19237,N_18713,N_18807);
nand U19238 (N_19238,N_19143,N_19142);
xor U19239 (N_19239,N_18818,N_19192);
nand U19240 (N_19240,N_18851,N_18796);
nand U19241 (N_19241,N_18673,N_18676);
and U19242 (N_19242,N_18948,N_19098);
nand U19243 (N_19243,N_18951,N_19128);
xnor U19244 (N_19244,N_19082,N_18911);
nor U19245 (N_19245,N_19198,N_19108);
nor U19246 (N_19246,N_19191,N_18762);
nand U19247 (N_19247,N_19075,N_18972);
nor U19248 (N_19248,N_18850,N_18652);
nor U19249 (N_19249,N_18924,N_19161);
nor U19250 (N_19250,N_18632,N_18929);
nor U19251 (N_19251,N_19110,N_19090);
and U19252 (N_19252,N_18692,N_18920);
and U19253 (N_19253,N_18960,N_18942);
nor U19254 (N_19254,N_18694,N_18615);
nor U19255 (N_19255,N_18827,N_19069);
xor U19256 (N_19256,N_18973,N_19015);
or U19257 (N_19257,N_19017,N_18889);
nand U19258 (N_19258,N_18976,N_19185);
and U19259 (N_19259,N_19056,N_18726);
or U19260 (N_19260,N_18742,N_18697);
or U19261 (N_19261,N_19112,N_18985);
nor U19262 (N_19262,N_18611,N_18639);
nor U19263 (N_19263,N_19005,N_18801);
nand U19264 (N_19264,N_18767,N_18871);
or U19265 (N_19265,N_19051,N_18980);
xor U19266 (N_19266,N_18719,N_18982);
or U19267 (N_19267,N_19134,N_19059);
nor U19268 (N_19268,N_18957,N_18787);
and U19269 (N_19269,N_18940,N_18688);
or U19270 (N_19270,N_18915,N_19107);
nand U19271 (N_19271,N_18802,N_19010);
nand U19272 (N_19272,N_18646,N_18682);
nand U19273 (N_19273,N_18991,N_18890);
and U19274 (N_19274,N_18804,N_18984);
xor U19275 (N_19275,N_18614,N_18702);
nor U19276 (N_19276,N_18774,N_18730);
nand U19277 (N_19277,N_18629,N_18710);
or U19278 (N_19278,N_18779,N_18723);
xnor U19279 (N_19279,N_19150,N_18927);
and U19280 (N_19280,N_18881,N_18620);
or U19281 (N_19281,N_18747,N_18873);
and U19282 (N_19282,N_18875,N_19077);
or U19283 (N_19283,N_18717,N_18908);
xor U19284 (N_19284,N_19086,N_18935);
xor U19285 (N_19285,N_19099,N_18653);
nor U19286 (N_19286,N_18609,N_18863);
or U19287 (N_19287,N_19095,N_19113);
or U19288 (N_19288,N_18853,N_19009);
xnor U19289 (N_19289,N_19153,N_19096);
xor U19290 (N_19290,N_18919,N_18758);
and U19291 (N_19291,N_19091,N_18902);
and U19292 (N_19292,N_18880,N_19123);
xor U19293 (N_19293,N_18877,N_19060);
or U19294 (N_19294,N_19116,N_19176);
and U19295 (N_19295,N_18635,N_18678);
or U19296 (N_19296,N_18885,N_19182);
and U19297 (N_19297,N_18975,N_19088);
or U19298 (N_19298,N_18843,N_18819);
nand U19299 (N_19299,N_18862,N_19001);
nor U19300 (N_19300,N_19035,N_19156);
xor U19301 (N_19301,N_18791,N_18823);
nor U19302 (N_19302,N_18763,N_18967);
nor U19303 (N_19303,N_18835,N_19043);
nand U19304 (N_19304,N_19158,N_18898);
and U19305 (N_19305,N_18749,N_19151);
and U19306 (N_19306,N_19124,N_18668);
xor U19307 (N_19307,N_18641,N_19171);
nor U19308 (N_19308,N_18687,N_19138);
and U19309 (N_19309,N_19031,N_19080);
xor U19310 (N_19310,N_19087,N_18669);
xnor U19311 (N_19311,N_18913,N_18868);
nand U19312 (N_19312,N_19014,N_18734);
xnor U19313 (N_19313,N_18794,N_19114);
or U19314 (N_19314,N_19132,N_18670);
nand U19315 (N_19315,N_19081,N_18636);
or U19316 (N_19316,N_18867,N_19190);
nand U19317 (N_19317,N_19078,N_19073);
nand U19318 (N_19318,N_18617,N_19149);
or U19319 (N_19319,N_18949,N_18683);
xor U19320 (N_19320,N_18786,N_18856);
nand U19321 (N_19321,N_19127,N_18921);
xnor U19322 (N_19322,N_18778,N_18813);
nor U19323 (N_19323,N_19029,N_19040);
nand U19324 (N_19324,N_18896,N_18983);
and U19325 (N_19325,N_18956,N_18816);
xor U19326 (N_19326,N_18809,N_19163);
nand U19327 (N_19327,N_18901,N_18644);
nor U19328 (N_19328,N_18612,N_18854);
nand U19329 (N_19329,N_18748,N_18701);
xor U19330 (N_19330,N_18781,N_18857);
xor U19331 (N_19331,N_18711,N_18760);
xor U19332 (N_19332,N_19135,N_19093);
nand U19333 (N_19333,N_19119,N_18729);
or U19334 (N_19334,N_19175,N_18798);
or U19335 (N_19335,N_19038,N_18696);
nor U19336 (N_19336,N_19018,N_18803);
xnor U19337 (N_19337,N_18712,N_18618);
or U19338 (N_19338,N_18680,N_19117);
or U19339 (N_19339,N_18663,N_18739);
nand U19340 (N_19340,N_19063,N_18977);
nand U19341 (N_19341,N_19102,N_18790);
nor U19342 (N_19342,N_18936,N_18756);
nor U19343 (N_19343,N_18780,N_18904);
xnor U19344 (N_19344,N_19126,N_19121);
xnor U19345 (N_19345,N_18876,N_19186);
nor U19346 (N_19346,N_18969,N_18754);
or U19347 (N_19347,N_18666,N_18736);
xnor U19348 (N_19348,N_19048,N_18662);
nor U19349 (N_19349,N_18811,N_18909);
nand U19350 (N_19350,N_18647,N_19061);
nand U19351 (N_19351,N_18814,N_18626);
xnor U19352 (N_19352,N_18933,N_18826);
and U19353 (N_19353,N_19194,N_18624);
nor U19354 (N_19354,N_18955,N_18751);
nor U19355 (N_19355,N_19178,N_18842);
nor U19356 (N_19356,N_18771,N_18943);
nor U19357 (N_19357,N_19118,N_18815);
and U19358 (N_19358,N_18950,N_18613);
nor U19359 (N_19359,N_19160,N_19196);
nand U19360 (N_19360,N_18848,N_18772);
nand U19361 (N_19361,N_19089,N_18892);
xor U19362 (N_19362,N_18681,N_18830);
and U19363 (N_19363,N_19168,N_18859);
xnor U19364 (N_19364,N_19197,N_19115);
nand U19365 (N_19365,N_19002,N_18986);
and U19366 (N_19366,N_19066,N_18634);
nand U19367 (N_19367,N_18705,N_18916);
and U19368 (N_19368,N_18601,N_19012);
and U19369 (N_19369,N_18770,N_19036);
nand U19370 (N_19370,N_19052,N_18822);
xnor U19371 (N_19371,N_19162,N_18743);
or U19372 (N_19372,N_19155,N_18718);
or U19373 (N_19373,N_18993,N_18788);
or U19374 (N_19374,N_18965,N_18628);
xor U19375 (N_19375,N_18608,N_19136);
or U19376 (N_19376,N_19104,N_19181);
nand U19377 (N_19377,N_18994,N_18905);
or U19378 (N_19378,N_18741,N_19125);
and U19379 (N_19379,N_19013,N_18700);
or U19380 (N_19380,N_18766,N_18939);
or U19381 (N_19381,N_18671,N_18891);
nand U19382 (N_19382,N_19021,N_19067);
or U19383 (N_19383,N_18797,N_19028);
or U19384 (N_19384,N_18661,N_18707);
and U19385 (N_19385,N_19147,N_19084);
nor U19386 (N_19386,N_19047,N_19189);
nand U19387 (N_19387,N_19146,N_18962);
xor U19388 (N_19388,N_19019,N_18727);
or U19389 (N_19389,N_19034,N_18709);
xnor U19390 (N_19390,N_18926,N_18878);
and U19391 (N_19391,N_18755,N_18855);
and U19392 (N_19392,N_18737,N_18996);
and U19393 (N_19393,N_18938,N_18793);
nand U19394 (N_19394,N_18789,N_19106);
nor U19395 (N_19395,N_18677,N_18954);
and U19396 (N_19396,N_18784,N_18844);
nand U19397 (N_19397,N_18746,N_18658);
nor U19398 (N_19398,N_18627,N_19195);
and U19399 (N_19399,N_18689,N_18978);
nand U19400 (N_19400,N_18997,N_18698);
nand U19401 (N_19401,N_18750,N_18998);
nor U19402 (N_19402,N_18820,N_19064);
nand U19403 (N_19403,N_19020,N_18769);
and U19404 (N_19404,N_18600,N_18721);
or U19405 (N_19405,N_19101,N_18637);
and U19406 (N_19406,N_19022,N_18733);
nand U19407 (N_19407,N_18879,N_19157);
and U19408 (N_19408,N_19164,N_18866);
and U19409 (N_19409,N_18900,N_18834);
xor U19410 (N_19410,N_19011,N_18937);
nor U19411 (N_19411,N_18765,N_18659);
or U19412 (N_19412,N_19167,N_18917);
xnor U19413 (N_19413,N_18964,N_18870);
xor U19414 (N_19414,N_18625,N_19025);
nor U19415 (N_19415,N_19042,N_19094);
xor U19416 (N_19416,N_19004,N_18970);
nand U19417 (N_19417,N_18651,N_18725);
nand U19418 (N_19418,N_18656,N_19054);
nand U19419 (N_19419,N_19023,N_18932);
nor U19420 (N_19420,N_18761,N_18861);
and U19421 (N_19421,N_19120,N_18987);
and U19422 (N_19422,N_19070,N_19188);
xor U19423 (N_19423,N_19174,N_18604);
nor U19424 (N_19424,N_19016,N_18650);
nand U19425 (N_19425,N_18914,N_18839);
or U19426 (N_19426,N_18806,N_19166);
nor U19427 (N_19427,N_18884,N_19148);
or U19428 (N_19428,N_19083,N_18716);
or U19429 (N_19429,N_19129,N_18773);
nor U19430 (N_19430,N_18740,N_18883);
or U19431 (N_19431,N_19026,N_18735);
nand U19432 (N_19432,N_19033,N_18708);
nand U19433 (N_19433,N_18699,N_19046);
and U19434 (N_19434,N_19057,N_18616);
or U19435 (N_19435,N_18812,N_19076);
nand U19436 (N_19436,N_19071,N_18831);
nor U19437 (N_19437,N_18640,N_18679);
xor U19438 (N_19438,N_19177,N_18603);
xor U19439 (N_19439,N_18849,N_18899);
and U19440 (N_19440,N_18777,N_18963);
or U19441 (N_19441,N_19058,N_18888);
nand U19442 (N_19442,N_18685,N_18783);
xor U19443 (N_19443,N_18672,N_19024);
or U19444 (N_19444,N_19139,N_18930);
nor U19445 (N_19445,N_18752,N_18958);
xor U19446 (N_19446,N_19068,N_19159);
and U19447 (N_19447,N_18858,N_18764);
nor U19448 (N_19448,N_18925,N_18805);
nand U19449 (N_19449,N_19065,N_18895);
xnor U19450 (N_19450,N_18953,N_18981);
nand U19451 (N_19451,N_19183,N_19062);
xor U19452 (N_19452,N_18995,N_19131);
nand U19453 (N_19453,N_18665,N_19154);
xnor U19454 (N_19454,N_18607,N_18989);
xor U19455 (N_19455,N_19027,N_18706);
xor U19456 (N_19456,N_18912,N_18808);
nor U19457 (N_19457,N_18645,N_18768);
and U19458 (N_19458,N_18887,N_19045);
nor U19459 (N_19459,N_18907,N_18825);
nand U19460 (N_19460,N_18934,N_19032);
nand U19461 (N_19461,N_18944,N_18810);
xnor U19462 (N_19462,N_18630,N_18845);
and U19463 (N_19463,N_18841,N_18821);
nor U19464 (N_19464,N_18693,N_19085);
nor U19465 (N_19465,N_18906,N_18633);
xnor U19466 (N_19466,N_18847,N_18655);
or U19467 (N_19467,N_18619,N_19187);
or U19468 (N_19468,N_18886,N_18753);
and U19469 (N_19469,N_18800,N_18836);
xor U19470 (N_19470,N_18648,N_18882);
or U19471 (N_19471,N_18846,N_18785);
nor U19472 (N_19472,N_18606,N_19074);
and U19473 (N_19473,N_18872,N_18928);
nand U19474 (N_19474,N_18795,N_18714);
xor U19475 (N_19475,N_18903,N_18695);
or U19476 (N_19476,N_19180,N_19184);
nand U19477 (N_19477,N_18894,N_18992);
nand U19478 (N_19478,N_18720,N_18910);
or U19479 (N_19479,N_19137,N_18674);
nand U19480 (N_19480,N_18893,N_19152);
nand U19481 (N_19481,N_19169,N_18968);
nor U19482 (N_19482,N_19041,N_19100);
and U19483 (N_19483,N_18631,N_18690);
xor U19484 (N_19484,N_18946,N_19130);
nand U19485 (N_19485,N_18722,N_19037);
and U19486 (N_19486,N_18621,N_19007);
xor U19487 (N_19487,N_19111,N_18691);
and U19488 (N_19488,N_18759,N_18610);
nor U19489 (N_19489,N_18776,N_18959);
nor U19490 (N_19490,N_18922,N_19097);
nand U19491 (N_19491,N_18792,N_18602);
or U19492 (N_19492,N_18918,N_19140);
nand U19493 (N_19493,N_19122,N_18605);
or U19494 (N_19494,N_19173,N_18869);
nor U19495 (N_19495,N_18966,N_18947);
nor U19496 (N_19496,N_18864,N_18684);
xor U19497 (N_19497,N_19008,N_18923);
nor U19498 (N_19498,N_18715,N_18660);
or U19499 (N_19499,N_18824,N_19079);
and U19500 (N_19500,N_18885,N_18708);
and U19501 (N_19501,N_19113,N_18774);
and U19502 (N_19502,N_18634,N_19079);
or U19503 (N_19503,N_18809,N_18874);
nand U19504 (N_19504,N_19060,N_18737);
nand U19505 (N_19505,N_18948,N_18757);
nand U19506 (N_19506,N_18860,N_18705);
nor U19507 (N_19507,N_18728,N_18910);
nor U19508 (N_19508,N_18953,N_18976);
or U19509 (N_19509,N_18948,N_18908);
xnor U19510 (N_19510,N_18827,N_18728);
or U19511 (N_19511,N_18753,N_18855);
xor U19512 (N_19512,N_19008,N_18892);
or U19513 (N_19513,N_18768,N_18716);
nand U19514 (N_19514,N_18854,N_18824);
xnor U19515 (N_19515,N_18683,N_18786);
or U19516 (N_19516,N_18745,N_19018);
nand U19517 (N_19517,N_18851,N_19041);
nor U19518 (N_19518,N_18634,N_18625);
nand U19519 (N_19519,N_18689,N_18769);
and U19520 (N_19520,N_18851,N_18738);
or U19521 (N_19521,N_18848,N_18986);
xor U19522 (N_19522,N_18679,N_18790);
nor U19523 (N_19523,N_18670,N_18705);
or U19524 (N_19524,N_18984,N_18767);
nand U19525 (N_19525,N_18956,N_18819);
or U19526 (N_19526,N_18934,N_18973);
and U19527 (N_19527,N_18651,N_18837);
nand U19528 (N_19528,N_18903,N_18767);
and U19529 (N_19529,N_18920,N_18848);
xnor U19530 (N_19530,N_19146,N_18756);
or U19531 (N_19531,N_18754,N_18953);
nor U19532 (N_19532,N_19141,N_19154);
and U19533 (N_19533,N_19078,N_18979);
xor U19534 (N_19534,N_18695,N_19163);
and U19535 (N_19535,N_18785,N_19008);
nand U19536 (N_19536,N_18696,N_18976);
nor U19537 (N_19537,N_19187,N_19151);
and U19538 (N_19538,N_18944,N_18720);
nor U19539 (N_19539,N_18994,N_18939);
nor U19540 (N_19540,N_19193,N_18787);
xnor U19541 (N_19541,N_18986,N_19186);
and U19542 (N_19542,N_19087,N_19039);
xor U19543 (N_19543,N_18957,N_18695);
or U19544 (N_19544,N_19111,N_18964);
xnor U19545 (N_19545,N_18759,N_19017);
nand U19546 (N_19546,N_19126,N_18811);
nand U19547 (N_19547,N_19025,N_18775);
nand U19548 (N_19548,N_19156,N_18698);
xor U19549 (N_19549,N_18834,N_18856);
nor U19550 (N_19550,N_18638,N_18741);
nor U19551 (N_19551,N_18641,N_19058);
or U19552 (N_19552,N_18784,N_18638);
xnor U19553 (N_19553,N_18662,N_18792);
nand U19554 (N_19554,N_18635,N_18673);
or U19555 (N_19555,N_18658,N_19111);
or U19556 (N_19556,N_18735,N_18794);
xor U19557 (N_19557,N_18658,N_19112);
xnor U19558 (N_19558,N_18754,N_18780);
xor U19559 (N_19559,N_18900,N_18838);
and U19560 (N_19560,N_18987,N_18845);
or U19561 (N_19561,N_18694,N_19014);
and U19562 (N_19562,N_18679,N_19069);
nor U19563 (N_19563,N_18861,N_18932);
and U19564 (N_19564,N_18932,N_18842);
or U19565 (N_19565,N_18639,N_18884);
nand U19566 (N_19566,N_18743,N_18693);
nand U19567 (N_19567,N_18934,N_18932);
nand U19568 (N_19568,N_18966,N_19035);
nand U19569 (N_19569,N_18679,N_18832);
xnor U19570 (N_19570,N_18900,N_18612);
nand U19571 (N_19571,N_18796,N_19197);
nand U19572 (N_19572,N_18678,N_18847);
or U19573 (N_19573,N_19023,N_18630);
or U19574 (N_19574,N_18873,N_19123);
nand U19575 (N_19575,N_18835,N_18828);
nand U19576 (N_19576,N_18767,N_18886);
nor U19577 (N_19577,N_18663,N_19098);
nor U19578 (N_19578,N_18935,N_19049);
nand U19579 (N_19579,N_18929,N_18903);
or U19580 (N_19580,N_19089,N_18886);
xnor U19581 (N_19581,N_18972,N_18832);
nand U19582 (N_19582,N_18729,N_18624);
and U19583 (N_19583,N_18901,N_19008);
and U19584 (N_19584,N_18718,N_19049);
xnor U19585 (N_19585,N_19012,N_19052);
and U19586 (N_19586,N_19026,N_19039);
nand U19587 (N_19587,N_18938,N_18904);
or U19588 (N_19588,N_18683,N_19037);
and U19589 (N_19589,N_19147,N_18961);
or U19590 (N_19590,N_19066,N_18877);
and U19591 (N_19591,N_19140,N_19081);
nor U19592 (N_19592,N_18999,N_19196);
nor U19593 (N_19593,N_18996,N_19001);
and U19594 (N_19594,N_18922,N_18710);
or U19595 (N_19595,N_19110,N_19153);
or U19596 (N_19596,N_18934,N_18855);
nor U19597 (N_19597,N_19003,N_19126);
or U19598 (N_19598,N_18777,N_19117);
nor U19599 (N_19599,N_18832,N_19014);
nand U19600 (N_19600,N_18829,N_18639);
nand U19601 (N_19601,N_18887,N_18875);
or U19602 (N_19602,N_18704,N_19080);
or U19603 (N_19603,N_18888,N_18777);
or U19604 (N_19604,N_19188,N_19106);
xnor U19605 (N_19605,N_18602,N_18775);
nand U19606 (N_19606,N_19132,N_19160);
nor U19607 (N_19607,N_19136,N_19029);
xnor U19608 (N_19608,N_18958,N_18887);
xor U19609 (N_19609,N_18949,N_18733);
xnor U19610 (N_19610,N_19071,N_18766);
nor U19611 (N_19611,N_18716,N_18679);
or U19612 (N_19612,N_18801,N_18715);
nand U19613 (N_19613,N_18987,N_18946);
nor U19614 (N_19614,N_19111,N_18631);
nand U19615 (N_19615,N_18825,N_18643);
xnor U19616 (N_19616,N_18609,N_19144);
or U19617 (N_19617,N_18792,N_18649);
or U19618 (N_19618,N_18701,N_18789);
xnor U19619 (N_19619,N_19148,N_19195);
nand U19620 (N_19620,N_19085,N_18835);
nand U19621 (N_19621,N_18853,N_18797);
nor U19622 (N_19622,N_18840,N_18743);
xor U19623 (N_19623,N_18846,N_19017);
and U19624 (N_19624,N_19136,N_18648);
xnor U19625 (N_19625,N_18875,N_19045);
nand U19626 (N_19626,N_18909,N_19119);
or U19627 (N_19627,N_18712,N_18695);
xnor U19628 (N_19628,N_18882,N_18888);
nor U19629 (N_19629,N_18941,N_18671);
nand U19630 (N_19630,N_18641,N_18722);
or U19631 (N_19631,N_18948,N_18737);
or U19632 (N_19632,N_18959,N_19139);
and U19633 (N_19633,N_18638,N_18758);
xor U19634 (N_19634,N_18956,N_18936);
and U19635 (N_19635,N_19149,N_19146);
nor U19636 (N_19636,N_19140,N_18937);
nand U19637 (N_19637,N_18614,N_18982);
or U19638 (N_19638,N_18754,N_18649);
or U19639 (N_19639,N_19159,N_18632);
nor U19640 (N_19640,N_19006,N_18827);
nor U19641 (N_19641,N_19149,N_18891);
nor U19642 (N_19642,N_18906,N_18988);
or U19643 (N_19643,N_19003,N_19113);
nor U19644 (N_19644,N_18748,N_18937);
nand U19645 (N_19645,N_18681,N_18723);
xnor U19646 (N_19646,N_19032,N_18968);
nand U19647 (N_19647,N_18948,N_18937);
nor U19648 (N_19648,N_18629,N_19140);
or U19649 (N_19649,N_18689,N_19070);
nand U19650 (N_19650,N_18673,N_18716);
nor U19651 (N_19651,N_19171,N_18986);
or U19652 (N_19652,N_18801,N_18655);
nor U19653 (N_19653,N_19180,N_18962);
or U19654 (N_19654,N_18965,N_19094);
xnor U19655 (N_19655,N_19119,N_18784);
and U19656 (N_19656,N_18686,N_18977);
nand U19657 (N_19657,N_18819,N_19049);
and U19658 (N_19658,N_18709,N_18957);
and U19659 (N_19659,N_19152,N_18892);
xor U19660 (N_19660,N_18960,N_18933);
and U19661 (N_19661,N_18972,N_19191);
or U19662 (N_19662,N_18758,N_18819);
xor U19663 (N_19663,N_18774,N_18806);
xor U19664 (N_19664,N_19076,N_19088);
xnor U19665 (N_19665,N_18701,N_18683);
xor U19666 (N_19666,N_18795,N_18994);
nor U19667 (N_19667,N_19015,N_18858);
nand U19668 (N_19668,N_18655,N_18677);
xnor U19669 (N_19669,N_18790,N_18820);
xnor U19670 (N_19670,N_18603,N_19126);
and U19671 (N_19671,N_18813,N_18986);
nand U19672 (N_19672,N_18895,N_19069);
xnor U19673 (N_19673,N_18700,N_18810);
and U19674 (N_19674,N_19153,N_18841);
nand U19675 (N_19675,N_18746,N_18667);
and U19676 (N_19676,N_19167,N_18888);
xor U19677 (N_19677,N_18724,N_19138);
and U19678 (N_19678,N_18607,N_18851);
and U19679 (N_19679,N_19186,N_18904);
nor U19680 (N_19680,N_19089,N_19110);
and U19681 (N_19681,N_19069,N_18639);
nor U19682 (N_19682,N_18876,N_18768);
and U19683 (N_19683,N_18813,N_18702);
and U19684 (N_19684,N_18941,N_18785);
xnor U19685 (N_19685,N_18747,N_18806);
nand U19686 (N_19686,N_18933,N_18741);
nand U19687 (N_19687,N_18657,N_19170);
or U19688 (N_19688,N_18759,N_18871);
nand U19689 (N_19689,N_19136,N_18763);
or U19690 (N_19690,N_19012,N_19064);
or U19691 (N_19691,N_18862,N_18649);
nor U19692 (N_19692,N_18969,N_18719);
and U19693 (N_19693,N_18840,N_18735);
or U19694 (N_19694,N_19186,N_18658);
nand U19695 (N_19695,N_19069,N_18682);
nand U19696 (N_19696,N_18751,N_18897);
xor U19697 (N_19697,N_18962,N_18990);
nor U19698 (N_19698,N_19196,N_19120);
nor U19699 (N_19699,N_19042,N_18870);
nor U19700 (N_19700,N_18923,N_18634);
nor U19701 (N_19701,N_18923,N_19196);
and U19702 (N_19702,N_18847,N_19034);
nand U19703 (N_19703,N_18983,N_18683);
nand U19704 (N_19704,N_18751,N_19099);
xnor U19705 (N_19705,N_18700,N_19023);
and U19706 (N_19706,N_18693,N_18657);
and U19707 (N_19707,N_18940,N_19112);
or U19708 (N_19708,N_19080,N_18727);
or U19709 (N_19709,N_18884,N_18799);
xor U19710 (N_19710,N_18941,N_18964);
xnor U19711 (N_19711,N_18854,N_18969);
xor U19712 (N_19712,N_19087,N_18816);
xnor U19713 (N_19713,N_18999,N_18605);
and U19714 (N_19714,N_19083,N_18710);
xnor U19715 (N_19715,N_18882,N_19134);
nand U19716 (N_19716,N_18713,N_18801);
or U19717 (N_19717,N_19010,N_19097);
or U19718 (N_19718,N_18725,N_18892);
xor U19719 (N_19719,N_18708,N_19081);
xor U19720 (N_19720,N_19123,N_19133);
xor U19721 (N_19721,N_18660,N_18825);
xnor U19722 (N_19722,N_18691,N_18852);
and U19723 (N_19723,N_18722,N_18653);
xnor U19724 (N_19724,N_18839,N_18702);
or U19725 (N_19725,N_19007,N_19139);
and U19726 (N_19726,N_18617,N_19181);
xor U19727 (N_19727,N_18644,N_18754);
nand U19728 (N_19728,N_19025,N_19119);
nor U19729 (N_19729,N_19141,N_18718);
nor U19730 (N_19730,N_18849,N_18613);
nor U19731 (N_19731,N_18806,N_18751);
and U19732 (N_19732,N_18629,N_18602);
nor U19733 (N_19733,N_18711,N_19094);
nand U19734 (N_19734,N_18705,N_18856);
or U19735 (N_19735,N_18752,N_18915);
or U19736 (N_19736,N_18970,N_18690);
nor U19737 (N_19737,N_18789,N_18840);
nand U19738 (N_19738,N_18702,N_19081);
or U19739 (N_19739,N_18773,N_18777);
nor U19740 (N_19740,N_18732,N_19014);
or U19741 (N_19741,N_18923,N_18919);
or U19742 (N_19742,N_19019,N_18988);
and U19743 (N_19743,N_19120,N_18868);
nor U19744 (N_19744,N_18956,N_18774);
nor U19745 (N_19745,N_18810,N_18892);
and U19746 (N_19746,N_18714,N_18726);
nand U19747 (N_19747,N_18883,N_18627);
and U19748 (N_19748,N_18600,N_19159);
xnor U19749 (N_19749,N_19167,N_19048);
and U19750 (N_19750,N_18741,N_18785);
or U19751 (N_19751,N_18692,N_19040);
nor U19752 (N_19752,N_18742,N_19193);
nand U19753 (N_19753,N_18966,N_19036);
xor U19754 (N_19754,N_19001,N_18968);
or U19755 (N_19755,N_18737,N_18867);
nor U19756 (N_19756,N_18635,N_18752);
or U19757 (N_19757,N_18923,N_18644);
xor U19758 (N_19758,N_18847,N_18731);
xnor U19759 (N_19759,N_18976,N_18886);
nor U19760 (N_19760,N_19020,N_18737);
and U19761 (N_19761,N_18949,N_18807);
nor U19762 (N_19762,N_19108,N_19148);
nor U19763 (N_19763,N_19099,N_19031);
or U19764 (N_19764,N_19040,N_18828);
xnor U19765 (N_19765,N_19062,N_18905);
xor U19766 (N_19766,N_19156,N_18613);
nor U19767 (N_19767,N_18753,N_19072);
nor U19768 (N_19768,N_18725,N_18637);
xor U19769 (N_19769,N_19147,N_18802);
and U19770 (N_19770,N_18957,N_19133);
nand U19771 (N_19771,N_19105,N_18898);
nor U19772 (N_19772,N_18940,N_19199);
or U19773 (N_19773,N_19044,N_18641);
xnor U19774 (N_19774,N_18878,N_19130);
and U19775 (N_19775,N_18855,N_18824);
or U19776 (N_19776,N_19128,N_18717);
xnor U19777 (N_19777,N_19152,N_18966);
or U19778 (N_19778,N_19018,N_18670);
xnor U19779 (N_19779,N_18828,N_19131);
nor U19780 (N_19780,N_18953,N_18957);
nor U19781 (N_19781,N_18726,N_18770);
nor U19782 (N_19782,N_19174,N_19095);
xor U19783 (N_19783,N_18937,N_18806);
or U19784 (N_19784,N_18885,N_19071);
xnor U19785 (N_19785,N_19107,N_19078);
nor U19786 (N_19786,N_18762,N_19120);
xor U19787 (N_19787,N_18698,N_19000);
or U19788 (N_19788,N_19016,N_18646);
nor U19789 (N_19789,N_18888,N_18928);
and U19790 (N_19790,N_19011,N_19099);
nor U19791 (N_19791,N_18636,N_19176);
xnor U19792 (N_19792,N_18647,N_19120);
nand U19793 (N_19793,N_18750,N_18965);
and U19794 (N_19794,N_18858,N_18973);
or U19795 (N_19795,N_19070,N_19105);
xor U19796 (N_19796,N_18668,N_18749);
or U19797 (N_19797,N_18737,N_18997);
and U19798 (N_19798,N_18745,N_18863);
and U19799 (N_19799,N_18630,N_19009);
xnor U19800 (N_19800,N_19511,N_19457);
xnor U19801 (N_19801,N_19697,N_19491);
nor U19802 (N_19802,N_19372,N_19402);
nand U19803 (N_19803,N_19753,N_19720);
or U19804 (N_19804,N_19740,N_19552);
and U19805 (N_19805,N_19713,N_19425);
xor U19806 (N_19806,N_19495,N_19761);
or U19807 (N_19807,N_19709,N_19238);
xor U19808 (N_19808,N_19261,N_19517);
nor U19809 (N_19809,N_19519,N_19514);
nor U19810 (N_19810,N_19437,N_19279);
nand U19811 (N_19811,N_19655,N_19695);
or U19812 (N_19812,N_19270,N_19274);
nand U19813 (N_19813,N_19742,N_19454);
and U19814 (N_19814,N_19275,N_19658);
nand U19815 (N_19815,N_19609,N_19217);
nand U19816 (N_19816,N_19555,N_19694);
nor U19817 (N_19817,N_19782,N_19232);
or U19818 (N_19818,N_19604,N_19775);
and U19819 (N_19819,N_19205,N_19470);
and U19820 (N_19820,N_19547,N_19717);
and U19821 (N_19821,N_19622,N_19605);
nand U19822 (N_19822,N_19202,N_19393);
xnor U19823 (N_19823,N_19318,N_19426);
nor U19824 (N_19824,N_19249,N_19591);
nand U19825 (N_19825,N_19749,N_19774);
xor U19826 (N_19826,N_19735,N_19567);
or U19827 (N_19827,N_19203,N_19421);
and U19828 (N_19828,N_19306,N_19209);
or U19829 (N_19829,N_19610,N_19502);
nand U19830 (N_19830,N_19583,N_19629);
and U19831 (N_19831,N_19588,N_19370);
nor U19832 (N_19832,N_19542,N_19452);
or U19833 (N_19833,N_19640,N_19615);
or U19834 (N_19834,N_19779,N_19710);
nand U19835 (N_19835,N_19660,N_19670);
and U19836 (N_19836,N_19215,N_19594);
xnor U19837 (N_19837,N_19265,N_19379);
or U19838 (N_19838,N_19330,N_19492);
xnor U19839 (N_19839,N_19763,N_19487);
and U19840 (N_19840,N_19561,N_19429);
nor U19841 (N_19841,N_19624,N_19786);
nor U19842 (N_19842,N_19407,N_19254);
xnor U19843 (N_19843,N_19651,N_19613);
and U19844 (N_19844,N_19500,N_19284);
and U19845 (N_19845,N_19637,N_19443);
xnor U19846 (N_19846,N_19439,N_19380);
and U19847 (N_19847,N_19549,N_19458);
xnor U19848 (N_19848,N_19332,N_19635);
xor U19849 (N_19849,N_19283,N_19724);
and U19850 (N_19850,N_19264,N_19718);
or U19851 (N_19851,N_19478,N_19577);
nor U19852 (N_19852,N_19490,N_19352);
nand U19853 (N_19853,N_19557,N_19772);
or U19854 (N_19854,N_19494,N_19391);
xnor U19855 (N_19855,N_19301,N_19731);
and U19856 (N_19856,N_19628,N_19516);
nor U19857 (N_19857,N_19218,N_19669);
nor U19858 (N_19858,N_19690,N_19676);
nor U19859 (N_19859,N_19785,N_19420);
xor U19860 (N_19860,N_19256,N_19445);
or U19861 (N_19861,N_19719,N_19755);
nand U19862 (N_19862,N_19553,N_19556);
xor U19863 (N_19863,N_19654,N_19367);
xor U19864 (N_19864,N_19508,N_19346);
nor U19865 (N_19865,N_19646,N_19444);
nand U19866 (N_19866,N_19705,N_19522);
or U19867 (N_19867,N_19277,N_19267);
xnor U19868 (N_19868,N_19228,N_19315);
xor U19869 (N_19869,N_19368,N_19224);
or U19870 (N_19870,N_19527,N_19608);
xnor U19871 (N_19871,N_19337,N_19585);
nand U19872 (N_19872,N_19392,N_19227);
xnor U19873 (N_19873,N_19754,N_19504);
nor U19874 (N_19874,N_19223,N_19533);
or U19875 (N_19875,N_19672,N_19349);
xor U19876 (N_19876,N_19448,N_19313);
nand U19877 (N_19877,N_19207,N_19276);
or U19878 (N_19878,N_19369,N_19258);
and U19879 (N_19879,N_19273,N_19331);
and U19880 (N_19880,N_19263,N_19317);
nor U19881 (N_19881,N_19463,N_19257);
nand U19882 (N_19882,N_19300,N_19278);
nor U19883 (N_19883,N_19399,N_19480);
or U19884 (N_19884,N_19663,N_19721);
nand U19885 (N_19885,N_19466,N_19353);
or U19886 (N_19886,N_19324,N_19680);
or U19887 (N_19887,N_19795,N_19506);
or U19888 (N_19888,N_19234,N_19389);
and U19889 (N_19889,N_19216,N_19348);
nand U19890 (N_19890,N_19736,N_19664);
nor U19891 (N_19891,N_19240,N_19312);
nand U19892 (N_19892,N_19387,N_19302);
and U19893 (N_19893,N_19250,N_19414);
nand U19894 (N_19894,N_19231,N_19418);
xnor U19895 (N_19895,N_19606,N_19411);
xnor U19896 (N_19896,N_19659,N_19638);
nand U19897 (N_19897,N_19550,N_19543);
or U19898 (N_19898,N_19416,N_19706);
nor U19899 (N_19899,N_19794,N_19206);
nor U19900 (N_19900,N_19639,N_19757);
and U19901 (N_19901,N_19350,N_19581);
nand U19902 (N_19902,N_19438,N_19599);
or U19903 (N_19903,N_19580,N_19469);
nand U19904 (N_19904,N_19220,N_19535);
nor U19905 (N_19905,N_19406,N_19509);
or U19906 (N_19906,N_19363,N_19376);
and U19907 (N_19907,N_19625,N_19771);
and U19908 (N_19908,N_19797,N_19401);
or U19909 (N_19909,N_19404,N_19489);
and U19910 (N_19910,N_19394,N_19518);
nor U19911 (N_19911,N_19688,N_19787);
nor U19912 (N_19912,N_19449,N_19326);
or U19913 (N_19913,N_19395,N_19684);
xor U19914 (N_19914,N_19462,N_19636);
xnor U19915 (N_19915,N_19356,N_19308);
nor U19916 (N_19916,N_19616,N_19582);
xor U19917 (N_19917,N_19481,N_19262);
xnor U19918 (N_19918,N_19311,N_19573);
xor U19919 (N_19919,N_19334,N_19653);
xnor U19920 (N_19920,N_19295,N_19722);
and U19921 (N_19921,N_19689,N_19623);
nor U19922 (N_19922,N_19716,N_19410);
xor U19923 (N_19923,N_19243,N_19540);
and U19924 (N_19924,N_19450,N_19428);
or U19925 (N_19925,N_19282,N_19575);
nor U19926 (N_19926,N_19687,N_19266);
nor U19927 (N_19927,N_19681,N_19351);
nand U19928 (N_19928,N_19596,N_19340);
and U19929 (N_19929,N_19385,N_19419);
nand U19930 (N_19930,N_19620,N_19560);
nor U19931 (N_19931,N_19280,N_19778);
or U19932 (N_19932,N_19298,N_19667);
xor U19933 (N_19933,N_19322,N_19335);
or U19934 (N_19934,N_19737,N_19403);
and U19935 (N_19935,N_19627,N_19378);
and U19936 (N_19936,N_19361,N_19612);
or U19937 (N_19937,N_19602,N_19345);
and U19938 (N_19938,N_19691,N_19729);
nand U19939 (N_19939,N_19255,N_19325);
xnor U19940 (N_19940,N_19472,N_19586);
xor U19941 (N_19941,N_19643,N_19661);
nand U19942 (N_19942,N_19656,N_19357);
or U19943 (N_19943,N_19631,N_19781);
or U19944 (N_19944,N_19520,N_19584);
nand U19945 (N_19945,N_19796,N_19388);
nand U19946 (N_19946,N_19479,N_19750);
or U19947 (N_19947,N_19513,N_19434);
or U19948 (N_19948,N_19532,N_19333);
nor U19949 (N_19949,N_19244,N_19601);
nand U19950 (N_19950,N_19728,N_19712);
xnor U19951 (N_19951,N_19734,N_19682);
xnor U19952 (N_19952,N_19521,N_19571);
and U19953 (N_19953,N_19748,N_19320);
and U19954 (N_19954,N_19590,N_19534);
nor U19955 (N_19955,N_19726,N_19446);
or U19956 (N_19956,N_19468,N_19642);
or U19957 (N_19957,N_19693,N_19292);
or U19958 (N_19958,N_19412,N_19536);
nand U19959 (N_19959,N_19679,N_19699);
and U19960 (N_19960,N_19291,N_19213);
nor U19961 (N_19961,N_19769,N_19529);
and U19962 (N_19962,N_19692,N_19537);
xnor U19963 (N_19963,N_19225,N_19751);
nand U19964 (N_19964,N_19743,N_19675);
or U19965 (N_19965,N_19593,N_19564);
and U19966 (N_19966,N_19386,N_19242);
and U19967 (N_19967,N_19526,N_19229);
nor U19968 (N_19968,N_19460,N_19245);
nor U19969 (N_19969,N_19666,N_19764);
nor U19970 (N_19970,N_19671,N_19545);
and U19971 (N_19971,N_19477,N_19467);
nor U19972 (N_19972,N_19396,N_19733);
and U19973 (N_19973,N_19436,N_19723);
nand U19974 (N_19974,N_19528,N_19600);
nand U19975 (N_19975,N_19465,N_19739);
nand U19976 (N_19976,N_19323,N_19607);
nor U19977 (N_19977,N_19503,N_19700);
nor U19978 (N_19978,N_19652,N_19569);
or U19979 (N_19979,N_19773,N_19711);
or U19980 (N_19980,N_19497,N_19461);
nor U19981 (N_19981,N_19767,N_19471);
nor U19982 (N_19982,N_19271,N_19548);
xor U19983 (N_19983,N_19515,N_19662);
xnor U19984 (N_19984,N_19563,N_19499);
nor U19985 (N_19985,N_19617,N_19630);
xnor U19986 (N_19986,N_19201,N_19741);
nor U19987 (N_19987,N_19756,N_19668);
xnor U19988 (N_19988,N_19762,N_19374);
nor U19989 (N_19989,N_19328,N_19725);
nor U19990 (N_19990,N_19214,N_19293);
and U19991 (N_19991,N_19373,N_19433);
and U19992 (N_19992,N_19568,N_19546);
and U19993 (N_19993,N_19641,N_19314);
nor U19994 (N_19994,N_19745,N_19704);
nand U19995 (N_19995,N_19299,N_19791);
nor U19996 (N_19996,N_19384,N_19336);
nand U19997 (N_19997,N_19305,N_19246);
nor U19998 (N_19998,N_19341,N_19377);
or U19999 (N_19999,N_19683,N_19297);
nor U20000 (N_20000,N_19342,N_19268);
xnor U20001 (N_20001,N_19677,N_19286);
nor U20002 (N_20002,N_19799,N_19765);
xnor U20003 (N_20003,N_19423,N_19365);
or U20004 (N_20004,N_19424,N_19674);
nand U20005 (N_20005,N_19714,N_19415);
xor U20006 (N_20006,N_19648,N_19747);
nor U20007 (N_20007,N_19304,N_19269);
and U20008 (N_20008,N_19746,N_19788);
and U20009 (N_20009,N_19212,N_19738);
nor U20010 (N_20010,N_19427,N_19432);
nor U20011 (N_20011,N_19364,N_19678);
and U20012 (N_20012,N_19290,N_19316);
or U20013 (N_20013,N_19633,N_19405);
nand U20014 (N_20014,N_19488,N_19760);
nor U20015 (N_20015,N_19707,N_19576);
and U20016 (N_20016,N_19589,N_19727);
nor U20017 (N_20017,N_19296,N_19210);
or U20018 (N_20018,N_19440,N_19559);
nand U20019 (N_20019,N_19579,N_19702);
nand U20020 (N_20020,N_19382,N_19598);
nand U20021 (N_20021,N_19338,N_19360);
nor U20022 (N_20022,N_19565,N_19759);
or U20023 (N_20023,N_19200,N_19241);
nand U20024 (N_20024,N_19701,N_19459);
or U20025 (N_20025,N_19456,N_19485);
and U20026 (N_20026,N_19474,N_19570);
and U20027 (N_20027,N_19248,N_19777);
nor U20028 (N_20028,N_19272,N_19219);
xor U20029 (N_20029,N_19347,N_19430);
nand U20030 (N_20030,N_19621,N_19222);
nand U20031 (N_20031,N_19447,N_19611);
or U20032 (N_20032,N_19650,N_19790);
xor U20033 (N_20033,N_19776,N_19355);
and U20034 (N_20034,N_19435,N_19233);
or U20035 (N_20035,N_19673,N_19507);
xnor U20036 (N_20036,N_19798,N_19783);
and U20037 (N_20037,N_19307,N_19685);
nand U20038 (N_20038,N_19319,N_19344);
and U20039 (N_20039,N_19732,N_19592);
nor U20040 (N_20040,N_19657,N_19285);
and U20041 (N_20041,N_19541,N_19758);
and U20042 (N_20042,N_19554,N_19486);
nand U20043 (N_20043,N_19383,N_19251);
nand U20044 (N_20044,N_19247,N_19789);
and U20045 (N_20045,N_19455,N_19398);
nand U20046 (N_20046,N_19354,N_19451);
xor U20047 (N_20047,N_19595,N_19371);
nand U20048 (N_20048,N_19343,N_19339);
or U20049 (N_20049,N_19260,N_19792);
or U20050 (N_20050,N_19366,N_19482);
xor U20051 (N_20051,N_19230,N_19259);
xor U20052 (N_20052,N_19730,N_19505);
nand U20053 (N_20053,N_19632,N_19498);
xnor U20054 (N_20054,N_19626,N_19686);
and U20055 (N_20055,N_19359,N_19597);
and U20056 (N_20056,N_19752,N_19551);
or U20057 (N_20057,N_19696,N_19390);
nand U20058 (N_20058,N_19362,N_19780);
and U20059 (N_20059,N_19281,N_19442);
xnor U20060 (N_20060,N_19523,N_19422);
and U20061 (N_20061,N_19310,N_19476);
xor U20062 (N_20062,N_19645,N_19539);
nor U20063 (N_20063,N_19558,N_19698);
nor U20064 (N_20064,N_19574,N_19634);
nor U20065 (N_20065,N_19400,N_19618);
nor U20066 (N_20066,N_19208,N_19397);
or U20067 (N_20067,N_19473,N_19289);
or U20068 (N_20068,N_19501,N_19484);
nor U20069 (N_20069,N_19744,N_19512);
or U20070 (N_20070,N_19409,N_19287);
or U20071 (N_20071,N_19294,N_19235);
xor U20072 (N_20072,N_19530,N_19309);
nand U20073 (N_20073,N_19793,N_19464);
nor U20074 (N_20074,N_19703,N_19572);
nor U20075 (N_20075,N_19538,N_19413);
or U20076 (N_20076,N_19578,N_19327);
or U20077 (N_20077,N_19562,N_19531);
xnor U20078 (N_20078,N_19239,N_19381);
nor U20079 (N_20079,N_19288,N_19544);
and U20080 (N_20080,N_19510,N_19766);
xnor U20081 (N_20081,N_19236,N_19603);
and U20082 (N_20082,N_19253,N_19375);
xnor U20083 (N_20083,N_19221,N_19358);
or U20084 (N_20084,N_19408,N_19715);
nand U20085 (N_20085,N_19252,N_19496);
xnor U20086 (N_20086,N_19784,N_19483);
and U20087 (N_20087,N_19770,N_19226);
or U20088 (N_20088,N_19665,N_19329);
or U20089 (N_20089,N_19644,N_19475);
nor U20090 (N_20090,N_19211,N_19525);
nor U20091 (N_20091,N_19647,N_19708);
or U20092 (N_20092,N_19431,N_19768);
nor U20093 (N_20093,N_19614,N_19524);
nand U20094 (N_20094,N_19493,N_19649);
or U20095 (N_20095,N_19619,N_19453);
nand U20096 (N_20096,N_19566,N_19303);
xor U20097 (N_20097,N_19321,N_19587);
xor U20098 (N_20098,N_19204,N_19237);
nor U20099 (N_20099,N_19417,N_19441);
nand U20100 (N_20100,N_19517,N_19231);
nor U20101 (N_20101,N_19638,N_19673);
nand U20102 (N_20102,N_19363,N_19763);
xor U20103 (N_20103,N_19453,N_19753);
and U20104 (N_20104,N_19309,N_19670);
xor U20105 (N_20105,N_19718,N_19311);
nand U20106 (N_20106,N_19610,N_19243);
xor U20107 (N_20107,N_19357,N_19326);
xnor U20108 (N_20108,N_19213,N_19614);
and U20109 (N_20109,N_19687,N_19607);
xor U20110 (N_20110,N_19720,N_19234);
or U20111 (N_20111,N_19265,N_19424);
and U20112 (N_20112,N_19201,N_19711);
nand U20113 (N_20113,N_19564,N_19531);
or U20114 (N_20114,N_19677,N_19325);
xor U20115 (N_20115,N_19554,N_19426);
or U20116 (N_20116,N_19560,N_19335);
and U20117 (N_20117,N_19246,N_19601);
xor U20118 (N_20118,N_19438,N_19653);
nand U20119 (N_20119,N_19584,N_19305);
and U20120 (N_20120,N_19236,N_19702);
or U20121 (N_20121,N_19284,N_19281);
or U20122 (N_20122,N_19463,N_19415);
and U20123 (N_20123,N_19669,N_19343);
and U20124 (N_20124,N_19517,N_19690);
nand U20125 (N_20125,N_19410,N_19549);
or U20126 (N_20126,N_19798,N_19444);
nor U20127 (N_20127,N_19400,N_19477);
and U20128 (N_20128,N_19306,N_19651);
or U20129 (N_20129,N_19336,N_19227);
and U20130 (N_20130,N_19347,N_19734);
and U20131 (N_20131,N_19315,N_19658);
or U20132 (N_20132,N_19697,N_19629);
or U20133 (N_20133,N_19284,N_19733);
and U20134 (N_20134,N_19235,N_19622);
xnor U20135 (N_20135,N_19261,N_19490);
nor U20136 (N_20136,N_19378,N_19448);
xor U20137 (N_20137,N_19593,N_19411);
and U20138 (N_20138,N_19426,N_19439);
or U20139 (N_20139,N_19772,N_19616);
xor U20140 (N_20140,N_19648,N_19532);
or U20141 (N_20141,N_19213,N_19602);
xnor U20142 (N_20142,N_19489,N_19730);
nand U20143 (N_20143,N_19576,N_19329);
nor U20144 (N_20144,N_19755,N_19589);
nor U20145 (N_20145,N_19638,N_19637);
nand U20146 (N_20146,N_19512,N_19442);
nor U20147 (N_20147,N_19316,N_19677);
xor U20148 (N_20148,N_19361,N_19724);
nor U20149 (N_20149,N_19675,N_19224);
nand U20150 (N_20150,N_19764,N_19418);
or U20151 (N_20151,N_19476,N_19716);
and U20152 (N_20152,N_19523,N_19671);
and U20153 (N_20153,N_19474,N_19383);
xnor U20154 (N_20154,N_19561,N_19458);
and U20155 (N_20155,N_19673,N_19593);
or U20156 (N_20156,N_19690,N_19696);
or U20157 (N_20157,N_19209,N_19693);
xor U20158 (N_20158,N_19636,N_19488);
and U20159 (N_20159,N_19381,N_19371);
xor U20160 (N_20160,N_19556,N_19566);
or U20161 (N_20161,N_19281,N_19472);
xor U20162 (N_20162,N_19362,N_19347);
and U20163 (N_20163,N_19648,N_19738);
or U20164 (N_20164,N_19557,N_19512);
nand U20165 (N_20165,N_19591,N_19437);
nor U20166 (N_20166,N_19654,N_19358);
and U20167 (N_20167,N_19480,N_19209);
nand U20168 (N_20168,N_19302,N_19581);
nand U20169 (N_20169,N_19464,N_19332);
and U20170 (N_20170,N_19479,N_19474);
or U20171 (N_20171,N_19728,N_19535);
nand U20172 (N_20172,N_19305,N_19520);
and U20173 (N_20173,N_19546,N_19773);
nand U20174 (N_20174,N_19442,N_19485);
and U20175 (N_20175,N_19592,N_19407);
or U20176 (N_20176,N_19406,N_19201);
and U20177 (N_20177,N_19581,N_19646);
nand U20178 (N_20178,N_19282,N_19256);
and U20179 (N_20179,N_19636,N_19448);
xor U20180 (N_20180,N_19372,N_19292);
nor U20181 (N_20181,N_19420,N_19742);
or U20182 (N_20182,N_19299,N_19214);
xor U20183 (N_20183,N_19527,N_19223);
nand U20184 (N_20184,N_19279,N_19413);
or U20185 (N_20185,N_19478,N_19633);
and U20186 (N_20186,N_19480,N_19343);
or U20187 (N_20187,N_19668,N_19339);
nor U20188 (N_20188,N_19208,N_19510);
nor U20189 (N_20189,N_19515,N_19346);
or U20190 (N_20190,N_19504,N_19524);
nand U20191 (N_20191,N_19290,N_19543);
or U20192 (N_20192,N_19515,N_19752);
nor U20193 (N_20193,N_19318,N_19591);
or U20194 (N_20194,N_19664,N_19546);
or U20195 (N_20195,N_19514,N_19532);
nand U20196 (N_20196,N_19418,N_19279);
and U20197 (N_20197,N_19707,N_19325);
nor U20198 (N_20198,N_19708,N_19465);
nor U20199 (N_20199,N_19560,N_19341);
nand U20200 (N_20200,N_19496,N_19509);
or U20201 (N_20201,N_19317,N_19426);
nor U20202 (N_20202,N_19769,N_19538);
or U20203 (N_20203,N_19794,N_19543);
or U20204 (N_20204,N_19516,N_19225);
and U20205 (N_20205,N_19204,N_19491);
nor U20206 (N_20206,N_19237,N_19416);
nand U20207 (N_20207,N_19358,N_19525);
nand U20208 (N_20208,N_19564,N_19348);
or U20209 (N_20209,N_19303,N_19250);
and U20210 (N_20210,N_19340,N_19469);
or U20211 (N_20211,N_19583,N_19404);
and U20212 (N_20212,N_19259,N_19386);
and U20213 (N_20213,N_19639,N_19398);
or U20214 (N_20214,N_19496,N_19711);
xor U20215 (N_20215,N_19239,N_19307);
nor U20216 (N_20216,N_19371,N_19786);
or U20217 (N_20217,N_19661,N_19610);
xor U20218 (N_20218,N_19227,N_19363);
nor U20219 (N_20219,N_19779,N_19673);
or U20220 (N_20220,N_19353,N_19798);
nor U20221 (N_20221,N_19466,N_19288);
and U20222 (N_20222,N_19425,N_19698);
and U20223 (N_20223,N_19634,N_19711);
or U20224 (N_20224,N_19332,N_19735);
nor U20225 (N_20225,N_19636,N_19505);
xor U20226 (N_20226,N_19560,N_19413);
nor U20227 (N_20227,N_19680,N_19443);
nor U20228 (N_20228,N_19562,N_19469);
nand U20229 (N_20229,N_19686,N_19442);
xor U20230 (N_20230,N_19437,N_19734);
xnor U20231 (N_20231,N_19735,N_19235);
or U20232 (N_20232,N_19254,N_19219);
nand U20233 (N_20233,N_19272,N_19542);
nor U20234 (N_20234,N_19232,N_19400);
xnor U20235 (N_20235,N_19546,N_19776);
nor U20236 (N_20236,N_19446,N_19496);
nand U20237 (N_20237,N_19776,N_19493);
nand U20238 (N_20238,N_19272,N_19635);
xor U20239 (N_20239,N_19787,N_19547);
nand U20240 (N_20240,N_19429,N_19347);
xor U20241 (N_20241,N_19618,N_19475);
nand U20242 (N_20242,N_19607,N_19582);
xor U20243 (N_20243,N_19613,N_19553);
and U20244 (N_20244,N_19413,N_19312);
or U20245 (N_20245,N_19644,N_19499);
xnor U20246 (N_20246,N_19625,N_19283);
xor U20247 (N_20247,N_19695,N_19629);
or U20248 (N_20248,N_19742,N_19388);
and U20249 (N_20249,N_19560,N_19751);
nor U20250 (N_20250,N_19611,N_19425);
nor U20251 (N_20251,N_19723,N_19509);
and U20252 (N_20252,N_19685,N_19261);
xor U20253 (N_20253,N_19635,N_19527);
nor U20254 (N_20254,N_19299,N_19730);
nand U20255 (N_20255,N_19446,N_19550);
xor U20256 (N_20256,N_19375,N_19232);
and U20257 (N_20257,N_19483,N_19393);
nand U20258 (N_20258,N_19359,N_19289);
and U20259 (N_20259,N_19266,N_19531);
and U20260 (N_20260,N_19387,N_19676);
or U20261 (N_20261,N_19433,N_19645);
or U20262 (N_20262,N_19752,N_19738);
xnor U20263 (N_20263,N_19776,N_19276);
and U20264 (N_20264,N_19453,N_19326);
nand U20265 (N_20265,N_19316,N_19634);
and U20266 (N_20266,N_19435,N_19539);
or U20267 (N_20267,N_19534,N_19206);
nor U20268 (N_20268,N_19269,N_19710);
nor U20269 (N_20269,N_19262,N_19799);
nand U20270 (N_20270,N_19250,N_19621);
xor U20271 (N_20271,N_19273,N_19619);
and U20272 (N_20272,N_19608,N_19681);
nor U20273 (N_20273,N_19386,N_19569);
and U20274 (N_20274,N_19437,N_19739);
and U20275 (N_20275,N_19746,N_19318);
nand U20276 (N_20276,N_19334,N_19491);
and U20277 (N_20277,N_19532,N_19201);
or U20278 (N_20278,N_19551,N_19334);
nor U20279 (N_20279,N_19283,N_19513);
nor U20280 (N_20280,N_19772,N_19319);
or U20281 (N_20281,N_19232,N_19667);
nor U20282 (N_20282,N_19219,N_19557);
and U20283 (N_20283,N_19490,N_19389);
xor U20284 (N_20284,N_19689,N_19584);
nor U20285 (N_20285,N_19204,N_19699);
nor U20286 (N_20286,N_19244,N_19428);
or U20287 (N_20287,N_19260,N_19278);
xnor U20288 (N_20288,N_19356,N_19741);
nor U20289 (N_20289,N_19397,N_19720);
xnor U20290 (N_20290,N_19666,N_19625);
and U20291 (N_20291,N_19719,N_19273);
nand U20292 (N_20292,N_19620,N_19602);
or U20293 (N_20293,N_19644,N_19431);
nor U20294 (N_20294,N_19508,N_19588);
xor U20295 (N_20295,N_19496,N_19793);
nand U20296 (N_20296,N_19342,N_19299);
and U20297 (N_20297,N_19363,N_19547);
or U20298 (N_20298,N_19672,N_19532);
or U20299 (N_20299,N_19279,N_19659);
xor U20300 (N_20300,N_19433,N_19222);
or U20301 (N_20301,N_19420,N_19331);
and U20302 (N_20302,N_19399,N_19386);
nor U20303 (N_20303,N_19433,N_19344);
or U20304 (N_20304,N_19464,N_19667);
nand U20305 (N_20305,N_19513,N_19278);
nand U20306 (N_20306,N_19282,N_19342);
nand U20307 (N_20307,N_19233,N_19758);
nand U20308 (N_20308,N_19205,N_19784);
or U20309 (N_20309,N_19308,N_19540);
nand U20310 (N_20310,N_19592,N_19329);
nand U20311 (N_20311,N_19611,N_19535);
and U20312 (N_20312,N_19764,N_19319);
nand U20313 (N_20313,N_19612,N_19582);
xor U20314 (N_20314,N_19322,N_19784);
nor U20315 (N_20315,N_19355,N_19634);
xor U20316 (N_20316,N_19461,N_19722);
nor U20317 (N_20317,N_19382,N_19634);
or U20318 (N_20318,N_19612,N_19784);
nor U20319 (N_20319,N_19463,N_19429);
nor U20320 (N_20320,N_19219,N_19338);
xor U20321 (N_20321,N_19292,N_19370);
and U20322 (N_20322,N_19582,N_19542);
xor U20323 (N_20323,N_19425,N_19637);
nand U20324 (N_20324,N_19563,N_19569);
and U20325 (N_20325,N_19266,N_19267);
or U20326 (N_20326,N_19254,N_19324);
xnor U20327 (N_20327,N_19607,N_19537);
xnor U20328 (N_20328,N_19620,N_19473);
or U20329 (N_20329,N_19343,N_19261);
nor U20330 (N_20330,N_19314,N_19289);
nand U20331 (N_20331,N_19786,N_19512);
xor U20332 (N_20332,N_19423,N_19503);
xnor U20333 (N_20333,N_19460,N_19691);
nor U20334 (N_20334,N_19366,N_19437);
nor U20335 (N_20335,N_19619,N_19612);
and U20336 (N_20336,N_19676,N_19694);
and U20337 (N_20337,N_19202,N_19713);
xnor U20338 (N_20338,N_19607,N_19755);
xnor U20339 (N_20339,N_19354,N_19226);
nor U20340 (N_20340,N_19297,N_19562);
nor U20341 (N_20341,N_19301,N_19365);
and U20342 (N_20342,N_19634,N_19413);
nand U20343 (N_20343,N_19648,N_19370);
and U20344 (N_20344,N_19669,N_19230);
or U20345 (N_20345,N_19362,N_19431);
or U20346 (N_20346,N_19714,N_19553);
nand U20347 (N_20347,N_19558,N_19702);
nand U20348 (N_20348,N_19393,N_19201);
and U20349 (N_20349,N_19201,N_19281);
and U20350 (N_20350,N_19210,N_19386);
xnor U20351 (N_20351,N_19210,N_19706);
nand U20352 (N_20352,N_19742,N_19413);
and U20353 (N_20353,N_19795,N_19410);
xnor U20354 (N_20354,N_19764,N_19393);
nand U20355 (N_20355,N_19432,N_19213);
nand U20356 (N_20356,N_19762,N_19306);
or U20357 (N_20357,N_19348,N_19780);
xnor U20358 (N_20358,N_19412,N_19251);
xor U20359 (N_20359,N_19550,N_19684);
nand U20360 (N_20360,N_19779,N_19258);
or U20361 (N_20361,N_19435,N_19494);
xor U20362 (N_20362,N_19417,N_19656);
nor U20363 (N_20363,N_19597,N_19444);
xnor U20364 (N_20364,N_19426,N_19289);
and U20365 (N_20365,N_19351,N_19385);
and U20366 (N_20366,N_19303,N_19588);
nor U20367 (N_20367,N_19493,N_19481);
nor U20368 (N_20368,N_19455,N_19777);
nand U20369 (N_20369,N_19756,N_19583);
and U20370 (N_20370,N_19718,N_19791);
and U20371 (N_20371,N_19334,N_19561);
xnor U20372 (N_20372,N_19415,N_19591);
or U20373 (N_20373,N_19580,N_19224);
nor U20374 (N_20374,N_19373,N_19331);
and U20375 (N_20375,N_19357,N_19548);
or U20376 (N_20376,N_19678,N_19592);
or U20377 (N_20377,N_19390,N_19619);
nand U20378 (N_20378,N_19449,N_19260);
or U20379 (N_20379,N_19513,N_19290);
nor U20380 (N_20380,N_19256,N_19237);
or U20381 (N_20381,N_19643,N_19427);
xnor U20382 (N_20382,N_19771,N_19248);
xor U20383 (N_20383,N_19797,N_19718);
nand U20384 (N_20384,N_19480,N_19239);
nand U20385 (N_20385,N_19698,N_19538);
or U20386 (N_20386,N_19292,N_19261);
nor U20387 (N_20387,N_19745,N_19215);
nand U20388 (N_20388,N_19598,N_19346);
or U20389 (N_20389,N_19686,N_19486);
nand U20390 (N_20390,N_19612,N_19237);
nand U20391 (N_20391,N_19698,N_19271);
and U20392 (N_20392,N_19774,N_19543);
nor U20393 (N_20393,N_19308,N_19452);
xnor U20394 (N_20394,N_19424,N_19439);
xnor U20395 (N_20395,N_19249,N_19505);
or U20396 (N_20396,N_19416,N_19618);
or U20397 (N_20397,N_19579,N_19615);
nand U20398 (N_20398,N_19308,N_19373);
xor U20399 (N_20399,N_19225,N_19549);
nand U20400 (N_20400,N_20353,N_20388);
xor U20401 (N_20401,N_20049,N_19913);
xnor U20402 (N_20402,N_20012,N_20072);
nor U20403 (N_20403,N_20390,N_19863);
nand U20404 (N_20404,N_20007,N_20392);
or U20405 (N_20405,N_19938,N_20336);
nand U20406 (N_20406,N_19847,N_19836);
nand U20407 (N_20407,N_20308,N_19823);
and U20408 (N_20408,N_19888,N_20151);
nand U20409 (N_20409,N_19957,N_20349);
nand U20410 (N_20410,N_20249,N_20378);
nand U20411 (N_20411,N_20071,N_19914);
and U20412 (N_20412,N_19831,N_20138);
or U20413 (N_20413,N_20347,N_19887);
and U20414 (N_20414,N_20203,N_19880);
nand U20415 (N_20415,N_20381,N_20396);
and U20416 (N_20416,N_20002,N_19993);
nor U20417 (N_20417,N_20316,N_20387);
and U20418 (N_20418,N_20334,N_19974);
or U20419 (N_20419,N_20332,N_19929);
and U20420 (N_20420,N_19967,N_19984);
xnor U20421 (N_20421,N_19804,N_20127);
and U20422 (N_20422,N_19899,N_20220);
nor U20423 (N_20423,N_19944,N_20222);
nor U20424 (N_20424,N_20078,N_20043);
nor U20425 (N_20425,N_20016,N_20257);
xor U20426 (N_20426,N_20196,N_20017);
nand U20427 (N_20427,N_19936,N_19969);
or U20428 (N_20428,N_19966,N_20258);
nor U20429 (N_20429,N_19864,N_20179);
nor U20430 (N_20430,N_20070,N_20094);
or U20431 (N_20431,N_20324,N_20097);
or U20432 (N_20432,N_20134,N_20194);
nand U20433 (N_20433,N_19833,N_20224);
nor U20434 (N_20434,N_19881,N_19801);
nor U20435 (N_20435,N_19932,N_20100);
xnor U20436 (N_20436,N_20109,N_19933);
xor U20437 (N_20437,N_20093,N_19806);
nor U20438 (N_20438,N_20310,N_19849);
nor U20439 (N_20439,N_20040,N_19965);
nor U20440 (N_20440,N_19991,N_19977);
nand U20441 (N_20441,N_19852,N_20338);
nand U20442 (N_20442,N_20216,N_20342);
and U20443 (N_20443,N_20162,N_19941);
nand U20444 (N_20444,N_20247,N_19908);
or U20445 (N_20445,N_20362,N_20340);
nor U20446 (N_20446,N_20176,N_20377);
nor U20447 (N_20447,N_19816,N_20372);
and U20448 (N_20448,N_20357,N_20114);
or U20449 (N_20449,N_20395,N_20294);
and U20450 (N_20450,N_20241,N_20158);
xnor U20451 (N_20451,N_19889,N_19937);
or U20452 (N_20452,N_20231,N_19988);
and U20453 (N_20453,N_20269,N_20025);
xnor U20454 (N_20454,N_20149,N_20036);
nor U20455 (N_20455,N_19999,N_19918);
or U20456 (N_20456,N_19963,N_20397);
or U20457 (N_20457,N_20175,N_19808);
and U20458 (N_20458,N_19825,N_19923);
nor U20459 (N_20459,N_20359,N_19939);
or U20460 (N_20460,N_20282,N_19931);
and U20461 (N_20461,N_20237,N_19903);
and U20462 (N_20462,N_19953,N_20370);
or U20463 (N_20463,N_19942,N_20126);
nor U20464 (N_20464,N_19878,N_20195);
or U20465 (N_20465,N_20321,N_20099);
and U20466 (N_20466,N_19870,N_19829);
xor U20467 (N_20467,N_20250,N_20183);
or U20468 (N_20468,N_20335,N_20329);
nor U20469 (N_20469,N_20364,N_20223);
or U20470 (N_20470,N_20302,N_20084);
or U20471 (N_20471,N_20000,N_19834);
and U20472 (N_20472,N_19990,N_19884);
xnor U20473 (N_20473,N_20004,N_20188);
xnor U20474 (N_20474,N_20339,N_20135);
nand U20475 (N_20475,N_20150,N_20037);
nand U20476 (N_20476,N_20119,N_20271);
xnor U20477 (N_20477,N_19983,N_20113);
and U20478 (N_20478,N_20356,N_20337);
xor U20479 (N_20479,N_19810,N_19869);
nand U20480 (N_20480,N_19827,N_19905);
nand U20481 (N_20481,N_19911,N_19940);
nand U20482 (N_20482,N_20140,N_20273);
nor U20483 (N_20483,N_20184,N_20058);
xnor U20484 (N_20484,N_20024,N_20199);
or U20485 (N_20485,N_20115,N_20023);
xnor U20486 (N_20486,N_19835,N_20259);
nor U20487 (N_20487,N_20173,N_19978);
or U20488 (N_20488,N_20219,N_19845);
and U20489 (N_20489,N_19982,N_20028);
and U20490 (N_20490,N_20276,N_19960);
or U20491 (N_20491,N_20108,N_19997);
and U20492 (N_20492,N_20101,N_20117);
nor U20493 (N_20493,N_20076,N_19925);
nand U20494 (N_20494,N_19964,N_20155);
and U20495 (N_20495,N_20112,N_20165);
xnor U20496 (N_20496,N_20105,N_20122);
and U20497 (N_20497,N_19976,N_20297);
xor U20498 (N_20498,N_20305,N_20055);
and U20499 (N_20499,N_20283,N_20146);
or U20500 (N_20500,N_20225,N_19853);
and U20501 (N_20501,N_20205,N_19865);
nor U20502 (N_20502,N_19901,N_19981);
nor U20503 (N_20503,N_20020,N_20299);
and U20504 (N_20504,N_20301,N_20379);
nor U20505 (N_20505,N_20064,N_20029);
nand U20506 (N_20506,N_20263,N_19876);
or U20507 (N_20507,N_20344,N_20075);
or U20508 (N_20508,N_19809,N_20198);
xnor U20509 (N_20509,N_20267,N_20256);
nor U20510 (N_20510,N_20345,N_20186);
and U20511 (N_20511,N_19951,N_20021);
nand U20512 (N_20512,N_20001,N_19874);
or U20513 (N_20513,N_19850,N_20323);
nand U20514 (N_20514,N_20048,N_19920);
xor U20515 (N_20515,N_19935,N_20069);
nand U20516 (N_20516,N_20209,N_20154);
xor U20517 (N_20517,N_19952,N_20272);
and U20518 (N_20518,N_19972,N_19821);
and U20519 (N_20519,N_20382,N_19996);
nand U20520 (N_20520,N_20130,N_20365);
nand U20521 (N_20521,N_19985,N_20252);
and U20522 (N_20522,N_20217,N_20110);
xor U20523 (N_20523,N_20202,N_19915);
nand U20524 (N_20524,N_20125,N_20383);
and U20525 (N_20525,N_20009,N_20062);
and U20526 (N_20526,N_20238,N_20380);
or U20527 (N_20527,N_19882,N_20330);
and U20528 (N_20528,N_19896,N_19954);
or U20529 (N_20529,N_20065,N_20056);
nor U20530 (N_20530,N_19818,N_20011);
and U20531 (N_20531,N_20348,N_20102);
nand U20532 (N_20532,N_19945,N_20088);
xor U20533 (N_20533,N_20170,N_20030);
nand U20534 (N_20534,N_20368,N_20264);
xnor U20535 (N_20535,N_19907,N_20228);
xor U20536 (N_20536,N_20248,N_20081);
nand U20537 (N_20537,N_20177,N_20018);
nand U20538 (N_20538,N_20089,N_20307);
or U20539 (N_20539,N_20235,N_19934);
nand U20540 (N_20540,N_19946,N_20240);
and U20541 (N_20541,N_20187,N_20211);
nand U20542 (N_20542,N_20006,N_19832);
or U20543 (N_20543,N_20193,N_20274);
nor U20544 (N_20544,N_19891,N_20287);
and U20545 (N_20545,N_20068,N_19839);
or U20546 (N_20546,N_20035,N_20019);
nor U20547 (N_20547,N_19838,N_20229);
or U20548 (N_20548,N_20346,N_20375);
nand U20549 (N_20549,N_20005,N_20083);
nand U20550 (N_20550,N_19987,N_20124);
xor U20551 (N_20551,N_20128,N_19958);
and U20552 (N_20552,N_20210,N_19830);
xor U20553 (N_20553,N_20373,N_20201);
xor U20554 (N_20554,N_19861,N_20369);
xnor U20555 (N_20555,N_20074,N_19851);
xnor U20556 (N_20556,N_20171,N_19860);
or U20557 (N_20557,N_19926,N_20098);
xor U20558 (N_20558,N_19854,N_19986);
xnor U20559 (N_20559,N_19924,N_20285);
nor U20560 (N_20560,N_20014,N_19970);
or U20561 (N_20561,N_19802,N_20277);
xor U20562 (N_20562,N_20385,N_20360);
nor U20563 (N_20563,N_19930,N_19877);
or U20564 (N_20564,N_20139,N_20057);
and U20565 (N_20565,N_19815,N_20262);
nand U20566 (N_20566,N_20157,N_20279);
nand U20567 (N_20567,N_20358,N_20161);
nor U20568 (N_20568,N_19900,N_20244);
xnor U20569 (N_20569,N_20137,N_19895);
xor U20570 (N_20570,N_20082,N_19968);
nand U20571 (N_20571,N_20166,N_20152);
nor U20572 (N_20572,N_20090,N_20280);
or U20573 (N_20573,N_20313,N_19959);
or U20574 (N_20574,N_20042,N_20221);
or U20575 (N_20575,N_20132,N_20092);
nand U20576 (N_20576,N_19826,N_19961);
nand U20577 (N_20577,N_20278,N_19928);
or U20578 (N_20578,N_20104,N_19943);
xnor U20579 (N_20579,N_20376,N_20164);
nand U20580 (N_20580,N_19846,N_19975);
and U20581 (N_20581,N_20296,N_20145);
nand U20582 (N_20582,N_20226,N_19822);
and U20583 (N_20583,N_20053,N_19948);
xnor U20584 (N_20584,N_20213,N_20087);
nor U20585 (N_20585,N_20207,N_20354);
and U20586 (N_20586,N_20163,N_20121);
xor U20587 (N_20587,N_20236,N_20169);
or U20588 (N_20588,N_20319,N_20208);
or U20589 (N_20589,N_19820,N_20077);
or U20590 (N_20590,N_20254,N_19885);
nor U20591 (N_20591,N_20003,N_20051);
nand U20592 (N_20592,N_19910,N_20391);
xnor U20593 (N_20593,N_20218,N_20026);
nor U20594 (N_20594,N_20041,N_20133);
and U20595 (N_20595,N_20059,N_20160);
nand U20596 (N_20596,N_20174,N_20239);
nor U20597 (N_20597,N_20034,N_20320);
or U20598 (N_20598,N_20111,N_19824);
nor U20599 (N_20599,N_20233,N_20144);
nor U20600 (N_20600,N_19902,N_20061);
and U20601 (N_20601,N_19921,N_20182);
nand U20602 (N_20602,N_20143,N_20047);
nand U20603 (N_20603,N_20118,N_20178);
nand U20604 (N_20604,N_19956,N_19916);
xnor U20605 (N_20605,N_20046,N_20107);
and U20606 (N_20606,N_20168,N_19909);
or U20607 (N_20607,N_19868,N_20243);
nand U20608 (N_20608,N_19859,N_20120);
or U20609 (N_20609,N_20331,N_20204);
nand U20610 (N_20610,N_20079,N_19904);
and U20611 (N_20611,N_20322,N_19980);
and U20612 (N_20612,N_19994,N_19867);
nor U20613 (N_20613,N_20350,N_20245);
nand U20614 (N_20614,N_19848,N_20291);
nand U20615 (N_20615,N_20399,N_20292);
nand U20616 (N_20616,N_20190,N_20015);
and U20617 (N_20617,N_20371,N_19893);
or U20618 (N_20618,N_19992,N_20141);
nand U20619 (N_20619,N_19947,N_20398);
xor U20620 (N_20620,N_20281,N_19883);
and U20621 (N_20621,N_19995,N_19949);
nand U20622 (N_20622,N_20333,N_19856);
nor U20623 (N_20623,N_20136,N_20284);
and U20624 (N_20624,N_19873,N_20214);
nand U20625 (N_20625,N_20032,N_20167);
nand U20626 (N_20626,N_20351,N_20343);
and U20627 (N_20627,N_20085,N_20159);
nor U20628 (N_20628,N_20010,N_20073);
nor U20629 (N_20629,N_19828,N_20095);
nor U20630 (N_20630,N_20363,N_19855);
nand U20631 (N_20631,N_19950,N_19927);
nor U20632 (N_20632,N_20008,N_20386);
and U20633 (N_20633,N_19955,N_20246);
nor U20634 (N_20634,N_20215,N_20148);
or U20635 (N_20635,N_19875,N_19858);
or U20636 (N_20636,N_20044,N_20289);
or U20637 (N_20637,N_19892,N_19998);
nor U20638 (N_20638,N_20227,N_20147);
nand U20639 (N_20639,N_20013,N_19971);
or U20640 (N_20640,N_20268,N_20066);
nor U20641 (N_20641,N_20086,N_20266);
nor U20642 (N_20642,N_20290,N_20315);
nor U20643 (N_20643,N_20131,N_20185);
xnor U20644 (N_20644,N_20311,N_20142);
or U20645 (N_20645,N_20096,N_19989);
and U20646 (N_20646,N_20116,N_20156);
nor U20647 (N_20647,N_20031,N_19843);
and U20648 (N_20648,N_19886,N_20050);
and U20649 (N_20649,N_19890,N_20123);
and U20650 (N_20650,N_20253,N_20341);
and U20651 (N_20651,N_20255,N_20038);
or U20652 (N_20652,N_20295,N_20197);
or U20653 (N_20653,N_19805,N_20033);
nand U20654 (N_20654,N_19894,N_19917);
and U20655 (N_20655,N_19879,N_20153);
or U20656 (N_20656,N_20293,N_19973);
xnor U20657 (N_20657,N_20327,N_20180);
nand U20658 (N_20658,N_19819,N_20027);
nor U20659 (N_20659,N_20103,N_20052);
nand U20660 (N_20660,N_20172,N_20304);
or U20661 (N_20661,N_20251,N_20181);
nor U20662 (N_20662,N_20384,N_20206);
and U20663 (N_20663,N_19862,N_19813);
nor U20664 (N_20664,N_20232,N_20200);
nand U20665 (N_20665,N_20192,N_19871);
or U20666 (N_20666,N_20063,N_20306);
and U20667 (N_20667,N_19979,N_20309);
and U20668 (N_20668,N_20234,N_20374);
or U20669 (N_20669,N_20328,N_20080);
nor U20670 (N_20670,N_20367,N_19817);
or U20671 (N_20671,N_20129,N_20260);
or U20672 (N_20672,N_19814,N_20298);
nand U20673 (N_20673,N_20230,N_20261);
or U20674 (N_20674,N_20286,N_20300);
and U20675 (N_20675,N_19800,N_20317);
xnor U20676 (N_20676,N_19807,N_19803);
or U20677 (N_20677,N_20242,N_20326);
nand U20678 (N_20678,N_20361,N_19857);
nor U20679 (N_20679,N_20106,N_19872);
nand U20680 (N_20680,N_20191,N_19898);
or U20681 (N_20681,N_20312,N_20045);
nor U20682 (N_20682,N_19812,N_19906);
xor U20683 (N_20683,N_19866,N_20288);
and U20684 (N_20684,N_20394,N_19919);
xnor U20685 (N_20685,N_20366,N_20022);
and U20686 (N_20686,N_19842,N_20054);
or U20687 (N_20687,N_20314,N_20325);
nor U20688 (N_20688,N_20091,N_20303);
and U20689 (N_20689,N_20060,N_20270);
and U20690 (N_20690,N_19912,N_20275);
xnor U20691 (N_20691,N_19962,N_19922);
or U20692 (N_20692,N_20393,N_19841);
nand U20693 (N_20693,N_19840,N_19837);
nand U20694 (N_20694,N_20067,N_20265);
xor U20695 (N_20695,N_20039,N_20355);
nor U20696 (N_20696,N_20352,N_20189);
xnor U20697 (N_20697,N_20318,N_19811);
or U20698 (N_20698,N_19897,N_20389);
and U20699 (N_20699,N_19844,N_20212);
nand U20700 (N_20700,N_20390,N_20204);
and U20701 (N_20701,N_20200,N_19963);
and U20702 (N_20702,N_20112,N_19940);
xor U20703 (N_20703,N_20340,N_20272);
nand U20704 (N_20704,N_19819,N_20297);
or U20705 (N_20705,N_20239,N_20220);
and U20706 (N_20706,N_19836,N_20012);
nand U20707 (N_20707,N_20007,N_20327);
and U20708 (N_20708,N_20378,N_20038);
xnor U20709 (N_20709,N_20297,N_20055);
or U20710 (N_20710,N_20216,N_20232);
xor U20711 (N_20711,N_20275,N_20130);
or U20712 (N_20712,N_20214,N_19825);
and U20713 (N_20713,N_20161,N_19829);
nor U20714 (N_20714,N_20056,N_20286);
or U20715 (N_20715,N_19899,N_19853);
xor U20716 (N_20716,N_20096,N_19884);
or U20717 (N_20717,N_20115,N_20390);
or U20718 (N_20718,N_20296,N_19895);
nand U20719 (N_20719,N_20266,N_20307);
nor U20720 (N_20720,N_20337,N_19964);
xor U20721 (N_20721,N_19930,N_20299);
nand U20722 (N_20722,N_19938,N_20267);
or U20723 (N_20723,N_19998,N_20311);
xor U20724 (N_20724,N_20166,N_20274);
or U20725 (N_20725,N_20087,N_20155);
nand U20726 (N_20726,N_20048,N_20172);
nor U20727 (N_20727,N_19831,N_19860);
nand U20728 (N_20728,N_20056,N_20084);
nand U20729 (N_20729,N_19974,N_20295);
xnor U20730 (N_20730,N_19837,N_20340);
or U20731 (N_20731,N_19895,N_19812);
xor U20732 (N_20732,N_20349,N_19808);
xor U20733 (N_20733,N_19831,N_20173);
nand U20734 (N_20734,N_20116,N_19801);
nand U20735 (N_20735,N_19858,N_20229);
nor U20736 (N_20736,N_20009,N_20057);
xor U20737 (N_20737,N_19938,N_20250);
and U20738 (N_20738,N_20113,N_19924);
or U20739 (N_20739,N_19844,N_20076);
nor U20740 (N_20740,N_20386,N_20094);
nand U20741 (N_20741,N_19826,N_20181);
nor U20742 (N_20742,N_20103,N_19946);
nor U20743 (N_20743,N_20169,N_19826);
or U20744 (N_20744,N_19901,N_20055);
and U20745 (N_20745,N_20377,N_19954);
or U20746 (N_20746,N_20206,N_19849);
or U20747 (N_20747,N_20107,N_20325);
and U20748 (N_20748,N_20052,N_19954);
or U20749 (N_20749,N_20318,N_20141);
xor U20750 (N_20750,N_20184,N_20389);
nor U20751 (N_20751,N_20000,N_20353);
nor U20752 (N_20752,N_20083,N_20357);
or U20753 (N_20753,N_20107,N_20062);
and U20754 (N_20754,N_19827,N_19816);
nand U20755 (N_20755,N_19887,N_20015);
or U20756 (N_20756,N_20396,N_19851);
nand U20757 (N_20757,N_20006,N_20073);
xor U20758 (N_20758,N_20356,N_20271);
and U20759 (N_20759,N_20066,N_20263);
nor U20760 (N_20760,N_20031,N_19987);
nand U20761 (N_20761,N_20140,N_19863);
nor U20762 (N_20762,N_19956,N_20260);
or U20763 (N_20763,N_20068,N_20202);
or U20764 (N_20764,N_20340,N_19969);
or U20765 (N_20765,N_19916,N_19875);
xor U20766 (N_20766,N_20055,N_19917);
xnor U20767 (N_20767,N_19855,N_20171);
or U20768 (N_20768,N_19934,N_20131);
or U20769 (N_20769,N_20389,N_19860);
and U20770 (N_20770,N_20302,N_19949);
or U20771 (N_20771,N_20101,N_20026);
and U20772 (N_20772,N_20266,N_20106);
and U20773 (N_20773,N_19940,N_20273);
xor U20774 (N_20774,N_19853,N_20266);
or U20775 (N_20775,N_20281,N_20256);
and U20776 (N_20776,N_20279,N_20051);
and U20777 (N_20777,N_19871,N_20098);
nand U20778 (N_20778,N_20323,N_20117);
xnor U20779 (N_20779,N_20231,N_19989);
and U20780 (N_20780,N_20196,N_20298);
nor U20781 (N_20781,N_19866,N_19817);
nor U20782 (N_20782,N_20370,N_20345);
nor U20783 (N_20783,N_20207,N_20223);
or U20784 (N_20784,N_20224,N_20074);
xor U20785 (N_20785,N_20352,N_20298);
and U20786 (N_20786,N_19837,N_20071);
nor U20787 (N_20787,N_20024,N_20094);
or U20788 (N_20788,N_20003,N_19995);
or U20789 (N_20789,N_20274,N_20264);
nand U20790 (N_20790,N_20257,N_19993);
and U20791 (N_20791,N_20217,N_20347);
or U20792 (N_20792,N_20357,N_20079);
or U20793 (N_20793,N_19936,N_20315);
nor U20794 (N_20794,N_20240,N_20101);
nand U20795 (N_20795,N_20317,N_20387);
nand U20796 (N_20796,N_20034,N_20101);
xnor U20797 (N_20797,N_19948,N_19952);
nor U20798 (N_20798,N_20353,N_20206);
nand U20799 (N_20799,N_19821,N_20305);
nor U20800 (N_20800,N_19956,N_20376);
or U20801 (N_20801,N_19931,N_20335);
nor U20802 (N_20802,N_20059,N_20116);
or U20803 (N_20803,N_19985,N_20249);
nor U20804 (N_20804,N_19871,N_20396);
and U20805 (N_20805,N_20000,N_20112);
xnor U20806 (N_20806,N_20326,N_19823);
and U20807 (N_20807,N_19935,N_19823);
nand U20808 (N_20808,N_19811,N_20192);
nand U20809 (N_20809,N_20375,N_20039);
and U20810 (N_20810,N_20063,N_19846);
xor U20811 (N_20811,N_20042,N_19907);
xor U20812 (N_20812,N_20342,N_19851);
and U20813 (N_20813,N_19859,N_19870);
and U20814 (N_20814,N_20066,N_20173);
or U20815 (N_20815,N_20354,N_19942);
or U20816 (N_20816,N_20027,N_19938);
xor U20817 (N_20817,N_19944,N_20066);
or U20818 (N_20818,N_19855,N_20365);
nor U20819 (N_20819,N_20130,N_19983);
or U20820 (N_20820,N_20068,N_20113);
and U20821 (N_20821,N_20231,N_20143);
xnor U20822 (N_20822,N_20278,N_20200);
xor U20823 (N_20823,N_20125,N_19877);
nor U20824 (N_20824,N_19959,N_20225);
nand U20825 (N_20825,N_20193,N_20084);
or U20826 (N_20826,N_20128,N_20316);
nor U20827 (N_20827,N_20122,N_19803);
nand U20828 (N_20828,N_19826,N_20324);
and U20829 (N_20829,N_20078,N_19918);
nand U20830 (N_20830,N_20351,N_20016);
xor U20831 (N_20831,N_20100,N_20315);
and U20832 (N_20832,N_20184,N_20355);
nand U20833 (N_20833,N_20029,N_20261);
or U20834 (N_20834,N_20226,N_20219);
nor U20835 (N_20835,N_20215,N_20176);
nor U20836 (N_20836,N_20276,N_19985);
or U20837 (N_20837,N_19848,N_20070);
nor U20838 (N_20838,N_20358,N_20314);
xor U20839 (N_20839,N_20037,N_20205);
nand U20840 (N_20840,N_19992,N_19803);
or U20841 (N_20841,N_20070,N_20384);
nor U20842 (N_20842,N_20012,N_20099);
and U20843 (N_20843,N_19985,N_19854);
or U20844 (N_20844,N_20163,N_20271);
nand U20845 (N_20845,N_20327,N_19841);
and U20846 (N_20846,N_20202,N_19925);
and U20847 (N_20847,N_19812,N_19893);
xor U20848 (N_20848,N_19866,N_19999);
xor U20849 (N_20849,N_20397,N_20263);
nand U20850 (N_20850,N_19931,N_20249);
and U20851 (N_20851,N_19858,N_19913);
and U20852 (N_20852,N_20281,N_20380);
nand U20853 (N_20853,N_20148,N_20203);
nor U20854 (N_20854,N_20116,N_19874);
nand U20855 (N_20855,N_20386,N_19877);
or U20856 (N_20856,N_20158,N_19999);
xor U20857 (N_20857,N_20388,N_20018);
nand U20858 (N_20858,N_20130,N_20055);
xnor U20859 (N_20859,N_20208,N_20138);
xnor U20860 (N_20860,N_20146,N_19972);
nor U20861 (N_20861,N_19862,N_20137);
or U20862 (N_20862,N_20368,N_20271);
nor U20863 (N_20863,N_19989,N_19853);
xnor U20864 (N_20864,N_20353,N_19825);
and U20865 (N_20865,N_20363,N_20061);
nand U20866 (N_20866,N_20231,N_19965);
nor U20867 (N_20867,N_20098,N_19896);
nor U20868 (N_20868,N_20049,N_20259);
or U20869 (N_20869,N_20239,N_20142);
nand U20870 (N_20870,N_20321,N_20259);
nor U20871 (N_20871,N_20049,N_20171);
nor U20872 (N_20872,N_19843,N_20235);
nand U20873 (N_20873,N_19822,N_20306);
or U20874 (N_20874,N_20092,N_20073);
nand U20875 (N_20875,N_20061,N_20230);
and U20876 (N_20876,N_19874,N_20238);
and U20877 (N_20877,N_20234,N_19985);
nor U20878 (N_20878,N_19883,N_20115);
nor U20879 (N_20879,N_19855,N_19935);
or U20880 (N_20880,N_20175,N_19852);
xor U20881 (N_20881,N_20333,N_20066);
xor U20882 (N_20882,N_19843,N_19861);
nand U20883 (N_20883,N_20337,N_19907);
nand U20884 (N_20884,N_20199,N_19881);
nor U20885 (N_20885,N_20198,N_20223);
and U20886 (N_20886,N_20139,N_19932);
and U20887 (N_20887,N_20205,N_20011);
nor U20888 (N_20888,N_20176,N_19976);
and U20889 (N_20889,N_20183,N_20135);
nor U20890 (N_20890,N_20245,N_20232);
nor U20891 (N_20891,N_20223,N_19837);
and U20892 (N_20892,N_20256,N_20003);
and U20893 (N_20893,N_20236,N_20248);
and U20894 (N_20894,N_20084,N_19869);
and U20895 (N_20895,N_20076,N_20207);
xnor U20896 (N_20896,N_20023,N_19865);
and U20897 (N_20897,N_19880,N_20157);
xor U20898 (N_20898,N_20001,N_20010);
xnor U20899 (N_20899,N_19813,N_19931);
nand U20900 (N_20900,N_20376,N_20165);
xor U20901 (N_20901,N_20002,N_19894);
or U20902 (N_20902,N_20101,N_19808);
or U20903 (N_20903,N_20070,N_20073);
or U20904 (N_20904,N_20357,N_20067);
and U20905 (N_20905,N_20205,N_20094);
nand U20906 (N_20906,N_19985,N_19951);
or U20907 (N_20907,N_20160,N_20030);
nand U20908 (N_20908,N_20245,N_19809);
xor U20909 (N_20909,N_19852,N_20036);
or U20910 (N_20910,N_20274,N_20090);
xnor U20911 (N_20911,N_20053,N_20340);
nand U20912 (N_20912,N_19898,N_20348);
or U20913 (N_20913,N_20185,N_19979);
nand U20914 (N_20914,N_20018,N_20029);
nor U20915 (N_20915,N_20250,N_20377);
and U20916 (N_20916,N_20130,N_20324);
nor U20917 (N_20917,N_20148,N_20118);
and U20918 (N_20918,N_19909,N_20320);
and U20919 (N_20919,N_19959,N_19863);
or U20920 (N_20920,N_20213,N_20316);
and U20921 (N_20921,N_20014,N_20173);
nor U20922 (N_20922,N_20270,N_19937);
nor U20923 (N_20923,N_20190,N_19937);
nand U20924 (N_20924,N_20051,N_20114);
xor U20925 (N_20925,N_20104,N_20383);
xor U20926 (N_20926,N_20376,N_19921);
or U20927 (N_20927,N_20396,N_20355);
nand U20928 (N_20928,N_19878,N_20005);
and U20929 (N_20929,N_19804,N_19974);
or U20930 (N_20930,N_20327,N_20345);
xnor U20931 (N_20931,N_20069,N_20346);
nand U20932 (N_20932,N_20272,N_19857);
nand U20933 (N_20933,N_20188,N_20011);
and U20934 (N_20934,N_19992,N_20168);
and U20935 (N_20935,N_20227,N_19855);
and U20936 (N_20936,N_20318,N_20194);
or U20937 (N_20937,N_20194,N_20263);
xor U20938 (N_20938,N_20186,N_20144);
and U20939 (N_20939,N_20233,N_20114);
and U20940 (N_20940,N_19943,N_20002);
or U20941 (N_20941,N_19975,N_20248);
nand U20942 (N_20942,N_19971,N_19863);
nand U20943 (N_20943,N_19850,N_20257);
or U20944 (N_20944,N_19998,N_20387);
nor U20945 (N_20945,N_20253,N_20194);
and U20946 (N_20946,N_19848,N_20243);
xor U20947 (N_20947,N_20185,N_20246);
or U20948 (N_20948,N_19997,N_20023);
xor U20949 (N_20949,N_20102,N_20136);
nand U20950 (N_20950,N_19966,N_20313);
nor U20951 (N_20951,N_20301,N_20332);
nor U20952 (N_20952,N_20185,N_20142);
nand U20953 (N_20953,N_20396,N_20177);
and U20954 (N_20954,N_20080,N_20156);
nor U20955 (N_20955,N_20071,N_20074);
nor U20956 (N_20956,N_20389,N_20022);
xnor U20957 (N_20957,N_19978,N_20082);
nor U20958 (N_20958,N_19825,N_20024);
nor U20959 (N_20959,N_19824,N_19934);
and U20960 (N_20960,N_19923,N_19857);
or U20961 (N_20961,N_20371,N_19970);
nand U20962 (N_20962,N_20322,N_19989);
and U20963 (N_20963,N_19834,N_20051);
and U20964 (N_20964,N_20010,N_20308);
nand U20965 (N_20965,N_20020,N_20389);
xnor U20966 (N_20966,N_19990,N_20257);
xor U20967 (N_20967,N_20057,N_20296);
and U20968 (N_20968,N_20036,N_19877);
or U20969 (N_20969,N_20107,N_20370);
and U20970 (N_20970,N_19840,N_20049);
nand U20971 (N_20971,N_20369,N_19983);
or U20972 (N_20972,N_20353,N_20054);
xnor U20973 (N_20973,N_19832,N_19947);
nand U20974 (N_20974,N_20243,N_20295);
xor U20975 (N_20975,N_19986,N_19909);
or U20976 (N_20976,N_20323,N_20218);
and U20977 (N_20977,N_19980,N_20372);
nand U20978 (N_20978,N_20062,N_20079);
xnor U20979 (N_20979,N_19927,N_19944);
xor U20980 (N_20980,N_20004,N_20328);
nand U20981 (N_20981,N_20018,N_19832);
nand U20982 (N_20982,N_20151,N_20281);
or U20983 (N_20983,N_20255,N_20057);
xor U20984 (N_20984,N_19894,N_20219);
or U20985 (N_20985,N_20306,N_20273);
nand U20986 (N_20986,N_20126,N_20287);
and U20987 (N_20987,N_20142,N_20399);
xnor U20988 (N_20988,N_19845,N_20006);
xnor U20989 (N_20989,N_20284,N_20011);
nor U20990 (N_20990,N_20223,N_20361);
nor U20991 (N_20991,N_20096,N_20080);
nor U20992 (N_20992,N_20378,N_20369);
nor U20993 (N_20993,N_20350,N_20371);
nor U20994 (N_20994,N_19865,N_20034);
or U20995 (N_20995,N_19859,N_19860);
xnor U20996 (N_20996,N_20207,N_19939);
or U20997 (N_20997,N_19947,N_20213);
nand U20998 (N_20998,N_20152,N_20346);
xor U20999 (N_20999,N_20290,N_20034);
nand U21000 (N_21000,N_20881,N_20600);
xor U21001 (N_21001,N_20448,N_20551);
and U21002 (N_21002,N_20896,N_20601);
nand U21003 (N_21003,N_20620,N_20756);
nand U21004 (N_21004,N_20466,N_20948);
or U21005 (N_21005,N_20415,N_20829);
or U21006 (N_21006,N_20979,N_20673);
nand U21007 (N_21007,N_20417,N_20694);
or U21008 (N_21008,N_20730,N_20405);
nor U21009 (N_21009,N_20739,N_20581);
and U21010 (N_21010,N_20828,N_20890);
nor U21011 (N_21011,N_20752,N_20850);
or U21012 (N_21012,N_20597,N_20479);
nand U21013 (N_21013,N_20903,N_20440);
xnor U21014 (N_21014,N_20592,N_20664);
and U21015 (N_21015,N_20871,N_20719);
or U21016 (N_21016,N_20461,N_20826);
nand U21017 (N_21017,N_20438,N_20681);
xor U21018 (N_21018,N_20671,N_20864);
nor U21019 (N_21019,N_20961,N_20988);
and U21020 (N_21020,N_20729,N_20552);
and U21021 (N_21021,N_20598,N_20678);
nand U21022 (N_21022,N_20542,N_20740);
and U21023 (N_21023,N_20793,N_20437);
xor U21024 (N_21024,N_20691,N_20843);
nor U21025 (N_21025,N_20804,N_20530);
xor U21026 (N_21026,N_20401,N_20974);
nor U21027 (N_21027,N_20540,N_20796);
or U21028 (N_21028,N_20699,N_20657);
nand U21029 (N_21029,N_20820,N_20870);
nand U21030 (N_21030,N_20546,N_20883);
and U21031 (N_21031,N_20888,N_20509);
or U21032 (N_21032,N_20989,N_20602);
xnor U21033 (N_21033,N_20934,N_20900);
nand U21034 (N_21034,N_20488,N_20875);
nor U21035 (N_21035,N_20460,N_20867);
nor U21036 (N_21036,N_20750,N_20483);
xor U21037 (N_21037,N_20901,N_20513);
and U21038 (N_21038,N_20630,N_20497);
or U21039 (N_21039,N_20762,N_20846);
nand U21040 (N_21040,N_20947,N_20824);
nand U21041 (N_21041,N_20527,N_20478);
or U21042 (N_21042,N_20915,N_20548);
xnor U21043 (N_21043,N_20679,N_20427);
and U21044 (N_21044,N_20410,N_20463);
and U21045 (N_21045,N_20932,N_20953);
nand U21046 (N_21046,N_20914,N_20480);
and U21047 (N_21047,N_20819,N_20442);
and U21048 (N_21048,N_20732,N_20672);
xor U21049 (N_21049,N_20590,N_20572);
nand U21050 (N_21050,N_20839,N_20666);
xor U21051 (N_21051,N_20521,N_20408);
xnor U21052 (N_21052,N_20971,N_20923);
or U21053 (N_21053,N_20507,N_20951);
and U21054 (N_21054,N_20702,N_20443);
nor U21055 (N_21055,N_20473,N_20860);
xor U21056 (N_21056,N_20959,N_20726);
or U21057 (N_21057,N_20921,N_20558);
and U21058 (N_21058,N_20591,N_20917);
nor U21059 (N_21059,N_20449,N_20859);
xor U21060 (N_21060,N_20698,N_20703);
or U21061 (N_21061,N_20919,N_20662);
and U21062 (N_21062,N_20557,N_20777);
and U21063 (N_21063,N_20676,N_20628);
or U21064 (N_21064,N_20603,N_20884);
xor U21065 (N_21065,N_20485,N_20701);
and U21066 (N_21066,N_20763,N_20553);
nor U21067 (N_21067,N_20781,N_20992);
nor U21068 (N_21068,N_20727,N_20541);
and U21069 (N_21069,N_20863,N_20754);
nor U21070 (N_21070,N_20432,N_20906);
or U21071 (N_21071,N_20852,N_20403);
nor U21072 (N_21072,N_20573,N_20728);
nand U21073 (N_21073,N_20798,N_20660);
nand U21074 (N_21074,N_20447,N_20543);
nor U21075 (N_21075,N_20584,N_20516);
nor U21076 (N_21076,N_20629,N_20813);
xor U21077 (N_21077,N_20986,N_20795);
nor U21078 (N_21078,N_20452,N_20471);
xor U21079 (N_21079,N_20769,N_20925);
nand U21080 (N_21080,N_20981,N_20505);
and U21081 (N_21081,N_20670,N_20773);
nand U21082 (N_21082,N_20619,N_20710);
nor U21083 (N_21083,N_20656,N_20807);
nor U21084 (N_21084,N_20642,N_20969);
nand U21085 (N_21085,N_20586,N_20840);
xnor U21086 (N_21086,N_20433,N_20425);
nor U21087 (N_21087,N_20588,N_20713);
and U21088 (N_21088,N_20685,N_20684);
xnor U21089 (N_21089,N_20537,N_20496);
xor U21090 (N_21090,N_20518,N_20686);
and U21091 (N_21091,N_20643,N_20411);
nand U21092 (N_21092,N_20880,N_20693);
xnor U21093 (N_21093,N_20476,N_20625);
or U21094 (N_21094,N_20930,N_20894);
nor U21095 (N_21095,N_20770,N_20823);
nand U21096 (N_21096,N_20578,N_20910);
and U21097 (N_21097,N_20922,N_20785);
xor U21098 (N_21098,N_20963,N_20465);
and U21099 (N_21099,N_20429,N_20851);
and U21100 (N_21100,N_20760,N_20717);
and U21101 (N_21101,N_20580,N_20982);
nor U21102 (N_21102,N_20531,N_20583);
nor U21103 (N_21103,N_20579,N_20831);
or U21104 (N_21104,N_20755,N_20658);
and U21105 (N_21105,N_20749,N_20997);
xnor U21106 (N_21106,N_20641,N_20617);
nor U21107 (N_21107,N_20806,N_20886);
or U21108 (N_21108,N_20690,N_20577);
nor U21109 (N_21109,N_20512,N_20544);
and U21110 (N_21110,N_20757,N_20802);
and U21111 (N_21111,N_20902,N_20955);
and U21112 (N_21112,N_20675,N_20822);
and U21113 (N_21113,N_20566,N_20495);
xor U21114 (N_21114,N_20524,N_20841);
nor U21115 (N_21115,N_20808,N_20593);
and U21116 (N_21116,N_20559,N_20941);
xor U21117 (N_21117,N_20523,N_20748);
xnor U21118 (N_21118,N_20651,N_20899);
nor U21119 (N_21119,N_20778,N_20874);
or U21120 (N_21120,N_20869,N_20956);
and U21121 (N_21121,N_20499,N_20797);
nand U21122 (N_21122,N_20789,N_20774);
xnor U21123 (N_21123,N_20611,N_20689);
nand U21124 (N_21124,N_20715,N_20990);
nor U21125 (N_21125,N_20721,N_20776);
and U21126 (N_21126,N_20878,N_20547);
and U21127 (N_21127,N_20599,N_20978);
xnor U21128 (N_21128,N_20810,N_20426);
nand U21129 (N_21129,N_20996,N_20674);
xnor U21130 (N_21130,N_20420,N_20842);
xnor U21131 (N_21131,N_20817,N_20450);
and U21132 (N_21132,N_20709,N_20957);
nor U21133 (N_21133,N_20825,N_20536);
xnor U21134 (N_21134,N_20920,N_20723);
nor U21135 (N_21135,N_20659,N_20434);
nand U21136 (N_21136,N_20938,N_20545);
nand U21137 (N_21137,N_20980,N_20646);
or U21138 (N_21138,N_20610,N_20409);
nor U21139 (N_21139,N_20983,N_20960);
nor U21140 (N_21140,N_20893,N_20467);
and U21141 (N_21141,N_20942,N_20435);
or U21142 (N_21142,N_20885,N_20812);
and U21143 (N_21143,N_20879,N_20428);
or U21144 (N_21144,N_20567,N_20718);
nand U21145 (N_21145,N_20794,N_20412);
xnor U21146 (N_21146,N_20407,N_20413);
and U21147 (N_21147,N_20764,N_20731);
xnor U21148 (N_21148,N_20845,N_20491);
nand U21149 (N_21149,N_20680,N_20775);
or U21150 (N_21150,N_20454,N_20984);
nor U21151 (N_21151,N_20766,N_20414);
nand U21152 (N_21152,N_20596,N_20761);
and U21153 (N_21153,N_20758,N_20652);
and U21154 (N_21154,N_20561,N_20973);
xor U21155 (N_21155,N_20844,N_20457);
xnor U21156 (N_21156,N_20668,N_20872);
nand U21157 (N_21157,N_20609,N_20622);
nor U21158 (N_21158,N_20882,N_20654);
nor U21159 (N_21159,N_20649,N_20555);
and U21160 (N_21160,N_20575,N_20783);
or U21161 (N_21161,N_20737,N_20400);
and U21162 (N_21162,N_20482,N_20431);
or U21163 (N_21163,N_20972,N_20605);
xnor U21164 (N_21164,N_20866,N_20614);
nor U21165 (N_21165,N_20967,N_20995);
nor U21166 (N_21166,N_20621,N_20464);
nand U21167 (N_21167,N_20430,N_20977);
nand U21168 (N_21168,N_20404,N_20522);
xor U21169 (N_21169,N_20929,N_20663);
xor U21170 (N_21170,N_20565,N_20626);
or U21171 (N_21171,N_20976,N_20631);
and U21172 (N_21172,N_20645,N_20539);
nor U21173 (N_21173,N_20486,N_20568);
xnor U21174 (N_21174,N_20792,N_20422);
nand U21175 (N_21175,N_20608,N_20991);
xor U21176 (N_21176,N_20607,N_20444);
or U21177 (N_21177,N_20868,N_20650);
nor U21178 (N_21178,N_20563,N_20459);
nor U21179 (N_21179,N_20742,N_20623);
and U21180 (N_21180,N_20470,N_20453);
and U21181 (N_21181,N_20943,N_20854);
nand U21182 (N_21182,N_20419,N_20576);
nand U21183 (N_21183,N_20833,N_20569);
nand U21184 (N_21184,N_20830,N_20954);
nand U21185 (N_21185,N_20744,N_20927);
or U21186 (N_21186,N_20618,N_20724);
and U21187 (N_21187,N_20911,N_20816);
nand U21188 (N_21188,N_20765,N_20469);
or U21189 (N_21189,N_20554,N_20891);
nor U21190 (N_21190,N_20661,N_20818);
xor U21191 (N_21191,N_20436,N_20582);
nor U21192 (N_21192,N_20604,N_20743);
nor U21193 (N_21193,N_20725,N_20423);
nand U21194 (N_21194,N_20987,N_20683);
nor U21195 (N_21195,N_20994,N_20418);
or U21196 (N_21196,N_20616,N_20735);
nor U21197 (N_21197,N_20708,N_20697);
nor U21198 (N_21198,N_20815,N_20722);
xor U21199 (N_21199,N_20615,N_20809);
or U21200 (N_21200,N_20918,N_20688);
or U21201 (N_21201,N_20790,N_20907);
xor U21202 (N_21202,N_20788,N_20692);
xor U21203 (N_21203,N_20862,N_20517);
nand U21204 (N_21204,N_20855,N_20791);
nand U21205 (N_21205,N_20514,N_20747);
and U21206 (N_21206,N_20638,N_20940);
and U21207 (N_21207,N_20639,N_20502);
xnor U21208 (N_21208,N_20771,N_20574);
nor U21209 (N_21209,N_20857,N_20711);
xor U21210 (N_21210,N_20472,N_20865);
xor U21211 (N_21211,N_20632,N_20767);
or U21212 (N_21212,N_20640,N_20475);
xnor U21213 (N_21213,N_20526,N_20926);
and U21214 (N_21214,N_20520,N_20564);
and U21215 (N_21215,N_20873,N_20944);
nor U21216 (N_21216,N_20474,N_20624);
and U21217 (N_21217,N_20462,N_20484);
or U21218 (N_21218,N_20669,N_20935);
xnor U21219 (N_21219,N_20647,N_20998);
or U21220 (N_21220,N_20655,N_20634);
xnor U21221 (N_21221,N_20494,N_20458);
xnor U21222 (N_21222,N_20751,N_20898);
xor U21223 (N_21223,N_20627,N_20912);
nand U21224 (N_21224,N_20421,N_20424);
nand U21225 (N_21225,N_20966,N_20635);
or U21226 (N_21226,N_20784,N_20667);
and U21227 (N_21227,N_20636,N_20847);
nor U21228 (N_21228,N_20928,N_20946);
nor U21229 (N_21229,N_20952,N_20993);
nor U21230 (N_21230,N_20876,N_20515);
xor U21231 (N_21231,N_20968,N_20779);
or U21232 (N_21232,N_20999,N_20538);
or U21233 (N_21233,N_20637,N_20533);
nand U21234 (N_21234,N_20803,N_20493);
and U21235 (N_21235,N_20549,N_20799);
nor U21236 (N_21236,N_20939,N_20805);
or U21237 (N_21237,N_20529,N_20481);
xor U21238 (N_21238,N_20498,N_20700);
or U21239 (N_21239,N_20931,N_20849);
xnor U21240 (N_21240,N_20402,N_20487);
nand U21241 (N_21241,N_20933,N_20519);
nand U21242 (N_21242,N_20741,N_20707);
or U21243 (N_21243,N_20595,N_20949);
nand U21244 (N_21244,N_20821,N_20511);
xor U21245 (N_21245,N_20492,N_20965);
nand U21246 (N_21246,N_20772,N_20644);
and U21247 (N_21247,N_20706,N_20687);
and U21248 (N_21248,N_20704,N_20682);
or U21249 (N_21249,N_20585,N_20633);
xnor U21250 (N_21250,N_20916,N_20525);
and U21251 (N_21251,N_20550,N_20653);
nand U21252 (N_21252,N_20837,N_20738);
nand U21253 (N_21253,N_20858,N_20853);
nor U21254 (N_21254,N_20446,N_20562);
nor U21255 (N_21255,N_20897,N_20500);
nor U21256 (N_21256,N_20856,N_20489);
nor U21257 (N_21257,N_20908,N_20455);
xnor U21258 (N_21258,N_20800,N_20836);
xor U21259 (N_21259,N_20456,N_20560);
nand U21260 (N_21260,N_20612,N_20451);
and U21261 (N_21261,N_20753,N_20503);
xnor U21262 (N_21262,N_20665,N_20508);
xnor U21263 (N_21263,N_20532,N_20913);
nor U21264 (N_21264,N_20501,N_20759);
nor U21265 (N_21265,N_20936,N_20909);
xnor U21266 (N_21266,N_20889,N_20746);
and U21267 (N_21267,N_20892,N_20648);
or U21268 (N_21268,N_20445,N_20677);
xnor U21269 (N_21269,N_20768,N_20504);
nor U21270 (N_21270,N_20835,N_20848);
nand U21271 (N_21271,N_20887,N_20827);
xor U21272 (N_21272,N_20801,N_20716);
nand U21273 (N_21273,N_20606,N_20734);
and U21274 (N_21274,N_20714,N_20811);
nand U21275 (N_21275,N_20964,N_20613);
or U21276 (N_21276,N_20787,N_20705);
nor U21277 (N_21277,N_20556,N_20468);
xnor U21278 (N_21278,N_20962,N_20937);
nor U21279 (N_21279,N_20570,N_20782);
nor U21280 (N_21280,N_20895,N_20904);
or U21281 (N_21281,N_20861,N_20510);
xnor U21282 (N_21282,N_20490,N_20733);
and U21283 (N_21283,N_20535,N_20736);
nor U21284 (N_21284,N_20985,N_20506);
or U21285 (N_21285,N_20712,N_20945);
and U21286 (N_21286,N_20477,N_20814);
and U21287 (N_21287,N_20589,N_20528);
nor U21288 (N_21288,N_20534,N_20877);
nand U21289 (N_21289,N_20832,N_20441);
and U21290 (N_21290,N_20834,N_20439);
nand U21291 (N_21291,N_20780,N_20587);
nor U21292 (N_21292,N_20745,N_20786);
xnor U21293 (N_21293,N_20970,N_20696);
nand U21294 (N_21294,N_20416,N_20720);
nor U21295 (N_21295,N_20975,N_20571);
nor U21296 (N_21296,N_20905,N_20838);
xnor U21297 (N_21297,N_20958,N_20406);
nor U21298 (N_21298,N_20950,N_20594);
xor U21299 (N_21299,N_20695,N_20924);
nor U21300 (N_21300,N_20659,N_20881);
or U21301 (N_21301,N_20928,N_20414);
and U21302 (N_21302,N_20871,N_20945);
xor U21303 (N_21303,N_20504,N_20748);
nor U21304 (N_21304,N_20571,N_20944);
nand U21305 (N_21305,N_20880,N_20456);
nand U21306 (N_21306,N_20903,N_20736);
nor U21307 (N_21307,N_20788,N_20615);
or U21308 (N_21308,N_20443,N_20791);
xnor U21309 (N_21309,N_20708,N_20422);
and U21310 (N_21310,N_20436,N_20536);
and U21311 (N_21311,N_20695,N_20709);
and U21312 (N_21312,N_20806,N_20808);
or U21313 (N_21313,N_20729,N_20741);
and U21314 (N_21314,N_20966,N_20871);
xor U21315 (N_21315,N_20829,N_20560);
nor U21316 (N_21316,N_20936,N_20902);
and U21317 (N_21317,N_20630,N_20590);
nor U21318 (N_21318,N_20518,N_20875);
xor U21319 (N_21319,N_20426,N_20747);
nor U21320 (N_21320,N_20522,N_20582);
nand U21321 (N_21321,N_20996,N_20784);
and U21322 (N_21322,N_20710,N_20773);
and U21323 (N_21323,N_20543,N_20979);
xnor U21324 (N_21324,N_20567,N_20515);
nor U21325 (N_21325,N_20473,N_20667);
xor U21326 (N_21326,N_20438,N_20554);
and U21327 (N_21327,N_20852,N_20976);
and U21328 (N_21328,N_20864,N_20570);
and U21329 (N_21329,N_20561,N_20958);
xor U21330 (N_21330,N_20569,N_20757);
nand U21331 (N_21331,N_20993,N_20708);
or U21332 (N_21332,N_20744,N_20563);
nand U21333 (N_21333,N_20579,N_20644);
or U21334 (N_21334,N_20813,N_20896);
nand U21335 (N_21335,N_20696,N_20853);
nor U21336 (N_21336,N_20528,N_20567);
nor U21337 (N_21337,N_20774,N_20937);
or U21338 (N_21338,N_20572,N_20475);
or U21339 (N_21339,N_20844,N_20640);
or U21340 (N_21340,N_20955,N_20784);
nand U21341 (N_21341,N_20507,N_20497);
or U21342 (N_21342,N_20976,N_20965);
or U21343 (N_21343,N_20940,N_20701);
nand U21344 (N_21344,N_20944,N_20559);
xor U21345 (N_21345,N_20811,N_20976);
xnor U21346 (N_21346,N_20830,N_20587);
xor U21347 (N_21347,N_20402,N_20597);
and U21348 (N_21348,N_20625,N_20582);
nand U21349 (N_21349,N_20518,N_20747);
nor U21350 (N_21350,N_20572,N_20629);
xnor U21351 (N_21351,N_20632,N_20576);
nand U21352 (N_21352,N_20702,N_20761);
xnor U21353 (N_21353,N_20522,N_20446);
nand U21354 (N_21354,N_20951,N_20974);
xor U21355 (N_21355,N_20938,N_20590);
nor U21356 (N_21356,N_20647,N_20831);
xnor U21357 (N_21357,N_20596,N_20559);
or U21358 (N_21358,N_20445,N_20497);
and U21359 (N_21359,N_20899,N_20823);
or U21360 (N_21360,N_20788,N_20965);
nand U21361 (N_21361,N_20786,N_20467);
and U21362 (N_21362,N_20493,N_20589);
or U21363 (N_21363,N_20945,N_20874);
and U21364 (N_21364,N_20534,N_20422);
xnor U21365 (N_21365,N_20412,N_20952);
nand U21366 (N_21366,N_20806,N_20483);
or U21367 (N_21367,N_20435,N_20951);
and U21368 (N_21368,N_20586,N_20972);
and U21369 (N_21369,N_20826,N_20671);
and U21370 (N_21370,N_20805,N_20591);
and U21371 (N_21371,N_20744,N_20968);
and U21372 (N_21372,N_20784,N_20499);
nand U21373 (N_21373,N_20789,N_20967);
nand U21374 (N_21374,N_20540,N_20829);
nor U21375 (N_21375,N_20739,N_20573);
and U21376 (N_21376,N_20736,N_20859);
xor U21377 (N_21377,N_20477,N_20766);
or U21378 (N_21378,N_20457,N_20557);
xnor U21379 (N_21379,N_20471,N_20411);
and U21380 (N_21380,N_20496,N_20452);
nand U21381 (N_21381,N_20918,N_20691);
nor U21382 (N_21382,N_20935,N_20817);
xor U21383 (N_21383,N_20740,N_20939);
xnor U21384 (N_21384,N_20844,N_20636);
and U21385 (N_21385,N_20596,N_20483);
or U21386 (N_21386,N_20452,N_20830);
xnor U21387 (N_21387,N_20451,N_20960);
or U21388 (N_21388,N_20772,N_20521);
or U21389 (N_21389,N_20578,N_20752);
xor U21390 (N_21390,N_20628,N_20511);
and U21391 (N_21391,N_20788,N_20709);
nand U21392 (N_21392,N_20947,N_20572);
xnor U21393 (N_21393,N_20766,N_20679);
or U21394 (N_21394,N_20607,N_20758);
xor U21395 (N_21395,N_20886,N_20998);
xor U21396 (N_21396,N_20685,N_20623);
xnor U21397 (N_21397,N_20449,N_20786);
nor U21398 (N_21398,N_20908,N_20445);
nor U21399 (N_21399,N_20585,N_20563);
xor U21400 (N_21400,N_20608,N_20639);
nor U21401 (N_21401,N_20881,N_20645);
or U21402 (N_21402,N_20834,N_20626);
and U21403 (N_21403,N_20922,N_20400);
nand U21404 (N_21404,N_20708,N_20714);
or U21405 (N_21405,N_20580,N_20520);
or U21406 (N_21406,N_20494,N_20789);
or U21407 (N_21407,N_20657,N_20761);
nor U21408 (N_21408,N_20417,N_20409);
nand U21409 (N_21409,N_20964,N_20445);
or U21410 (N_21410,N_20567,N_20455);
xor U21411 (N_21411,N_20916,N_20892);
nand U21412 (N_21412,N_20703,N_20631);
or U21413 (N_21413,N_20708,N_20628);
nor U21414 (N_21414,N_20934,N_20565);
xnor U21415 (N_21415,N_20474,N_20412);
or U21416 (N_21416,N_20528,N_20888);
or U21417 (N_21417,N_20942,N_20873);
xnor U21418 (N_21418,N_20894,N_20585);
and U21419 (N_21419,N_20420,N_20521);
xor U21420 (N_21420,N_20828,N_20425);
and U21421 (N_21421,N_20685,N_20726);
nand U21422 (N_21422,N_20536,N_20539);
nor U21423 (N_21423,N_20658,N_20465);
and U21424 (N_21424,N_20781,N_20818);
xor U21425 (N_21425,N_20974,N_20597);
or U21426 (N_21426,N_20958,N_20461);
nor U21427 (N_21427,N_20830,N_20709);
and U21428 (N_21428,N_20822,N_20700);
nand U21429 (N_21429,N_20930,N_20799);
or U21430 (N_21430,N_20875,N_20761);
xor U21431 (N_21431,N_20413,N_20998);
xnor U21432 (N_21432,N_20547,N_20735);
nand U21433 (N_21433,N_20790,N_20914);
and U21434 (N_21434,N_20660,N_20445);
nor U21435 (N_21435,N_20826,N_20433);
or U21436 (N_21436,N_20616,N_20529);
nor U21437 (N_21437,N_20970,N_20716);
nor U21438 (N_21438,N_20655,N_20725);
and U21439 (N_21439,N_20581,N_20745);
or U21440 (N_21440,N_20548,N_20623);
nor U21441 (N_21441,N_20696,N_20491);
nand U21442 (N_21442,N_20871,N_20838);
or U21443 (N_21443,N_20848,N_20957);
or U21444 (N_21444,N_20913,N_20423);
nor U21445 (N_21445,N_20958,N_20570);
xnor U21446 (N_21446,N_20562,N_20489);
and U21447 (N_21447,N_20987,N_20701);
nor U21448 (N_21448,N_20625,N_20596);
xnor U21449 (N_21449,N_20657,N_20760);
xor U21450 (N_21450,N_20820,N_20985);
xor U21451 (N_21451,N_20843,N_20722);
nor U21452 (N_21452,N_20671,N_20850);
xnor U21453 (N_21453,N_20855,N_20417);
and U21454 (N_21454,N_20541,N_20638);
or U21455 (N_21455,N_20835,N_20744);
or U21456 (N_21456,N_20468,N_20626);
and U21457 (N_21457,N_20863,N_20716);
or U21458 (N_21458,N_20625,N_20577);
nor U21459 (N_21459,N_20403,N_20722);
and U21460 (N_21460,N_20817,N_20631);
or U21461 (N_21461,N_20866,N_20509);
or U21462 (N_21462,N_20525,N_20590);
xor U21463 (N_21463,N_20486,N_20928);
or U21464 (N_21464,N_20431,N_20508);
nand U21465 (N_21465,N_20572,N_20428);
nand U21466 (N_21466,N_20894,N_20924);
nor U21467 (N_21467,N_20842,N_20702);
nor U21468 (N_21468,N_20433,N_20421);
nor U21469 (N_21469,N_20475,N_20889);
and U21470 (N_21470,N_20721,N_20554);
nand U21471 (N_21471,N_20638,N_20532);
and U21472 (N_21472,N_20712,N_20706);
and U21473 (N_21473,N_20458,N_20651);
or U21474 (N_21474,N_20645,N_20756);
or U21475 (N_21475,N_20521,N_20960);
nand U21476 (N_21476,N_20785,N_20864);
nor U21477 (N_21477,N_20755,N_20501);
nand U21478 (N_21478,N_20781,N_20712);
or U21479 (N_21479,N_20625,N_20517);
xnor U21480 (N_21480,N_20974,N_20530);
nand U21481 (N_21481,N_20438,N_20844);
xnor U21482 (N_21482,N_20873,N_20683);
nor U21483 (N_21483,N_20776,N_20902);
nand U21484 (N_21484,N_20693,N_20417);
nand U21485 (N_21485,N_20882,N_20935);
nand U21486 (N_21486,N_20835,N_20407);
and U21487 (N_21487,N_20914,N_20729);
or U21488 (N_21488,N_20502,N_20631);
nor U21489 (N_21489,N_20500,N_20994);
xor U21490 (N_21490,N_20880,N_20430);
or U21491 (N_21491,N_20576,N_20927);
xor U21492 (N_21492,N_20614,N_20864);
nor U21493 (N_21493,N_20552,N_20793);
xor U21494 (N_21494,N_20863,N_20703);
xnor U21495 (N_21495,N_20616,N_20959);
and U21496 (N_21496,N_20441,N_20678);
nor U21497 (N_21497,N_20754,N_20915);
and U21498 (N_21498,N_20733,N_20705);
xnor U21499 (N_21499,N_20466,N_20584);
nor U21500 (N_21500,N_20673,N_20647);
nor U21501 (N_21501,N_20485,N_20787);
or U21502 (N_21502,N_20686,N_20510);
and U21503 (N_21503,N_20433,N_20781);
nor U21504 (N_21504,N_20940,N_20599);
nand U21505 (N_21505,N_20921,N_20739);
and U21506 (N_21506,N_20836,N_20665);
nor U21507 (N_21507,N_20625,N_20924);
and U21508 (N_21508,N_20752,N_20520);
xnor U21509 (N_21509,N_20842,N_20874);
nand U21510 (N_21510,N_20517,N_20538);
nand U21511 (N_21511,N_20796,N_20892);
or U21512 (N_21512,N_20468,N_20661);
nand U21513 (N_21513,N_20661,N_20700);
nand U21514 (N_21514,N_20563,N_20710);
xor U21515 (N_21515,N_20768,N_20914);
xor U21516 (N_21516,N_20730,N_20728);
nor U21517 (N_21517,N_20965,N_20527);
or U21518 (N_21518,N_20722,N_20490);
nand U21519 (N_21519,N_20935,N_20649);
nand U21520 (N_21520,N_20519,N_20702);
or U21521 (N_21521,N_20866,N_20710);
nand U21522 (N_21522,N_20418,N_20885);
and U21523 (N_21523,N_20739,N_20811);
nor U21524 (N_21524,N_20748,N_20793);
and U21525 (N_21525,N_20941,N_20858);
nand U21526 (N_21526,N_20829,N_20642);
nand U21527 (N_21527,N_20965,N_20405);
xor U21528 (N_21528,N_20526,N_20758);
nor U21529 (N_21529,N_20504,N_20839);
nand U21530 (N_21530,N_20903,N_20428);
nand U21531 (N_21531,N_20701,N_20689);
nor U21532 (N_21532,N_20495,N_20616);
xor U21533 (N_21533,N_20761,N_20527);
nand U21534 (N_21534,N_20820,N_20774);
or U21535 (N_21535,N_20821,N_20515);
or U21536 (N_21536,N_20658,N_20588);
or U21537 (N_21537,N_20921,N_20542);
or U21538 (N_21538,N_20690,N_20836);
or U21539 (N_21539,N_20914,N_20423);
nor U21540 (N_21540,N_20781,N_20813);
nor U21541 (N_21541,N_20446,N_20555);
xor U21542 (N_21542,N_20439,N_20727);
nand U21543 (N_21543,N_20575,N_20999);
and U21544 (N_21544,N_20635,N_20947);
and U21545 (N_21545,N_20874,N_20825);
nor U21546 (N_21546,N_20696,N_20550);
xnor U21547 (N_21547,N_20735,N_20532);
xnor U21548 (N_21548,N_20742,N_20694);
nor U21549 (N_21549,N_20626,N_20999);
nor U21550 (N_21550,N_20778,N_20594);
nor U21551 (N_21551,N_20532,N_20930);
nand U21552 (N_21552,N_20512,N_20542);
or U21553 (N_21553,N_20421,N_20885);
and U21554 (N_21554,N_20835,N_20865);
xnor U21555 (N_21555,N_20740,N_20647);
and U21556 (N_21556,N_20842,N_20546);
xnor U21557 (N_21557,N_20433,N_20575);
or U21558 (N_21558,N_20771,N_20410);
nor U21559 (N_21559,N_20752,N_20538);
nor U21560 (N_21560,N_20744,N_20809);
and U21561 (N_21561,N_20707,N_20548);
nor U21562 (N_21562,N_20726,N_20732);
xnor U21563 (N_21563,N_20545,N_20694);
and U21564 (N_21564,N_20537,N_20913);
and U21565 (N_21565,N_20971,N_20617);
xor U21566 (N_21566,N_20699,N_20483);
or U21567 (N_21567,N_20958,N_20850);
and U21568 (N_21568,N_20530,N_20770);
nand U21569 (N_21569,N_20405,N_20430);
nand U21570 (N_21570,N_20898,N_20640);
nor U21571 (N_21571,N_20881,N_20787);
xor U21572 (N_21572,N_20977,N_20638);
or U21573 (N_21573,N_20997,N_20747);
xor U21574 (N_21574,N_20928,N_20995);
and U21575 (N_21575,N_20612,N_20678);
nor U21576 (N_21576,N_20572,N_20424);
nand U21577 (N_21577,N_20856,N_20497);
and U21578 (N_21578,N_20673,N_20799);
or U21579 (N_21579,N_20741,N_20932);
nand U21580 (N_21580,N_20859,N_20683);
nand U21581 (N_21581,N_20992,N_20796);
nor U21582 (N_21582,N_20678,N_20759);
or U21583 (N_21583,N_20491,N_20931);
nand U21584 (N_21584,N_20523,N_20643);
or U21585 (N_21585,N_20496,N_20728);
xor U21586 (N_21586,N_20693,N_20871);
and U21587 (N_21587,N_20436,N_20835);
nand U21588 (N_21588,N_20758,N_20746);
nor U21589 (N_21589,N_20687,N_20881);
nand U21590 (N_21590,N_20870,N_20950);
nand U21591 (N_21591,N_20808,N_20972);
or U21592 (N_21592,N_20626,N_20701);
xnor U21593 (N_21593,N_20760,N_20547);
and U21594 (N_21594,N_20660,N_20429);
xnor U21595 (N_21595,N_20810,N_20934);
nor U21596 (N_21596,N_20823,N_20776);
or U21597 (N_21597,N_20903,N_20480);
xor U21598 (N_21598,N_20962,N_20711);
xnor U21599 (N_21599,N_20612,N_20706);
nor U21600 (N_21600,N_21217,N_21365);
or U21601 (N_21601,N_21209,N_21269);
nand U21602 (N_21602,N_21525,N_21399);
xnor U21603 (N_21603,N_21099,N_21549);
nand U21604 (N_21604,N_21366,N_21530);
xnor U21605 (N_21605,N_21281,N_21285);
xor U21606 (N_21606,N_21489,N_21221);
nand U21607 (N_21607,N_21149,N_21581);
xor U21608 (N_21608,N_21477,N_21522);
xor U21609 (N_21609,N_21352,N_21174);
or U21610 (N_21610,N_21331,N_21214);
nor U21611 (N_21611,N_21015,N_21293);
nand U21612 (N_21612,N_21491,N_21077);
nor U21613 (N_21613,N_21304,N_21047);
and U21614 (N_21614,N_21026,N_21559);
nand U21615 (N_21615,N_21327,N_21248);
nor U21616 (N_21616,N_21592,N_21146);
and U21617 (N_21617,N_21247,N_21424);
or U21618 (N_21618,N_21091,N_21230);
xnor U21619 (N_21619,N_21268,N_21594);
nor U21620 (N_21620,N_21396,N_21052);
xnor U21621 (N_21621,N_21140,N_21188);
nor U21622 (N_21622,N_21419,N_21449);
nand U21623 (N_21623,N_21351,N_21289);
and U21624 (N_21624,N_21120,N_21429);
nor U21625 (N_21625,N_21215,N_21505);
xor U21626 (N_21626,N_21046,N_21595);
nand U21627 (N_21627,N_21073,N_21179);
nand U21628 (N_21628,N_21196,N_21253);
nand U21629 (N_21629,N_21361,N_21017);
xnor U21630 (N_21630,N_21133,N_21459);
nor U21631 (N_21631,N_21451,N_21488);
nor U21632 (N_21632,N_21078,N_21490);
nor U21633 (N_21633,N_21264,N_21409);
nand U21634 (N_21634,N_21598,N_21193);
nor U21635 (N_21635,N_21271,N_21212);
nor U21636 (N_21636,N_21266,N_21506);
or U21637 (N_21637,N_21296,N_21464);
nor U21638 (N_21638,N_21083,N_21108);
nand U21639 (N_21639,N_21245,N_21323);
and U21640 (N_21640,N_21080,N_21340);
xnor U21641 (N_21641,N_21104,N_21139);
nand U21642 (N_21642,N_21486,N_21313);
or U21643 (N_21643,N_21460,N_21481);
xor U21644 (N_21644,N_21030,N_21238);
nand U21645 (N_21645,N_21210,N_21584);
xnor U21646 (N_21646,N_21317,N_21412);
and U21647 (N_21647,N_21225,N_21154);
or U21648 (N_21648,N_21265,N_21569);
nor U21649 (N_21649,N_21256,N_21144);
nor U21650 (N_21650,N_21555,N_21158);
nor U21651 (N_21651,N_21336,N_21575);
nand U21652 (N_21652,N_21448,N_21462);
or U21653 (N_21653,N_21012,N_21004);
nor U21654 (N_21654,N_21413,N_21369);
nand U21655 (N_21655,N_21148,N_21276);
nand U21656 (N_21656,N_21498,N_21223);
nor U21657 (N_21657,N_21386,N_21586);
or U21658 (N_21658,N_21123,N_21367);
or U21659 (N_21659,N_21470,N_21437);
nand U21660 (N_21660,N_21025,N_21573);
or U21661 (N_21661,N_21392,N_21234);
nor U21662 (N_21662,N_21346,N_21049);
or U21663 (N_21663,N_21321,N_21356);
or U21664 (N_21664,N_21360,N_21492);
or U21665 (N_21665,N_21425,N_21391);
or U21666 (N_21666,N_21294,N_21385);
nor U21667 (N_21667,N_21041,N_21539);
and U21668 (N_21668,N_21572,N_21226);
nor U21669 (N_21669,N_21354,N_21087);
and U21670 (N_21670,N_21267,N_21095);
nand U21671 (N_21671,N_21301,N_21185);
xor U21672 (N_21672,N_21428,N_21009);
nor U21673 (N_21673,N_21348,N_21187);
xnor U21674 (N_21674,N_21329,N_21447);
or U21675 (N_21675,N_21473,N_21454);
or U21676 (N_21676,N_21241,N_21507);
and U21677 (N_21677,N_21560,N_21283);
or U21678 (N_21678,N_21275,N_21090);
nor U21679 (N_21679,N_21445,N_21007);
xor U21680 (N_21680,N_21084,N_21224);
or U21681 (N_21681,N_21307,N_21444);
nor U21682 (N_21682,N_21547,N_21337);
xnor U21683 (N_21683,N_21053,N_21054);
and U21684 (N_21684,N_21173,N_21517);
nor U21685 (N_21685,N_21551,N_21159);
or U21686 (N_21686,N_21531,N_21011);
nand U21687 (N_21687,N_21231,N_21190);
nand U21688 (N_21688,N_21119,N_21504);
and U21689 (N_21689,N_21060,N_21115);
or U21690 (N_21690,N_21161,N_21599);
xor U21691 (N_21691,N_21527,N_21420);
and U21692 (N_21692,N_21236,N_21567);
or U21693 (N_21693,N_21389,N_21455);
xnor U21694 (N_21694,N_21561,N_21254);
nand U21695 (N_21695,N_21545,N_21502);
nand U21696 (N_21696,N_21516,N_21178);
nor U21697 (N_21697,N_21111,N_21397);
or U21698 (N_21698,N_21362,N_21082);
or U21699 (N_21699,N_21280,N_21135);
and U21700 (N_21700,N_21151,N_21568);
xor U21701 (N_21701,N_21086,N_21045);
and U21702 (N_21702,N_21417,N_21203);
nor U21703 (N_21703,N_21192,N_21006);
xor U21704 (N_21704,N_21028,N_21353);
nor U21705 (N_21705,N_21194,N_21079);
or U21706 (N_21706,N_21003,N_21593);
and U21707 (N_21707,N_21503,N_21295);
and U21708 (N_21708,N_21242,N_21169);
or U21709 (N_21709,N_21411,N_21302);
xor U21710 (N_21710,N_21316,N_21358);
nand U21711 (N_21711,N_21122,N_21495);
nor U21712 (N_21712,N_21379,N_21333);
nor U21713 (N_21713,N_21483,N_21515);
xnor U21714 (N_21714,N_21533,N_21044);
and U21715 (N_21715,N_21363,N_21374);
nor U21716 (N_21716,N_21398,N_21128);
nor U21717 (N_21717,N_21322,N_21508);
or U21718 (N_21718,N_21163,N_21407);
and U21719 (N_21719,N_21220,N_21553);
or U21720 (N_21720,N_21585,N_21400);
or U21721 (N_21721,N_21463,N_21408);
or U21722 (N_21722,N_21040,N_21423);
and U21723 (N_21723,N_21499,N_21213);
xnor U21724 (N_21724,N_21309,N_21116);
nand U21725 (N_21725,N_21270,N_21450);
nor U21726 (N_21726,N_21556,N_21018);
nor U21727 (N_21727,N_21278,N_21075);
nor U21728 (N_21728,N_21570,N_21579);
nor U21729 (N_21729,N_21465,N_21546);
nor U21730 (N_21730,N_21421,N_21359);
and U21731 (N_21731,N_21021,N_21166);
and U21732 (N_21732,N_21022,N_21114);
nor U21733 (N_21733,N_21103,N_21482);
nor U21734 (N_21734,N_21291,N_21059);
and U21735 (N_21735,N_21107,N_21131);
nand U21736 (N_21736,N_21355,N_21055);
nor U21737 (N_21737,N_21211,N_21339);
xnor U21738 (N_21738,N_21132,N_21002);
or U21739 (N_21739,N_21577,N_21521);
nand U21740 (N_21740,N_21070,N_21514);
xor U21741 (N_21741,N_21534,N_21442);
xor U21742 (N_21742,N_21314,N_21582);
and U21743 (N_21743,N_21510,N_21526);
and U21744 (N_21744,N_21344,N_21023);
or U21745 (N_21745,N_21142,N_21176);
and U21746 (N_21746,N_21260,N_21479);
nor U21747 (N_21747,N_21251,N_21320);
and U21748 (N_21748,N_21427,N_21165);
or U21749 (N_21749,N_21298,N_21167);
and U21750 (N_21750,N_21402,N_21338);
nand U21751 (N_21751,N_21198,N_21162);
nor U21752 (N_21752,N_21164,N_21288);
nor U21753 (N_21753,N_21257,N_21147);
and U21754 (N_21754,N_21287,N_21117);
and U21755 (N_21755,N_21032,N_21019);
nor U21756 (N_21756,N_21461,N_21388);
xnor U21757 (N_21757,N_21284,N_21098);
xor U21758 (N_21758,N_21074,N_21175);
or U21759 (N_21759,N_21375,N_21529);
or U21760 (N_21760,N_21458,N_21347);
nor U21761 (N_21761,N_21239,N_21102);
nor U21762 (N_21762,N_21204,N_21171);
and U21763 (N_21763,N_21106,N_21118);
nor U21764 (N_21764,N_21562,N_21250);
nand U21765 (N_21765,N_21299,N_21141);
nand U21766 (N_21766,N_21010,N_21509);
or U21767 (N_21767,N_21031,N_21076);
nand U21768 (N_21768,N_21540,N_21100);
and U21769 (N_21769,N_21308,N_21172);
and U21770 (N_21770,N_21438,N_21050);
nand U21771 (N_21771,N_21195,N_21237);
and U21772 (N_21772,N_21382,N_21160);
and U21773 (N_21773,N_21168,N_21277);
or U21774 (N_21774,N_21094,N_21469);
nor U21775 (N_21775,N_21229,N_21512);
xnor U21776 (N_21776,N_21519,N_21487);
and U21777 (N_21777,N_21286,N_21152);
xnor U21778 (N_21778,N_21414,N_21051);
and U21779 (N_21779,N_21156,N_21043);
and U21780 (N_21780,N_21415,N_21186);
and U21781 (N_21781,N_21472,N_21484);
nand U21782 (N_21782,N_21564,N_21387);
nor U21783 (N_21783,N_21014,N_21008);
nor U21784 (N_21784,N_21112,N_21282);
xor U21785 (N_21785,N_21068,N_21441);
nand U21786 (N_21786,N_21199,N_21101);
xor U21787 (N_21787,N_21528,N_21452);
or U21788 (N_21788,N_21541,N_21588);
or U21789 (N_21789,N_21218,N_21081);
or U21790 (N_21790,N_21134,N_21071);
nor U21791 (N_21791,N_21467,N_21170);
xor U21792 (N_21792,N_21542,N_21453);
or U21793 (N_21793,N_21378,N_21093);
and U21794 (N_21794,N_21113,N_21088);
or U21795 (N_21795,N_21036,N_21001);
and U21796 (N_21796,N_21089,N_21349);
nor U21797 (N_21797,N_21532,N_21246);
nand U21798 (N_21798,N_21550,N_21207);
nand U21799 (N_21799,N_21129,N_21233);
and U21800 (N_21800,N_21303,N_21377);
or U21801 (N_21801,N_21216,N_21262);
and U21802 (N_21802,N_21205,N_21261);
or U21803 (N_21803,N_21566,N_21240);
nand U21804 (N_21804,N_21183,N_21056);
xnor U21805 (N_21805,N_21042,N_21381);
xnor U21806 (N_21806,N_21232,N_21370);
and U21807 (N_21807,N_21342,N_21350);
nand U21808 (N_21808,N_21235,N_21496);
nand U21809 (N_21809,N_21466,N_21290);
xor U21810 (N_21810,N_21145,N_21476);
nor U21811 (N_21811,N_21109,N_21580);
and U21812 (N_21812,N_21493,N_21252);
and U21813 (N_21813,N_21305,N_21578);
and U21814 (N_21814,N_21373,N_21371);
or U21815 (N_21815,N_21554,N_21124);
or U21816 (N_21816,N_21535,N_21180);
xnor U21817 (N_21817,N_21137,N_21596);
nor U21818 (N_21818,N_21039,N_21279);
xor U21819 (N_21819,N_21273,N_21368);
xor U21820 (N_21820,N_21272,N_21153);
xor U21821 (N_21821,N_21405,N_21474);
xnor U21822 (N_21822,N_21416,N_21155);
and U21823 (N_21823,N_21332,N_21064);
nand U21824 (N_21824,N_21538,N_21457);
nor U21825 (N_21825,N_21058,N_21244);
nor U21826 (N_21826,N_21544,N_21263);
and U21827 (N_21827,N_21105,N_21468);
or U21828 (N_21828,N_21523,N_21557);
xor U21829 (N_21829,N_21182,N_21548);
and U21830 (N_21830,N_21430,N_21418);
or U21831 (N_21831,N_21587,N_21027);
nor U21832 (N_21832,N_21552,N_21243);
nor U21833 (N_21833,N_21357,N_21334);
nor U21834 (N_21834,N_21406,N_21292);
or U21835 (N_21835,N_21583,N_21311);
xor U21836 (N_21836,N_21063,N_21315);
nor U21837 (N_21837,N_21364,N_21037);
nor U21838 (N_21838,N_21067,N_21020);
or U21839 (N_21839,N_21258,N_21536);
xnor U21840 (N_21840,N_21069,N_21410);
or U21841 (N_21841,N_21033,N_21208);
xnor U21842 (N_21842,N_21395,N_21383);
nor U21843 (N_21843,N_21440,N_21434);
nor U21844 (N_21844,N_21048,N_21274);
nand U21845 (N_21845,N_21125,N_21376);
or U21846 (N_21846,N_21590,N_21439);
or U21847 (N_21847,N_21057,N_21576);
and U21848 (N_21848,N_21335,N_21518);
and U21849 (N_21849,N_21494,N_21571);
or U21850 (N_21850,N_21431,N_21543);
and U21851 (N_21851,N_21558,N_21456);
xnor U21852 (N_21852,N_21497,N_21034);
or U21853 (N_21853,N_21306,N_21197);
nor U21854 (N_21854,N_21478,N_21443);
nand U21855 (N_21855,N_21005,N_21157);
nand U21856 (N_21856,N_21259,N_21136);
nand U21857 (N_21857,N_21390,N_21181);
nor U21858 (N_21858,N_21227,N_21249);
or U21859 (N_21859,N_21061,N_21372);
and U21860 (N_21860,N_21511,N_21597);
xor U21861 (N_21861,N_21065,N_21085);
or U21862 (N_21862,N_21013,N_21480);
and U21863 (N_21863,N_21016,N_21485);
nor U21864 (N_21864,N_21435,N_21038);
xnor U21865 (N_21865,N_21401,N_21228);
or U21866 (N_21866,N_21130,N_21343);
nand U21867 (N_21867,N_21029,N_21121);
xor U21868 (N_21868,N_21426,N_21471);
and U21869 (N_21869,N_21150,N_21345);
and U21870 (N_21870,N_21110,N_21319);
nand U21871 (N_21871,N_21446,N_21189);
nand U21872 (N_21872,N_21436,N_21310);
xnor U21873 (N_21873,N_21330,N_21206);
nand U21874 (N_21874,N_21312,N_21324);
nor U21875 (N_21875,N_21066,N_21024);
xnor U21876 (N_21876,N_21404,N_21328);
and U21877 (N_21877,N_21341,N_21191);
xnor U21878 (N_21878,N_21325,N_21062);
and U21879 (N_21879,N_21138,N_21565);
nor U21880 (N_21880,N_21563,N_21184);
or U21881 (N_21881,N_21393,N_21500);
xor U21882 (N_21882,N_21520,N_21219);
nand U21883 (N_21883,N_21127,N_21326);
xnor U21884 (N_21884,N_21318,N_21297);
nor U21885 (N_21885,N_21384,N_21574);
nor U21886 (N_21886,N_21475,N_21000);
nor U21887 (N_21887,N_21537,N_21202);
or U21888 (N_21888,N_21177,N_21097);
nor U21889 (N_21889,N_21200,N_21072);
nor U21890 (N_21890,N_21403,N_21432);
xor U21891 (N_21891,N_21591,N_21433);
or U21892 (N_21892,N_21035,N_21143);
xnor U21893 (N_21893,N_21092,N_21222);
nor U21894 (N_21894,N_21096,N_21524);
nand U21895 (N_21895,N_21300,N_21201);
and U21896 (N_21896,N_21501,N_21380);
nand U21897 (N_21897,N_21422,N_21126);
nor U21898 (N_21898,N_21589,N_21255);
or U21899 (N_21899,N_21394,N_21513);
nand U21900 (N_21900,N_21348,N_21350);
or U21901 (N_21901,N_21513,N_21205);
nor U21902 (N_21902,N_21115,N_21192);
xor U21903 (N_21903,N_21054,N_21212);
nor U21904 (N_21904,N_21422,N_21377);
and U21905 (N_21905,N_21397,N_21078);
nor U21906 (N_21906,N_21254,N_21029);
xor U21907 (N_21907,N_21286,N_21093);
nor U21908 (N_21908,N_21499,N_21290);
and U21909 (N_21909,N_21055,N_21251);
and U21910 (N_21910,N_21282,N_21532);
xnor U21911 (N_21911,N_21179,N_21595);
nor U21912 (N_21912,N_21200,N_21301);
nand U21913 (N_21913,N_21237,N_21226);
and U21914 (N_21914,N_21024,N_21002);
or U21915 (N_21915,N_21330,N_21491);
or U21916 (N_21916,N_21380,N_21349);
nor U21917 (N_21917,N_21131,N_21565);
xnor U21918 (N_21918,N_21089,N_21314);
nor U21919 (N_21919,N_21080,N_21425);
nor U21920 (N_21920,N_21091,N_21503);
or U21921 (N_21921,N_21490,N_21246);
nand U21922 (N_21922,N_21480,N_21492);
or U21923 (N_21923,N_21089,N_21023);
nand U21924 (N_21924,N_21151,N_21150);
and U21925 (N_21925,N_21533,N_21342);
xnor U21926 (N_21926,N_21104,N_21058);
and U21927 (N_21927,N_21374,N_21569);
or U21928 (N_21928,N_21370,N_21320);
or U21929 (N_21929,N_21097,N_21455);
xnor U21930 (N_21930,N_21379,N_21502);
nand U21931 (N_21931,N_21119,N_21390);
nand U21932 (N_21932,N_21413,N_21491);
or U21933 (N_21933,N_21210,N_21595);
and U21934 (N_21934,N_21253,N_21481);
or U21935 (N_21935,N_21150,N_21171);
nand U21936 (N_21936,N_21535,N_21475);
and U21937 (N_21937,N_21438,N_21484);
and U21938 (N_21938,N_21033,N_21329);
nor U21939 (N_21939,N_21289,N_21369);
nand U21940 (N_21940,N_21439,N_21214);
nand U21941 (N_21941,N_21040,N_21186);
nand U21942 (N_21942,N_21275,N_21591);
nor U21943 (N_21943,N_21060,N_21429);
xor U21944 (N_21944,N_21020,N_21389);
nand U21945 (N_21945,N_21343,N_21297);
or U21946 (N_21946,N_21016,N_21057);
or U21947 (N_21947,N_21192,N_21432);
or U21948 (N_21948,N_21478,N_21531);
xor U21949 (N_21949,N_21460,N_21444);
and U21950 (N_21950,N_21289,N_21125);
and U21951 (N_21951,N_21505,N_21495);
nor U21952 (N_21952,N_21238,N_21553);
nor U21953 (N_21953,N_21158,N_21432);
and U21954 (N_21954,N_21563,N_21361);
or U21955 (N_21955,N_21212,N_21080);
xnor U21956 (N_21956,N_21509,N_21004);
nor U21957 (N_21957,N_21184,N_21000);
nor U21958 (N_21958,N_21299,N_21103);
or U21959 (N_21959,N_21256,N_21479);
nand U21960 (N_21960,N_21116,N_21265);
and U21961 (N_21961,N_21059,N_21384);
nor U21962 (N_21962,N_21273,N_21367);
or U21963 (N_21963,N_21170,N_21062);
nand U21964 (N_21964,N_21305,N_21434);
nor U21965 (N_21965,N_21207,N_21551);
nor U21966 (N_21966,N_21021,N_21281);
nand U21967 (N_21967,N_21351,N_21196);
nand U21968 (N_21968,N_21135,N_21074);
or U21969 (N_21969,N_21222,N_21471);
or U21970 (N_21970,N_21092,N_21525);
xor U21971 (N_21971,N_21388,N_21550);
nand U21972 (N_21972,N_21487,N_21473);
or U21973 (N_21973,N_21567,N_21202);
xor U21974 (N_21974,N_21422,N_21375);
nand U21975 (N_21975,N_21508,N_21468);
nand U21976 (N_21976,N_21267,N_21553);
xor U21977 (N_21977,N_21251,N_21166);
and U21978 (N_21978,N_21505,N_21582);
xor U21979 (N_21979,N_21190,N_21504);
or U21980 (N_21980,N_21364,N_21327);
nand U21981 (N_21981,N_21452,N_21390);
and U21982 (N_21982,N_21357,N_21175);
xnor U21983 (N_21983,N_21121,N_21562);
nand U21984 (N_21984,N_21571,N_21058);
nor U21985 (N_21985,N_21518,N_21198);
and U21986 (N_21986,N_21465,N_21318);
nor U21987 (N_21987,N_21555,N_21557);
and U21988 (N_21988,N_21302,N_21585);
nand U21989 (N_21989,N_21108,N_21564);
or U21990 (N_21990,N_21442,N_21443);
or U21991 (N_21991,N_21431,N_21538);
nor U21992 (N_21992,N_21142,N_21274);
and U21993 (N_21993,N_21166,N_21534);
or U21994 (N_21994,N_21056,N_21224);
and U21995 (N_21995,N_21177,N_21457);
nand U21996 (N_21996,N_21247,N_21567);
or U21997 (N_21997,N_21201,N_21241);
nand U21998 (N_21998,N_21427,N_21441);
nor U21999 (N_21999,N_21498,N_21537);
or U22000 (N_22000,N_21180,N_21383);
nor U22001 (N_22001,N_21462,N_21101);
and U22002 (N_22002,N_21501,N_21307);
or U22003 (N_22003,N_21205,N_21191);
or U22004 (N_22004,N_21495,N_21178);
nor U22005 (N_22005,N_21316,N_21367);
xor U22006 (N_22006,N_21131,N_21591);
or U22007 (N_22007,N_21155,N_21000);
nor U22008 (N_22008,N_21483,N_21584);
nor U22009 (N_22009,N_21253,N_21102);
nor U22010 (N_22010,N_21072,N_21136);
nand U22011 (N_22011,N_21587,N_21242);
xnor U22012 (N_22012,N_21589,N_21121);
and U22013 (N_22013,N_21053,N_21327);
and U22014 (N_22014,N_21413,N_21140);
and U22015 (N_22015,N_21472,N_21322);
and U22016 (N_22016,N_21545,N_21005);
or U22017 (N_22017,N_21150,N_21311);
nor U22018 (N_22018,N_21402,N_21156);
or U22019 (N_22019,N_21438,N_21153);
and U22020 (N_22020,N_21381,N_21040);
nand U22021 (N_22021,N_21357,N_21054);
or U22022 (N_22022,N_21206,N_21103);
or U22023 (N_22023,N_21290,N_21010);
and U22024 (N_22024,N_21029,N_21387);
xnor U22025 (N_22025,N_21215,N_21132);
nor U22026 (N_22026,N_21331,N_21537);
and U22027 (N_22027,N_21113,N_21433);
xnor U22028 (N_22028,N_21002,N_21514);
nor U22029 (N_22029,N_21340,N_21093);
and U22030 (N_22030,N_21106,N_21417);
nand U22031 (N_22031,N_21189,N_21012);
and U22032 (N_22032,N_21187,N_21231);
or U22033 (N_22033,N_21394,N_21156);
xor U22034 (N_22034,N_21208,N_21472);
nor U22035 (N_22035,N_21537,N_21309);
xnor U22036 (N_22036,N_21149,N_21349);
or U22037 (N_22037,N_21006,N_21081);
nor U22038 (N_22038,N_21392,N_21393);
or U22039 (N_22039,N_21510,N_21048);
or U22040 (N_22040,N_21342,N_21559);
xor U22041 (N_22041,N_21519,N_21513);
nor U22042 (N_22042,N_21001,N_21364);
or U22043 (N_22043,N_21307,N_21176);
and U22044 (N_22044,N_21039,N_21489);
or U22045 (N_22045,N_21578,N_21423);
nor U22046 (N_22046,N_21368,N_21143);
xnor U22047 (N_22047,N_21178,N_21330);
nand U22048 (N_22048,N_21254,N_21275);
xor U22049 (N_22049,N_21397,N_21254);
or U22050 (N_22050,N_21403,N_21338);
or U22051 (N_22051,N_21232,N_21208);
or U22052 (N_22052,N_21494,N_21402);
and U22053 (N_22053,N_21247,N_21147);
and U22054 (N_22054,N_21207,N_21150);
or U22055 (N_22055,N_21528,N_21136);
and U22056 (N_22056,N_21125,N_21377);
or U22057 (N_22057,N_21033,N_21504);
xor U22058 (N_22058,N_21063,N_21599);
xnor U22059 (N_22059,N_21160,N_21364);
xor U22060 (N_22060,N_21227,N_21291);
or U22061 (N_22061,N_21500,N_21375);
xnor U22062 (N_22062,N_21402,N_21382);
xor U22063 (N_22063,N_21192,N_21220);
xnor U22064 (N_22064,N_21592,N_21536);
or U22065 (N_22065,N_21571,N_21000);
nor U22066 (N_22066,N_21583,N_21083);
nor U22067 (N_22067,N_21585,N_21088);
and U22068 (N_22068,N_21108,N_21551);
or U22069 (N_22069,N_21093,N_21064);
or U22070 (N_22070,N_21119,N_21538);
or U22071 (N_22071,N_21134,N_21102);
or U22072 (N_22072,N_21490,N_21100);
nor U22073 (N_22073,N_21488,N_21031);
xor U22074 (N_22074,N_21587,N_21147);
nor U22075 (N_22075,N_21570,N_21282);
and U22076 (N_22076,N_21497,N_21067);
nand U22077 (N_22077,N_21551,N_21483);
xor U22078 (N_22078,N_21367,N_21371);
xnor U22079 (N_22079,N_21585,N_21589);
and U22080 (N_22080,N_21456,N_21512);
xnor U22081 (N_22081,N_21546,N_21332);
xnor U22082 (N_22082,N_21207,N_21381);
nand U22083 (N_22083,N_21166,N_21344);
or U22084 (N_22084,N_21182,N_21301);
and U22085 (N_22085,N_21243,N_21287);
or U22086 (N_22086,N_21369,N_21533);
or U22087 (N_22087,N_21587,N_21382);
xor U22088 (N_22088,N_21458,N_21281);
and U22089 (N_22089,N_21103,N_21339);
and U22090 (N_22090,N_21050,N_21373);
xnor U22091 (N_22091,N_21385,N_21522);
nor U22092 (N_22092,N_21458,N_21287);
nand U22093 (N_22093,N_21159,N_21105);
nor U22094 (N_22094,N_21040,N_21561);
nor U22095 (N_22095,N_21555,N_21050);
or U22096 (N_22096,N_21129,N_21230);
nor U22097 (N_22097,N_21019,N_21359);
and U22098 (N_22098,N_21297,N_21278);
nor U22099 (N_22099,N_21142,N_21158);
nor U22100 (N_22100,N_21357,N_21231);
xnor U22101 (N_22101,N_21429,N_21573);
and U22102 (N_22102,N_21348,N_21443);
nand U22103 (N_22103,N_21244,N_21582);
or U22104 (N_22104,N_21203,N_21070);
xor U22105 (N_22105,N_21174,N_21228);
xnor U22106 (N_22106,N_21325,N_21215);
nand U22107 (N_22107,N_21275,N_21213);
nand U22108 (N_22108,N_21238,N_21215);
nor U22109 (N_22109,N_21404,N_21210);
and U22110 (N_22110,N_21200,N_21041);
or U22111 (N_22111,N_21021,N_21574);
and U22112 (N_22112,N_21447,N_21232);
or U22113 (N_22113,N_21328,N_21351);
and U22114 (N_22114,N_21347,N_21563);
nand U22115 (N_22115,N_21141,N_21504);
xor U22116 (N_22116,N_21122,N_21144);
and U22117 (N_22117,N_21170,N_21294);
xnor U22118 (N_22118,N_21006,N_21546);
and U22119 (N_22119,N_21436,N_21362);
and U22120 (N_22120,N_21397,N_21417);
nand U22121 (N_22121,N_21124,N_21241);
and U22122 (N_22122,N_21197,N_21288);
xor U22123 (N_22123,N_21110,N_21364);
xor U22124 (N_22124,N_21299,N_21497);
or U22125 (N_22125,N_21050,N_21428);
nor U22126 (N_22126,N_21280,N_21470);
or U22127 (N_22127,N_21427,N_21288);
nand U22128 (N_22128,N_21252,N_21464);
nor U22129 (N_22129,N_21482,N_21039);
or U22130 (N_22130,N_21447,N_21519);
nand U22131 (N_22131,N_21248,N_21433);
nand U22132 (N_22132,N_21026,N_21583);
or U22133 (N_22133,N_21168,N_21094);
or U22134 (N_22134,N_21462,N_21495);
and U22135 (N_22135,N_21277,N_21478);
or U22136 (N_22136,N_21424,N_21302);
and U22137 (N_22137,N_21279,N_21241);
or U22138 (N_22138,N_21050,N_21366);
xnor U22139 (N_22139,N_21470,N_21584);
and U22140 (N_22140,N_21283,N_21175);
and U22141 (N_22141,N_21534,N_21585);
or U22142 (N_22142,N_21079,N_21471);
nor U22143 (N_22143,N_21507,N_21302);
or U22144 (N_22144,N_21005,N_21252);
xor U22145 (N_22145,N_21100,N_21047);
and U22146 (N_22146,N_21055,N_21235);
and U22147 (N_22147,N_21303,N_21368);
nand U22148 (N_22148,N_21032,N_21003);
nor U22149 (N_22149,N_21157,N_21096);
xor U22150 (N_22150,N_21011,N_21115);
nor U22151 (N_22151,N_21035,N_21480);
and U22152 (N_22152,N_21327,N_21352);
and U22153 (N_22153,N_21469,N_21482);
or U22154 (N_22154,N_21492,N_21039);
and U22155 (N_22155,N_21232,N_21130);
nand U22156 (N_22156,N_21127,N_21053);
nand U22157 (N_22157,N_21157,N_21067);
or U22158 (N_22158,N_21523,N_21353);
or U22159 (N_22159,N_21146,N_21022);
nand U22160 (N_22160,N_21365,N_21209);
and U22161 (N_22161,N_21527,N_21214);
or U22162 (N_22162,N_21409,N_21498);
xor U22163 (N_22163,N_21062,N_21493);
nand U22164 (N_22164,N_21148,N_21560);
or U22165 (N_22165,N_21488,N_21128);
nand U22166 (N_22166,N_21578,N_21080);
xnor U22167 (N_22167,N_21216,N_21492);
and U22168 (N_22168,N_21280,N_21483);
nor U22169 (N_22169,N_21212,N_21342);
and U22170 (N_22170,N_21461,N_21143);
nand U22171 (N_22171,N_21308,N_21147);
or U22172 (N_22172,N_21119,N_21599);
nand U22173 (N_22173,N_21163,N_21046);
nor U22174 (N_22174,N_21186,N_21220);
and U22175 (N_22175,N_21010,N_21107);
xnor U22176 (N_22176,N_21392,N_21002);
and U22177 (N_22177,N_21483,N_21399);
and U22178 (N_22178,N_21537,N_21501);
nor U22179 (N_22179,N_21382,N_21381);
or U22180 (N_22180,N_21074,N_21516);
xnor U22181 (N_22181,N_21043,N_21589);
nand U22182 (N_22182,N_21576,N_21350);
or U22183 (N_22183,N_21137,N_21274);
xor U22184 (N_22184,N_21516,N_21028);
and U22185 (N_22185,N_21017,N_21575);
nand U22186 (N_22186,N_21417,N_21558);
xnor U22187 (N_22187,N_21056,N_21384);
or U22188 (N_22188,N_21501,N_21403);
or U22189 (N_22189,N_21266,N_21243);
or U22190 (N_22190,N_21584,N_21169);
nand U22191 (N_22191,N_21536,N_21144);
nor U22192 (N_22192,N_21491,N_21376);
nand U22193 (N_22193,N_21196,N_21431);
or U22194 (N_22194,N_21564,N_21113);
or U22195 (N_22195,N_21470,N_21255);
and U22196 (N_22196,N_21028,N_21196);
nand U22197 (N_22197,N_21200,N_21052);
and U22198 (N_22198,N_21323,N_21304);
and U22199 (N_22199,N_21306,N_21561);
nor U22200 (N_22200,N_21611,N_21857);
and U22201 (N_22201,N_21657,N_22016);
and U22202 (N_22202,N_21850,N_22027);
nand U22203 (N_22203,N_21854,N_21874);
nor U22204 (N_22204,N_21767,N_21921);
nand U22205 (N_22205,N_21714,N_22086);
nor U22206 (N_22206,N_21839,N_21630);
xnor U22207 (N_22207,N_22190,N_22067);
nand U22208 (N_22208,N_21965,N_22178);
nand U22209 (N_22209,N_21866,N_21710);
xnor U22210 (N_22210,N_21761,N_21875);
or U22211 (N_22211,N_21898,N_22182);
xor U22212 (N_22212,N_22117,N_22012);
and U22213 (N_22213,N_21820,N_21750);
or U22214 (N_22214,N_21703,N_22163);
nand U22215 (N_22215,N_21887,N_21787);
nor U22216 (N_22216,N_22164,N_21963);
and U22217 (N_22217,N_21769,N_22015);
and U22218 (N_22218,N_22127,N_22056);
or U22219 (N_22219,N_21666,N_22156);
xnor U22220 (N_22220,N_21958,N_21731);
nand U22221 (N_22221,N_22011,N_21999);
nand U22222 (N_22222,N_21735,N_22158);
nor U22223 (N_22223,N_22186,N_22151);
nor U22224 (N_22224,N_21723,N_22169);
and U22225 (N_22225,N_21784,N_22116);
nand U22226 (N_22226,N_21929,N_22106);
nand U22227 (N_22227,N_22013,N_21834);
or U22228 (N_22228,N_22197,N_21986);
or U22229 (N_22229,N_21851,N_21702);
xor U22230 (N_22230,N_22179,N_22032);
xor U22231 (N_22231,N_21924,N_21638);
or U22232 (N_22232,N_21847,N_21737);
xor U22233 (N_22233,N_21890,N_21892);
and U22234 (N_22234,N_22039,N_22193);
or U22235 (N_22235,N_21619,N_21713);
xnor U22236 (N_22236,N_21604,N_21828);
and U22237 (N_22237,N_21726,N_22189);
and U22238 (N_22238,N_21815,N_22148);
and U22239 (N_22239,N_21936,N_21801);
or U22240 (N_22240,N_21848,N_21639);
or U22241 (N_22241,N_22129,N_22160);
xor U22242 (N_22242,N_22187,N_21774);
and U22243 (N_22243,N_22074,N_21602);
xnor U22244 (N_22244,N_22022,N_22131);
or U22245 (N_22245,N_21669,N_22119);
nand U22246 (N_22246,N_21880,N_21681);
nor U22247 (N_22247,N_21653,N_22143);
nor U22248 (N_22248,N_22034,N_22084);
or U22249 (N_22249,N_22052,N_22043);
xnor U22250 (N_22250,N_21660,N_21625);
nand U22251 (N_22251,N_21860,N_22089);
xnor U22252 (N_22252,N_21951,N_22007);
xnor U22253 (N_22253,N_22088,N_22159);
nand U22254 (N_22254,N_21684,N_21891);
nand U22255 (N_22255,N_21606,N_21833);
xor U22256 (N_22256,N_22188,N_21682);
nand U22257 (N_22257,N_21800,N_22018);
nand U22258 (N_22258,N_21778,N_22114);
nand U22259 (N_22259,N_21786,N_22110);
and U22260 (N_22260,N_21843,N_21781);
and U22261 (N_22261,N_21996,N_22126);
xor U22262 (N_22262,N_21941,N_22028);
nand U22263 (N_22263,N_21841,N_21937);
nand U22264 (N_22264,N_21728,N_21616);
or U22265 (N_22265,N_21867,N_22140);
and U22266 (N_22266,N_21915,N_21830);
nor U22267 (N_22267,N_22181,N_21837);
nor U22268 (N_22268,N_21995,N_21722);
xnor U22269 (N_22269,N_22055,N_22115);
and U22270 (N_22270,N_22132,N_21642);
or U22271 (N_22271,N_21945,N_21708);
nor U22272 (N_22272,N_21683,N_22167);
or U22273 (N_22273,N_21641,N_21677);
and U22274 (N_22274,N_21897,N_21966);
and U22275 (N_22275,N_21738,N_21791);
xor U22276 (N_22276,N_21690,N_21975);
and U22277 (N_22277,N_21615,N_21698);
nor U22278 (N_22278,N_21705,N_22014);
xor U22279 (N_22279,N_22057,N_21893);
nor U22280 (N_22280,N_21836,N_21755);
xnor U22281 (N_22281,N_21845,N_21699);
and U22282 (N_22282,N_21647,N_22085);
and U22283 (N_22283,N_21931,N_22105);
nor U22284 (N_22284,N_21785,N_21668);
or U22285 (N_22285,N_22079,N_21852);
nand U22286 (N_22286,N_21600,N_21656);
or U22287 (N_22287,N_21869,N_21806);
nor U22288 (N_22288,N_22196,N_22121);
nand U22289 (N_22289,N_21825,N_21691);
or U22290 (N_22290,N_21959,N_22162);
nand U22291 (N_22291,N_21745,N_21706);
or U22292 (N_22292,N_21911,N_21829);
xor U22293 (N_22293,N_22120,N_22113);
or U22294 (N_22294,N_21992,N_21650);
nor U22295 (N_22295,N_22112,N_22104);
xor U22296 (N_22296,N_22198,N_21694);
nand U22297 (N_22297,N_21909,N_21809);
nor U22298 (N_22298,N_21918,N_22049);
and U22299 (N_22299,N_21980,N_21700);
nor U22300 (N_22300,N_22137,N_22036);
and U22301 (N_22301,N_22175,N_21917);
or U22302 (N_22302,N_22058,N_21881);
xnor U22303 (N_22303,N_21969,N_21664);
nand U22304 (N_22304,N_21832,N_22145);
and U22305 (N_22305,N_21756,N_22176);
or U22306 (N_22306,N_22122,N_21620);
nand U22307 (N_22307,N_22184,N_21676);
and U22308 (N_22308,N_22069,N_21842);
and U22309 (N_22309,N_21824,N_21725);
and U22310 (N_22310,N_21923,N_21793);
or U22311 (N_22311,N_21811,N_21776);
nand U22312 (N_22312,N_21766,N_21943);
and U22313 (N_22313,N_21822,N_21721);
and U22314 (N_22314,N_22053,N_21888);
nor U22315 (N_22315,N_21622,N_21973);
xor U22316 (N_22316,N_21695,N_22083);
or U22317 (N_22317,N_21686,N_21868);
and U22318 (N_22318,N_21910,N_21991);
and U22319 (N_22319,N_21914,N_21982);
nor U22320 (N_22320,N_21783,N_21763);
xor U22321 (N_22321,N_21944,N_21974);
xor U22322 (N_22322,N_22020,N_21771);
xnor U22323 (N_22323,N_22098,N_22174);
or U22324 (N_22324,N_21905,N_21717);
or U22325 (N_22325,N_21729,N_22109);
nand U22326 (N_22326,N_21614,N_21633);
nor U22327 (N_22327,N_21777,N_21961);
or U22328 (N_22328,N_21817,N_21696);
xor U22329 (N_22329,N_21697,N_21605);
xnor U22330 (N_22330,N_22153,N_21716);
and U22331 (N_22331,N_21758,N_22050);
and U22332 (N_22332,N_21707,N_22030);
or U22333 (N_22333,N_21799,N_22038);
nand U22334 (N_22334,N_21997,N_21925);
nor U22335 (N_22335,N_21912,N_21913);
or U22336 (N_22336,N_21636,N_22044);
nor U22337 (N_22337,N_22173,N_21709);
nor U22338 (N_22338,N_22063,N_21687);
nor U22339 (N_22339,N_21648,N_21727);
nor U22340 (N_22340,N_21952,N_22177);
nor U22341 (N_22341,N_22191,N_22047);
xor U22342 (N_22342,N_21661,N_21818);
nor U22343 (N_22343,N_21623,N_21916);
or U22344 (N_22344,N_21688,N_21775);
nand U22345 (N_22345,N_21994,N_21844);
or U22346 (N_22346,N_21928,N_21645);
and U22347 (N_22347,N_21862,N_22138);
nor U22348 (N_22348,N_21835,N_21603);
nand U22349 (N_22349,N_21972,N_21896);
nor U22350 (N_22350,N_21654,N_22144);
and U22351 (N_22351,N_21878,N_22005);
and U22352 (N_22352,N_21797,N_21938);
and U22353 (N_22353,N_21990,N_22170);
or U22354 (N_22354,N_21689,N_22006);
nand U22355 (N_22355,N_21627,N_21617);
nand U22356 (N_22356,N_22054,N_22192);
xor U22357 (N_22357,N_21930,N_22024);
xor U22358 (N_22358,N_21629,N_21858);
nand U22359 (N_22359,N_21855,N_21672);
nand U22360 (N_22360,N_21673,N_21987);
and U22361 (N_22361,N_22070,N_21864);
xnor U22362 (N_22362,N_21838,N_21655);
and U22363 (N_22363,N_21652,N_22108);
and U22364 (N_22364,N_22072,N_22095);
nand U22365 (N_22365,N_22097,N_21610);
and U22366 (N_22366,N_21821,N_22107);
xor U22367 (N_22367,N_21704,N_22017);
and U22368 (N_22368,N_21747,N_21635);
and U22369 (N_22369,N_22139,N_22092);
and U22370 (N_22370,N_21871,N_21979);
or U22371 (N_22371,N_22009,N_21612);
and U22372 (N_22372,N_21993,N_21876);
nand U22373 (N_22373,N_21927,N_21662);
and U22374 (N_22374,N_22155,N_21624);
xnor U22375 (N_22375,N_21663,N_21746);
or U22376 (N_22376,N_21906,N_22029);
nor U22377 (N_22377,N_22080,N_21877);
nand U22378 (N_22378,N_21794,N_21601);
nand U22379 (N_22379,N_21649,N_22035);
or U22380 (N_22380,N_21609,N_21718);
nand U22381 (N_22381,N_21751,N_22099);
and U22382 (N_22382,N_22041,N_22147);
or U22383 (N_22383,N_21935,N_21957);
or U22384 (N_22384,N_21953,N_21949);
nand U22385 (N_22385,N_21846,N_22076);
or U22386 (N_22386,N_22118,N_21765);
nand U22387 (N_22387,N_21651,N_21680);
xor U22388 (N_22388,N_22135,N_22002);
nand U22389 (N_22389,N_21863,N_22051);
xor U22390 (N_22390,N_22031,N_21643);
and U22391 (N_22391,N_21886,N_21740);
nand U22392 (N_22392,N_21899,N_22165);
and U22393 (N_22393,N_21637,N_22059);
and U22394 (N_22394,N_22141,N_21968);
and U22395 (N_22395,N_21970,N_22185);
and U22396 (N_22396,N_21849,N_21805);
or U22397 (N_22397,N_21724,N_21967);
and U22398 (N_22398,N_22171,N_22096);
or U22399 (N_22399,N_21632,N_21895);
nand U22400 (N_22400,N_21932,N_21856);
nand U22401 (N_22401,N_21613,N_21960);
or U22402 (N_22402,N_22021,N_21883);
nand U22403 (N_22403,N_21762,N_21807);
nand U22404 (N_22404,N_22068,N_22061);
and U22405 (N_22405,N_21901,N_22195);
xnor U22406 (N_22406,N_21665,N_21978);
nor U22407 (N_22407,N_21768,N_22172);
xor U22408 (N_22408,N_21940,N_22037);
nand U22409 (N_22409,N_21808,N_21942);
or U22410 (N_22410,N_21667,N_21872);
nand U22411 (N_22411,N_22183,N_21674);
or U22412 (N_22412,N_22046,N_21865);
nor U22413 (N_22413,N_22103,N_21810);
nand U22414 (N_22414,N_21964,N_22136);
xor U22415 (N_22415,N_22154,N_22128);
or U22416 (N_22416,N_21802,N_21922);
nand U22417 (N_22417,N_22142,N_21983);
nand U22418 (N_22418,N_22008,N_21628);
or U22419 (N_22419,N_22146,N_21788);
xor U22420 (N_22420,N_21780,N_21903);
and U22421 (N_22421,N_22010,N_21753);
and U22422 (N_22422,N_21692,N_22000);
xor U22423 (N_22423,N_21671,N_21889);
nand U22424 (N_22424,N_21823,N_21947);
nor U22425 (N_22425,N_22075,N_22025);
nor U22426 (N_22426,N_21946,N_21744);
or U22427 (N_22427,N_21962,N_21926);
or U22428 (N_22428,N_21840,N_22199);
or U22429 (N_22429,N_21646,N_21779);
xor U22430 (N_22430,N_21908,N_22123);
or U22431 (N_22431,N_21748,N_22161);
or U22432 (N_22432,N_22111,N_21827);
or U22433 (N_22433,N_21782,N_21796);
nand U22434 (N_22434,N_21773,N_21741);
xnor U22435 (N_22435,N_22033,N_21658);
xor U22436 (N_22436,N_21789,N_21770);
xor U22437 (N_22437,N_22060,N_21733);
nand U22438 (N_22438,N_21772,N_21795);
and U22439 (N_22439,N_21988,N_21920);
nor U22440 (N_22440,N_22082,N_21985);
and U22441 (N_22441,N_22157,N_21948);
nand U22442 (N_22442,N_21732,N_21826);
nor U22443 (N_22443,N_21607,N_22062);
nor U22444 (N_22444,N_21739,N_21644);
xor U22445 (N_22445,N_21950,N_21907);
xnor U22446 (N_22446,N_21618,N_22042);
and U22447 (N_22447,N_21879,N_21870);
nor U22448 (N_22448,N_21812,N_21933);
nor U22449 (N_22449,N_22134,N_21720);
and U22450 (N_22450,N_21659,N_21885);
or U22451 (N_22451,N_21873,N_21956);
and U22452 (N_22452,N_21955,N_22149);
or U22453 (N_22453,N_22066,N_22004);
nor U22454 (N_22454,N_21814,N_21631);
nor U22455 (N_22455,N_22077,N_21831);
and U22456 (N_22456,N_21989,N_22023);
nand U22457 (N_22457,N_21904,N_21884);
or U22458 (N_22458,N_21900,N_21749);
or U22459 (N_22459,N_21813,N_21971);
and U22460 (N_22460,N_21790,N_21736);
or U22461 (N_22461,N_22090,N_21804);
and U22462 (N_22462,N_21608,N_22003);
and U22463 (N_22463,N_22166,N_22133);
or U22464 (N_22464,N_22087,N_21894);
xnor U22465 (N_22465,N_22065,N_21757);
and U22466 (N_22466,N_22026,N_21977);
nor U22467 (N_22467,N_22168,N_22001);
or U22468 (N_22468,N_21853,N_21816);
xnor U22469 (N_22469,N_21939,N_22094);
or U22470 (N_22470,N_21712,N_22019);
nor U22471 (N_22471,N_21752,N_22150);
or U22472 (N_22472,N_21754,N_22100);
nand U22473 (N_22473,N_21719,N_21634);
and U22474 (N_22474,N_22078,N_21760);
or U22475 (N_22475,N_21819,N_21859);
or U22476 (N_22476,N_21679,N_22130);
nand U22477 (N_22477,N_22093,N_21626);
and U22478 (N_22478,N_21743,N_21730);
or U22479 (N_22479,N_22071,N_21902);
nand U22480 (N_22480,N_21792,N_22102);
nand U22481 (N_22481,N_21798,N_21711);
nor U22482 (N_22482,N_21764,N_21861);
nand U22483 (N_22483,N_21670,N_22064);
nand U22484 (N_22484,N_21640,N_21882);
nand U22485 (N_22485,N_22091,N_22040);
or U22486 (N_22486,N_21919,N_21734);
and U22487 (N_22487,N_21715,N_21984);
nand U22488 (N_22488,N_21742,N_22048);
xnor U22489 (N_22489,N_21934,N_22101);
and U22490 (N_22490,N_21976,N_21678);
or U22491 (N_22491,N_21759,N_22152);
and U22492 (N_22492,N_21675,N_22073);
xnor U22493 (N_22493,N_21621,N_21981);
and U22494 (N_22494,N_22045,N_22180);
nand U22495 (N_22495,N_21954,N_22081);
or U22496 (N_22496,N_21685,N_21693);
nand U22497 (N_22497,N_21803,N_22125);
nor U22498 (N_22498,N_21998,N_22124);
xor U22499 (N_22499,N_22194,N_21701);
nor U22500 (N_22500,N_21766,N_22099);
xor U22501 (N_22501,N_21774,N_21847);
nand U22502 (N_22502,N_22169,N_21622);
nor U22503 (N_22503,N_21742,N_21897);
or U22504 (N_22504,N_21644,N_21965);
and U22505 (N_22505,N_22097,N_21829);
and U22506 (N_22506,N_22127,N_22125);
nand U22507 (N_22507,N_21813,N_21795);
or U22508 (N_22508,N_21767,N_22199);
nor U22509 (N_22509,N_21973,N_21724);
nand U22510 (N_22510,N_21957,N_21761);
nand U22511 (N_22511,N_22056,N_22025);
nand U22512 (N_22512,N_21651,N_21770);
nor U22513 (N_22513,N_22124,N_21793);
nand U22514 (N_22514,N_22157,N_21871);
nor U22515 (N_22515,N_21868,N_22068);
nor U22516 (N_22516,N_21879,N_22174);
and U22517 (N_22517,N_22176,N_22125);
nand U22518 (N_22518,N_21866,N_21638);
and U22519 (N_22519,N_21616,N_22001);
or U22520 (N_22520,N_21864,N_21706);
nand U22521 (N_22521,N_22037,N_22144);
or U22522 (N_22522,N_21662,N_21634);
xnor U22523 (N_22523,N_21765,N_22029);
nand U22524 (N_22524,N_21618,N_21819);
or U22525 (N_22525,N_21878,N_22164);
nor U22526 (N_22526,N_21930,N_21992);
nand U22527 (N_22527,N_21684,N_21857);
nand U22528 (N_22528,N_21922,N_21981);
xor U22529 (N_22529,N_21978,N_22025);
nand U22530 (N_22530,N_22052,N_22088);
nor U22531 (N_22531,N_22156,N_22134);
xnor U22532 (N_22532,N_21996,N_21768);
nand U22533 (N_22533,N_21821,N_21675);
nor U22534 (N_22534,N_22097,N_21944);
xnor U22535 (N_22535,N_21999,N_22031);
nand U22536 (N_22536,N_21655,N_21704);
nand U22537 (N_22537,N_22195,N_22001);
nand U22538 (N_22538,N_21848,N_22171);
xor U22539 (N_22539,N_21951,N_21993);
xor U22540 (N_22540,N_21767,N_22063);
nand U22541 (N_22541,N_21657,N_21609);
and U22542 (N_22542,N_22082,N_21786);
xnor U22543 (N_22543,N_21665,N_22021);
nand U22544 (N_22544,N_21613,N_21672);
xor U22545 (N_22545,N_21613,N_22120);
nand U22546 (N_22546,N_22191,N_22115);
nor U22547 (N_22547,N_21957,N_21839);
or U22548 (N_22548,N_21716,N_21834);
or U22549 (N_22549,N_21822,N_22131);
and U22550 (N_22550,N_21769,N_21662);
nor U22551 (N_22551,N_21944,N_21798);
xnor U22552 (N_22552,N_21921,N_21664);
and U22553 (N_22553,N_21671,N_22018);
nor U22554 (N_22554,N_21726,N_21770);
nor U22555 (N_22555,N_22176,N_22004);
xor U22556 (N_22556,N_22193,N_21953);
nand U22557 (N_22557,N_21950,N_22102);
xor U22558 (N_22558,N_21904,N_21816);
and U22559 (N_22559,N_21679,N_21828);
xor U22560 (N_22560,N_21881,N_21946);
nor U22561 (N_22561,N_21912,N_21600);
nand U22562 (N_22562,N_21701,N_21828);
or U22563 (N_22563,N_21625,N_21810);
nand U22564 (N_22564,N_21672,N_21956);
nor U22565 (N_22565,N_21985,N_21643);
or U22566 (N_22566,N_21990,N_21755);
nand U22567 (N_22567,N_21917,N_21699);
nand U22568 (N_22568,N_21882,N_21676);
and U22569 (N_22569,N_21964,N_21688);
nor U22570 (N_22570,N_21981,N_21609);
nor U22571 (N_22571,N_22057,N_22181);
xor U22572 (N_22572,N_21615,N_21839);
nand U22573 (N_22573,N_21840,N_22176);
xnor U22574 (N_22574,N_21649,N_21736);
nor U22575 (N_22575,N_22186,N_21820);
xnor U22576 (N_22576,N_21620,N_21684);
and U22577 (N_22577,N_21906,N_22034);
xor U22578 (N_22578,N_21768,N_21739);
nand U22579 (N_22579,N_21856,N_21850);
nand U22580 (N_22580,N_22037,N_21941);
nand U22581 (N_22581,N_21770,N_21867);
and U22582 (N_22582,N_21647,N_22199);
nor U22583 (N_22583,N_21893,N_22180);
and U22584 (N_22584,N_21863,N_21921);
xnor U22585 (N_22585,N_21872,N_21892);
xor U22586 (N_22586,N_21651,N_21769);
or U22587 (N_22587,N_22002,N_22180);
or U22588 (N_22588,N_21687,N_21776);
nand U22589 (N_22589,N_22105,N_21656);
nand U22590 (N_22590,N_22147,N_22032);
nor U22591 (N_22591,N_22109,N_21986);
and U22592 (N_22592,N_21947,N_21946);
nor U22593 (N_22593,N_22099,N_21630);
nand U22594 (N_22594,N_22057,N_22135);
xnor U22595 (N_22595,N_21762,N_21702);
or U22596 (N_22596,N_21847,N_22135);
and U22597 (N_22597,N_21724,N_22074);
nand U22598 (N_22598,N_21973,N_21606);
xor U22599 (N_22599,N_21664,N_21707);
nand U22600 (N_22600,N_22085,N_21985);
xnor U22601 (N_22601,N_21747,N_22141);
nand U22602 (N_22602,N_21753,N_21966);
and U22603 (N_22603,N_21796,N_21633);
nand U22604 (N_22604,N_21950,N_21760);
or U22605 (N_22605,N_21639,N_21679);
or U22606 (N_22606,N_21962,N_21886);
and U22607 (N_22607,N_21704,N_21971);
and U22608 (N_22608,N_22096,N_21839);
or U22609 (N_22609,N_21708,N_21884);
nor U22610 (N_22610,N_22154,N_22020);
nor U22611 (N_22611,N_21924,N_22114);
nor U22612 (N_22612,N_21885,N_21752);
xnor U22613 (N_22613,N_21716,N_22173);
nor U22614 (N_22614,N_21961,N_21707);
or U22615 (N_22615,N_22021,N_22176);
xnor U22616 (N_22616,N_22034,N_21765);
or U22617 (N_22617,N_21663,N_21951);
xnor U22618 (N_22618,N_22027,N_21780);
xor U22619 (N_22619,N_22073,N_22174);
and U22620 (N_22620,N_22196,N_21690);
nand U22621 (N_22621,N_22166,N_21883);
or U22622 (N_22622,N_21705,N_22114);
and U22623 (N_22623,N_21818,N_21875);
or U22624 (N_22624,N_22190,N_22043);
or U22625 (N_22625,N_21876,N_22138);
and U22626 (N_22626,N_21835,N_22067);
nand U22627 (N_22627,N_22015,N_22148);
or U22628 (N_22628,N_22174,N_22058);
and U22629 (N_22629,N_21780,N_21700);
or U22630 (N_22630,N_22138,N_21819);
nor U22631 (N_22631,N_22082,N_22124);
and U22632 (N_22632,N_21822,N_21645);
nor U22633 (N_22633,N_21940,N_22138);
nor U22634 (N_22634,N_21877,N_21612);
or U22635 (N_22635,N_21824,N_22004);
nand U22636 (N_22636,N_22076,N_21836);
xnor U22637 (N_22637,N_21996,N_21741);
xnor U22638 (N_22638,N_21760,N_22044);
nor U22639 (N_22639,N_22105,N_21854);
or U22640 (N_22640,N_21834,N_21699);
xnor U22641 (N_22641,N_21983,N_21663);
nor U22642 (N_22642,N_21745,N_21868);
and U22643 (N_22643,N_21798,N_21934);
xor U22644 (N_22644,N_21748,N_21659);
or U22645 (N_22645,N_21912,N_21909);
nor U22646 (N_22646,N_21854,N_21696);
and U22647 (N_22647,N_21923,N_21615);
xnor U22648 (N_22648,N_21840,N_21631);
nand U22649 (N_22649,N_21641,N_22030);
xnor U22650 (N_22650,N_21776,N_21927);
nor U22651 (N_22651,N_22192,N_21991);
or U22652 (N_22652,N_22193,N_21661);
and U22653 (N_22653,N_21929,N_21624);
or U22654 (N_22654,N_22028,N_22032);
and U22655 (N_22655,N_22080,N_21804);
xor U22656 (N_22656,N_21859,N_21884);
and U22657 (N_22657,N_22023,N_21673);
nor U22658 (N_22658,N_22133,N_21664);
xor U22659 (N_22659,N_22080,N_21630);
and U22660 (N_22660,N_21803,N_22199);
or U22661 (N_22661,N_22041,N_21779);
nor U22662 (N_22662,N_22198,N_22146);
nor U22663 (N_22663,N_22170,N_22073);
and U22664 (N_22664,N_22016,N_22001);
xor U22665 (N_22665,N_21896,N_21868);
and U22666 (N_22666,N_21812,N_21905);
nand U22667 (N_22667,N_21673,N_21763);
or U22668 (N_22668,N_21851,N_21866);
and U22669 (N_22669,N_22167,N_21644);
xor U22670 (N_22670,N_22033,N_21682);
nand U22671 (N_22671,N_21676,N_22176);
or U22672 (N_22672,N_21634,N_21887);
nand U22673 (N_22673,N_21838,N_22198);
nor U22674 (N_22674,N_21666,N_22148);
nand U22675 (N_22675,N_22091,N_21961);
and U22676 (N_22676,N_21774,N_21953);
xor U22677 (N_22677,N_21803,N_21639);
nor U22678 (N_22678,N_21690,N_21770);
xor U22679 (N_22679,N_22093,N_21706);
xor U22680 (N_22680,N_21829,N_21711);
xnor U22681 (N_22681,N_22003,N_22061);
or U22682 (N_22682,N_21709,N_21613);
or U22683 (N_22683,N_21856,N_22149);
or U22684 (N_22684,N_21756,N_21742);
nor U22685 (N_22685,N_22145,N_21896);
or U22686 (N_22686,N_21753,N_21831);
xnor U22687 (N_22687,N_22066,N_21821);
and U22688 (N_22688,N_21891,N_22070);
nand U22689 (N_22689,N_21867,N_21885);
xor U22690 (N_22690,N_22036,N_21924);
nor U22691 (N_22691,N_21884,N_21943);
and U22692 (N_22692,N_21854,N_22043);
or U22693 (N_22693,N_22080,N_21984);
nand U22694 (N_22694,N_21773,N_21748);
xor U22695 (N_22695,N_21752,N_21935);
or U22696 (N_22696,N_21781,N_21890);
xnor U22697 (N_22697,N_21711,N_22143);
xnor U22698 (N_22698,N_22192,N_22072);
xor U22699 (N_22699,N_22121,N_21941);
nand U22700 (N_22700,N_22176,N_22092);
nand U22701 (N_22701,N_22172,N_21667);
xnor U22702 (N_22702,N_21754,N_22159);
nand U22703 (N_22703,N_22005,N_21909);
or U22704 (N_22704,N_22010,N_22025);
xnor U22705 (N_22705,N_21746,N_21686);
xnor U22706 (N_22706,N_21846,N_22003);
and U22707 (N_22707,N_21807,N_21883);
xnor U22708 (N_22708,N_22184,N_21923);
or U22709 (N_22709,N_21891,N_21900);
or U22710 (N_22710,N_21662,N_21685);
or U22711 (N_22711,N_22105,N_21679);
nor U22712 (N_22712,N_21773,N_21934);
or U22713 (N_22713,N_21939,N_21813);
nand U22714 (N_22714,N_21868,N_22150);
xor U22715 (N_22715,N_22150,N_21866);
and U22716 (N_22716,N_21923,N_21896);
nor U22717 (N_22717,N_22099,N_21945);
and U22718 (N_22718,N_21887,N_21867);
nor U22719 (N_22719,N_21620,N_21973);
and U22720 (N_22720,N_21653,N_22119);
nor U22721 (N_22721,N_21975,N_22022);
nand U22722 (N_22722,N_21854,N_21698);
xnor U22723 (N_22723,N_22043,N_22123);
and U22724 (N_22724,N_22124,N_21966);
or U22725 (N_22725,N_21639,N_22047);
nand U22726 (N_22726,N_21885,N_21988);
xor U22727 (N_22727,N_21634,N_21669);
or U22728 (N_22728,N_22053,N_22028);
or U22729 (N_22729,N_21989,N_21698);
nor U22730 (N_22730,N_21771,N_21632);
xor U22731 (N_22731,N_21815,N_21915);
and U22732 (N_22732,N_21745,N_21820);
nand U22733 (N_22733,N_22022,N_21711);
or U22734 (N_22734,N_21964,N_21681);
nand U22735 (N_22735,N_21727,N_21855);
xor U22736 (N_22736,N_21675,N_22177);
nor U22737 (N_22737,N_21661,N_21685);
and U22738 (N_22738,N_22183,N_22100);
xor U22739 (N_22739,N_21752,N_22091);
or U22740 (N_22740,N_21844,N_21865);
nand U22741 (N_22741,N_22086,N_21835);
xnor U22742 (N_22742,N_22031,N_22186);
nor U22743 (N_22743,N_21755,N_21720);
and U22744 (N_22744,N_22174,N_21907);
nor U22745 (N_22745,N_21992,N_21779);
nand U22746 (N_22746,N_22084,N_22057);
xor U22747 (N_22747,N_21731,N_21695);
and U22748 (N_22748,N_21963,N_21738);
nor U22749 (N_22749,N_21850,N_22013);
or U22750 (N_22750,N_21952,N_21911);
xor U22751 (N_22751,N_22051,N_21777);
or U22752 (N_22752,N_21969,N_22100);
and U22753 (N_22753,N_21646,N_21920);
nand U22754 (N_22754,N_21616,N_21665);
nor U22755 (N_22755,N_22167,N_21934);
nand U22756 (N_22756,N_21700,N_22076);
or U22757 (N_22757,N_21868,N_21690);
and U22758 (N_22758,N_21977,N_22080);
or U22759 (N_22759,N_21677,N_22172);
nand U22760 (N_22760,N_21800,N_21942);
nand U22761 (N_22761,N_21689,N_21710);
nor U22762 (N_22762,N_21932,N_21604);
nand U22763 (N_22763,N_22104,N_21857);
and U22764 (N_22764,N_21855,N_22070);
and U22765 (N_22765,N_21938,N_22123);
xnor U22766 (N_22766,N_22138,N_22049);
xor U22767 (N_22767,N_22158,N_22144);
and U22768 (N_22768,N_21621,N_21810);
or U22769 (N_22769,N_22114,N_21850);
nand U22770 (N_22770,N_21987,N_21684);
nand U22771 (N_22771,N_22156,N_21614);
nand U22772 (N_22772,N_21839,N_21857);
nor U22773 (N_22773,N_21976,N_21763);
and U22774 (N_22774,N_21602,N_22159);
nand U22775 (N_22775,N_21787,N_21981);
nand U22776 (N_22776,N_21774,N_21872);
xor U22777 (N_22777,N_21637,N_21946);
or U22778 (N_22778,N_21880,N_21656);
xor U22779 (N_22779,N_22090,N_21802);
nor U22780 (N_22780,N_21927,N_21795);
nand U22781 (N_22781,N_22092,N_22185);
or U22782 (N_22782,N_21804,N_22038);
nor U22783 (N_22783,N_21681,N_21932);
nand U22784 (N_22784,N_21730,N_21935);
or U22785 (N_22785,N_21964,N_21905);
xnor U22786 (N_22786,N_21613,N_21918);
nor U22787 (N_22787,N_21824,N_21694);
or U22788 (N_22788,N_22062,N_21744);
nor U22789 (N_22789,N_21883,N_22062);
xnor U22790 (N_22790,N_21918,N_21989);
or U22791 (N_22791,N_22154,N_22066);
or U22792 (N_22792,N_21684,N_22081);
and U22793 (N_22793,N_22118,N_21724);
and U22794 (N_22794,N_21629,N_21971);
and U22795 (N_22795,N_22042,N_21739);
nor U22796 (N_22796,N_21840,N_22124);
nor U22797 (N_22797,N_21747,N_21732);
xor U22798 (N_22798,N_21669,N_21769);
xnor U22799 (N_22799,N_21940,N_21790);
xnor U22800 (N_22800,N_22433,N_22455);
or U22801 (N_22801,N_22325,N_22722);
xor U22802 (N_22802,N_22292,N_22390);
or U22803 (N_22803,N_22756,N_22226);
or U22804 (N_22804,N_22478,N_22426);
or U22805 (N_22805,N_22514,N_22662);
nor U22806 (N_22806,N_22754,N_22439);
xnor U22807 (N_22807,N_22472,N_22264);
xor U22808 (N_22808,N_22427,N_22412);
or U22809 (N_22809,N_22644,N_22725);
xnor U22810 (N_22810,N_22459,N_22270);
nand U22811 (N_22811,N_22527,N_22741);
nor U22812 (N_22812,N_22232,N_22288);
nor U22813 (N_22813,N_22667,N_22386);
and U22814 (N_22814,N_22685,N_22551);
and U22815 (N_22815,N_22457,N_22387);
nor U22816 (N_22816,N_22327,N_22733);
xnor U22817 (N_22817,N_22425,N_22770);
xor U22818 (N_22818,N_22613,N_22734);
or U22819 (N_22819,N_22240,N_22561);
nor U22820 (N_22820,N_22592,N_22587);
or U22821 (N_22821,N_22569,N_22661);
and U22822 (N_22822,N_22748,N_22278);
nor U22823 (N_22823,N_22300,N_22250);
or U22824 (N_22824,N_22638,N_22217);
xor U22825 (N_22825,N_22747,N_22678);
and U22826 (N_22826,N_22351,N_22394);
xor U22827 (N_22827,N_22724,N_22378);
nand U22828 (N_22828,N_22467,N_22577);
xor U22829 (N_22829,N_22711,N_22749);
xnor U22830 (N_22830,N_22333,N_22784);
nand U22831 (N_22831,N_22256,N_22323);
or U22832 (N_22832,N_22714,N_22218);
nand U22833 (N_22833,N_22437,N_22589);
nor U22834 (N_22834,N_22694,N_22380);
nand U22835 (N_22835,N_22744,N_22225);
xnor U22836 (N_22836,N_22600,N_22706);
and U22837 (N_22837,N_22778,N_22388);
or U22838 (N_22838,N_22556,N_22564);
nor U22839 (N_22839,N_22237,N_22681);
xor U22840 (N_22840,N_22374,N_22486);
and U22841 (N_22841,N_22448,N_22285);
or U22842 (N_22842,N_22214,N_22657);
xnor U22843 (N_22843,N_22316,N_22654);
xnor U22844 (N_22844,N_22652,N_22313);
xnor U22845 (N_22845,N_22261,N_22347);
nand U22846 (N_22846,N_22328,N_22690);
nor U22847 (N_22847,N_22541,N_22293);
xnor U22848 (N_22848,N_22758,N_22428);
nor U22849 (N_22849,N_22759,N_22408);
or U22850 (N_22850,N_22583,N_22373);
xnor U22851 (N_22851,N_22721,N_22717);
xor U22852 (N_22852,N_22421,N_22399);
or U22853 (N_22853,N_22696,N_22555);
or U22854 (N_22854,N_22306,N_22231);
or U22855 (N_22855,N_22496,N_22783);
nor U22856 (N_22856,N_22477,N_22247);
nand U22857 (N_22857,N_22775,N_22346);
xnor U22858 (N_22858,N_22698,N_22487);
and U22859 (N_22859,N_22660,N_22672);
or U22860 (N_22860,N_22618,N_22201);
and U22861 (N_22861,N_22671,N_22311);
xor U22862 (N_22862,N_22286,N_22326);
xnor U22863 (N_22863,N_22382,N_22463);
or U22864 (N_22864,N_22760,N_22401);
nand U22865 (N_22865,N_22720,N_22728);
or U22866 (N_22866,N_22623,N_22650);
nand U22867 (N_22867,N_22376,N_22547);
or U22868 (N_22868,N_22621,N_22359);
xor U22869 (N_22869,N_22416,N_22210);
xnor U22870 (N_22870,N_22367,N_22515);
or U22871 (N_22871,N_22682,N_22277);
and U22872 (N_22872,N_22742,N_22458);
and U22873 (N_22873,N_22490,N_22567);
or U22874 (N_22874,N_22361,N_22279);
and U22875 (N_22875,N_22389,N_22369);
nor U22876 (N_22876,N_22712,N_22764);
nand U22877 (N_22877,N_22317,N_22795);
or U22878 (N_22878,N_22637,N_22509);
or U22879 (N_22879,N_22640,N_22691);
nor U22880 (N_22880,N_22499,N_22588);
and U22881 (N_22881,N_22565,N_22796);
nand U22882 (N_22882,N_22263,N_22350);
nor U22883 (N_22883,N_22449,N_22417);
nand U22884 (N_22884,N_22655,N_22493);
or U22885 (N_22885,N_22665,N_22236);
nand U22886 (N_22886,N_22715,N_22651);
and U22887 (N_22887,N_22420,N_22597);
nand U22888 (N_22888,N_22546,N_22705);
or U22889 (N_22889,N_22702,N_22594);
xnor U22890 (N_22890,N_22701,N_22372);
nor U22891 (N_22891,N_22379,N_22465);
or U22892 (N_22892,N_22513,N_22550);
nand U22893 (N_22893,N_22686,N_22666);
nand U22894 (N_22894,N_22442,N_22745);
and U22895 (N_22895,N_22572,N_22568);
and U22896 (N_22896,N_22602,N_22614);
nand U22897 (N_22897,N_22771,N_22357);
and U22898 (N_22898,N_22700,N_22582);
and U22899 (N_22899,N_22522,N_22785);
or U22900 (N_22900,N_22731,N_22345);
or U22901 (N_22901,N_22438,N_22593);
and U22902 (N_22902,N_22675,N_22776);
or U22903 (N_22903,N_22633,N_22719);
or U22904 (N_22904,N_22708,N_22730);
and U22905 (N_22905,N_22268,N_22538);
nand U22906 (N_22906,N_22500,N_22331);
and U22907 (N_22907,N_22519,N_22689);
or U22908 (N_22908,N_22646,N_22520);
and U22909 (N_22909,N_22392,N_22343);
or U22910 (N_22910,N_22301,N_22777);
and U22911 (N_22911,N_22322,N_22607);
and U22912 (N_22912,N_22707,N_22419);
nand U22913 (N_22913,N_22510,N_22338);
nor U22914 (N_22914,N_22781,N_22406);
xnor U22915 (N_22915,N_22571,N_22391);
xor U22916 (N_22916,N_22239,N_22549);
nor U22917 (N_22917,N_22533,N_22634);
xor U22918 (N_22918,N_22273,N_22503);
or U22919 (N_22919,N_22619,N_22530);
nand U22920 (N_22920,N_22548,N_22334);
or U22921 (N_22921,N_22601,N_22352);
xor U22922 (N_22922,N_22488,N_22475);
nand U22923 (N_22923,N_22625,N_22215);
or U22924 (N_22924,N_22265,N_22304);
xor U22925 (N_22925,N_22431,N_22308);
and U22926 (N_22926,N_22570,N_22251);
nor U22927 (N_22927,N_22511,N_22337);
or U22928 (N_22928,N_22212,N_22456);
nand U22929 (N_22929,N_22255,N_22558);
nand U22930 (N_22930,N_22751,N_22245);
xnor U22931 (N_22931,N_22676,N_22553);
and U22932 (N_22932,N_22603,N_22710);
or U22933 (N_22933,N_22639,N_22750);
nor U22934 (N_22934,N_22375,N_22642);
or U22935 (N_22935,N_22544,N_22377);
or U22936 (N_22936,N_22444,N_22409);
nand U22937 (N_22937,N_22729,N_22435);
nor U22938 (N_22938,N_22483,N_22769);
nand U22939 (N_22939,N_22606,N_22418);
nand U22940 (N_22940,N_22470,N_22274);
nand U22941 (N_22941,N_22441,N_22506);
or U22942 (N_22942,N_22414,N_22363);
or U22943 (N_22943,N_22295,N_22446);
and U22944 (N_22944,N_22653,N_22318);
nand U22945 (N_22945,N_22238,N_22224);
and U22946 (N_22946,N_22739,N_22280);
xor U22947 (N_22947,N_22562,N_22407);
nor U22948 (N_22948,N_22339,N_22608);
or U22949 (N_22949,N_22221,N_22732);
and U22950 (N_22950,N_22452,N_22434);
nor U22951 (N_22951,N_22340,N_22709);
or U22952 (N_22952,N_22688,N_22257);
xnor U22953 (N_22953,N_22755,N_22680);
or U22954 (N_22954,N_22566,N_22205);
nand U22955 (N_22955,N_22529,N_22782);
xnor U22956 (N_22956,N_22223,N_22315);
or U22957 (N_22957,N_22779,N_22559);
nand U22958 (N_22958,N_22780,N_22504);
or U22959 (N_22959,N_22267,N_22489);
or U22960 (N_22960,N_22684,N_22332);
nand U22961 (N_22961,N_22494,N_22604);
nand U22962 (N_22962,N_22716,N_22299);
nand U22963 (N_22963,N_22726,N_22479);
or U22964 (N_22964,N_22788,N_22629);
nor U22965 (N_22965,N_22355,N_22248);
nor U22966 (N_22966,N_22669,N_22537);
nor U22967 (N_22967,N_22360,N_22440);
nor U22968 (N_22968,N_22584,N_22396);
nor U22969 (N_22969,N_22249,N_22517);
nand U22970 (N_22970,N_22628,N_22560);
nor U22971 (N_22971,N_22737,N_22259);
or U22972 (N_22972,N_22402,N_22356);
and U22973 (N_22973,N_22471,N_22348);
or U22974 (N_22974,N_22234,N_22424);
nand U22975 (N_22975,N_22574,N_22289);
and U22976 (N_22976,N_22746,N_22242);
nor U22977 (N_22977,N_22397,N_22206);
and U22978 (N_22978,N_22349,N_22579);
or U22979 (N_22979,N_22523,N_22241);
nand U22980 (N_22980,N_22799,N_22481);
xor U22981 (N_22981,N_22723,N_22595);
or U22982 (N_22982,N_22753,N_22491);
nor U22983 (N_22983,N_22664,N_22235);
and U22984 (N_22984,N_22297,N_22366);
xnor U22985 (N_22985,N_22791,N_22429);
nand U22986 (N_22986,N_22230,N_22736);
and U22987 (N_22987,N_22545,N_22631);
nand U22988 (N_22988,N_22395,N_22430);
xnor U22989 (N_22989,N_22518,N_22269);
and U22990 (N_22990,N_22445,N_22468);
or U22991 (N_22991,N_22580,N_22659);
nor U22992 (N_22992,N_22258,N_22599);
and U22993 (N_22993,N_22365,N_22789);
nor U22994 (N_22994,N_22704,N_22647);
nor U22995 (N_22995,N_22658,N_22581);
nor U22996 (N_22996,N_22516,N_22798);
xor U22997 (N_22997,N_22461,N_22495);
nand U22998 (N_22998,N_22735,N_22703);
nand U22999 (N_22999,N_22648,N_22786);
nand U23000 (N_23000,N_22532,N_22320);
xnor U23001 (N_23001,N_22586,N_22498);
or U23002 (N_23002,N_22632,N_22793);
nand U23003 (N_23003,N_22324,N_22370);
nand U23004 (N_23004,N_22693,N_22443);
nor U23005 (N_23005,N_22609,N_22415);
xor U23006 (N_23006,N_22563,N_22266);
nand U23007 (N_23007,N_22413,N_22229);
nand U23008 (N_23008,N_22466,N_22436);
or U23009 (N_23009,N_22670,N_22344);
nand U23010 (N_23010,N_22697,N_22319);
nor U23011 (N_23011,N_22204,N_22752);
nor U23012 (N_23012,N_22228,N_22740);
nor U23013 (N_23013,N_22610,N_22384);
or U23014 (N_23014,N_22773,N_22512);
xnor U23015 (N_23015,N_22636,N_22643);
and U23016 (N_23016,N_22573,N_22695);
or U23017 (N_23017,N_22552,N_22207);
nor U23018 (N_23018,N_22282,N_22718);
or U23019 (N_23019,N_22476,N_22526);
nand U23020 (N_23020,N_22687,N_22462);
or U23021 (N_23021,N_22284,N_22208);
or U23022 (N_23022,N_22649,N_22321);
xnor U23023 (N_23023,N_22611,N_22453);
xnor U23024 (N_23024,N_22576,N_22617);
and U23025 (N_23025,N_22227,N_22287);
nand U23026 (N_23026,N_22209,N_22738);
nand U23027 (N_23027,N_22505,N_22674);
xor U23028 (N_23028,N_22612,N_22341);
or U23029 (N_23029,N_22294,N_22244);
nor U23030 (N_23030,N_22310,N_22296);
and U23031 (N_23031,N_22787,N_22598);
nor U23032 (N_23032,N_22535,N_22626);
nor U23033 (N_23033,N_22590,N_22335);
nor U23034 (N_23034,N_22246,N_22303);
nor U23035 (N_23035,N_22216,N_22497);
or U23036 (N_23036,N_22554,N_22450);
or U23037 (N_23037,N_22305,N_22615);
nand U23038 (N_23038,N_22404,N_22772);
or U23039 (N_23039,N_22213,N_22485);
and U23040 (N_23040,N_22381,N_22400);
nor U23041 (N_23041,N_22200,N_22307);
xnor U23042 (N_23042,N_22507,N_22358);
nand U23043 (N_23043,N_22743,N_22302);
or U23044 (N_23044,N_22578,N_22219);
or U23045 (N_23045,N_22540,N_22330);
nor U23046 (N_23046,N_22620,N_22591);
or U23047 (N_23047,N_22474,N_22627);
and U23048 (N_23048,N_22243,N_22596);
or U23049 (N_23049,N_22482,N_22525);
and U23050 (N_23050,N_22790,N_22679);
or U23051 (N_23051,N_22403,N_22543);
nand U23052 (N_23052,N_22534,N_22766);
and U23053 (N_23053,N_22797,N_22276);
or U23054 (N_23054,N_22309,N_22368);
and U23055 (N_23055,N_22524,N_22492);
or U23056 (N_23056,N_22423,N_22656);
and U23057 (N_23057,N_22262,N_22254);
xnor U23058 (N_23058,N_22762,N_22281);
nor U23059 (N_23059,N_22641,N_22410);
and U23060 (N_23060,N_22792,N_22645);
or U23061 (N_23061,N_22398,N_22447);
or U23062 (N_23062,N_22575,N_22767);
nor U23063 (N_23063,N_22393,N_22616);
or U23064 (N_23064,N_22405,N_22291);
and U23065 (N_23065,N_22342,N_22312);
or U23066 (N_23066,N_22761,N_22354);
nor U23067 (N_23067,N_22364,N_22683);
xor U23068 (N_23068,N_22692,N_22464);
nor U23069 (N_23069,N_22314,N_22329);
nor U23070 (N_23070,N_22727,N_22774);
nand U23071 (N_23071,N_22202,N_22668);
nor U23072 (N_23072,N_22271,N_22283);
and U23073 (N_23073,N_22203,N_22422);
nand U23074 (N_23074,N_22765,N_22480);
nor U23075 (N_23075,N_22605,N_22794);
or U23076 (N_23076,N_22635,N_22411);
nor U23077 (N_23077,N_22539,N_22371);
nand U23078 (N_23078,N_22211,N_22275);
xnor U23079 (N_23079,N_22298,N_22385);
or U23080 (N_23080,N_22451,N_22233);
xor U23081 (N_23081,N_22624,N_22460);
nor U23082 (N_23082,N_22673,N_22622);
or U23083 (N_23083,N_22336,N_22531);
and U23084 (N_23084,N_22272,N_22757);
xor U23085 (N_23085,N_22528,N_22502);
and U23086 (N_23086,N_22473,N_22699);
nor U23087 (N_23087,N_22454,N_22469);
and U23088 (N_23088,N_22557,N_22663);
xor U23089 (N_23089,N_22220,N_22290);
or U23090 (N_23090,N_22542,N_22383);
xnor U23091 (N_23091,N_22713,N_22484);
nand U23092 (N_23092,N_22521,N_22585);
nand U23093 (N_23093,N_22768,N_22252);
nand U23094 (N_23094,N_22501,N_22508);
nand U23095 (N_23095,N_22260,N_22362);
nand U23096 (N_23096,N_22536,N_22253);
or U23097 (N_23097,N_22432,N_22630);
nand U23098 (N_23098,N_22353,N_22222);
nor U23099 (N_23099,N_22763,N_22677);
and U23100 (N_23100,N_22555,N_22288);
nor U23101 (N_23101,N_22635,N_22485);
and U23102 (N_23102,N_22698,N_22497);
or U23103 (N_23103,N_22554,N_22454);
xnor U23104 (N_23104,N_22248,N_22764);
xor U23105 (N_23105,N_22285,N_22268);
xor U23106 (N_23106,N_22569,N_22268);
or U23107 (N_23107,N_22218,N_22725);
nor U23108 (N_23108,N_22737,N_22509);
nand U23109 (N_23109,N_22268,N_22383);
and U23110 (N_23110,N_22268,N_22322);
nor U23111 (N_23111,N_22637,N_22599);
or U23112 (N_23112,N_22402,N_22697);
xnor U23113 (N_23113,N_22691,N_22718);
xor U23114 (N_23114,N_22333,N_22646);
or U23115 (N_23115,N_22420,N_22232);
and U23116 (N_23116,N_22354,N_22353);
xor U23117 (N_23117,N_22249,N_22732);
and U23118 (N_23118,N_22459,N_22299);
nor U23119 (N_23119,N_22560,N_22349);
or U23120 (N_23120,N_22325,N_22459);
and U23121 (N_23121,N_22626,N_22532);
or U23122 (N_23122,N_22310,N_22533);
and U23123 (N_23123,N_22233,N_22717);
or U23124 (N_23124,N_22517,N_22450);
xor U23125 (N_23125,N_22677,N_22476);
nand U23126 (N_23126,N_22486,N_22351);
or U23127 (N_23127,N_22421,N_22213);
nand U23128 (N_23128,N_22429,N_22263);
xnor U23129 (N_23129,N_22375,N_22393);
and U23130 (N_23130,N_22655,N_22394);
nor U23131 (N_23131,N_22261,N_22233);
and U23132 (N_23132,N_22310,N_22761);
nor U23133 (N_23133,N_22672,N_22493);
and U23134 (N_23134,N_22611,N_22579);
and U23135 (N_23135,N_22462,N_22465);
and U23136 (N_23136,N_22229,N_22331);
or U23137 (N_23137,N_22291,N_22223);
xor U23138 (N_23138,N_22335,N_22707);
xnor U23139 (N_23139,N_22297,N_22721);
and U23140 (N_23140,N_22426,N_22706);
xor U23141 (N_23141,N_22297,N_22378);
or U23142 (N_23142,N_22385,N_22637);
nand U23143 (N_23143,N_22383,N_22435);
or U23144 (N_23144,N_22257,N_22674);
nand U23145 (N_23145,N_22386,N_22269);
and U23146 (N_23146,N_22681,N_22459);
or U23147 (N_23147,N_22290,N_22249);
nand U23148 (N_23148,N_22398,N_22710);
or U23149 (N_23149,N_22759,N_22299);
nand U23150 (N_23150,N_22317,N_22566);
nor U23151 (N_23151,N_22507,N_22458);
nand U23152 (N_23152,N_22509,N_22289);
or U23153 (N_23153,N_22455,N_22414);
nor U23154 (N_23154,N_22750,N_22232);
or U23155 (N_23155,N_22309,N_22695);
nand U23156 (N_23156,N_22312,N_22460);
or U23157 (N_23157,N_22431,N_22718);
nand U23158 (N_23158,N_22312,N_22562);
nor U23159 (N_23159,N_22569,N_22604);
nand U23160 (N_23160,N_22549,N_22451);
xor U23161 (N_23161,N_22458,N_22731);
or U23162 (N_23162,N_22653,N_22266);
nor U23163 (N_23163,N_22321,N_22590);
nand U23164 (N_23164,N_22661,N_22746);
nor U23165 (N_23165,N_22338,N_22669);
nand U23166 (N_23166,N_22278,N_22253);
or U23167 (N_23167,N_22382,N_22776);
nor U23168 (N_23168,N_22603,N_22615);
and U23169 (N_23169,N_22640,N_22749);
xnor U23170 (N_23170,N_22479,N_22296);
xor U23171 (N_23171,N_22577,N_22666);
xnor U23172 (N_23172,N_22635,N_22341);
nor U23173 (N_23173,N_22574,N_22327);
and U23174 (N_23174,N_22624,N_22622);
or U23175 (N_23175,N_22784,N_22717);
or U23176 (N_23176,N_22614,N_22522);
xnor U23177 (N_23177,N_22289,N_22611);
nor U23178 (N_23178,N_22605,N_22214);
nor U23179 (N_23179,N_22713,N_22572);
nor U23180 (N_23180,N_22577,N_22558);
xor U23181 (N_23181,N_22700,N_22697);
xnor U23182 (N_23182,N_22325,N_22397);
or U23183 (N_23183,N_22428,N_22587);
nor U23184 (N_23184,N_22384,N_22266);
nor U23185 (N_23185,N_22552,N_22250);
and U23186 (N_23186,N_22280,N_22388);
xnor U23187 (N_23187,N_22333,N_22501);
xnor U23188 (N_23188,N_22205,N_22335);
xor U23189 (N_23189,N_22669,N_22257);
or U23190 (N_23190,N_22461,N_22496);
and U23191 (N_23191,N_22240,N_22479);
nor U23192 (N_23192,N_22563,N_22726);
nor U23193 (N_23193,N_22316,N_22381);
nand U23194 (N_23194,N_22613,N_22641);
or U23195 (N_23195,N_22597,N_22487);
xor U23196 (N_23196,N_22468,N_22643);
nand U23197 (N_23197,N_22789,N_22619);
and U23198 (N_23198,N_22566,N_22336);
nand U23199 (N_23199,N_22229,N_22785);
xnor U23200 (N_23200,N_22441,N_22261);
or U23201 (N_23201,N_22462,N_22719);
and U23202 (N_23202,N_22743,N_22636);
nor U23203 (N_23203,N_22383,N_22424);
nor U23204 (N_23204,N_22510,N_22675);
xnor U23205 (N_23205,N_22596,N_22616);
nor U23206 (N_23206,N_22278,N_22641);
and U23207 (N_23207,N_22355,N_22445);
nor U23208 (N_23208,N_22465,N_22531);
xnor U23209 (N_23209,N_22525,N_22766);
xnor U23210 (N_23210,N_22526,N_22355);
or U23211 (N_23211,N_22623,N_22697);
xnor U23212 (N_23212,N_22419,N_22251);
xor U23213 (N_23213,N_22388,N_22446);
and U23214 (N_23214,N_22235,N_22395);
nand U23215 (N_23215,N_22439,N_22509);
nand U23216 (N_23216,N_22327,N_22296);
nand U23217 (N_23217,N_22294,N_22641);
nor U23218 (N_23218,N_22602,N_22374);
xor U23219 (N_23219,N_22581,N_22797);
nand U23220 (N_23220,N_22625,N_22282);
and U23221 (N_23221,N_22609,N_22326);
xor U23222 (N_23222,N_22583,N_22707);
xnor U23223 (N_23223,N_22653,N_22764);
nand U23224 (N_23224,N_22326,N_22365);
or U23225 (N_23225,N_22564,N_22416);
xor U23226 (N_23226,N_22467,N_22707);
xor U23227 (N_23227,N_22442,N_22593);
xnor U23228 (N_23228,N_22711,N_22241);
nand U23229 (N_23229,N_22211,N_22787);
xnor U23230 (N_23230,N_22240,N_22544);
nand U23231 (N_23231,N_22275,N_22593);
and U23232 (N_23232,N_22512,N_22589);
xnor U23233 (N_23233,N_22447,N_22248);
nor U23234 (N_23234,N_22530,N_22763);
nand U23235 (N_23235,N_22394,N_22320);
or U23236 (N_23236,N_22391,N_22626);
and U23237 (N_23237,N_22737,N_22733);
and U23238 (N_23238,N_22245,N_22769);
xnor U23239 (N_23239,N_22370,N_22427);
and U23240 (N_23240,N_22736,N_22318);
and U23241 (N_23241,N_22334,N_22514);
and U23242 (N_23242,N_22444,N_22442);
nand U23243 (N_23243,N_22335,N_22408);
xor U23244 (N_23244,N_22389,N_22356);
nand U23245 (N_23245,N_22592,N_22289);
nor U23246 (N_23246,N_22562,N_22368);
xnor U23247 (N_23247,N_22445,N_22769);
and U23248 (N_23248,N_22429,N_22430);
xor U23249 (N_23249,N_22428,N_22423);
xor U23250 (N_23250,N_22516,N_22768);
nand U23251 (N_23251,N_22458,N_22669);
or U23252 (N_23252,N_22675,N_22757);
and U23253 (N_23253,N_22362,N_22361);
xnor U23254 (N_23254,N_22567,N_22493);
xnor U23255 (N_23255,N_22459,N_22286);
xnor U23256 (N_23256,N_22608,N_22466);
nor U23257 (N_23257,N_22733,N_22744);
nor U23258 (N_23258,N_22517,N_22482);
or U23259 (N_23259,N_22795,N_22694);
or U23260 (N_23260,N_22369,N_22224);
or U23261 (N_23261,N_22641,N_22472);
or U23262 (N_23262,N_22360,N_22457);
or U23263 (N_23263,N_22227,N_22450);
nand U23264 (N_23264,N_22736,N_22237);
nand U23265 (N_23265,N_22486,N_22660);
or U23266 (N_23266,N_22302,N_22608);
or U23267 (N_23267,N_22349,N_22287);
nand U23268 (N_23268,N_22269,N_22625);
xor U23269 (N_23269,N_22481,N_22732);
nor U23270 (N_23270,N_22451,N_22359);
and U23271 (N_23271,N_22283,N_22504);
xnor U23272 (N_23272,N_22254,N_22782);
and U23273 (N_23273,N_22535,N_22389);
nor U23274 (N_23274,N_22381,N_22235);
nor U23275 (N_23275,N_22653,N_22400);
nor U23276 (N_23276,N_22779,N_22473);
nor U23277 (N_23277,N_22503,N_22716);
xnor U23278 (N_23278,N_22798,N_22342);
or U23279 (N_23279,N_22275,N_22675);
and U23280 (N_23280,N_22258,N_22524);
xnor U23281 (N_23281,N_22451,N_22544);
nor U23282 (N_23282,N_22654,N_22441);
nor U23283 (N_23283,N_22408,N_22359);
and U23284 (N_23284,N_22618,N_22407);
and U23285 (N_23285,N_22366,N_22541);
or U23286 (N_23286,N_22430,N_22547);
or U23287 (N_23287,N_22631,N_22383);
nor U23288 (N_23288,N_22307,N_22693);
xor U23289 (N_23289,N_22397,N_22395);
nand U23290 (N_23290,N_22387,N_22506);
or U23291 (N_23291,N_22691,N_22334);
nor U23292 (N_23292,N_22602,N_22514);
or U23293 (N_23293,N_22464,N_22459);
and U23294 (N_23294,N_22377,N_22382);
xor U23295 (N_23295,N_22363,N_22264);
nand U23296 (N_23296,N_22391,N_22206);
nor U23297 (N_23297,N_22736,N_22324);
nor U23298 (N_23298,N_22525,N_22279);
nor U23299 (N_23299,N_22475,N_22711);
xnor U23300 (N_23300,N_22557,N_22300);
and U23301 (N_23301,N_22765,N_22764);
and U23302 (N_23302,N_22394,N_22762);
nor U23303 (N_23303,N_22656,N_22316);
nand U23304 (N_23304,N_22234,N_22381);
nor U23305 (N_23305,N_22353,N_22266);
xnor U23306 (N_23306,N_22380,N_22718);
nand U23307 (N_23307,N_22764,N_22224);
nand U23308 (N_23308,N_22260,N_22438);
and U23309 (N_23309,N_22582,N_22397);
xor U23310 (N_23310,N_22322,N_22685);
xnor U23311 (N_23311,N_22786,N_22667);
and U23312 (N_23312,N_22225,N_22524);
xor U23313 (N_23313,N_22527,N_22605);
or U23314 (N_23314,N_22307,N_22388);
nor U23315 (N_23315,N_22253,N_22733);
and U23316 (N_23316,N_22479,N_22454);
xnor U23317 (N_23317,N_22527,N_22759);
nand U23318 (N_23318,N_22545,N_22349);
nor U23319 (N_23319,N_22407,N_22233);
xor U23320 (N_23320,N_22424,N_22468);
and U23321 (N_23321,N_22579,N_22769);
or U23322 (N_23322,N_22469,N_22472);
and U23323 (N_23323,N_22643,N_22269);
nor U23324 (N_23324,N_22209,N_22489);
nor U23325 (N_23325,N_22471,N_22410);
nor U23326 (N_23326,N_22585,N_22663);
nand U23327 (N_23327,N_22599,N_22591);
and U23328 (N_23328,N_22296,N_22307);
or U23329 (N_23329,N_22665,N_22734);
xor U23330 (N_23330,N_22546,N_22590);
or U23331 (N_23331,N_22559,N_22299);
xor U23332 (N_23332,N_22641,N_22764);
or U23333 (N_23333,N_22377,N_22361);
or U23334 (N_23334,N_22604,N_22656);
nor U23335 (N_23335,N_22447,N_22623);
xnor U23336 (N_23336,N_22495,N_22594);
nor U23337 (N_23337,N_22203,N_22443);
or U23338 (N_23338,N_22612,N_22212);
and U23339 (N_23339,N_22446,N_22606);
or U23340 (N_23340,N_22688,N_22584);
nand U23341 (N_23341,N_22521,N_22318);
nand U23342 (N_23342,N_22702,N_22274);
xor U23343 (N_23343,N_22608,N_22796);
or U23344 (N_23344,N_22526,N_22752);
or U23345 (N_23345,N_22594,N_22682);
and U23346 (N_23346,N_22316,N_22683);
xnor U23347 (N_23347,N_22422,N_22760);
or U23348 (N_23348,N_22369,N_22548);
xnor U23349 (N_23349,N_22312,N_22202);
xnor U23350 (N_23350,N_22258,N_22321);
xor U23351 (N_23351,N_22202,N_22437);
xnor U23352 (N_23352,N_22723,N_22630);
or U23353 (N_23353,N_22723,N_22694);
or U23354 (N_23354,N_22229,N_22641);
nand U23355 (N_23355,N_22646,N_22594);
nor U23356 (N_23356,N_22333,N_22582);
xnor U23357 (N_23357,N_22490,N_22411);
xor U23358 (N_23358,N_22347,N_22793);
xor U23359 (N_23359,N_22522,N_22314);
and U23360 (N_23360,N_22428,N_22535);
nand U23361 (N_23361,N_22602,N_22558);
nor U23362 (N_23362,N_22272,N_22771);
nand U23363 (N_23363,N_22399,N_22747);
or U23364 (N_23364,N_22729,N_22376);
or U23365 (N_23365,N_22318,N_22334);
xor U23366 (N_23366,N_22282,N_22300);
nor U23367 (N_23367,N_22687,N_22595);
xor U23368 (N_23368,N_22240,N_22208);
and U23369 (N_23369,N_22258,N_22739);
nand U23370 (N_23370,N_22661,N_22778);
or U23371 (N_23371,N_22434,N_22343);
nand U23372 (N_23372,N_22491,N_22496);
or U23373 (N_23373,N_22297,N_22372);
nor U23374 (N_23374,N_22347,N_22269);
or U23375 (N_23375,N_22439,N_22575);
nor U23376 (N_23376,N_22423,N_22450);
xor U23377 (N_23377,N_22525,N_22578);
and U23378 (N_23378,N_22529,N_22255);
nand U23379 (N_23379,N_22507,N_22273);
nand U23380 (N_23380,N_22441,N_22269);
nand U23381 (N_23381,N_22530,N_22731);
nand U23382 (N_23382,N_22727,N_22514);
or U23383 (N_23383,N_22556,N_22689);
or U23384 (N_23384,N_22715,N_22382);
nor U23385 (N_23385,N_22630,N_22329);
and U23386 (N_23386,N_22360,N_22537);
nor U23387 (N_23387,N_22702,N_22351);
or U23388 (N_23388,N_22491,N_22561);
nand U23389 (N_23389,N_22685,N_22385);
nand U23390 (N_23390,N_22688,N_22633);
or U23391 (N_23391,N_22233,N_22577);
or U23392 (N_23392,N_22567,N_22395);
and U23393 (N_23393,N_22312,N_22626);
nand U23394 (N_23394,N_22248,N_22512);
nand U23395 (N_23395,N_22280,N_22585);
or U23396 (N_23396,N_22597,N_22274);
and U23397 (N_23397,N_22353,N_22449);
and U23398 (N_23398,N_22562,N_22425);
or U23399 (N_23399,N_22497,N_22411);
nor U23400 (N_23400,N_23332,N_23140);
or U23401 (N_23401,N_22985,N_23183);
nand U23402 (N_23402,N_22931,N_23367);
xnor U23403 (N_23403,N_22924,N_23311);
nand U23404 (N_23404,N_23250,N_23156);
or U23405 (N_23405,N_23347,N_23087);
or U23406 (N_23406,N_23081,N_22903);
or U23407 (N_23407,N_23319,N_23068);
nand U23408 (N_23408,N_23126,N_22982);
nand U23409 (N_23409,N_22919,N_22997);
nand U23410 (N_23410,N_22943,N_23276);
nand U23411 (N_23411,N_23294,N_23322);
xnor U23412 (N_23412,N_23037,N_23162);
nor U23413 (N_23413,N_23038,N_23091);
xor U23414 (N_23414,N_22901,N_23242);
nand U23415 (N_23415,N_22980,N_23122);
nand U23416 (N_23416,N_22959,N_23317);
nor U23417 (N_23417,N_23172,N_23358);
and U23418 (N_23418,N_23348,N_23269);
and U23419 (N_23419,N_23168,N_22979);
nor U23420 (N_23420,N_23115,N_23053);
xnor U23421 (N_23421,N_22887,N_23079);
and U23422 (N_23422,N_23147,N_23229);
nand U23423 (N_23423,N_23137,N_23143);
and U23424 (N_23424,N_23362,N_22905);
xor U23425 (N_23425,N_22821,N_23372);
or U23426 (N_23426,N_22845,N_23336);
nand U23427 (N_23427,N_23135,N_22954);
nand U23428 (N_23428,N_23000,N_22899);
nand U23429 (N_23429,N_23393,N_23164);
and U23430 (N_23430,N_23234,N_23200);
or U23431 (N_23431,N_22806,N_22925);
xnor U23432 (N_23432,N_23128,N_22850);
nor U23433 (N_23433,N_23369,N_23099);
xor U23434 (N_23434,N_22998,N_23342);
xnor U23435 (N_23435,N_22842,N_23152);
or U23436 (N_23436,N_23290,N_22862);
nor U23437 (N_23437,N_23257,N_23016);
or U23438 (N_23438,N_23142,N_23330);
nand U23439 (N_23439,N_22993,N_23092);
nor U23440 (N_23440,N_22817,N_23205);
nor U23441 (N_23441,N_23343,N_23378);
nand U23442 (N_23442,N_23195,N_23356);
xor U23443 (N_23443,N_23299,N_23289);
and U23444 (N_23444,N_22824,N_23161);
xor U23445 (N_23445,N_23111,N_23063);
nand U23446 (N_23446,N_23320,N_22836);
nand U23447 (N_23447,N_22804,N_23387);
nor U23448 (N_23448,N_22946,N_22975);
and U23449 (N_23449,N_23208,N_23117);
nor U23450 (N_23450,N_22964,N_22840);
and U23451 (N_23451,N_22861,N_23007);
nand U23452 (N_23452,N_23240,N_23009);
and U23453 (N_23453,N_23003,N_22874);
or U23454 (N_23454,N_23024,N_22889);
and U23455 (N_23455,N_22971,N_23192);
nor U23456 (N_23456,N_23145,N_22927);
xor U23457 (N_23457,N_23020,N_23374);
xnor U23458 (N_23458,N_23293,N_22801);
xor U23459 (N_23459,N_23207,N_23069);
nand U23460 (N_23460,N_22855,N_23057);
nor U23461 (N_23461,N_22955,N_23101);
and U23462 (N_23462,N_22894,N_23224);
and U23463 (N_23463,N_22870,N_23325);
and U23464 (N_23464,N_22911,N_23329);
and U23465 (N_23465,N_23338,N_22922);
nor U23466 (N_23466,N_22920,N_23231);
and U23467 (N_23467,N_23216,N_23246);
and U23468 (N_23468,N_22841,N_22973);
nor U23469 (N_23469,N_23389,N_23061);
or U23470 (N_23470,N_23353,N_22953);
nand U23471 (N_23471,N_22968,N_23165);
or U23472 (N_23472,N_23095,N_22983);
or U23473 (N_23473,N_23002,N_23153);
and U23474 (N_23474,N_23112,N_23113);
nor U23475 (N_23475,N_23260,N_22984);
nor U23476 (N_23476,N_23073,N_23071);
nor U23477 (N_23477,N_23151,N_22871);
or U23478 (N_23478,N_22858,N_23194);
and U23479 (N_23479,N_22978,N_23265);
or U23480 (N_23480,N_23340,N_23108);
nor U23481 (N_23481,N_23005,N_23059);
or U23482 (N_23482,N_23187,N_23222);
xnor U23483 (N_23483,N_23304,N_23093);
or U23484 (N_23484,N_22947,N_23077);
nor U23485 (N_23485,N_23188,N_23076);
xnor U23486 (N_23486,N_22992,N_23055);
nor U23487 (N_23487,N_23104,N_23345);
xor U23488 (N_23488,N_23282,N_22849);
nor U23489 (N_23489,N_23217,N_23014);
and U23490 (N_23490,N_23110,N_22988);
or U23491 (N_23491,N_23255,N_22825);
or U23492 (N_23492,N_23316,N_23237);
nand U23493 (N_23493,N_23243,N_23043);
xor U23494 (N_23494,N_22891,N_23158);
nor U23495 (N_23495,N_23377,N_22933);
and U23496 (N_23496,N_23106,N_23127);
nor U23497 (N_23497,N_22950,N_23021);
nor U23498 (N_23498,N_22910,N_23365);
and U23499 (N_23499,N_23333,N_23350);
xor U23500 (N_23500,N_23254,N_22819);
or U23501 (N_23501,N_23303,N_22852);
nor U23502 (N_23502,N_23180,N_23198);
xnor U23503 (N_23503,N_23241,N_22923);
or U23504 (N_23504,N_23213,N_22869);
xor U23505 (N_23505,N_23399,N_23261);
nor U23506 (N_23506,N_23373,N_23041);
and U23507 (N_23507,N_22865,N_22989);
nand U23508 (N_23508,N_23049,N_22814);
and U23509 (N_23509,N_23176,N_22827);
nor U23510 (N_23510,N_22913,N_23100);
or U23511 (N_23511,N_23228,N_22876);
nand U23512 (N_23512,N_23349,N_23048);
nor U23513 (N_23513,N_22990,N_22812);
nor U23514 (N_23514,N_22914,N_22890);
xor U23515 (N_23515,N_22936,N_22906);
nor U23516 (N_23516,N_22999,N_22823);
and U23517 (N_23517,N_22873,N_23086);
nor U23518 (N_23518,N_23235,N_23191);
or U23519 (N_23519,N_23163,N_23313);
and U23520 (N_23520,N_23083,N_23141);
xnor U23521 (N_23521,N_22864,N_23326);
nor U23522 (N_23522,N_23244,N_23097);
xnor U23523 (N_23523,N_23042,N_23075);
nor U23524 (N_23524,N_23285,N_23098);
nand U23525 (N_23525,N_22863,N_23144);
xnor U23526 (N_23526,N_23186,N_22826);
nor U23527 (N_23527,N_22972,N_23036);
and U23528 (N_23528,N_23114,N_22857);
nand U23529 (N_23529,N_23088,N_23050);
nand U23530 (N_23530,N_22929,N_23392);
nand U23531 (N_23531,N_23232,N_23105);
or U23532 (N_23532,N_23305,N_23226);
and U23533 (N_23533,N_23096,N_22844);
or U23534 (N_23534,N_22810,N_22854);
xnor U23535 (N_23535,N_22856,N_23258);
nand U23536 (N_23536,N_23175,N_22888);
xor U23537 (N_23537,N_23150,N_22877);
and U23538 (N_23538,N_23357,N_22860);
xnor U23539 (N_23539,N_23125,N_23376);
and U23540 (N_23540,N_23171,N_22872);
nand U23541 (N_23541,N_22867,N_22941);
and U23542 (N_23542,N_23394,N_23028);
nand U23543 (N_23543,N_23017,N_23045);
or U23544 (N_23544,N_22951,N_23090);
nand U23545 (N_23545,N_23359,N_22944);
nand U23546 (N_23546,N_23056,N_22886);
xnor U23547 (N_23547,N_23287,N_22960);
nor U23548 (N_23548,N_23245,N_23291);
xnor U23549 (N_23549,N_23341,N_23065);
xnor U23550 (N_23550,N_22909,N_23263);
or U23551 (N_23551,N_22962,N_23102);
or U23552 (N_23552,N_23133,N_23278);
nor U23553 (N_23553,N_23344,N_23174);
and U23554 (N_23554,N_22918,N_23302);
nor U23555 (N_23555,N_23157,N_23268);
nor U23556 (N_23556,N_23170,N_23085);
nand U23557 (N_23557,N_22987,N_23084);
nor U23558 (N_23558,N_22974,N_23351);
nand U23559 (N_23559,N_23391,N_23366);
or U23560 (N_23560,N_23027,N_22948);
and U23561 (N_23561,N_22934,N_23247);
and U23562 (N_23562,N_23146,N_23080);
xnor U23563 (N_23563,N_23310,N_22938);
xnor U23564 (N_23564,N_22896,N_22847);
or U23565 (N_23565,N_22994,N_22900);
nand U23566 (N_23566,N_22868,N_23361);
xor U23567 (N_23567,N_23190,N_23306);
nand U23568 (N_23568,N_23339,N_23390);
xnor U23569 (N_23569,N_22834,N_22815);
xor U23570 (N_23570,N_23398,N_22986);
nand U23571 (N_23571,N_22970,N_23018);
xor U23572 (N_23572,N_22880,N_23199);
and U23573 (N_23573,N_22831,N_23368);
nor U23574 (N_23574,N_23236,N_23030);
nor U23575 (N_23575,N_23355,N_22800);
nand U23576 (N_23576,N_23215,N_22928);
nor U23577 (N_23577,N_23248,N_23169);
or U23578 (N_23578,N_22912,N_22915);
and U23579 (N_23579,N_23138,N_23107);
nor U23580 (N_23580,N_23252,N_22939);
or U23581 (N_23581,N_23301,N_23040);
xnor U23582 (N_23582,N_23166,N_23010);
and U23583 (N_23583,N_23277,N_23202);
nor U23584 (N_23584,N_23283,N_23382);
nand U23585 (N_23585,N_23315,N_23292);
nor U23586 (N_23586,N_23067,N_23379);
or U23587 (N_23587,N_23214,N_22843);
or U23588 (N_23588,N_22884,N_23173);
xnor U23589 (N_23589,N_23380,N_23318);
or U23590 (N_23590,N_23121,N_22803);
xnor U23591 (N_23591,N_23267,N_23223);
or U23592 (N_23592,N_23033,N_23381);
or U23593 (N_23593,N_23388,N_22963);
or U23594 (N_23594,N_23060,N_23286);
nor U23595 (N_23595,N_23279,N_22976);
xor U23596 (N_23596,N_22822,N_23072);
nand U23597 (N_23597,N_23044,N_22904);
nand U23598 (N_23598,N_22932,N_23274);
xnor U23599 (N_23599,N_23204,N_23203);
or U23600 (N_23600,N_23004,N_22908);
nor U23601 (N_23601,N_23062,N_22885);
nand U23602 (N_23602,N_23066,N_23239);
nand U23603 (N_23603,N_22882,N_23177);
xor U23604 (N_23604,N_23120,N_23078);
xor U23605 (N_23605,N_23262,N_22921);
nor U23606 (N_23606,N_23070,N_22935);
and U23607 (N_23607,N_22813,N_22811);
nor U23608 (N_23608,N_23312,N_23307);
or U23609 (N_23609,N_23346,N_22866);
or U23610 (N_23610,N_22859,N_22961);
and U23611 (N_23611,N_23026,N_23058);
or U23612 (N_23612,N_22995,N_23227);
and U23613 (N_23613,N_23012,N_23185);
nor U23614 (N_23614,N_22828,N_23370);
nor U23615 (N_23615,N_22878,N_22875);
xnor U23616 (N_23616,N_23280,N_22881);
xnor U23617 (N_23617,N_23211,N_23284);
or U23618 (N_23618,N_23022,N_23238);
and U23619 (N_23619,N_23259,N_23360);
nand U23620 (N_23620,N_23189,N_22952);
nand U23621 (N_23621,N_22820,N_23103);
or U23622 (N_23622,N_22892,N_23335);
or U23623 (N_23623,N_22956,N_23013);
nor U23624 (N_23624,N_22851,N_22846);
nand U23625 (N_23625,N_23251,N_23034);
and U23626 (N_23626,N_22916,N_23288);
nand U23627 (N_23627,N_22830,N_23015);
nand U23628 (N_23628,N_23155,N_23118);
xnor U23629 (N_23629,N_23201,N_23383);
nor U23630 (N_23630,N_23298,N_23212);
nor U23631 (N_23631,N_23025,N_23300);
xnor U23632 (N_23632,N_23193,N_23148);
and U23633 (N_23633,N_23295,N_22833);
nand U23634 (N_23634,N_23160,N_23130);
xor U23635 (N_23635,N_23396,N_23132);
nor U23636 (N_23636,N_22966,N_23220);
nor U23637 (N_23637,N_23337,N_23327);
xnor U23638 (N_23638,N_23039,N_23124);
nand U23639 (N_23639,N_22942,N_22805);
nor U23640 (N_23640,N_23046,N_23385);
nand U23641 (N_23641,N_23272,N_22839);
nor U23642 (N_23642,N_22895,N_23264);
and U23643 (N_23643,N_22981,N_23011);
xnor U23644 (N_23644,N_22829,N_23363);
or U23645 (N_23645,N_23321,N_23273);
and U23646 (N_23646,N_23197,N_22996);
nor U23647 (N_23647,N_23397,N_23064);
xor U23648 (N_23648,N_22917,N_22807);
xnor U23649 (N_23649,N_23219,N_23116);
nand U23650 (N_23650,N_23082,N_23136);
nor U23651 (N_23651,N_23386,N_23123);
xor U23652 (N_23652,N_23308,N_23328);
nand U23653 (N_23653,N_23221,N_23249);
xor U23654 (N_23654,N_22965,N_23266);
and U23655 (N_23655,N_23109,N_23323);
and U23656 (N_23656,N_23129,N_23051);
or U23657 (N_23657,N_22848,N_23314);
or U23658 (N_23658,N_23352,N_22879);
or U23659 (N_23659,N_22907,N_23233);
or U23660 (N_23660,N_22838,N_23031);
nand U23661 (N_23661,N_23364,N_23006);
nor U23662 (N_23662,N_23275,N_23296);
nor U23663 (N_23663,N_23154,N_22853);
or U23664 (N_23664,N_23270,N_22832);
xnor U23665 (N_23665,N_22958,N_23309);
xnor U23666 (N_23666,N_22883,N_23253);
nor U23667 (N_23667,N_22940,N_23054);
and U23668 (N_23668,N_23375,N_23371);
nor U23669 (N_23669,N_23139,N_23395);
xnor U23670 (N_23670,N_22802,N_23271);
nor U23671 (N_23671,N_23008,N_22898);
xnor U23672 (N_23672,N_22816,N_23032);
nor U23673 (N_23673,N_23023,N_22991);
xnor U23674 (N_23674,N_23331,N_23354);
or U23675 (N_23675,N_23019,N_22893);
and U23676 (N_23676,N_23167,N_23256);
and U23677 (N_23677,N_23119,N_23196);
xor U23678 (N_23678,N_22977,N_22902);
or U23679 (N_23679,N_23179,N_23230);
and U23680 (N_23680,N_22957,N_23218);
nand U23681 (N_23681,N_22926,N_23074);
or U23682 (N_23682,N_23384,N_22837);
nand U23683 (N_23683,N_22967,N_23149);
nand U23684 (N_23684,N_22945,N_23035);
or U23685 (N_23685,N_23184,N_22949);
nor U23686 (N_23686,N_22809,N_22818);
nor U23687 (N_23687,N_23001,N_22835);
and U23688 (N_23688,N_23225,N_23281);
or U23689 (N_23689,N_23209,N_22808);
nand U23690 (N_23690,N_23029,N_22930);
xor U23691 (N_23691,N_23297,N_23178);
nand U23692 (N_23692,N_23324,N_22897);
nor U23693 (N_23693,N_23089,N_23052);
xnor U23694 (N_23694,N_22969,N_23134);
and U23695 (N_23695,N_23206,N_23334);
nor U23696 (N_23696,N_22937,N_23181);
xnor U23697 (N_23697,N_23094,N_23210);
or U23698 (N_23698,N_23182,N_23047);
nand U23699 (N_23699,N_23159,N_23131);
or U23700 (N_23700,N_22866,N_22948);
nand U23701 (N_23701,N_22948,N_23399);
and U23702 (N_23702,N_23396,N_22985);
nor U23703 (N_23703,N_23093,N_23279);
and U23704 (N_23704,N_23229,N_23296);
and U23705 (N_23705,N_23391,N_22963);
xnor U23706 (N_23706,N_22917,N_23338);
nand U23707 (N_23707,N_23007,N_22870);
nor U23708 (N_23708,N_22832,N_23187);
nor U23709 (N_23709,N_22890,N_23238);
or U23710 (N_23710,N_23169,N_23252);
nand U23711 (N_23711,N_23102,N_23194);
or U23712 (N_23712,N_23305,N_22920);
xnor U23713 (N_23713,N_23051,N_22847);
xor U23714 (N_23714,N_23104,N_23341);
nand U23715 (N_23715,N_23340,N_23195);
nand U23716 (N_23716,N_23237,N_23179);
nor U23717 (N_23717,N_23321,N_23285);
and U23718 (N_23718,N_23009,N_22912);
and U23719 (N_23719,N_23034,N_22829);
or U23720 (N_23720,N_23398,N_23375);
and U23721 (N_23721,N_22835,N_22995);
xnor U23722 (N_23722,N_22820,N_22867);
nand U23723 (N_23723,N_23034,N_23024);
xnor U23724 (N_23724,N_23037,N_23299);
nor U23725 (N_23725,N_23314,N_22993);
and U23726 (N_23726,N_23363,N_23219);
nand U23727 (N_23727,N_23359,N_22889);
nor U23728 (N_23728,N_22870,N_22865);
or U23729 (N_23729,N_23247,N_23379);
and U23730 (N_23730,N_23265,N_23122);
nand U23731 (N_23731,N_22817,N_22947);
and U23732 (N_23732,N_23012,N_23299);
nand U23733 (N_23733,N_23150,N_22912);
xor U23734 (N_23734,N_23258,N_23250);
xor U23735 (N_23735,N_23096,N_22995);
or U23736 (N_23736,N_23053,N_22960);
and U23737 (N_23737,N_23066,N_22898);
or U23738 (N_23738,N_23084,N_22909);
nand U23739 (N_23739,N_23177,N_23115);
or U23740 (N_23740,N_23366,N_22840);
nand U23741 (N_23741,N_23006,N_23043);
nand U23742 (N_23742,N_23027,N_22844);
nor U23743 (N_23743,N_23149,N_22853);
or U23744 (N_23744,N_23199,N_23379);
nor U23745 (N_23745,N_22978,N_23047);
nor U23746 (N_23746,N_23089,N_22814);
nand U23747 (N_23747,N_23003,N_22997);
or U23748 (N_23748,N_23287,N_22866);
xor U23749 (N_23749,N_23131,N_23168);
and U23750 (N_23750,N_22984,N_22909);
nor U23751 (N_23751,N_22884,N_22967);
nor U23752 (N_23752,N_22958,N_22943);
xor U23753 (N_23753,N_22987,N_23338);
or U23754 (N_23754,N_23166,N_23370);
xnor U23755 (N_23755,N_22854,N_22952);
nand U23756 (N_23756,N_23174,N_22900);
nand U23757 (N_23757,N_23351,N_22943);
and U23758 (N_23758,N_23180,N_23156);
and U23759 (N_23759,N_23383,N_22983);
nor U23760 (N_23760,N_22892,N_22867);
nor U23761 (N_23761,N_23050,N_23019);
nor U23762 (N_23762,N_23132,N_23051);
nor U23763 (N_23763,N_23091,N_22885);
nor U23764 (N_23764,N_23203,N_23277);
and U23765 (N_23765,N_23132,N_22847);
nor U23766 (N_23766,N_22831,N_23396);
xor U23767 (N_23767,N_23033,N_23037);
or U23768 (N_23768,N_22884,N_23326);
nor U23769 (N_23769,N_23321,N_22885);
or U23770 (N_23770,N_23230,N_22877);
nor U23771 (N_23771,N_23395,N_23359);
nand U23772 (N_23772,N_23256,N_22887);
nor U23773 (N_23773,N_23060,N_23214);
and U23774 (N_23774,N_22994,N_23068);
xnor U23775 (N_23775,N_23296,N_23228);
and U23776 (N_23776,N_22865,N_23313);
nor U23777 (N_23777,N_23008,N_22885);
xor U23778 (N_23778,N_22916,N_23030);
and U23779 (N_23779,N_23309,N_22880);
or U23780 (N_23780,N_23388,N_23280);
nor U23781 (N_23781,N_23109,N_23330);
and U23782 (N_23782,N_22856,N_22939);
xnor U23783 (N_23783,N_22861,N_22935);
nor U23784 (N_23784,N_22934,N_22895);
and U23785 (N_23785,N_23199,N_23176);
xnor U23786 (N_23786,N_23141,N_23014);
or U23787 (N_23787,N_23174,N_23153);
nand U23788 (N_23788,N_23366,N_23142);
nand U23789 (N_23789,N_23148,N_23270);
nand U23790 (N_23790,N_22973,N_23289);
and U23791 (N_23791,N_22803,N_23272);
nor U23792 (N_23792,N_23379,N_23389);
nand U23793 (N_23793,N_22813,N_23100);
or U23794 (N_23794,N_22992,N_22901);
or U23795 (N_23795,N_23389,N_23142);
xor U23796 (N_23796,N_23282,N_23333);
nor U23797 (N_23797,N_23065,N_22857);
xor U23798 (N_23798,N_22964,N_23053);
and U23799 (N_23799,N_23034,N_23195);
or U23800 (N_23800,N_23034,N_23351);
nor U23801 (N_23801,N_23069,N_23131);
or U23802 (N_23802,N_23040,N_23229);
or U23803 (N_23803,N_22970,N_23228);
or U23804 (N_23804,N_22956,N_22947);
nand U23805 (N_23805,N_22884,N_23393);
xnor U23806 (N_23806,N_23096,N_23124);
xor U23807 (N_23807,N_23237,N_23307);
nand U23808 (N_23808,N_23058,N_23179);
and U23809 (N_23809,N_22983,N_23000);
or U23810 (N_23810,N_23022,N_22844);
nor U23811 (N_23811,N_23150,N_23199);
xor U23812 (N_23812,N_22994,N_23043);
or U23813 (N_23813,N_22886,N_23273);
xnor U23814 (N_23814,N_23219,N_23103);
nand U23815 (N_23815,N_23099,N_23184);
or U23816 (N_23816,N_23051,N_23240);
and U23817 (N_23817,N_22952,N_23208);
or U23818 (N_23818,N_23011,N_22837);
xnor U23819 (N_23819,N_23184,N_23237);
xnor U23820 (N_23820,N_23146,N_22943);
or U23821 (N_23821,N_22893,N_23264);
and U23822 (N_23822,N_23021,N_23055);
or U23823 (N_23823,N_23189,N_23025);
xnor U23824 (N_23824,N_23248,N_22933);
nor U23825 (N_23825,N_23103,N_23248);
nand U23826 (N_23826,N_22913,N_23200);
and U23827 (N_23827,N_23061,N_23356);
or U23828 (N_23828,N_23286,N_23173);
xnor U23829 (N_23829,N_23095,N_22849);
nor U23830 (N_23830,N_22886,N_22983);
nor U23831 (N_23831,N_23183,N_23188);
nor U23832 (N_23832,N_23016,N_23348);
nand U23833 (N_23833,N_23305,N_23043);
and U23834 (N_23834,N_22967,N_23044);
or U23835 (N_23835,N_22820,N_23080);
nor U23836 (N_23836,N_22862,N_23180);
xnor U23837 (N_23837,N_23148,N_22838);
xor U23838 (N_23838,N_23163,N_23249);
nor U23839 (N_23839,N_23020,N_22834);
and U23840 (N_23840,N_23392,N_22914);
nand U23841 (N_23841,N_23126,N_23207);
nand U23842 (N_23842,N_22999,N_22939);
or U23843 (N_23843,N_23271,N_22883);
or U23844 (N_23844,N_23394,N_23058);
nor U23845 (N_23845,N_23216,N_23102);
and U23846 (N_23846,N_23059,N_23324);
xnor U23847 (N_23847,N_23152,N_22894);
xor U23848 (N_23848,N_23247,N_22959);
xnor U23849 (N_23849,N_23271,N_22926);
nor U23850 (N_23850,N_23145,N_23359);
nor U23851 (N_23851,N_22948,N_23151);
or U23852 (N_23852,N_23151,N_23155);
nand U23853 (N_23853,N_23382,N_23065);
or U23854 (N_23854,N_23241,N_23161);
or U23855 (N_23855,N_23160,N_23129);
nor U23856 (N_23856,N_23121,N_23300);
nor U23857 (N_23857,N_23153,N_23022);
nor U23858 (N_23858,N_23368,N_22861);
and U23859 (N_23859,N_23030,N_23072);
or U23860 (N_23860,N_23189,N_22892);
xnor U23861 (N_23861,N_23220,N_22814);
xor U23862 (N_23862,N_23180,N_23373);
xor U23863 (N_23863,N_23368,N_23290);
nand U23864 (N_23864,N_22902,N_23335);
xor U23865 (N_23865,N_23156,N_22919);
and U23866 (N_23866,N_23178,N_22988);
and U23867 (N_23867,N_22834,N_22903);
and U23868 (N_23868,N_23067,N_23141);
and U23869 (N_23869,N_23357,N_23268);
nor U23870 (N_23870,N_22999,N_23351);
or U23871 (N_23871,N_23370,N_23052);
or U23872 (N_23872,N_23060,N_23336);
xor U23873 (N_23873,N_23189,N_23064);
and U23874 (N_23874,N_22847,N_22968);
or U23875 (N_23875,N_23347,N_23289);
xor U23876 (N_23876,N_23003,N_23044);
and U23877 (N_23877,N_23261,N_22838);
xor U23878 (N_23878,N_23297,N_22938);
and U23879 (N_23879,N_23035,N_22823);
nand U23880 (N_23880,N_22999,N_23313);
and U23881 (N_23881,N_23293,N_23053);
and U23882 (N_23882,N_23344,N_22905);
nand U23883 (N_23883,N_23260,N_23273);
or U23884 (N_23884,N_23216,N_22824);
nor U23885 (N_23885,N_22991,N_23197);
xor U23886 (N_23886,N_22867,N_23219);
or U23887 (N_23887,N_22963,N_23100);
nor U23888 (N_23888,N_23317,N_22807);
nand U23889 (N_23889,N_23017,N_23118);
nand U23890 (N_23890,N_23327,N_22901);
nor U23891 (N_23891,N_22901,N_22994);
xor U23892 (N_23892,N_23279,N_23078);
nand U23893 (N_23893,N_22888,N_23337);
nor U23894 (N_23894,N_23300,N_23304);
nand U23895 (N_23895,N_23258,N_23291);
nor U23896 (N_23896,N_23206,N_23168);
xnor U23897 (N_23897,N_23129,N_22980);
xor U23898 (N_23898,N_22954,N_22890);
or U23899 (N_23899,N_23352,N_22871);
xor U23900 (N_23900,N_22887,N_23096);
nand U23901 (N_23901,N_22853,N_22863);
xor U23902 (N_23902,N_23306,N_22861);
and U23903 (N_23903,N_22990,N_23153);
nor U23904 (N_23904,N_23205,N_23382);
nor U23905 (N_23905,N_22857,N_23287);
or U23906 (N_23906,N_23330,N_22806);
xnor U23907 (N_23907,N_22936,N_23184);
and U23908 (N_23908,N_22963,N_23353);
nand U23909 (N_23909,N_23220,N_22891);
or U23910 (N_23910,N_22866,N_23285);
or U23911 (N_23911,N_23142,N_22801);
and U23912 (N_23912,N_23325,N_23292);
xor U23913 (N_23913,N_23034,N_23067);
nand U23914 (N_23914,N_23075,N_23397);
xnor U23915 (N_23915,N_22991,N_23260);
nor U23916 (N_23916,N_23012,N_23110);
nand U23917 (N_23917,N_23189,N_23187);
and U23918 (N_23918,N_22896,N_23231);
nor U23919 (N_23919,N_22949,N_23002);
nor U23920 (N_23920,N_23385,N_22907);
and U23921 (N_23921,N_22892,N_23018);
nand U23922 (N_23922,N_23391,N_23208);
or U23923 (N_23923,N_22975,N_23232);
nor U23924 (N_23924,N_22915,N_23275);
xor U23925 (N_23925,N_23393,N_22945);
or U23926 (N_23926,N_22909,N_23336);
nor U23927 (N_23927,N_22835,N_22932);
nor U23928 (N_23928,N_23334,N_22911);
nor U23929 (N_23929,N_23242,N_23225);
xor U23930 (N_23930,N_23021,N_22946);
xor U23931 (N_23931,N_23313,N_23195);
nor U23932 (N_23932,N_22825,N_23347);
nand U23933 (N_23933,N_22844,N_22864);
nor U23934 (N_23934,N_23291,N_23207);
nor U23935 (N_23935,N_23000,N_23265);
nor U23936 (N_23936,N_23056,N_23364);
or U23937 (N_23937,N_23304,N_23270);
or U23938 (N_23938,N_23184,N_23047);
or U23939 (N_23939,N_23021,N_22963);
and U23940 (N_23940,N_23147,N_23023);
and U23941 (N_23941,N_23024,N_23187);
and U23942 (N_23942,N_23364,N_23010);
and U23943 (N_23943,N_22845,N_22800);
or U23944 (N_23944,N_22919,N_23375);
or U23945 (N_23945,N_23184,N_23271);
or U23946 (N_23946,N_22864,N_23056);
and U23947 (N_23947,N_22859,N_23117);
nand U23948 (N_23948,N_23118,N_23133);
and U23949 (N_23949,N_22866,N_22846);
xnor U23950 (N_23950,N_22885,N_23270);
or U23951 (N_23951,N_22816,N_22912);
or U23952 (N_23952,N_23203,N_22898);
nor U23953 (N_23953,N_23033,N_23147);
nor U23954 (N_23954,N_22980,N_23049);
nor U23955 (N_23955,N_22925,N_23048);
and U23956 (N_23956,N_22908,N_22941);
or U23957 (N_23957,N_23168,N_23393);
or U23958 (N_23958,N_23397,N_23135);
nand U23959 (N_23959,N_23350,N_23090);
xnor U23960 (N_23960,N_23052,N_23245);
and U23961 (N_23961,N_23298,N_23044);
nor U23962 (N_23962,N_23073,N_22869);
or U23963 (N_23963,N_22864,N_23181);
or U23964 (N_23964,N_23241,N_23320);
or U23965 (N_23965,N_23104,N_22815);
and U23966 (N_23966,N_23184,N_23364);
nor U23967 (N_23967,N_23353,N_22937);
nor U23968 (N_23968,N_22848,N_22954);
nor U23969 (N_23969,N_23372,N_23039);
or U23970 (N_23970,N_23136,N_22851);
xor U23971 (N_23971,N_23125,N_23315);
nor U23972 (N_23972,N_23181,N_23061);
or U23973 (N_23973,N_23128,N_23005);
xor U23974 (N_23974,N_23094,N_23379);
xor U23975 (N_23975,N_23122,N_23234);
nor U23976 (N_23976,N_22968,N_23294);
nor U23977 (N_23977,N_23235,N_22955);
and U23978 (N_23978,N_22910,N_23187);
nor U23979 (N_23979,N_23296,N_22878);
and U23980 (N_23980,N_23276,N_22851);
and U23981 (N_23981,N_22962,N_23219);
and U23982 (N_23982,N_22929,N_23258);
and U23983 (N_23983,N_22839,N_23328);
and U23984 (N_23984,N_22967,N_22852);
and U23985 (N_23985,N_22837,N_23261);
or U23986 (N_23986,N_22880,N_23335);
nand U23987 (N_23987,N_22868,N_23233);
nand U23988 (N_23988,N_23178,N_22933);
or U23989 (N_23989,N_22820,N_23138);
nor U23990 (N_23990,N_23209,N_23306);
nand U23991 (N_23991,N_23039,N_22908);
or U23992 (N_23992,N_23155,N_22888);
xor U23993 (N_23993,N_23023,N_22867);
xnor U23994 (N_23994,N_23282,N_22960);
or U23995 (N_23995,N_23184,N_23149);
nor U23996 (N_23996,N_23137,N_23177);
xnor U23997 (N_23997,N_23142,N_22814);
nor U23998 (N_23998,N_23299,N_23338);
xor U23999 (N_23999,N_22872,N_22802);
and U24000 (N_24000,N_23792,N_23851);
xnor U24001 (N_24001,N_23667,N_23848);
or U24002 (N_24002,N_23646,N_23766);
xnor U24003 (N_24003,N_23659,N_23897);
and U24004 (N_24004,N_23807,N_23689);
nand U24005 (N_24005,N_23534,N_23495);
nor U24006 (N_24006,N_23912,N_23533);
or U24007 (N_24007,N_23625,N_23428);
nand U24008 (N_24008,N_23862,N_23571);
nand U24009 (N_24009,N_23749,N_23902);
and U24010 (N_24010,N_23997,N_23604);
or U24011 (N_24011,N_23596,N_23471);
xnor U24012 (N_24012,N_23413,N_23568);
nor U24013 (N_24013,N_23401,N_23884);
and U24014 (N_24014,N_23705,N_23589);
nand U24015 (N_24015,N_23765,N_23810);
xor U24016 (N_24016,N_23979,N_23900);
and U24017 (N_24017,N_23719,N_23984);
xor U24018 (N_24018,N_23639,N_23505);
or U24019 (N_24019,N_23592,N_23929);
or U24020 (N_24020,N_23799,N_23951);
xor U24021 (N_24021,N_23905,N_23873);
or U24022 (N_24022,N_23891,N_23725);
and U24023 (N_24023,N_23650,N_23866);
nor U24024 (N_24024,N_23886,N_23797);
xnor U24025 (N_24025,N_23861,N_23580);
nor U24026 (N_24026,N_23594,N_23536);
or U24027 (N_24027,N_23586,N_23924);
and U24028 (N_24028,N_23809,N_23709);
nor U24029 (N_24029,N_23971,N_23754);
nor U24030 (N_24030,N_23697,N_23598);
nor U24031 (N_24031,N_23467,N_23635);
nor U24032 (N_24032,N_23478,N_23508);
nor U24033 (N_24033,N_23856,N_23877);
and U24034 (N_24034,N_23823,N_23785);
xnor U24035 (N_24035,N_23423,N_23842);
nand U24036 (N_24036,N_23717,N_23612);
and U24037 (N_24037,N_23798,N_23411);
and U24038 (N_24038,N_23437,N_23665);
and U24039 (N_24039,N_23706,N_23913);
xnor U24040 (N_24040,N_23822,N_23811);
xnor U24041 (N_24041,N_23521,N_23513);
xnor U24042 (N_24042,N_23472,N_23552);
nand U24043 (N_24043,N_23400,N_23640);
nor U24044 (N_24044,N_23998,N_23479);
nor U24045 (N_24045,N_23915,N_23663);
or U24046 (N_24046,N_23961,N_23948);
or U24047 (N_24047,N_23932,N_23776);
xor U24048 (N_24048,N_23444,N_23456);
or U24049 (N_24049,N_23492,N_23645);
nand U24050 (N_24050,N_23581,N_23933);
and U24051 (N_24051,N_23484,N_23517);
xnor U24052 (N_24052,N_23519,N_23488);
and U24053 (N_24053,N_23840,N_23599);
nand U24054 (N_24054,N_23652,N_23853);
xor U24055 (N_24055,N_23416,N_23942);
or U24056 (N_24056,N_23977,N_23660);
nor U24057 (N_24057,N_23728,N_23629);
nand U24058 (N_24058,N_23607,N_23542);
nand U24059 (N_24059,N_23459,N_23541);
nor U24060 (N_24060,N_23889,N_23618);
xor U24061 (N_24061,N_23720,N_23623);
or U24062 (N_24062,N_23457,N_23914);
and U24063 (N_24063,N_23516,N_23414);
and U24064 (N_24064,N_23672,N_23812);
nand U24065 (N_24065,N_23554,N_23608);
nand U24066 (N_24066,N_23702,N_23895);
xor U24067 (N_24067,N_23434,N_23491);
nand U24068 (N_24068,N_23818,N_23701);
xnor U24069 (N_24069,N_23990,N_23758);
and U24070 (N_24070,N_23455,N_23600);
nand U24071 (N_24071,N_23616,N_23547);
xor U24072 (N_24072,N_23863,N_23801);
nor U24073 (N_24073,N_23800,N_23966);
and U24074 (N_24074,N_23772,N_23871);
xor U24075 (N_24075,N_23538,N_23458);
or U24076 (N_24076,N_23675,N_23658);
or U24077 (N_24077,N_23838,N_23831);
and U24078 (N_24078,N_23826,N_23733);
nand U24079 (N_24079,N_23920,N_23903);
xnor U24080 (N_24080,N_23816,N_23908);
or U24081 (N_24081,N_23893,N_23576);
nor U24082 (N_24082,N_23806,N_23967);
xor U24083 (N_24083,N_23734,N_23627);
xnor U24084 (N_24084,N_23885,N_23588);
or U24085 (N_24085,N_23653,N_23408);
nand U24086 (N_24086,N_23759,N_23703);
nand U24087 (N_24087,N_23503,N_23969);
nor U24088 (N_24088,N_23791,N_23779);
nor U24089 (N_24089,N_23959,N_23614);
nand U24090 (N_24090,N_23683,N_23922);
xor U24091 (N_24091,N_23539,N_23795);
and U24092 (N_24092,N_23778,N_23518);
and U24093 (N_24093,N_23497,N_23919);
or U24094 (N_24094,N_23679,N_23910);
nor U24095 (N_24095,N_23960,N_23739);
and U24096 (N_24096,N_23845,N_23832);
xor U24097 (N_24097,N_23502,N_23407);
nor U24098 (N_24098,N_23964,N_23954);
xor U24099 (N_24099,N_23436,N_23514);
or U24100 (N_24100,N_23859,N_23753);
nor U24101 (N_24101,N_23546,N_23664);
nor U24102 (N_24102,N_23936,N_23412);
and U24103 (N_24103,N_23545,N_23881);
and U24104 (N_24104,N_23661,N_23402);
nand U24105 (N_24105,N_23793,N_23973);
or U24106 (N_24106,N_23738,N_23473);
nand U24107 (N_24107,N_23420,N_23763);
xor U24108 (N_24108,N_23712,N_23707);
and U24109 (N_24109,N_23633,N_23926);
xnor U24110 (N_24110,N_23958,N_23626);
nor U24111 (N_24111,N_23642,N_23982);
nor U24112 (N_24112,N_23510,N_23916);
xnor U24113 (N_24113,N_23846,N_23480);
nor U24114 (N_24114,N_23943,N_23424);
xor U24115 (N_24115,N_23737,N_23898);
or U24116 (N_24116,N_23708,N_23606);
nor U24117 (N_24117,N_23711,N_23621);
nor U24118 (N_24118,N_23965,N_23449);
and U24119 (N_24119,N_23777,N_23418);
nor U24120 (N_24120,N_23637,N_23446);
nand U24121 (N_24121,N_23493,N_23744);
xnor U24122 (N_24122,N_23764,N_23427);
nor U24123 (N_24123,N_23590,N_23980);
nand U24124 (N_24124,N_23573,N_23462);
nand U24125 (N_24125,N_23406,N_23988);
nor U24126 (N_24126,N_23403,N_23947);
or U24127 (N_24127,N_23894,N_23433);
and U24128 (N_24128,N_23559,N_23578);
nand U24129 (N_24129,N_23722,N_23788);
nand U24130 (N_24130,N_23803,N_23551);
nand U24131 (N_24131,N_23487,N_23426);
xor U24132 (N_24132,N_23574,N_23431);
and U24133 (N_24133,N_23666,N_23847);
or U24134 (N_24134,N_23858,N_23579);
nand U24135 (N_24135,N_23419,N_23532);
or U24136 (N_24136,N_23745,N_23986);
xnor U24137 (N_24137,N_23756,N_23714);
or U24138 (N_24138,N_23972,N_23904);
or U24139 (N_24139,N_23976,N_23565);
or U24140 (N_24140,N_23481,N_23544);
nand U24141 (N_24141,N_23781,N_23691);
nor U24142 (N_24142,N_23981,N_23819);
and U24143 (N_24143,N_23483,N_23991);
or U24144 (N_24144,N_23624,N_23918);
and U24145 (N_24145,N_23655,N_23743);
nand U24146 (N_24146,N_23435,N_23970);
nor U24147 (N_24147,N_23887,N_23732);
and U24148 (N_24148,N_23713,N_23515);
nor U24149 (N_24149,N_23556,N_23787);
nor U24150 (N_24150,N_23582,N_23489);
nand U24151 (N_24151,N_23775,N_23553);
nand U24152 (N_24152,N_23825,N_23726);
and U24153 (N_24153,N_23501,N_23693);
nor U24154 (N_24154,N_23802,N_23453);
or U24155 (N_24155,N_23724,N_23525);
and U24156 (N_24156,N_23685,N_23888);
xnor U24157 (N_24157,N_23794,N_23837);
nor U24158 (N_24158,N_23439,N_23716);
and U24159 (N_24159,N_23448,N_23486);
or U24160 (N_24160,N_23469,N_23432);
xnor U24161 (N_24161,N_23610,N_23657);
and U24162 (N_24162,N_23855,N_23928);
and U24163 (N_24163,N_23442,N_23696);
and U24164 (N_24164,N_23727,N_23796);
nor U24165 (N_24165,N_23975,N_23814);
and U24166 (N_24166,N_23784,N_23499);
or U24167 (N_24167,N_23482,N_23773);
or U24168 (N_24168,N_23690,N_23562);
xor U24169 (N_24169,N_23937,N_23949);
and U24170 (N_24170,N_23561,N_23874);
nor U24171 (N_24171,N_23901,N_23537);
nand U24172 (N_24172,N_23741,N_23694);
or U24173 (N_24173,N_23995,N_23867);
nor U24174 (N_24174,N_23549,N_23835);
and U24175 (N_24175,N_23992,N_23834);
nand U24176 (N_24176,N_23445,N_23931);
nand U24177 (N_24177,N_23944,N_23595);
and U24178 (N_24178,N_23630,N_23836);
or U24179 (N_24179,N_23490,N_23939);
and U24180 (N_24180,N_23715,N_23955);
or U24181 (N_24181,N_23723,N_23421);
or U24182 (N_24182,N_23555,N_23450);
and U24183 (N_24183,N_23742,N_23882);
nand U24184 (N_24184,N_23934,N_23828);
nor U24185 (N_24185,N_23425,N_23429);
xnor U24186 (N_24186,N_23447,N_23570);
or U24187 (N_24187,N_23940,N_23619);
nand U24188 (N_24188,N_23978,N_23466);
or U24189 (N_24189,N_23524,N_23643);
and U24190 (N_24190,N_23470,N_23527);
nand U24191 (N_24191,N_23464,N_23774);
or U24192 (N_24192,N_23875,N_23746);
xnor U24193 (N_24193,N_23617,N_23632);
nand U24194 (N_24194,N_23747,N_23415);
and U24195 (N_24195,N_23654,N_23682);
nand U24196 (N_24196,N_23849,N_23935);
and U24197 (N_24197,N_23963,N_23730);
nand U24198 (N_24198,N_23656,N_23852);
nand U24199 (N_24199,N_23647,N_23460);
xnor U24200 (N_24200,N_23587,N_23671);
or U24201 (N_24201,N_23463,N_23631);
xnor U24202 (N_24202,N_23535,N_23648);
and U24203 (N_24203,N_23699,N_23644);
and U24204 (N_24204,N_23824,N_23560);
nor U24205 (N_24205,N_23504,N_23974);
xor U24206 (N_24206,N_23520,N_23477);
nor U24207 (N_24207,N_23996,N_23899);
and U24208 (N_24208,N_23540,N_23569);
or U24209 (N_24209,N_23805,N_23748);
nor U24210 (N_24210,N_23718,N_23770);
and U24211 (N_24211,N_23443,N_23669);
nor U24212 (N_24212,N_23827,N_23622);
xor U24213 (N_24213,N_23465,N_23789);
xnor U24214 (N_24214,N_23755,N_23839);
nand U24215 (N_24215,N_23417,N_23687);
or U24216 (N_24216,N_23760,N_23957);
nor U24217 (N_24217,N_23767,N_23678);
or U24218 (N_24218,N_23968,N_23662);
or U24219 (N_24219,N_23509,N_23485);
nor U24220 (N_24220,N_23896,N_23651);
or U24221 (N_24221,N_23989,N_23609);
nor U24222 (N_24222,N_23602,N_23768);
and U24223 (N_24223,N_23451,N_23790);
nor U24224 (N_24224,N_23557,N_23761);
or U24225 (N_24225,N_23577,N_23771);
nor U24226 (N_24226,N_23751,N_23528);
xor U24227 (N_24227,N_23636,N_23952);
nor U24228 (N_24228,N_23878,N_23870);
nand U24229 (N_24229,N_23860,N_23422);
nor U24230 (N_24230,N_23808,N_23620);
nor U24231 (N_24231,N_23543,N_23649);
nand U24232 (N_24232,N_23454,N_23410);
xnor U24233 (N_24233,N_23677,N_23605);
xnor U24234 (N_24234,N_23476,N_23813);
and U24235 (N_24235,N_23925,N_23927);
nor U24236 (N_24236,N_23868,N_23531);
nand U24237 (N_24237,N_23404,N_23731);
and U24238 (N_24238,N_23548,N_23597);
xnor U24239 (N_24239,N_23880,N_23945);
and U24240 (N_24240,N_23566,N_23953);
or U24241 (N_24241,N_23686,N_23729);
and U24242 (N_24242,N_23591,N_23750);
xnor U24243 (N_24243,N_23634,N_23804);
nor U24244 (N_24244,N_23833,N_23841);
nor U24245 (N_24245,N_23704,N_23550);
nand U24246 (N_24246,N_23921,N_23430);
and U24247 (N_24247,N_23879,N_23830);
nand U24248 (N_24248,N_23983,N_23909);
and U24249 (N_24249,N_23684,N_23769);
nor U24250 (N_24250,N_23680,N_23780);
nand U24251 (N_24251,N_23611,N_23613);
and U24252 (N_24252,N_23530,N_23512);
nor U24253 (N_24253,N_23815,N_23821);
or U24254 (N_24254,N_23500,N_23872);
nor U24255 (N_24255,N_23917,N_23681);
nor U24256 (N_24256,N_23615,N_23529);
xor U24257 (N_24257,N_23567,N_23695);
or U24258 (N_24258,N_23883,N_23564);
xor U24259 (N_24259,N_23911,N_23628);
and U24260 (N_24260,N_23593,N_23907);
and U24261 (N_24261,N_23710,N_23993);
or U24262 (N_24262,N_23946,N_23494);
xor U24263 (N_24263,N_23850,N_23923);
and U24264 (N_24264,N_23994,N_23575);
or U24265 (N_24265,N_23585,N_23956);
nand U24266 (N_24266,N_23721,N_23857);
nor U24267 (N_24267,N_23438,N_23890);
or U24268 (N_24268,N_23999,N_23700);
nand U24269 (N_24269,N_23752,N_23475);
nor U24270 (N_24270,N_23762,N_23817);
nand U24271 (N_24271,N_23962,N_23865);
xor U24272 (N_24272,N_23820,N_23930);
or U24273 (N_24273,N_23498,N_23735);
nor U24274 (N_24274,N_23941,N_23583);
nor U24275 (N_24275,N_23938,N_23572);
nand U24276 (N_24276,N_23496,N_23698);
nand U24277 (N_24277,N_23876,N_23526);
nand U24278 (N_24278,N_23783,N_23786);
or U24279 (N_24279,N_23692,N_23603);
or U24280 (N_24280,N_23522,N_23452);
nor U24281 (N_24281,N_23674,N_23740);
nor U24282 (N_24282,N_23782,N_23673);
nand U24283 (N_24283,N_23950,N_23468);
and U24284 (N_24284,N_23638,N_23736);
xor U24285 (N_24285,N_23854,N_23474);
nand U24286 (N_24286,N_23688,N_23869);
xnor U24287 (N_24287,N_23892,N_23843);
or U24288 (N_24288,N_23563,N_23985);
nand U24289 (N_24289,N_23641,N_23405);
and U24290 (N_24290,N_23757,N_23584);
and U24291 (N_24291,N_23461,N_23511);
and U24292 (N_24292,N_23676,N_23441);
nand U24293 (N_24293,N_23906,N_23507);
or U24294 (N_24294,N_23558,N_23844);
nor U24295 (N_24295,N_23523,N_23506);
nor U24296 (N_24296,N_23409,N_23440);
nor U24297 (N_24297,N_23601,N_23670);
xor U24298 (N_24298,N_23864,N_23829);
and U24299 (N_24299,N_23987,N_23668);
nand U24300 (N_24300,N_23691,N_23547);
nand U24301 (N_24301,N_23895,N_23807);
or U24302 (N_24302,N_23525,N_23766);
and U24303 (N_24303,N_23592,N_23506);
xnor U24304 (N_24304,N_23664,N_23620);
or U24305 (N_24305,N_23924,N_23468);
nor U24306 (N_24306,N_23970,N_23904);
xor U24307 (N_24307,N_23698,N_23634);
or U24308 (N_24308,N_23507,N_23415);
xor U24309 (N_24309,N_23500,N_23658);
xnor U24310 (N_24310,N_23819,N_23590);
or U24311 (N_24311,N_23923,N_23771);
nand U24312 (N_24312,N_23928,N_23644);
nand U24313 (N_24313,N_23466,N_23936);
nand U24314 (N_24314,N_23978,N_23736);
or U24315 (N_24315,N_23838,N_23475);
or U24316 (N_24316,N_23972,N_23569);
nor U24317 (N_24317,N_23476,N_23662);
nor U24318 (N_24318,N_23744,N_23774);
and U24319 (N_24319,N_23461,N_23827);
or U24320 (N_24320,N_23830,N_23484);
or U24321 (N_24321,N_23987,N_23908);
nand U24322 (N_24322,N_23918,N_23419);
nand U24323 (N_24323,N_23683,N_23650);
nor U24324 (N_24324,N_23824,N_23920);
xnor U24325 (N_24325,N_23472,N_23415);
or U24326 (N_24326,N_23743,N_23855);
nor U24327 (N_24327,N_23620,N_23579);
and U24328 (N_24328,N_23841,N_23870);
nand U24329 (N_24329,N_23454,N_23847);
nor U24330 (N_24330,N_23860,N_23527);
xnor U24331 (N_24331,N_23845,N_23822);
xor U24332 (N_24332,N_23713,N_23944);
nor U24333 (N_24333,N_23623,N_23859);
or U24334 (N_24334,N_23864,N_23679);
and U24335 (N_24335,N_23799,N_23800);
nor U24336 (N_24336,N_23517,N_23537);
xnor U24337 (N_24337,N_23594,N_23592);
nor U24338 (N_24338,N_23425,N_23758);
nand U24339 (N_24339,N_23906,N_23739);
or U24340 (N_24340,N_23439,N_23621);
or U24341 (N_24341,N_23647,N_23578);
and U24342 (N_24342,N_23700,N_23951);
nor U24343 (N_24343,N_23853,N_23468);
nand U24344 (N_24344,N_23771,N_23547);
xor U24345 (N_24345,N_23967,N_23956);
nor U24346 (N_24346,N_23764,N_23697);
xor U24347 (N_24347,N_23403,N_23651);
xnor U24348 (N_24348,N_23807,N_23475);
nand U24349 (N_24349,N_23906,N_23498);
or U24350 (N_24350,N_23528,N_23718);
and U24351 (N_24351,N_23944,N_23937);
nor U24352 (N_24352,N_23882,N_23871);
nor U24353 (N_24353,N_23931,N_23703);
and U24354 (N_24354,N_23576,N_23574);
xnor U24355 (N_24355,N_23919,N_23520);
xor U24356 (N_24356,N_23899,N_23841);
nand U24357 (N_24357,N_23950,N_23934);
nand U24358 (N_24358,N_23655,N_23770);
or U24359 (N_24359,N_23871,N_23978);
xnor U24360 (N_24360,N_23597,N_23668);
nor U24361 (N_24361,N_23736,N_23840);
xor U24362 (N_24362,N_23586,N_23708);
xnor U24363 (N_24363,N_23497,N_23440);
xnor U24364 (N_24364,N_23464,N_23486);
nor U24365 (N_24365,N_23465,N_23943);
xnor U24366 (N_24366,N_23476,N_23745);
nor U24367 (N_24367,N_23418,N_23431);
and U24368 (N_24368,N_23889,N_23977);
or U24369 (N_24369,N_23626,N_23871);
and U24370 (N_24370,N_23428,N_23896);
nor U24371 (N_24371,N_23543,N_23591);
nand U24372 (N_24372,N_23852,N_23750);
and U24373 (N_24373,N_23853,N_23496);
and U24374 (N_24374,N_23755,N_23868);
and U24375 (N_24375,N_23592,N_23595);
nor U24376 (N_24376,N_23903,N_23833);
and U24377 (N_24377,N_23741,N_23852);
xnor U24378 (N_24378,N_23893,N_23548);
nand U24379 (N_24379,N_23974,N_23701);
and U24380 (N_24380,N_23412,N_23792);
nor U24381 (N_24381,N_23904,N_23570);
xnor U24382 (N_24382,N_23454,N_23515);
xor U24383 (N_24383,N_23662,N_23933);
nand U24384 (N_24384,N_23978,N_23825);
or U24385 (N_24385,N_23930,N_23556);
nand U24386 (N_24386,N_23922,N_23887);
xnor U24387 (N_24387,N_23731,N_23824);
or U24388 (N_24388,N_23534,N_23639);
xor U24389 (N_24389,N_23709,N_23839);
xnor U24390 (N_24390,N_23788,N_23932);
and U24391 (N_24391,N_23735,N_23613);
xnor U24392 (N_24392,N_23447,N_23682);
xnor U24393 (N_24393,N_23725,N_23994);
nand U24394 (N_24394,N_23470,N_23860);
and U24395 (N_24395,N_23829,N_23411);
nor U24396 (N_24396,N_23903,N_23968);
nand U24397 (N_24397,N_23402,N_23646);
xnor U24398 (N_24398,N_23881,N_23937);
nand U24399 (N_24399,N_23559,N_23647);
or U24400 (N_24400,N_23403,N_23622);
xor U24401 (N_24401,N_23547,N_23742);
or U24402 (N_24402,N_23847,N_23818);
xor U24403 (N_24403,N_23872,N_23697);
or U24404 (N_24404,N_23944,N_23493);
and U24405 (N_24405,N_23727,N_23473);
and U24406 (N_24406,N_23681,N_23543);
nor U24407 (N_24407,N_23626,N_23963);
and U24408 (N_24408,N_23525,N_23739);
nor U24409 (N_24409,N_23517,N_23905);
xnor U24410 (N_24410,N_23683,N_23743);
nor U24411 (N_24411,N_23406,N_23698);
xnor U24412 (N_24412,N_23437,N_23475);
xnor U24413 (N_24413,N_23533,N_23766);
and U24414 (N_24414,N_23972,N_23450);
xor U24415 (N_24415,N_23893,N_23666);
nor U24416 (N_24416,N_23845,N_23952);
nor U24417 (N_24417,N_23475,N_23820);
or U24418 (N_24418,N_23704,N_23682);
nor U24419 (N_24419,N_23401,N_23745);
nor U24420 (N_24420,N_23811,N_23833);
or U24421 (N_24421,N_23669,N_23401);
or U24422 (N_24422,N_23669,N_23573);
nand U24423 (N_24423,N_23427,N_23853);
and U24424 (N_24424,N_23855,N_23724);
and U24425 (N_24425,N_23641,N_23680);
nand U24426 (N_24426,N_23403,N_23460);
or U24427 (N_24427,N_23535,N_23571);
nand U24428 (N_24428,N_23444,N_23683);
nand U24429 (N_24429,N_23999,N_23591);
nor U24430 (N_24430,N_23822,N_23643);
or U24431 (N_24431,N_23616,N_23447);
nor U24432 (N_24432,N_23830,N_23574);
and U24433 (N_24433,N_23970,N_23746);
or U24434 (N_24434,N_23913,N_23922);
nor U24435 (N_24435,N_23415,N_23863);
and U24436 (N_24436,N_23455,N_23465);
and U24437 (N_24437,N_23621,N_23663);
nor U24438 (N_24438,N_23537,N_23868);
nand U24439 (N_24439,N_23771,N_23402);
or U24440 (N_24440,N_23848,N_23640);
xor U24441 (N_24441,N_23478,N_23894);
nor U24442 (N_24442,N_23658,N_23460);
nor U24443 (N_24443,N_23464,N_23974);
and U24444 (N_24444,N_23776,N_23438);
or U24445 (N_24445,N_23779,N_23796);
xor U24446 (N_24446,N_23854,N_23620);
nand U24447 (N_24447,N_23830,N_23593);
nand U24448 (N_24448,N_23854,N_23806);
nor U24449 (N_24449,N_23918,N_23572);
nor U24450 (N_24450,N_23470,N_23483);
nand U24451 (N_24451,N_23758,N_23706);
or U24452 (N_24452,N_23594,N_23506);
nand U24453 (N_24453,N_23856,N_23901);
nor U24454 (N_24454,N_23494,N_23815);
nand U24455 (N_24455,N_23880,N_23787);
xor U24456 (N_24456,N_23978,N_23810);
nor U24457 (N_24457,N_23716,N_23579);
nand U24458 (N_24458,N_23916,N_23943);
nor U24459 (N_24459,N_23495,N_23450);
or U24460 (N_24460,N_23637,N_23496);
nor U24461 (N_24461,N_23937,N_23821);
and U24462 (N_24462,N_23583,N_23515);
or U24463 (N_24463,N_23831,N_23882);
xor U24464 (N_24464,N_23982,N_23600);
xor U24465 (N_24465,N_23902,N_23987);
nor U24466 (N_24466,N_23859,N_23599);
or U24467 (N_24467,N_23831,N_23698);
or U24468 (N_24468,N_23537,N_23404);
and U24469 (N_24469,N_23679,N_23811);
or U24470 (N_24470,N_23635,N_23834);
nand U24471 (N_24471,N_23591,N_23790);
and U24472 (N_24472,N_23933,N_23615);
nor U24473 (N_24473,N_23638,N_23802);
xnor U24474 (N_24474,N_23659,N_23641);
nor U24475 (N_24475,N_23499,N_23899);
nand U24476 (N_24476,N_23929,N_23992);
nand U24477 (N_24477,N_23806,N_23658);
nor U24478 (N_24478,N_23663,N_23999);
and U24479 (N_24479,N_23646,N_23768);
xor U24480 (N_24480,N_23907,N_23668);
or U24481 (N_24481,N_23676,N_23926);
and U24482 (N_24482,N_23882,N_23907);
or U24483 (N_24483,N_23648,N_23794);
or U24484 (N_24484,N_23774,N_23843);
nor U24485 (N_24485,N_23582,N_23477);
nand U24486 (N_24486,N_23821,N_23555);
nand U24487 (N_24487,N_23822,N_23549);
nor U24488 (N_24488,N_23453,N_23841);
or U24489 (N_24489,N_23788,N_23756);
nor U24490 (N_24490,N_23790,N_23771);
or U24491 (N_24491,N_23530,N_23729);
and U24492 (N_24492,N_23797,N_23564);
nor U24493 (N_24493,N_23686,N_23634);
xor U24494 (N_24494,N_23546,N_23997);
and U24495 (N_24495,N_23557,N_23671);
or U24496 (N_24496,N_23574,N_23929);
or U24497 (N_24497,N_23676,N_23448);
nand U24498 (N_24498,N_23700,N_23666);
nor U24499 (N_24499,N_23616,N_23851);
or U24500 (N_24500,N_23411,N_23891);
and U24501 (N_24501,N_23589,N_23448);
nand U24502 (N_24502,N_23778,N_23835);
nor U24503 (N_24503,N_23849,N_23605);
and U24504 (N_24504,N_23598,N_23699);
or U24505 (N_24505,N_23735,N_23908);
nand U24506 (N_24506,N_23939,N_23786);
xor U24507 (N_24507,N_23783,N_23861);
nor U24508 (N_24508,N_23723,N_23948);
and U24509 (N_24509,N_23939,N_23555);
and U24510 (N_24510,N_23997,N_23787);
or U24511 (N_24511,N_23544,N_23717);
xor U24512 (N_24512,N_23793,N_23677);
and U24513 (N_24513,N_23465,N_23858);
nand U24514 (N_24514,N_23407,N_23996);
or U24515 (N_24515,N_23423,N_23511);
nand U24516 (N_24516,N_23408,N_23442);
and U24517 (N_24517,N_23803,N_23871);
or U24518 (N_24518,N_23673,N_23404);
nand U24519 (N_24519,N_23597,N_23549);
nor U24520 (N_24520,N_23828,N_23805);
or U24521 (N_24521,N_23690,N_23407);
nand U24522 (N_24522,N_23618,N_23599);
nand U24523 (N_24523,N_23797,N_23711);
and U24524 (N_24524,N_23882,N_23415);
or U24525 (N_24525,N_23955,N_23450);
xnor U24526 (N_24526,N_23680,N_23560);
and U24527 (N_24527,N_23720,N_23894);
nor U24528 (N_24528,N_23814,N_23825);
xnor U24529 (N_24529,N_23724,N_23479);
nor U24530 (N_24530,N_23659,N_23830);
nand U24531 (N_24531,N_23742,N_23864);
xnor U24532 (N_24532,N_23716,N_23979);
xor U24533 (N_24533,N_23913,N_23934);
nand U24534 (N_24534,N_23965,N_23801);
nor U24535 (N_24535,N_23651,N_23839);
and U24536 (N_24536,N_23736,N_23990);
or U24537 (N_24537,N_23437,N_23822);
or U24538 (N_24538,N_23956,N_23799);
xor U24539 (N_24539,N_23455,N_23862);
xor U24540 (N_24540,N_23605,N_23779);
nor U24541 (N_24541,N_23677,N_23508);
nor U24542 (N_24542,N_23626,N_23708);
xnor U24543 (N_24543,N_23627,N_23591);
nor U24544 (N_24544,N_23719,N_23982);
nor U24545 (N_24545,N_23915,N_23638);
nand U24546 (N_24546,N_23913,N_23838);
xnor U24547 (N_24547,N_23498,N_23835);
and U24548 (N_24548,N_23839,N_23473);
nand U24549 (N_24549,N_23427,N_23842);
and U24550 (N_24550,N_23813,N_23964);
and U24551 (N_24551,N_23825,N_23807);
and U24552 (N_24552,N_23609,N_23585);
nor U24553 (N_24553,N_23775,N_23459);
and U24554 (N_24554,N_23462,N_23472);
nand U24555 (N_24555,N_23656,N_23558);
xnor U24556 (N_24556,N_23478,N_23402);
nor U24557 (N_24557,N_23628,N_23712);
nand U24558 (N_24558,N_23987,N_23666);
xor U24559 (N_24559,N_23904,N_23683);
or U24560 (N_24560,N_23487,N_23513);
nand U24561 (N_24561,N_23917,N_23750);
xor U24562 (N_24562,N_23826,N_23827);
or U24563 (N_24563,N_23711,N_23474);
nand U24564 (N_24564,N_23608,N_23963);
and U24565 (N_24565,N_23830,N_23670);
xnor U24566 (N_24566,N_23402,N_23818);
nand U24567 (N_24567,N_23625,N_23527);
nor U24568 (N_24568,N_23694,N_23449);
nor U24569 (N_24569,N_23653,N_23416);
nand U24570 (N_24570,N_23774,N_23840);
xnor U24571 (N_24571,N_23505,N_23975);
nand U24572 (N_24572,N_23575,N_23750);
xor U24573 (N_24573,N_23684,N_23412);
and U24574 (N_24574,N_23765,N_23965);
nor U24575 (N_24575,N_23668,N_23672);
or U24576 (N_24576,N_23790,N_23627);
nor U24577 (N_24577,N_23603,N_23754);
and U24578 (N_24578,N_23713,N_23525);
xor U24579 (N_24579,N_23523,N_23410);
or U24580 (N_24580,N_23627,N_23722);
and U24581 (N_24581,N_23668,N_23594);
and U24582 (N_24582,N_23995,N_23668);
nand U24583 (N_24583,N_23964,N_23796);
xnor U24584 (N_24584,N_23582,N_23444);
or U24585 (N_24585,N_23945,N_23636);
xnor U24586 (N_24586,N_23616,N_23943);
and U24587 (N_24587,N_23718,N_23617);
and U24588 (N_24588,N_23730,N_23552);
xor U24589 (N_24589,N_23712,N_23975);
nor U24590 (N_24590,N_23793,N_23607);
xnor U24591 (N_24591,N_23816,N_23907);
and U24592 (N_24592,N_23881,N_23678);
xnor U24593 (N_24593,N_23667,N_23592);
nor U24594 (N_24594,N_23674,N_23739);
nand U24595 (N_24595,N_23820,N_23437);
nand U24596 (N_24596,N_23643,N_23909);
nand U24597 (N_24597,N_23876,N_23604);
or U24598 (N_24598,N_23775,N_23859);
nand U24599 (N_24599,N_23661,N_23965);
nand U24600 (N_24600,N_24420,N_24352);
xor U24601 (N_24601,N_24528,N_24300);
nand U24602 (N_24602,N_24366,N_24084);
and U24603 (N_24603,N_24510,N_24560);
nand U24604 (N_24604,N_24068,N_24421);
or U24605 (N_24605,N_24122,N_24441);
and U24606 (N_24606,N_24478,N_24156);
nor U24607 (N_24607,N_24577,N_24148);
nand U24608 (N_24608,N_24470,N_24091);
xnor U24609 (N_24609,N_24503,N_24354);
or U24610 (N_24610,N_24162,N_24115);
or U24611 (N_24611,N_24015,N_24059);
nor U24612 (N_24612,N_24297,N_24306);
nand U24613 (N_24613,N_24062,N_24022);
nand U24614 (N_24614,N_24449,N_24096);
nor U24615 (N_24615,N_24128,N_24439);
xor U24616 (N_24616,N_24320,N_24427);
or U24617 (N_24617,N_24559,N_24295);
and U24618 (N_24618,N_24269,N_24255);
or U24619 (N_24619,N_24339,N_24363);
nand U24620 (N_24620,N_24280,N_24271);
and U24621 (N_24621,N_24337,N_24580);
or U24622 (N_24622,N_24322,N_24292);
or U24623 (N_24623,N_24053,N_24565);
nand U24624 (N_24624,N_24511,N_24374);
or U24625 (N_24625,N_24395,N_24074);
or U24626 (N_24626,N_24129,N_24316);
nand U24627 (N_24627,N_24512,N_24442);
or U24628 (N_24628,N_24391,N_24151);
or U24629 (N_24629,N_24561,N_24536);
xor U24630 (N_24630,N_24153,N_24026);
or U24631 (N_24631,N_24370,N_24481);
or U24632 (N_24632,N_24276,N_24576);
nor U24633 (N_24633,N_24457,N_24033);
nor U24634 (N_24634,N_24000,N_24139);
xnor U24635 (N_24635,N_24309,N_24010);
nand U24636 (N_24636,N_24226,N_24400);
xnor U24637 (N_24637,N_24246,N_24112);
nand U24638 (N_24638,N_24546,N_24557);
nor U24639 (N_24639,N_24168,N_24463);
or U24640 (N_24640,N_24164,N_24399);
nand U24641 (N_24641,N_24278,N_24249);
nand U24642 (N_24642,N_24046,N_24023);
xor U24643 (N_24643,N_24516,N_24406);
and U24644 (N_24644,N_24458,N_24008);
xor U24645 (N_24645,N_24252,N_24445);
nor U24646 (N_24646,N_24346,N_24462);
and U24647 (N_24647,N_24248,N_24082);
and U24648 (N_24648,N_24054,N_24013);
or U24649 (N_24649,N_24019,N_24012);
and U24650 (N_24650,N_24069,N_24042);
nor U24651 (N_24651,N_24403,N_24589);
or U24652 (N_24652,N_24283,N_24152);
xnor U24653 (N_24653,N_24087,N_24055);
xnor U24654 (N_24654,N_24212,N_24450);
and U24655 (N_24655,N_24509,N_24459);
and U24656 (N_24656,N_24253,N_24437);
xnor U24657 (N_24657,N_24564,N_24174);
or U24658 (N_24658,N_24480,N_24104);
or U24659 (N_24659,N_24483,N_24235);
nand U24660 (N_24660,N_24185,N_24296);
and U24661 (N_24661,N_24359,N_24382);
or U24662 (N_24662,N_24380,N_24034);
or U24663 (N_24663,N_24488,N_24551);
nand U24664 (N_24664,N_24425,N_24251);
nor U24665 (N_24665,N_24085,N_24132);
or U24666 (N_24666,N_24213,N_24083);
and U24667 (N_24667,N_24570,N_24304);
and U24668 (N_24668,N_24529,N_24256);
xor U24669 (N_24669,N_24543,N_24250);
xnor U24670 (N_24670,N_24145,N_24274);
or U24671 (N_24671,N_24196,N_24094);
nand U24672 (N_24672,N_24279,N_24259);
or U24673 (N_24673,N_24195,N_24114);
nand U24674 (N_24674,N_24065,N_24461);
nor U24675 (N_24675,N_24327,N_24313);
or U24676 (N_24676,N_24206,N_24474);
nand U24677 (N_24677,N_24335,N_24429);
or U24678 (N_24678,N_24149,N_24171);
and U24679 (N_24679,N_24095,N_24435);
and U24680 (N_24680,N_24574,N_24314);
and U24681 (N_24681,N_24107,N_24507);
nand U24682 (N_24682,N_24423,N_24203);
and U24683 (N_24683,N_24092,N_24229);
xnor U24684 (N_24684,N_24569,N_24018);
or U24685 (N_24685,N_24179,N_24125);
and U24686 (N_24686,N_24016,N_24336);
nand U24687 (N_24687,N_24411,N_24245);
xnor U24688 (N_24688,N_24410,N_24358);
nor U24689 (N_24689,N_24475,N_24303);
nor U24690 (N_24690,N_24355,N_24590);
xnor U24691 (N_24691,N_24531,N_24290);
or U24692 (N_24692,N_24440,N_24538);
or U24693 (N_24693,N_24263,N_24289);
and U24694 (N_24694,N_24298,N_24581);
nor U24695 (N_24695,N_24455,N_24238);
nor U24696 (N_24696,N_24247,N_24090);
nand U24697 (N_24697,N_24323,N_24049);
xnor U24698 (N_24698,N_24479,N_24392);
nor U24699 (N_24699,N_24052,N_24522);
nor U24700 (N_24700,N_24077,N_24535);
nand U24701 (N_24701,N_24540,N_24446);
xor U24702 (N_24702,N_24430,N_24230);
and U24703 (N_24703,N_24341,N_24201);
xor U24704 (N_24704,N_24113,N_24556);
nor U24705 (N_24705,N_24039,N_24264);
nand U24706 (N_24706,N_24524,N_24121);
nor U24707 (N_24707,N_24072,N_24521);
nand U24708 (N_24708,N_24379,N_24209);
xnor U24709 (N_24709,N_24351,N_24050);
nand U24710 (N_24710,N_24386,N_24007);
and U24711 (N_24711,N_24527,N_24473);
nor U24712 (N_24712,N_24242,N_24599);
nor U24713 (N_24713,N_24377,N_24293);
nand U24714 (N_24714,N_24554,N_24431);
xnor U24715 (N_24715,N_24011,N_24378);
nand U24716 (N_24716,N_24312,N_24004);
nor U24717 (N_24717,N_24387,N_24542);
nand U24718 (N_24718,N_24040,N_24534);
or U24719 (N_24719,N_24286,N_24585);
nand U24720 (N_24720,N_24071,N_24166);
or U24721 (N_24721,N_24109,N_24070);
and U24722 (N_24722,N_24281,N_24329);
nor U24723 (N_24723,N_24262,N_24558);
nor U24724 (N_24724,N_24258,N_24003);
nor U24725 (N_24725,N_24191,N_24552);
and U24726 (N_24726,N_24364,N_24482);
nor U24727 (N_24727,N_24302,N_24595);
and U24728 (N_24728,N_24525,N_24273);
nand U24729 (N_24729,N_24267,N_24402);
or U24730 (N_24730,N_24566,N_24224);
and U24731 (N_24731,N_24343,N_24284);
and U24732 (N_24732,N_24257,N_24562);
xor U24733 (N_24733,N_24150,N_24079);
nor U24734 (N_24734,N_24424,N_24240);
nand U24735 (N_24735,N_24357,N_24194);
and U24736 (N_24736,N_24025,N_24385);
nor U24737 (N_24737,N_24118,N_24147);
xor U24738 (N_24738,N_24029,N_24088);
nand U24739 (N_24739,N_24078,N_24447);
or U24740 (N_24740,N_24130,N_24157);
or U24741 (N_24741,N_24197,N_24381);
nor U24742 (N_24742,N_24494,N_24367);
nand U24743 (N_24743,N_24066,N_24591);
xor U24744 (N_24744,N_24338,N_24567);
and U24745 (N_24745,N_24575,N_24161);
or U24746 (N_24746,N_24178,N_24321);
nand U24747 (N_24747,N_24319,N_24513);
nor U24748 (N_24748,N_24434,N_24448);
nand U24749 (N_24749,N_24127,N_24124);
nor U24750 (N_24750,N_24371,N_24519);
nand U24751 (N_24751,N_24523,N_24460);
nor U24752 (N_24752,N_24412,N_24444);
xor U24753 (N_24753,N_24108,N_24270);
xnor U24754 (N_24754,N_24307,N_24135);
or U24755 (N_24755,N_24187,N_24080);
xor U24756 (N_24756,N_24549,N_24202);
and U24757 (N_24757,N_24433,N_24426);
nor U24758 (N_24758,N_24176,N_24453);
nand U24759 (N_24759,N_24117,N_24227);
and U24760 (N_24760,N_24401,N_24582);
or U24761 (N_24761,N_24517,N_24443);
or U24762 (N_24762,N_24515,N_24225);
nand U24763 (N_24763,N_24404,N_24597);
or U24764 (N_24764,N_24553,N_24001);
nor U24765 (N_24765,N_24190,N_24102);
and U24766 (N_24766,N_24594,N_24484);
xor U24767 (N_24767,N_24324,N_24291);
and U24768 (N_24768,N_24368,N_24486);
nand U24769 (N_24769,N_24372,N_24548);
xnor U24770 (N_24770,N_24490,N_24530);
nor U24771 (N_24771,N_24045,N_24106);
or U24772 (N_24772,N_24317,N_24219);
or U24773 (N_24773,N_24428,N_24350);
and U24774 (N_24774,N_24330,N_24331);
and U24775 (N_24775,N_24119,N_24504);
and U24776 (N_24776,N_24237,N_24360);
nor U24777 (N_24777,N_24183,N_24211);
or U24778 (N_24778,N_24032,N_24485);
xnor U24779 (N_24779,N_24514,N_24310);
xor U24780 (N_24780,N_24159,N_24353);
and U24781 (N_24781,N_24277,N_24345);
nor U24782 (N_24782,N_24394,N_24221);
or U24783 (N_24783,N_24188,N_24141);
and U24784 (N_24784,N_24586,N_24027);
nand U24785 (N_24785,N_24089,N_24199);
or U24786 (N_24786,N_24285,N_24305);
and U24787 (N_24787,N_24573,N_24223);
nand U24788 (N_24788,N_24154,N_24389);
or U24789 (N_24789,N_24432,N_24398);
xnor U24790 (N_24790,N_24487,N_24163);
and U24791 (N_24791,N_24058,N_24105);
nand U24792 (N_24792,N_24550,N_24451);
nor U24793 (N_24793,N_24028,N_24210);
nand U24794 (N_24794,N_24100,N_24265);
and U24795 (N_24795,N_24489,N_24217);
nor U24796 (N_24796,N_24344,N_24233);
and U24797 (N_24797,N_24408,N_24332);
xnor U24798 (N_24798,N_24299,N_24340);
or U24799 (N_24799,N_24361,N_24583);
or U24800 (N_24800,N_24181,N_24021);
nand U24801 (N_24801,N_24593,N_24467);
nor U24802 (N_24802,N_24405,N_24193);
xor U24803 (N_24803,N_24035,N_24547);
xor U24804 (N_24804,N_24288,N_24452);
or U24805 (N_24805,N_24020,N_24198);
or U24806 (N_24806,N_24137,N_24333);
nor U24807 (N_24807,N_24063,N_24076);
nor U24808 (N_24808,N_24241,N_24017);
or U24809 (N_24809,N_24097,N_24180);
xnor U24810 (N_24810,N_24328,N_24311);
nor U24811 (N_24811,N_24496,N_24234);
nand U24812 (N_24812,N_24144,N_24587);
nand U24813 (N_24813,N_24413,N_24347);
nand U24814 (N_24814,N_24545,N_24172);
nand U24815 (N_24815,N_24061,N_24365);
nand U24816 (N_24816,N_24030,N_24031);
nand U24817 (N_24817,N_24348,N_24584);
nor U24818 (N_24818,N_24282,N_24454);
xor U24819 (N_24819,N_24498,N_24167);
or U24820 (N_24820,N_24006,N_24131);
nor U24821 (N_24821,N_24390,N_24067);
or U24822 (N_24822,N_24579,N_24133);
nor U24823 (N_24823,N_24578,N_24060);
nand U24824 (N_24824,N_24177,N_24120);
nor U24825 (N_24825,N_24056,N_24436);
or U24826 (N_24826,N_24146,N_24173);
or U24827 (N_24827,N_24471,N_24533);
xnor U24828 (N_24828,N_24207,N_24537);
nand U24829 (N_24829,N_24477,N_24170);
nor U24830 (N_24830,N_24093,N_24138);
and U24831 (N_24831,N_24111,N_24266);
nor U24832 (N_24832,N_24228,N_24081);
xnor U24833 (N_24833,N_24236,N_24472);
or U24834 (N_24834,N_24588,N_24465);
or U24835 (N_24835,N_24469,N_24438);
nand U24836 (N_24836,N_24243,N_24064);
nor U24837 (N_24837,N_24476,N_24362);
nand U24838 (N_24838,N_24409,N_24222);
xor U24839 (N_24839,N_24499,N_24175);
and U24840 (N_24840,N_24369,N_24216);
nor U24841 (N_24841,N_24526,N_24415);
nor U24842 (N_24842,N_24397,N_24541);
xnor U24843 (N_24843,N_24005,N_24532);
nor U24844 (N_24844,N_24272,N_24110);
nor U24845 (N_24845,N_24598,N_24356);
nor U24846 (N_24846,N_24342,N_24375);
xor U24847 (N_24847,N_24036,N_24116);
nor U24848 (N_24848,N_24407,N_24126);
or U24849 (N_24849,N_24205,N_24261);
nor U24850 (N_24850,N_24393,N_24568);
or U24851 (N_24851,N_24098,N_24134);
nand U24852 (N_24852,N_24215,N_24037);
nor U24853 (N_24853,N_24254,N_24231);
nor U24854 (N_24854,N_24464,N_24555);
nor U24855 (N_24855,N_24075,N_24155);
nor U24856 (N_24856,N_24334,N_24572);
nand U24857 (N_24857,N_24396,N_24260);
nand U24858 (N_24858,N_24239,N_24419);
xor U24859 (N_24859,N_24038,N_24294);
or U24860 (N_24860,N_24466,N_24544);
nand U24861 (N_24861,N_24520,N_24204);
xnor U24862 (N_24862,N_24502,N_24057);
and U24863 (N_24863,N_24184,N_24165);
xnor U24864 (N_24864,N_24142,N_24101);
nor U24865 (N_24865,N_24220,N_24268);
nand U24866 (N_24866,N_24208,N_24418);
or U24867 (N_24867,N_24014,N_24244);
nand U24868 (N_24868,N_24596,N_24495);
xnor U24869 (N_24869,N_24493,N_24497);
nor U24870 (N_24870,N_24416,N_24325);
xnor U24871 (N_24871,N_24318,N_24326);
nor U24872 (N_24872,N_24086,N_24123);
nand U24873 (N_24873,N_24468,N_24592);
xor U24874 (N_24874,N_24047,N_24044);
xnor U24875 (N_24875,N_24143,N_24287);
and U24876 (N_24876,N_24491,N_24508);
xnor U24877 (N_24877,N_24160,N_24518);
nor U24878 (N_24878,N_24383,N_24308);
nor U24879 (N_24879,N_24563,N_24505);
or U24880 (N_24880,N_24414,N_24024);
nor U24881 (N_24881,N_24422,N_24189);
nand U24882 (N_24882,N_24200,N_24140);
nand U24883 (N_24883,N_24376,N_24099);
and U24884 (N_24884,N_24051,N_24501);
xnor U24885 (N_24885,N_24506,N_24384);
nor U24886 (N_24886,N_24182,N_24073);
xor U24887 (N_24887,N_24009,N_24275);
or U24888 (N_24888,N_24041,N_24417);
nor U24889 (N_24889,N_24315,N_24492);
xnor U24890 (N_24890,N_24002,N_24373);
xor U24891 (N_24891,N_24539,N_24192);
or U24892 (N_24892,N_24158,N_24571);
nand U24893 (N_24893,N_24301,N_24456);
nor U24894 (N_24894,N_24232,N_24218);
xor U24895 (N_24895,N_24048,N_24500);
and U24896 (N_24896,N_24388,N_24169);
and U24897 (N_24897,N_24103,N_24136);
nand U24898 (N_24898,N_24043,N_24214);
xor U24899 (N_24899,N_24186,N_24349);
and U24900 (N_24900,N_24407,N_24403);
and U24901 (N_24901,N_24319,N_24087);
or U24902 (N_24902,N_24160,N_24488);
nand U24903 (N_24903,N_24082,N_24465);
and U24904 (N_24904,N_24084,N_24257);
nand U24905 (N_24905,N_24419,N_24442);
nand U24906 (N_24906,N_24562,N_24338);
nand U24907 (N_24907,N_24387,N_24141);
and U24908 (N_24908,N_24089,N_24309);
or U24909 (N_24909,N_24207,N_24108);
nand U24910 (N_24910,N_24040,N_24533);
and U24911 (N_24911,N_24094,N_24220);
nand U24912 (N_24912,N_24212,N_24514);
or U24913 (N_24913,N_24595,N_24563);
nand U24914 (N_24914,N_24194,N_24498);
and U24915 (N_24915,N_24408,N_24480);
nor U24916 (N_24916,N_24499,N_24246);
or U24917 (N_24917,N_24549,N_24216);
nor U24918 (N_24918,N_24221,N_24561);
or U24919 (N_24919,N_24367,N_24135);
xnor U24920 (N_24920,N_24268,N_24125);
nor U24921 (N_24921,N_24339,N_24366);
nand U24922 (N_24922,N_24591,N_24099);
xor U24923 (N_24923,N_24088,N_24007);
or U24924 (N_24924,N_24529,N_24286);
or U24925 (N_24925,N_24241,N_24327);
nand U24926 (N_24926,N_24165,N_24001);
xnor U24927 (N_24927,N_24251,N_24401);
nand U24928 (N_24928,N_24352,N_24001);
xor U24929 (N_24929,N_24301,N_24371);
xnor U24930 (N_24930,N_24025,N_24496);
nor U24931 (N_24931,N_24570,N_24112);
or U24932 (N_24932,N_24427,N_24011);
nor U24933 (N_24933,N_24074,N_24551);
or U24934 (N_24934,N_24100,N_24385);
or U24935 (N_24935,N_24593,N_24085);
nor U24936 (N_24936,N_24035,N_24490);
nor U24937 (N_24937,N_24327,N_24212);
or U24938 (N_24938,N_24379,N_24594);
nand U24939 (N_24939,N_24188,N_24115);
xnor U24940 (N_24940,N_24281,N_24320);
xor U24941 (N_24941,N_24283,N_24356);
or U24942 (N_24942,N_24166,N_24331);
nand U24943 (N_24943,N_24351,N_24364);
nand U24944 (N_24944,N_24296,N_24381);
nor U24945 (N_24945,N_24306,N_24211);
and U24946 (N_24946,N_24373,N_24237);
and U24947 (N_24947,N_24074,N_24243);
and U24948 (N_24948,N_24233,N_24508);
and U24949 (N_24949,N_24228,N_24052);
and U24950 (N_24950,N_24500,N_24454);
and U24951 (N_24951,N_24327,N_24540);
xnor U24952 (N_24952,N_24151,N_24044);
or U24953 (N_24953,N_24196,N_24206);
or U24954 (N_24954,N_24080,N_24188);
and U24955 (N_24955,N_24335,N_24246);
xor U24956 (N_24956,N_24203,N_24412);
or U24957 (N_24957,N_24477,N_24400);
nand U24958 (N_24958,N_24532,N_24389);
xor U24959 (N_24959,N_24494,N_24386);
and U24960 (N_24960,N_24334,N_24543);
and U24961 (N_24961,N_24147,N_24481);
nor U24962 (N_24962,N_24072,N_24391);
nor U24963 (N_24963,N_24221,N_24408);
or U24964 (N_24964,N_24226,N_24019);
nand U24965 (N_24965,N_24455,N_24237);
or U24966 (N_24966,N_24217,N_24417);
nand U24967 (N_24967,N_24211,N_24421);
or U24968 (N_24968,N_24186,N_24374);
nand U24969 (N_24969,N_24317,N_24326);
or U24970 (N_24970,N_24535,N_24439);
nand U24971 (N_24971,N_24015,N_24503);
nand U24972 (N_24972,N_24527,N_24080);
and U24973 (N_24973,N_24516,N_24463);
xor U24974 (N_24974,N_24381,N_24044);
and U24975 (N_24975,N_24346,N_24189);
xor U24976 (N_24976,N_24420,N_24100);
xnor U24977 (N_24977,N_24224,N_24377);
and U24978 (N_24978,N_24428,N_24554);
nor U24979 (N_24979,N_24284,N_24578);
xor U24980 (N_24980,N_24510,N_24219);
or U24981 (N_24981,N_24464,N_24429);
nand U24982 (N_24982,N_24299,N_24288);
nand U24983 (N_24983,N_24326,N_24569);
nand U24984 (N_24984,N_24135,N_24145);
or U24985 (N_24985,N_24374,N_24206);
xor U24986 (N_24986,N_24277,N_24067);
or U24987 (N_24987,N_24268,N_24017);
and U24988 (N_24988,N_24305,N_24045);
nand U24989 (N_24989,N_24347,N_24436);
xor U24990 (N_24990,N_24528,N_24532);
and U24991 (N_24991,N_24094,N_24018);
xnor U24992 (N_24992,N_24047,N_24099);
xnor U24993 (N_24993,N_24284,N_24421);
or U24994 (N_24994,N_24594,N_24034);
and U24995 (N_24995,N_24185,N_24449);
xnor U24996 (N_24996,N_24015,N_24336);
or U24997 (N_24997,N_24598,N_24411);
and U24998 (N_24998,N_24075,N_24442);
xor U24999 (N_24999,N_24565,N_24507);
and U25000 (N_25000,N_24184,N_24063);
xor U25001 (N_25001,N_24382,N_24400);
xnor U25002 (N_25002,N_24070,N_24374);
xor U25003 (N_25003,N_24007,N_24328);
and U25004 (N_25004,N_24417,N_24228);
nand U25005 (N_25005,N_24178,N_24458);
nand U25006 (N_25006,N_24237,N_24106);
nand U25007 (N_25007,N_24242,N_24339);
and U25008 (N_25008,N_24360,N_24344);
or U25009 (N_25009,N_24479,N_24394);
or U25010 (N_25010,N_24454,N_24309);
xnor U25011 (N_25011,N_24488,N_24231);
xor U25012 (N_25012,N_24226,N_24410);
nor U25013 (N_25013,N_24386,N_24472);
nor U25014 (N_25014,N_24472,N_24218);
or U25015 (N_25015,N_24565,N_24281);
xor U25016 (N_25016,N_24376,N_24378);
nand U25017 (N_25017,N_24303,N_24068);
nor U25018 (N_25018,N_24462,N_24461);
or U25019 (N_25019,N_24106,N_24498);
and U25020 (N_25020,N_24110,N_24075);
and U25021 (N_25021,N_24471,N_24182);
xnor U25022 (N_25022,N_24424,N_24162);
nor U25023 (N_25023,N_24084,N_24356);
nand U25024 (N_25024,N_24316,N_24140);
nor U25025 (N_25025,N_24297,N_24547);
nor U25026 (N_25026,N_24189,N_24238);
xor U25027 (N_25027,N_24052,N_24363);
and U25028 (N_25028,N_24227,N_24104);
nand U25029 (N_25029,N_24399,N_24448);
nand U25030 (N_25030,N_24546,N_24397);
and U25031 (N_25031,N_24035,N_24034);
nand U25032 (N_25032,N_24220,N_24339);
nor U25033 (N_25033,N_24591,N_24364);
and U25034 (N_25034,N_24225,N_24357);
nand U25035 (N_25035,N_24291,N_24243);
nor U25036 (N_25036,N_24178,N_24078);
xnor U25037 (N_25037,N_24329,N_24518);
or U25038 (N_25038,N_24314,N_24021);
nor U25039 (N_25039,N_24410,N_24258);
nor U25040 (N_25040,N_24121,N_24327);
nor U25041 (N_25041,N_24024,N_24538);
and U25042 (N_25042,N_24279,N_24025);
xor U25043 (N_25043,N_24011,N_24018);
xnor U25044 (N_25044,N_24328,N_24096);
and U25045 (N_25045,N_24524,N_24248);
and U25046 (N_25046,N_24244,N_24549);
and U25047 (N_25047,N_24177,N_24574);
nor U25048 (N_25048,N_24578,N_24254);
nand U25049 (N_25049,N_24509,N_24189);
and U25050 (N_25050,N_24370,N_24354);
nor U25051 (N_25051,N_24092,N_24049);
and U25052 (N_25052,N_24239,N_24010);
nor U25053 (N_25053,N_24088,N_24312);
nor U25054 (N_25054,N_24519,N_24530);
nor U25055 (N_25055,N_24244,N_24440);
nor U25056 (N_25056,N_24132,N_24415);
xor U25057 (N_25057,N_24149,N_24477);
and U25058 (N_25058,N_24120,N_24465);
or U25059 (N_25059,N_24501,N_24117);
nand U25060 (N_25060,N_24420,N_24150);
xnor U25061 (N_25061,N_24396,N_24174);
xor U25062 (N_25062,N_24333,N_24082);
or U25063 (N_25063,N_24417,N_24528);
and U25064 (N_25064,N_24596,N_24557);
nand U25065 (N_25065,N_24160,N_24366);
or U25066 (N_25066,N_24487,N_24309);
or U25067 (N_25067,N_24479,N_24057);
and U25068 (N_25068,N_24207,N_24490);
nor U25069 (N_25069,N_24326,N_24510);
xor U25070 (N_25070,N_24041,N_24093);
nor U25071 (N_25071,N_24529,N_24206);
nand U25072 (N_25072,N_24029,N_24317);
and U25073 (N_25073,N_24202,N_24434);
nor U25074 (N_25074,N_24058,N_24253);
xnor U25075 (N_25075,N_24436,N_24071);
nor U25076 (N_25076,N_24356,N_24168);
nand U25077 (N_25077,N_24497,N_24389);
and U25078 (N_25078,N_24366,N_24154);
and U25079 (N_25079,N_24134,N_24036);
nor U25080 (N_25080,N_24151,N_24244);
nor U25081 (N_25081,N_24326,N_24359);
xor U25082 (N_25082,N_24216,N_24201);
nand U25083 (N_25083,N_24296,N_24542);
nand U25084 (N_25084,N_24169,N_24341);
or U25085 (N_25085,N_24546,N_24336);
or U25086 (N_25086,N_24490,N_24465);
nor U25087 (N_25087,N_24271,N_24240);
and U25088 (N_25088,N_24079,N_24053);
nor U25089 (N_25089,N_24521,N_24302);
nand U25090 (N_25090,N_24501,N_24394);
nand U25091 (N_25091,N_24083,N_24556);
or U25092 (N_25092,N_24591,N_24386);
xor U25093 (N_25093,N_24137,N_24274);
nor U25094 (N_25094,N_24026,N_24585);
and U25095 (N_25095,N_24527,N_24538);
nand U25096 (N_25096,N_24169,N_24567);
and U25097 (N_25097,N_24160,N_24410);
xnor U25098 (N_25098,N_24000,N_24053);
xnor U25099 (N_25099,N_24145,N_24151);
xnor U25100 (N_25100,N_24308,N_24481);
or U25101 (N_25101,N_24007,N_24122);
nor U25102 (N_25102,N_24145,N_24085);
nand U25103 (N_25103,N_24479,N_24329);
or U25104 (N_25104,N_24360,N_24200);
or U25105 (N_25105,N_24079,N_24178);
nor U25106 (N_25106,N_24403,N_24108);
xor U25107 (N_25107,N_24115,N_24260);
nor U25108 (N_25108,N_24391,N_24000);
nor U25109 (N_25109,N_24237,N_24047);
xnor U25110 (N_25110,N_24535,N_24105);
and U25111 (N_25111,N_24131,N_24411);
and U25112 (N_25112,N_24270,N_24423);
xor U25113 (N_25113,N_24492,N_24159);
nor U25114 (N_25114,N_24383,N_24194);
nand U25115 (N_25115,N_24297,N_24592);
nor U25116 (N_25116,N_24455,N_24340);
xnor U25117 (N_25117,N_24115,N_24598);
xor U25118 (N_25118,N_24329,N_24355);
nand U25119 (N_25119,N_24428,N_24361);
nand U25120 (N_25120,N_24513,N_24532);
nor U25121 (N_25121,N_24595,N_24478);
xnor U25122 (N_25122,N_24408,N_24326);
or U25123 (N_25123,N_24109,N_24316);
xor U25124 (N_25124,N_24092,N_24132);
or U25125 (N_25125,N_24368,N_24323);
xnor U25126 (N_25126,N_24415,N_24340);
and U25127 (N_25127,N_24325,N_24333);
nand U25128 (N_25128,N_24420,N_24396);
nor U25129 (N_25129,N_24365,N_24431);
or U25130 (N_25130,N_24445,N_24424);
and U25131 (N_25131,N_24556,N_24333);
nor U25132 (N_25132,N_24373,N_24503);
or U25133 (N_25133,N_24543,N_24056);
or U25134 (N_25134,N_24044,N_24476);
or U25135 (N_25135,N_24271,N_24244);
xor U25136 (N_25136,N_24107,N_24382);
nor U25137 (N_25137,N_24311,N_24326);
xnor U25138 (N_25138,N_24516,N_24069);
xnor U25139 (N_25139,N_24216,N_24270);
or U25140 (N_25140,N_24284,N_24218);
and U25141 (N_25141,N_24420,N_24033);
xor U25142 (N_25142,N_24567,N_24204);
nand U25143 (N_25143,N_24059,N_24338);
and U25144 (N_25144,N_24181,N_24341);
nand U25145 (N_25145,N_24121,N_24036);
or U25146 (N_25146,N_24551,N_24220);
xnor U25147 (N_25147,N_24127,N_24368);
nand U25148 (N_25148,N_24322,N_24249);
and U25149 (N_25149,N_24076,N_24582);
nor U25150 (N_25150,N_24396,N_24118);
xnor U25151 (N_25151,N_24195,N_24135);
nand U25152 (N_25152,N_24449,N_24194);
or U25153 (N_25153,N_24397,N_24491);
xnor U25154 (N_25154,N_24233,N_24253);
xnor U25155 (N_25155,N_24338,N_24560);
and U25156 (N_25156,N_24154,N_24045);
and U25157 (N_25157,N_24105,N_24468);
and U25158 (N_25158,N_24096,N_24204);
nor U25159 (N_25159,N_24155,N_24144);
or U25160 (N_25160,N_24320,N_24491);
and U25161 (N_25161,N_24366,N_24179);
nor U25162 (N_25162,N_24181,N_24314);
nand U25163 (N_25163,N_24319,N_24269);
nor U25164 (N_25164,N_24306,N_24551);
and U25165 (N_25165,N_24007,N_24323);
nand U25166 (N_25166,N_24385,N_24019);
and U25167 (N_25167,N_24014,N_24004);
and U25168 (N_25168,N_24532,N_24138);
nor U25169 (N_25169,N_24508,N_24410);
nor U25170 (N_25170,N_24236,N_24517);
and U25171 (N_25171,N_24052,N_24044);
nor U25172 (N_25172,N_24446,N_24584);
xor U25173 (N_25173,N_24583,N_24109);
and U25174 (N_25174,N_24401,N_24100);
nor U25175 (N_25175,N_24436,N_24099);
and U25176 (N_25176,N_24077,N_24307);
and U25177 (N_25177,N_24327,N_24329);
nand U25178 (N_25178,N_24183,N_24100);
nand U25179 (N_25179,N_24409,N_24270);
nor U25180 (N_25180,N_24495,N_24090);
nand U25181 (N_25181,N_24518,N_24041);
nor U25182 (N_25182,N_24556,N_24541);
xnor U25183 (N_25183,N_24526,N_24051);
and U25184 (N_25184,N_24213,N_24363);
nand U25185 (N_25185,N_24428,N_24038);
nand U25186 (N_25186,N_24021,N_24151);
nand U25187 (N_25187,N_24589,N_24155);
and U25188 (N_25188,N_24571,N_24273);
and U25189 (N_25189,N_24291,N_24203);
nor U25190 (N_25190,N_24106,N_24249);
and U25191 (N_25191,N_24554,N_24409);
nand U25192 (N_25192,N_24081,N_24364);
and U25193 (N_25193,N_24034,N_24093);
or U25194 (N_25194,N_24206,N_24174);
or U25195 (N_25195,N_24204,N_24338);
nand U25196 (N_25196,N_24168,N_24279);
or U25197 (N_25197,N_24411,N_24082);
xnor U25198 (N_25198,N_24424,N_24150);
and U25199 (N_25199,N_24222,N_24344);
or U25200 (N_25200,N_25066,N_24619);
nor U25201 (N_25201,N_25037,N_24663);
or U25202 (N_25202,N_25070,N_25079);
nand U25203 (N_25203,N_24734,N_24904);
or U25204 (N_25204,N_24882,N_24810);
and U25205 (N_25205,N_25198,N_24608);
nor U25206 (N_25206,N_24961,N_24789);
xnor U25207 (N_25207,N_25188,N_25185);
nor U25208 (N_25208,N_25102,N_25101);
nor U25209 (N_25209,N_24714,N_25116);
xor U25210 (N_25210,N_24696,N_25058);
or U25211 (N_25211,N_24707,N_25056);
and U25212 (N_25212,N_24912,N_24960);
xor U25213 (N_25213,N_25089,N_24713);
nand U25214 (N_25214,N_24623,N_25153);
nor U25215 (N_25215,N_24809,N_25014);
nand U25216 (N_25216,N_24895,N_24824);
xor U25217 (N_25217,N_25197,N_24800);
xor U25218 (N_25218,N_24692,N_24931);
or U25219 (N_25219,N_24651,N_24614);
nor U25220 (N_25220,N_25118,N_24637);
or U25221 (N_25221,N_24954,N_25146);
nor U25222 (N_25222,N_24851,N_24730);
or U25223 (N_25223,N_25176,N_25168);
nor U25224 (N_25224,N_24698,N_24990);
xnor U25225 (N_25225,N_24673,N_24924);
and U25226 (N_25226,N_24729,N_24820);
or U25227 (N_25227,N_24903,N_25020);
and U25228 (N_25228,N_24976,N_25167);
or U25229 (N_25229,N_24836,N_24963);
nand U25230 (N_25230,N_25055,N_25155);
or U25231 (N_25231,N_24622,N_24975);
xor U25232 (N_25232,N_25039,N_24926);
or U25233 (N_25233,N_24704,N_24878);
nand U25234 (N_25234,N_24909,N_24812);
nor U25235 (N_25235,N_24712,N_24934);
xor U25236 (N_25236,N_24965,N_25002);
nand U25237 (N_25237,N_24756,N_24879);
and U25238 (N_25238,N_25011,N_24833);
nor U25239 (N_25239,N_25027,N_24765);
xnor U25240 (N_25240,N_25144,N_25163);
xor U25241 (N_25241,N_24877,N_24773);
or U25242 (N_25242,N_25162,N_24735);
xnor U25243 (N_25243,N_25126,N_24847);
nor U25244 (N_25244,N_25145,N_24936);
or U25245 (N_25245,N_24659,N_24636);
or U25246 (N_25246,N_24641,N_25080);
xor U25247 (N_25247,N_25022,N_24604);
and U25248 (N_25248,N_24726,N_25179);
nand U25249 (N_25249,N_24840,N_24950);
nor U25250 (N_25250,N_24980,N_24806);
xnor U25251 (N_25251,N_25125,N_24617);
and U25252 (N_25252,N_24937,N_25029);
or U25253 (N_25253,N_24690,N_24889);
xnor U25254 (N_25254,N_24921,N_24603);
nand U25255 (N_25255,N_24817,N_24791);
nor U25256 (N_25256,N_24630,N_24670);
and U25257 (N_25257,N_24660,N_25184);
nor U25258 (N_25258,N_24830,N_25105);
or U25259 (N_25259,N_24941,N_24816);
nand U25260 (N_25260,N_24994,N_24664);
and U25261 (N_25261,N_25087,N_24741);
nand U25262 (N_25262,N_24762,N_24688);
or U25263 (N_25263,N_25030,N_24635);
or U25264 (N_25264,N_24891,N_24790);
nand U25265 (N_25265,N_25062,N_24991);
nand U25266 (N_25266,N_24866,N_25104);
nand U25267 (N_25267,N_25128,N_25034);
and U25268 (N_25268,N_24613,N_24780);
and U25269 (N_25269,N_24881,N_24600);
and U25270 (N_25270,N_25000,N_24747);
nor U25271 (N_25271,N_24658,N_24985);
or U25272 (N_25272,N_24753,N_24802);
or U25273 (N_25273,N_24843,N_24986);
or U25274 (N_25274,N_25007,N_25004);
nor U25275 (N_25275,N_24988,N_24621);
or U25276 (N_25276,N_25041,N_24942);
or U25277 (N_25277,N_24971,N_24788);
nand U25278 (N_25278,N_24702,N_25068);
nor U25279 (N_25279,N_25161,N_25077);
nand U25280 (N_25280,N_24770,N_25067);
and U25281 (N_25281,N_24952,N_25152);
nor U25282 (N_25282,N_24998,N_24737);
or U25283 (N_25283,N_24957,N_24871);
nand U25284 (N_25284,N_25107,N_24855);
or U25285 (N_25285,N_24606,N_25008);
xnor U25286 (N_25286,N_25016,N_25012);
and U25287 (N_25287,N_24811,N_25138);
nand U25288 (N_25288,N_25129,N_24846);
or U25289 (N_25289,N_24913,N_24687);
xnor U25290 (N_25290,N_25042,N_24757);
nor U25291 (N_25291,N_24739,N_24805);
nor U25292 (N_25292,N_25098,N_24849);
or U25293 (N_25293,N_24798,N_24629);
and U25294 (N_25294,N_24911,N_25090);
nor U25295 (N_25295,N_25048,N_24727);
nor U25296 (N_25296,N_24640,N_24672);
nor U25297 (N_25297,N_24873,N_24825);
xnor U25298 (N_25298,N_24697,N_25114);
nor U25299 (N_25299,N_24869,N_24939);
xor U25300 (N_25300,N_24905,N_24923);
xor U25301 (N_25301,N_24888,N_24868);
xor U25302 (N_25302,N_25151,N_24933);
or U25303 (N_25303,N_24894,N_24793);
nand U25304 (N_25304,N_25021,N_25033);
nand U25305 (N_25305,N_24804,N_24943);
or U25306 (N_25306,N_25172,N_25137);
nor U25307 (N_25307,N_24842,N_24738);
nand U25308 (N_25308,N_25071,N_24815);
nor U25309 (N_25309,N_25109,N_24981);
nand U25310 (N_25310,N_24918,N_25018);
and U25311 (N_25311,N_24654,N_24951);
or U25312 (N_25312,N_25001,N_25143);
and U25313 (N_25313,N_25028,N_24979);
nand U25314 (N_25314,N_25149,N_24611);
nand U25315 (N_25315,N_25133,N_24758);
or U25316 (N_25316,N_25053,N_24845);
or U25317 (N_25317,N_24661,N_24844);
xor U25318 (N_25318,N_25113,N_25178);
or U25319 (N_25319,N_24930,N_24643);
nor U25320 (N_25320,N_24677,N_24656);
nor U25321 (N_25321,N_24982,N_24748);
or U25322 (N_25322,N_24970,N_24625);
xnor U25323 (N_25323,N_24801,N_24733);
or U25324 (N_25324,N_25026,N_24813);
nor U25325 (N_25325,N_24919,N_25106);
nor U25326 (N_25326,N_24665,N_25192);
nand U25327 (N_25327,N_24745,N_25078);
xnor U25328 (N_25328,N_24620,N_25032);
nor U25329 (N_25329,N_24647,N_25196);
nand U25330 (N_25330,N_24685,N_25040);
nand U25331 (N_25331,N_25047,N_24728);
or U25332 (N_25332,N_24646,N_25072);
nor U25333 (N_25333,N_25199,N_24794);
nor U25334 (N_25334,N_25023,N_25076);
xnor U25335 (N_25335,N_24666,N_24967);
and U25336 (N_25336,N_24995,N_24610);
nand U25337 (N_25337,N_25009,N_24964);
nor U25338 (N_25338,N_24870,N_24779);
nand U25339 (N_25339,N_24837,N_24675);
or U25340 (N_25340,N_24819,N_24821);
xnor U25341 (N_25341,N_24972,N_24947);
nand U25342 (N_25342,N_24917,N_24907);
nand U25343 (N_25343,N_25132,N_24955);
xnor U25344 (N_25344,N_25181,N_25157);
or U25345 (N_25345,N_24743,N_25139);
nor U25346 (N_25346,N_25038,N_24683);
nand U25347 (N_25347,N_25054,N_25006);
xnor U25348 (N_25348,N_25065,N_24774);
and U25349 (N_25349,N_24694,N_25124);
nand U25350 (N_25350,N_25097,N_24814);
or U25351 (N_25351,N_24865,N_25010);
nand U25352 (N_25352,N_24719,N_24875);
xnor U25353 (N_25353,N_25088,N_24996);
or U25354 (N_25354,N_24902,N_24703);
xor U25355 (N_25355,N_24959,N_25131);
nor U25356 (N_25356,N_24786,N_24962);
xor U25357 (N_25357,N_24674,N_24874);
nand U25358 (N_25358,N_25050,N_25121);
nor U25359 (N_25359,N_24898,N_24772);
nand U25360 (N_25360,N_25082,N_25142);
nand U25361 (N_25361,N_25059,N_24648);
nand U25362 (N_25362,N_24792,N_24601);
nand U25363 (N_25363,N_24850,N_25094);
nor U25364 (N_25364,N_24668,N_24899);
and U25365 (N_25365,N_24634,N_25134);
nand U25366 (N_25366,N_24657,N_24910);
nand U25367 (N_25367,N_24796,N_25120);
nand U25368 (N_25368,N_25140,N_24827);
and U25369 (N_25369,N_25085,N_25069);
nor U25370 (N_25370,N_25110,N_24944);
or U25371 (N_25371,N_25193,N_24838);
or U25372 (N_25372,N_24607,N_25003);
xor U25373 (N_25373,N_25046,N_24626);
nand U25374 (N_25374,N_24859,N_25186);
or U25375 (N_25375,N_25074,N_24624);
and U25376 (N_25376,N_24858,N_24721);
nor U25377 (N_25377,N_24715,N_24771);
nand U25378 (N_25378,N_24615,N_25189);
or U25379 (N_25379,N_24750,N_25112);
nor U25380 (N_25380,N_24984,N_24890);
and U25381 (N_25381,N_24605,N_24686);
and U25382 (N_25382,N_25005,N_24983);
nor U25383 (N_25383,N_24612,N_24669);
and U25384 (N_25384,N_25130,N_25017);
and U25385 (N_25385,N_24808,N_25166);
or U25386 (N_25386,N_24650,N_25043);
and U25387 (N_25387,N_24725,N_24631);
or U25388 (N_25388,N_25063,N_24680);
nand U25389 (N_25389,N_24776,N_24736);
xnor U25390 (N_25390,N_24940,N_24928);
and U25391 (N_25391,N_24916,N_24681);
or U25392 (N_25392,N_24749,N_25064);
xnor U25393 (N_25393,N_25061,N_24723);
or U25394 (N_25394,N_24717,N_24992);
or U25395 (N_25395,N_24828,N_25148);
nand U25396 (N_25396,N_24925,N_24699);
xor U25397 (N_25397,N_24787,N_24627);
nor U25398 (N_25398,N_25092,N_24906);
xnor U25399 (N_25399,N_24766,N_24863);
nand U25400 (N_25400,N_25147,N_25180);
and U25401 (N_25401,N_25174,N_25191);
and U25402 (N_25402,N_24908,N_24807);
and U25403 (N_25403,N_24768,N_25057);
or U25404 (N_25404,N_25100,N_24989);
or U25405 (N_25405,N_25170,N_25159);
or U25406 (N_25406,N_24755,N_24900);
or U25407 (N_25407,N_25103,N_24977);
nor U25408 (N_25408,N_24958,N_25091);
or U25409 (N_25409,N_24649,N_24709);
nand U25410 (N_25410,N_24968,N_25171);
nand U25411 (N_25411,N_25177,N_24701);
nor U25412 (N_25412,N_24662,N_24775);
or U25413 (N_25413,N_24705,N_25084);
nand U25414 (N_25414,N_25035,N_24653);
or U25415 (N_25415,N_24782,N_24731);
xor U25416 (N_25416,N_24978,N_25169);
xor U25417 (N_25417,N_25096,N_25183);
nand U25418 (N_25418,N_24710,N_24880);
xnor U25419 (N_25419,N_24922,N_24896);
nor U25420 (N_25420,N_24915,N_24784);
nor U25421 (N_25421,N_24700,N_24974);
xor U25422 (N_25422,N_24831,N_24679);
xnor U25423 (N_25423,N_24883,N_24823);
xnor U25424 (N_25424,N_24632,N_24720);
nand U25425 (N_25425,N_24803,N_24876);
nor U25426 (N_25426,N_24864,N_25182);
and U25427 (N_25427,N_25086,N_24785);
xor U25428 (N_25428,N_25051,N_25013);
or U25429 (N_25429,N_25060,N_25164);
xnor U25430 (N_25430,N_24886,N_24693);
xnor U25431 (N_25431,N_24861,N_24832);
or U25432 (N_25432,N_24993,N_24752);
nand U25433 (N_25433,N_24848,N_24732);
nand U25434 (N_25434,N_24997,N_25025);
nand U25435 (N_25435,N_24781,N_25135);
nand U25436 (N_25436,N_24938,N_24602);
xnor U25437 (N_25437,N_24671,N_24638);
nor U25438 (N_25438,N_24763,N_24740);
nand U25439 (N_25439,N_25044,N_25127);
nand U25440 (N_25440,N_24724,N_24711);
nand U25441 (N_25441,N_24856,N_24744);
nand U25442 (N_25442,N_24797,N_24949);
xnor U25443 (N_25443,N_25175,N_24945);
and U25444 (N_25444,N_24678,N_24754);
nand U25445 (N_25445,N_24642,N_24948);
nor U25446 (N_25446,N_25052,N_24914);
nand U25447 (N_25447,N_24853,N_24872);
and U25448 (N_25448,N_24857,N_24822);
nand U25449 (N_25449,N_24682,N_25160);
or U25450 (N_25450,N_24655,N_24644);
or U25451 (N_25451,N_25108,N_24969);
nand U25452 (N_25452,N_24973,N_24718);
or U25453 (N_25453,N_24708,N_24778);
xor U25454 (N_25454,N_24829,N_24818);
or U25455 (N_25455,N_24893,N_24826);
xnor U25456 (N_25456,N_24633,N_24920);
nor U25457 (N_25457,N_24722,N_24783);
or U25458 (N_25458,N_24932,N_24751);
nand U25459 (N_25459,N_24764,N_25165);
and U25460 (N_25460,N_24706,N_24689);
nor U25461 (N_25461,N_24884,N_25117);
and U25462 (N_25462,N_24799,N_24953);
nor U25463 (N_25463,N_25075,N_24761);
nor U25464 (N_25464,N_24645,N_25036);
nor U25465 (N_25465,N_24862,N_24684);
or U25466 (N_25466,N_25154,N_24885);
xor U25467 (N_25467,N_25123,N_24927);
xnor U25468 (N_25468,N_24839,N_24854);
nand U25469 (N_25469,N_24652,N_24777);
and U25470 (N_25470,N_24795,N_24628);
xor U25471 (N_25471,N_24639,N_25115);
nand U25472 (N_25472,N_24691,N_24852);
and U25473 (N_25473,N_25031,N_25081);
or U25474 (N_25474,N_24746,N_25141);
nor U25475 (N_25475,N_24966,N_24860);
nand U25476 (N_25476,N_25095,N_25187);
and U25477 (N_25477,N_25019,N_24695);
nor U25478 (N_25478,N_24867,N_24892);
nor U25479 (N_25479,N_24716,N_24999);
and U25480 (N_25480,N_25111,N_25099);
or U25481 (N_25481,N_24667,N_24609);
xnor U25482 (N_25482,N_24956,N_24759);
nand U25483 (N_25483,N_25045,N_25015);
and U25484 (N_25484,N_24769,N_25093);
and U25485 (N_25485,N_25156,N_24834);
nor U25486 (N_25486,N_24616,N_25158);
or U25487 (N_25487,N_24742,N_24760);
nor U25488 (N_25488,N_25194,N_24767);
nor U25489 (N_25489,N_25073,N_24935);
or U25490 (N_25490,N_25049,N_24946);
or U25491 (N_25491,N_25122,N_25150);
and U25492 (N_25492,N_25024,N_24835);
and U25493 (N_25493,N_25190,N_24897);
nor U25494 (N_25494,N_25119,N_24618);
and U25495 (N_25495,N_24929,N_24887);
nor U25496 (N_25496,N_25083,N_24676);
nand U25497 (N_25497,N_24901,N_24987);
and U25498 (N_25498,N_24841,N_25173);
nand U25499 (N_25499,N_25195,N_25136);
xnor U25500 (N_25500,N_25179,N_24668);
and U25501 (N_25501,N_24968,N_24773);
or U25502 (N_25502,N_25172,N_24797);
xnor U25503 (N_25503,N_24615,N_25142);
xor U25504 (N_25504,N_25092,N_25115);
or U25505 (N_25505,N_24720,N_24608);
nand U25506 (N_25506,N_25017,N_25195);
or U25507 (N_25507,N_24951,N_24647);
nand U25508 (N_25508,N_24750,N_24749);
and U25509 (N_25509,N_24615,N_24678);
nor U25510 (N_25510,N_25065,N_25156);
xnor U25511 (N_25511,N_24953,N_24797);
and U25512 (N_25512,N_24929,N_25097);
xnor U25513 (N_25513,N_24755,N_25081);
or U25514 (N_25514,N_24780,N_24771);
xor U25515 (N_25515,N_24691,N_24896);
and U25516 (N_25516,N_25168,N_24792);
or U25517 (N_25517,N_25067,N_24806);
nor U25518 (N_25518,N_25007,N_24753);
and U25519 (N_25519,N_25077,N_24785);
xnor U25520 (N_25520,N_24879,N_24823);
and U25521 (N_25521,N_24962,N_24782);
nand U25522 (N_25522,N_24649,N_24853);
nor U25523 (N_25523,N_25012,N_24614);
and U25524 (N_25524,N_25138,N_24889);
nor U25525 (N_25525,N_24973,N_24830);
nor U25526 (N_25526,N_24968,N_25167);
or U25527 (N_25527,N_24800,N_24911);
nor U25528 (N_25528,N_24965,N_24981);
nor U25529 (N_25529,N_24609,N_24627);
xnor U25530 (N_25530,N_25088,N_24768);
and U25531 (N_25531,N_24916,N_24868);
or U25532 (N_25532,N_24646,N_24940);
nand U25533 (N_25533,N_24626,N_24854);
nor U25534 (N_25534,N_24933,N_24911);
xor U25535 (N_25535,N_24787,N_24836);
nor U25536 (N_25536,N_24659,N_25018);
or U25537 (N_25537,N_25065,N_25154);
nor U25538 (N_25538,N_25068,N_24686);
nand U25539 (N_25539,N_24603,N_25021);
xnor U25540 (N_25540,N_25086,N_24960);
and U25541 (N_25541,N_24635,N_25094);
nand U25542 (N_25542,N_25135,N_24653);
and U25543 (N_25543,N_24813,N_25028);
or U25544 (N_25544,N_24677,N_25050);
xnor U25545 (N_25545,N_24650,N_25153);
or U25546 (N_25546,N_25009,N_25186);
or U25547 (N_25547,N_24983,N_24666);
nor U25548 (N_25548,N_24969,N_24777);
nand U25549 (N_25549,N_25102,N_24620);
nand U25550 (N_25550,N_24669,N_24883);
or U25551 (N_25551,N_25025,N_24712);
xnor U25552 (N_25552,N_25012,N_24653);
nand U25553 (N_25553,N_25046,N_24680);
nand U25554 (N_25554,N_24638,N_24933);
or U25555 (N_25555,N_24723,N_24972);
xor U25556 (N_25556,N_24878,N_24967);
nand U25557 (N_25557,N_24823,N_24959);
or U25558 (N_25558,N_25135,N_25199);
or U25559 (N_25559,N_25193,N_25122);
nor U25560 (N_25560,N_25074,N_24726);
and U25561 (N_25561,N_24815,N_25085);
nor U25562 (N_25562,N_25007,N_25138);
nand U25563 (N_25563,N_24707,N_25052);
nor U25564 (N_25564,N_25145,N_24989);
xnor U25565 (N_25565,N_24729,N_24891);
or U25566 (N_25566,N_24813,N_25113);
nand U25567 (N_25567,N_24743,N_24982);
and U25568 (N_25568,N_25078,N_24961);
or U25569 (N_25569,N_24874,N_25173);
nand U25570 (N_25570,N_24729,N_25053);
nor U25571 (N_25571,N_24756,N_25144);
and U25572 (N_25572,N_24993,N_24687);
or U25573 (N_25573,N_24747,N_25106);
and U25574 (N_25574,N_24757,N_25013);
nand U25575 (N_25575,N_24849,N_24781);
nor U25576 (N_25576,N_24836,N_24732);
nand U25577 (N_25577,N_25141,N_24924);
nor U25578 (N_25578,N_24903,N_24671);
or U25579 (N_25579,N_24652,N_25007);
nor U25580 (N_25580,N_24919,N_25169);
nand U25581 (N_25581,N_24836,N_24617);
nand U25582 (N_25582,N_25051,N_24878);
nand U25583 (N_25583,N_24868,N_24650);
nand U25584 (N_25584,N_24759,N_24959);
xnor U25585 (N_25585,N_24897,N_25021);
xnor U25586 (N_25586,N_24796,N_24768);
nor U25587 (N_25587,N_25094,N_24735);
and U25588 (N_25588,N_24874,N_24826);
nor U25589 (N_25589,N_25014,N_24942);
nor U25590 (N_25590,N_24980,N_24669);
or U25591 (N_25591,N_25156,N_24912);
nand U25592 (N_25592,N_24640,N_24652);
nor U25593 (N_25593,N_24761,N_24723);
nor U25594 (N_25594,N_24724,N_25119);
or U25595 (N_25595,N_24678,N_24898);
and U25596 (N_25596,N_24807,N_24799);
nand U25597 (N_25597,N_24917,N_24830);
and U25598 (N_25598,N_25015,N_24731);
xor U25599 (N_25599,N_24724,N_24747);
nor U25600 (N_25600,N_24907,N_24799);
or U25601 (N_25601,N_24898,N_24846);
xor U25602 (N_25602,N_24786,N_24658);
xor U25603 (N_25603,N_24703,N_24942);
nor U25604 (N_25604,N_24655,N_24950);
xor U25605 (N_25605,N_24671,N_24705);
xnor U25606 (N_25606,N_24706,N_24787);
and U25607 (N_25607,N_25082,N_25137);
nor U25608 (N_25608,N_25006,N_25166);
and U25609 (N_25609,N_24860,N_24742);
and U25610 (N_25610,N_24641,N_25124);
xnor U25611 (N_25611,N_24950,N_24860);
nor U25612 (N_25612,N_25165,N_25022);
xor U25613 (N_25613,N_24938,N_25118);
nor U25614 (N_25614,N_24727,N_24621);
and U25615 (N_25615,N_25163,N_24652);
and U25616 (N_25616,N_24810,N_25199);
or U25617 (N_25617,N_24806,N_24772);
nand U25618 (N_25618,N_24738,N_24998);
and U25619 (N_25619,N_25006,N_24671);
and U25620 (N_25620,N_24967,N_25185);
xor U25621 (N_25621,N_24778,N_24709);
nand U25622 (N_25622,N_24952,N_25141);
or U25623 (N_25623,N_24899,N_25196);
nand U25624 (N_25624,N_24777,N_24885);
or U25625 (N_25625,N_24783,N_24601);
and U25626 (N_25626,N_24641,N_24873);
nand U25627 (N_25627,N_24622,N_24646);
xnor U25628 (N_25628,N_24620,N_24856);
or U25629 (N_25629,N_24991,N_24961);
or U25630 (N_25630,N_25180,N_24909);
nor U25631 (N_25631,N_25176,N_25040);
or U25632 (N_25632,N_25175,N_24908);
nand U25633 (N_25633,N_25178,N_25148);
and U25634 (N_25634,N_24832,N_25116);
and U25635 (N_25635,N_24694,N_24753);
and U25636 (N_25636,N_24740,N_24673);
or U25637 (N_25637,N_25124,N_24820);
nor U25638 (N_25638,N_25172,N_24823);
xor U25639 (N_25639,N_24780,N_25187);
and U25640 (N_25640,N_25053,N_24826);
or U25641 (N_25641,N_24949,N_24693);
nand U25642 (N_25642,N_24885,N_24816);
nor U25643 (N_25643,N_24746,N_25014);
nand U25644 (N_25644,N_24621,N_24923);
nand U25645 (N_25645,N_25024,N_25100);
nor U25646 (N_25646,N_24705,N_24644);
nor U25647 (N_25647,N_24709,N_24895);
or U25648 (N_25648,N_24848,N_24730);
and U25649 (N_25649,N_24792,N_24670);
nor U25650 (N_25650,N_24937,N_25039);
nor U25651 (N_25651,N_24723,N_24602);
or U25652 (N_25652,N_24662,N_24851);
and U25653 (N_25653,N_24679,N_25108);
xnor U25654 (N_25654,N_24613,N_24755);
xnor U25655 (N_25655,N_25130,N_24725);
nand U25656 (N_25656,N_24790,N_25020);
xor U25657 (N_25657,N_24636,N_24804);
nor U25658 (N_25658,N_25083,N_25041);
or U25659 (N_25659,N_24860,N_24969);
and U25660 (N_25660,N_24995,N_24979);
xor U25661 (N_25661,N_25064,N_24858);
nand U25662 (N_25662,N_24990,N_24702);
xnor U25663 (N_25663,N_24793,N_25058);
or U25664 (N_25664,N_24705,N_24953);
nand U25665 (N_25665,N_24866,N_24853);
nand U25666 (N_25666,N_24894,N_24647);
or U25667 (N_25667,N_24664,N_25019);
nand U25668 (N_25668,N_24759,N_24734);
nor U25669 (N_25669,N_24646,N_24790);
and U25670 (N_25670,N_24645,N_24630);
nor U25671 (N_25671,N_24788,N_25097);
or U25672 (N_25672,N_24637,N_24639);
or U25673 (N_25673,N_24641,N_24883);
or U25674 (N_25674,N_24742,N_24735);
and U25675 (N_25675,N_24853,N_25090);
and U25676 (N_25676,N_24750,N_25062);
and U25677 (N_25677,N_24658,N_24825);
and U25678 (N_25678,N_24775,N_25057);
and U25679 (N_25679,N_25045,N_24786);
nand U25680 (N_25680,N_24755,N_24790);
nand U25681 (N_25681,N_24882,N_25135);
or U25682 (N_25682,N_25074,N_25007);
nand U25683 (N_25683,N_24882,N_24846);
xnor U25684 (N_25684,N_25103,N_24838);
and U25685 (N_25685,N_24722,N_24704);
nand U25686 (N_25686,N_24643,N_24892);
or U25687 (N_25687,N_25055,N_24979);
and U25688 (N_25688,N_25003,N_24968);
xor U25689 (N_25689,N_24719,N_24972);
or U25690 (N_25690,N_24892,N_25102);
and U25691 (N_25691,N_24850,N_25010);
xor U25692 (N_25692,N_24981,N_24985);
nor U25693 (N_25693,N_24820,N_24928);
xor U25694 (N_25694,N_24716,N_25027);
or U25695 (N_25695,N_24814,N_25172);
and U25696 (N_25696,N_24728,N_24681);
xor U25697 (N_25697,N_24652,N_24712);
nand U25698 (N_25698,N_25180,N_24772);
nor U25699 (N_25699,N_24868,N_24636);
or U25700 (N_25700,N_24858,N_25073);
or U25701 (N_25701,N_24949,N_24787);
nor U25702 (N_25702,N_24737,N_25132);
or U25703 (N_25703,N_24846,N_24943);
nor U25704 (N_25704,N_24903,N_24851);
and U25705 (N_25705,N_25054,N_25110);
or U25706 (N_25706,N_24936,N_24713);
nor U25707 (N_25707,N_24747,N_24693);
or U25708 (N_25708,N_24935,N_24640);
and U25709 (N_25709,N_24718,N_24925);
xnor U25710 (N_25710,N_24845,N_24639);
nand U25711 (N_25711,N_24795,N_24717);
xor U25712 (N_25712,N_24684,N_24985);
or U25713 (N_25713,N_25104,N_24876);
nor U25714 (N_25714,N_24629,N_24747);
and U25715 (N_25715,N_24858,N_24868);
and U25716 (N_25716,N_24761,N_24603);
xnor U25717 (N_25717,N_24732,N_24703);
and U25718 (N_25718,N_24934,N_24844);
nand U25719 (N_25719,N_24901,N_24897);
or U25720 (N_25720,N_25147,N_24739);
xor U25721 (N_25721,N_24894,N_24877);
and U25722 (N_25722,N_25010,N_24699);
nand U25723 (N_25723,N_24908,N_24637);
nand U25724 (N_25724,N_25104,N_24853);
nor U25725 (N_25725,N_24701,N_25030);
nor U25726 (N_25726,N_25106,N_25119);
and U25727 (N_25727,N_25060,N_24736);
or U25728 (N_25728,N_24848,N_24955);
xor U25729 (N_25729,N_24846,N_24865);
or U25730 (N_25730,N_25114,N_25060);
or U25731 (N_25731,N_25141,N_24717);
nand U25732 (N_25732,N_24959,N_25094);
or U25733 (N_25733,N_25011,N_24868);
or U25734 (N_25734,N_24955,N_24711);
or U25735 (N_25735,N_24775,N_25077);
and U25736 (N_25736,N_24977,N_24897);
and U25737 (N_25737,N_24618,N_24742);
xnor U25738 (N_25738,N_24983,N_25139);
nor U25739 (N_25739,N_24721,N_24914);
or U25740 (N_25740,N_24924,N_24868);
or U25741 (N_25741,N_24925,N_24967);
nor U25742 (N_25742,N_24722,N_24675);
or U25743 (N_25743,N_25135,N_24648);
and U25744 (N_25744,N_24897,N_25048);
nor U25745 (N_25745,N_24982,N_25124);
nor U25746 (N_25746,N_24607,N_25114);
nand U25747 (N_25747,N_25165,N_25028);
and U25748 (N_25748,N_24648,N_24712);
and U25749 (N_25749,N_25048,N_25005);
and U25750 (N_25750,N_24732,N_24795);
nor U25751 (N_25751,N_24779,N_24962);
nand U25752 (N_25752,N_24866,N_24870);
nand U25753 (N_25753,N_25012,N_24984);
nand U25754 (N_25754,N_25151,N_24963);
xnor U25755 (N_25755,N_24644,N_24715);
nor U25756 (N_25756,N_24854,N_25130);
or U25757 (N_25757,N_24785,N_25040);
nand U25758 (N_25758,N_24769,N_24823);
nand U25759 (N_25759,N_24785,N_24846);
nand U25760 (N_25760,N_24705,N_24769);
nor U25761 (N_25761,N_25161,N_24869);
xnor U25762 (N_25762,N_25067,N_24650);
nand U25763 (N_25763,N_24923,N_24890);
or U25764 (N_25764,N_25169,N_25031);
or U25765 (N_25765,N_24603,N_24706);
and U25766 (N_25766,N_24820,N_24793);
nand U25767 (N_25767,N_24608,N_24780);
or U25768 (N_25768,N_25017,N_24722);
and U25769 (N_25769,N_25174,N_24711);
nor U25770 (N_25770,N_25095,N_24656);
xor U25771 (N_25771,N_24866,N_24633);
or U25772 (N_25772,N_24776,N_25126);
xnor U25773 (N_25773,N_24918,N_24889);
nand U25774 (N_25774,N_24658,N_25175);
or U25775 (N_25775,N_24792,N_25187);
xor U25776 (N_25776,N_25124,N_24876);
nand U25777 (N_25777,N_24950,N_24790);
and U25778 (N_25778,N_25071,N_24708);
and U25779 (N_25779,N_25147,N_25028);
nor U25780 (N_25780,N_25159,N_25114);
xor U25781 (N_25781,N_24672,N_24838);
and U25782 (N_25782,N_24929,N_24943);
and U25783 (N_25783,N_24866,N_25169);
or U25784 (N_25784,N_24807,N_24772);
xor U25785 (N_25785,N_24757,N_24936);
nor U25786 (N_25786,N_24893,N_24987);
and U25787 (N_25787,N_25001,N_25044);
or U25788 (N_25788,N_24935,N_24855);
nor U25789 (N_25789,N_24969,N_24867);
nor U25790 (N_25790,N_24808,N_25034);
and U25791 (N_25791,N_25028,N_24714);
or U25792 (N_25792,N_24651,N_24605);
nand U25793 (N_25793,N_25028,N_25094);
nand U25794 (N_25794,N_24953,N_24823);
nand U25795 (N_25795,N_25079,N_24916);
xor U25796 (N_25796,N_24777,N_24979);
and U25797 (N_25797,N_24715,N_24600);
and U25798 (N_25798,N_25123,N_25075);
xnor U25799 (N_25799,N_24883,N_24961);
xnor U25800 (N_25800,N_25354,N_25566);
and U25801 (N_25801,N_25383,N_25734);
xnor U25802 (N_25802,N_25272,N_25765);
xor U25803 (N_25803,N_25224,N_25527);
nand U25804 (N_25804,N_25664,N_25449);
nand U25805 (N_25805,N_25523,N_25200);
or U25806 (N_25806,N_25248,N_25752);
xnor U25807 (N_25807,N_25508,N_25243);
and U25808 (N_25808,N_25301,N_25751);
xor U25809 (N_25809,N_25220,N_25334);
xor U25810 (N_25810,N_25533,N_25766);
nor U25811 (N_25811,N_25281,N_25551);
nor U25812 (N_25812,N_25614,N_25625);
xor U25813 (N_25813,N_25704,N_25588);
or U25814 (N_25814,N_25306,N_25548);
nor U25815 (N_25815,N_25363,N_25410);
xnor U25816 (N_25816,N_25439,N_25634);
nor U25817 (N_25817,N_25484,N_25789);
xor U25818 (N_25818,N_25794,N_25706);
or U25819 (N_25819,N_25405,N_25639);
and U25820 (N_25820,N_25576,N_25416);
or U25821 (N_25821,N_25320,N_25528);
or U25822 (N_25822,N_25387,N_25604);
nor U25823 (N_25823,N_25650,N_25225);
nand U25824 (N_25824,N_25519,N_25744);
nand U25825 (N_25825,N_25412,N_25295);
nor U25826 (N_25826,N_25244,N_25502);
or U25827 (N_25827,N_25441,N_25228);
nand U25828 (N_25828,N_25382,N_25635);
or U25829 (N_25829,N_25356,N_25379);
xnor U25830 (N_25830,N_25791,N_25785);
and U25831 (N_25831,N_25471,N_25307);
and U25832 (N_25832,N_25649,N_25414);
and U25833 (N_25833,N_25485,N_25345);
xor U25834 (N_25834,N_25573,N_25761);
xor U25835 (N_25835,N_25384,N_25518);
or U25836 (N_25836,N_25556,N_25788);
and U25837 (N_25837,N_25386,N_25458);
and U25838 (N_25838,N_25696,N_25633);
or U25839 (N_25839,N_25343,N_25495);
xor U25840 (N_25840,N_25456,N_25310);
nor U25841 (N_25841,N_25487,N_25401);
xor U25842 (N_25842,N_25514,N_25593);
nand U25843 (N_25843,N_25462,N_25474);
nor U25844 (N_25844,N_25772,N_25698);
or U25845 (N_25845,N_25489,N_25231);
and U25846 (N_25846,N_25426,N_25715);
and U25847 (N_25847,N_25505,N_25746);
nand U25848 (N_25848,N_25669,N_25433);
xor U25849 (N_25849,N_25777,N_25648);
and U25850 (N_25850,N_25442,N_25799);
or U25851 (N_25851,N_25641,N_25452);
or U25852 (N_25852,N_25663,N_25233);
xnor U25853 (N_25853,N_25720,N_25685);
or U25854 (N_25854,N_25239,N_25705);
and U25855 (N_25855,N_25780,N_25718);
xnor U25856 (N_25856,N_25292,N_25303);
nor U25857 (N_25857,N_25795,N_25603);
nor U25858 (N_25858,N_25652,N_25411);
xnor U25859 (N_25859,N_25304,N_25376);
and U25860 (N_25860,N_25674,N_25309);
or U25861 (N_25861,N_25290,N_25355);
or U25862 (N_25862,N_25690,N_25438);
and U25863 (N_25863,N_25773,N_25755);
and U25864 (N_25864,N_25529,N_25672);
xor U25865 (N_25865,N_25359,N_25675);
xnor U25866 (N_25866,N_25557,N_25629);
xnor U25867 (N_25867,N_25268,N_25740);
nor U25868 (N_25868,N_25403,N_25291);
nand U25869 (N_25869,N_25296,N_25782);
nor U25870 (N_25870,N_25700,N_25432);
xor U25871 (N_25871,N_25476,N_25346);
or U25872 (N_25872,N_25217,N_25575);
and U25873 (N_25873,N_25367,N_25499);
nor U25874 (N_25874,N_25493,N_25360);
or U25875 (N_25875,N_25246,N_25400);
xor U25876 (N_25876,N_25714,N_25445);
nand U25877 (N_25877,N_25678,N_25455);
xnor U25878 (N_25878,N_25477,N_25627);
nor U25879 (N_25879,N_25786,N_25587);
or U25880 (N_25880,N_25257,N_25294);
nor U25881 (N_25881,N_25541,N_25424);
nor U25882 (N_25882,N_25347,N_25284);
xnor U25883 (N_25883,N_25707,N_25327);
nor U25884 (N_25884,N_25394,N_25776);
or U25885 (N_25885,N_25247,N_25375);
and U25886 (N_25886,N_25745,N_25601);
nand U25887 (N_25887,N_25270,N_25554);
nand U25888 (N_25888,N_25372,N_25645);
or U25889 (N_25889,N_25626,N_25380);
xnor U25890 (N_25890,N_25261,N_25699);
nand U25891 (N_25891,N_25723,N_25643);
or U25892 (N_25892,N_25368,N_25733);
or U25893 (N_25893,N_25205,N_25610);
or U25894 (N_25894,N_25646,N_25753);
nand U25895 (N_25895,N_25687,N_25222);
and U25896 (N_25896,N_25506,N_25511);
and U25897 (N_25897,N_25223,N_25275);
xnor U25898 (N_25898,N_25616,N_25313);
or U25899 (N_25899,N_25538,N_25448);
nor U25900 (N_25900,N_25407,N_25447);
nor U25901 (N_25901,N_25461,N_25336);
nand U25902 (N_25902,N_25312,N_25507);
nor U25903 (N_25903,N_25258,N_25749);
or U25904 (N_25904,N_25737,N_25622);
nand U25905 (N_25905,N_25662,N_25762);
or U25906 (N_25906,N_25280,N_25615);
nor U25907 (N_25907,N_25395,N_25774);
and U25908 (N_25908,N_25348,N_25337);
nand U25909 (N_25909,N_25708,N_25726);
and U25910 (N_25910,N_25206,N_25532);
or U25911 (N_25911,N_25605,N_25287);
nor U25912 (N_25912,N_25201,N_25742);
or U25913 (N_25913,N_25719,N_25311);
nand U25914 (N_25914,N_25586,N_25612);
and U25915 (N_25915,N_25637,N_25568);
and U25916 (N_25916,N_25415,N_25227);
xor U25917 (N_25917,N_25654,N_25567);
nand U25918 (N_25918,N_25325,N_25350);
or U25919 (N_25919,N_25323,N_25388);
nand U25920 (N_25920,N_25389,N_25322);
and U25921 (N_25921,N_25620,N_25249);
nand U25922 (N_25922,N_25565,N_25716);
or U25923 (N_25923,N_25450,N_25778);
nor U25924 (N_25924,N_25333,N_25743);
and U25925 (N_25925,N_25366,N_25331);
or U25926 (N_25926,N_25491,N_25202);
or U25927 (N_25927,N_25328,N_25624);
and U25928 (N_25928,N_25709,N_25404);
xnor U25929 (N_25929,N_25535,N_25465);
nand U25930 (N_25930,N_25259,N_25293);
nor U25931 (N_25931,N_25725,N_25245);
nor U25932 (N_25932,N_25209,N_25531);
nor U25933 (N_25933,N_25362,N_25278);
or U25934 (N_25934,N_25264,N_25392);
xnor U25935 (N_25935,N_25212,N_25621);
and U25936 (N_25936,N_25361,N_25315);
and U25937 (N_25937,N_25510,N_25552);
xor U25938 (N_25938,N_25607,N_25580);
and U25939 (N_25939,N_25764,N_25435);
or U25940 (N_25940,N_25473,N_25314);
or U25941 (N_25941,N_25539,N_25494);
nor U25942 (N_25942,N_25521,N_25747);
nand U25943 (N_25943,N_25653,N_25750);
and U25944 (N_25944,N_25429,N_25235);
nor U25945 (N_25945,N_25358,N_25561);
or U25946 (N_25946,N_25436,N_25781);
and U25947 (N_25947,N_25691,N_25501);
nand U25948 (N_25948,N_25598,N_25644);
nor U25949 (N_25949,N_25480,N_25570);
or U25950 (N_25950,N_25421,N_25546);
and U25951 (N_25951,N_25798,N_25694);
nand U25952 (N_25952,N_25673,N_25592);
xnor U25953 (N_25953,N_25730,N_25513);
xnor U25954 (N_25954,N_25783,N_25695);
nor U25955 (N_25955,N_25594,N_25210);
or U25956 (N_25956,N_25482,N_25251);
nor U25957 (N_25957,N_25682,N_25451);
nand U25958 (N_25958,N_25378,N_25796);
and U25959 (N_25959,N_25440,N_25767);
nand U25960 (N_25960,N_25736,N_25324);
nand U25961 (N_25961,N_25717,N_25738);
xor U25962 (N_25962,N_25671,N_25692);
nand U25963 (N_25963,N_25229,N_25769);
or U25964 (N_25964,N_25319,N_25374);
and U25965 (N_25965,N_25265,N_25656);
nor U25966 (N_25966,N_25710,N_25219);
or U25967 (N_25967,N_25397,N_25599);
xor U25968 (N_25968,N_25266,N_25677);
xor U25969 (N_25969,N_25763,N_25298);
xor U25970 (N_25970,N_25509,N_25775);
nor U25971 (N_25971,N_25263,N_25520);
nand U25972 (N_25972,N_25686,N_25431);
xor U25973 (N_25973,N_25544,N_25215);
nor U25974 (N_25974,N_25406,N_25443);
nand U25975 (N_25975,N_25420,N_25269);
nand U25976 (N_25976,N_25681,N_25326);
nand U25977 (N_25977,N_25467,N_25665);
and U25978 (N_25978,N_25793,N_25732);
and U25979 (N_25979,N_25797,N_25537);
xor U25980 (N_25980,N_25545,N_25475);
nand U25981 (N_25981,N_25211,N_25208);
and U25982 (N_25982,N_25391,N_25623);
nor U25983 (N_25983,N_25305,N_25697);
xnor U25984 (N_25984,N_25398,N_25759);
nor U25985 (N_25985,N_25596,N_25370);
and U25986 (N_25986,N_25413,N_25279);
xor U25987 (N_25987,N_25329,N_25418);
nor U25988 (N_25988,N_25600,N_25446);
nor U25989 (N_25989,N_25640,N_25542);
nand U25990 (N_25990,N_25430,N_25504);
nand U25991 (N_25991,N_25254,N_25748);
or U25992 (N_25992,N_25524,N_25369);
nand U25993 (N_25993,N_25676,N_25549);
nand U25994 (N_25994,N_25344,N_25632);
nand U25995 (N_25995,N_25666,N_25417);
and U25996 (N_25996,N_25457,N_25760);
nand U25997 (N_25997,N_25574,N_25735);
nor U25998 (N_25998,N_25582,N_25739);
nor U25999 (N_25999,N_25792,N_25218);
nor U26000 (N_26000,N_25617,N_25670);
nand U26001 (N_26001,N_25498,N_25659);
xor U26002 (N_26002,N_25779,N_25352);
xnor U26003 (N_26003,N_25606,N_25332);
and U26004 (N_26004,N_25300,N_25230);
nor U26005 (N_26005,N_25299,N_25741);
or U26006 (N_26006,N_25536,N_25727);
or U26007 (N_26007,N_25425,N_25252);
and U26008 (N_26008,N_25468,N_25583);
or U26009 (N_26009,N_25558,N_25619);
or U26010 (N_26010,N_25241,N_25428);
xnor U26011 (N_26011,N_25559,N_25340);
xnor U26012 (N_26012,N_25381,N_25630);
nor U26013 (N_26013,N_25771,N_25402);
nor U26014 (N_26014,N_25553,N_25683);
and U26015 (N_26015,N_25547,N_25486);
or U26016 (N_26016,N_25479,N_25490);
nor U26017 (N_26017,N_25351,N_25453);
nand U26018 (N_26018,N_25658,N_25492);
or U26019 (N_26019,N_25285,N_25562);
and U26020 (N_26020,N_25688,N_25464);
xor U26021 (N_26021,N_25585,N_25540);
nand U26022 (N_26022,N_25399,N_25226);
nand U26023 (N_26023,N_25722,N_25602);
nand U26024 (N_26024,N_25419,N_25271);
and U26025 (N_26025,N_25595,N_25262);
nor U26026 (N_26026,N_25500,N_25579);
nand U26027 (N_26027,N_25371,N_25638);
and U26028 (N_26028,N_25297,N_25423);
or U26029 (N_26029,N_25512,N_25385);
nor U26030 (N_26030,N_25661,N_25597);
nand U26031 (N_26031,N_25283,N_25422);
xor U26032 (N_26032,N_25338,N_25481);
and U26033 (N_26033,N_25668,N_25240);
xnor U26034 (N_26034,N_25255,N_25790);
and U26035 (N_26035,N_25689,N_25483);
xnor U26036 (N_26036,N_25444,N_25636);
nor U26037 (N_26037,N_25768,N_25427);
nand U26038 (N_26038,N_25702,N_25408);
xnor U26039 (N_26039,N_25581,N_25353);
xnor U26040 (N_26040,N_25274,N_25530);
nor U26041 (N_26041,N_25591,N_25260);
and U26042 (N_26042,N_25667,N_25232);
or U26043 (N_26043,N_25684,N_25357);
nor U26044 (N_26044,N_25341,N_25463);
nand U26045 (N_26045,N_25373,N_25724);
or U26046 (N_26046,N_25288,N_25515);
and U26047 (N_26047,N_25470,N_25611);
nor U26048 (N_26048,N_25390,N_25631);
xnor U26049 (N_26049,N_25393,N_25365);
nor U26050 (N_26050,N_25655,N_25563);
and U26051 (N_26051,N_25216,N_25526);
and U26052 (N_26052,N_25618,N_25497);
and U26053 (N_26053,N_25469,N_25349);
and U26054 (N_26054,N_25286,N_25238);
nand U26055 (N_26055,N_25321,N_25628);
xnor U26056 (N_26056,N_25267,N_25787);
xnor U26057 (N_26057,N_25472,N_25728);
nor U26058 (N_26058,N_25434,N_25534);
xor U26059 (N_26059,N_25204,N_25693);
xor U26060 (N_26060,N_25555,N_25608);
nor U26061 (N_26061,N_25330,N_25517);
or U26062 (N_26062,N_25731,N_25282);
and U26063 (N_26063,N_25589,N_25317);
and U26064 (N_26064,N_25647,N_25459);
xor U26065 (N_26065,N_25770,N_25214);
or U26066 (N_26066,N_25364,N_25577);
xor U26067 (N_26067,N_25756,N_25578);
nand U26068 (N_26068,N_25316,N_25572);
nand U26069 (N_26069,N_25318,N_25522);
nor U26070 (N_26070,N_25250,N_25496);
nor U26071 (N_26071,N_25213,N_25754);
nand U26072 (N_26072,N_25651,N_25571);
xnor U26073 (N_26073,N_25339,N_25237);
nand U26074 (N_26074,N_25757,N_25680);
nor U26075 (N_26075,N_25560,N_25543);
nand U26076 (N_26076,N_25308,N_25525);
nor U26077 (N_26077,N_25550,N_25711);
nand U26078 (N_26078,N_25342,N_25516);
xnor U26079 (N_26079,N_25679,N_25253);
nand U26080 (N_26080,N_25460,N_25335);
and U26081 (N_26081,N_25454,N_25488);
and U26082 (N_26082,N_25221,N_25721);
xor U26083 (N_26083,N_25276,N_25503);
nor U26084 (N_26084,N_25242,N_25273);
nand U26085 (N_26085,N_25642,N_25713);
nand U26086 (N_26086,N_25289,N_25590);
nand U26087 (N_26087,N_25657,N_25758);
xnor U26088 (N_26088,N_25409,N_25277);
and U26089 (N_26089,N_25256,N_25236);
and U26090 (N_26090,N_25784,N_25377);
nor U26091 (N_26091,N_25613,N_25701);
and U26092 (N_26092,N_25660,N_25207);
and U26093 (N_26093,N_25703,N_25437);
nor U26094 (N_26094,N_25584,N_25729);
or U26095 (N_26095,N_25396,N_25569);
nor U26096 (N_26096,N_25466,N_25564);
and U26097 (N_26097,N_25234,N_25609);
nor U26098 (N_26098,N_25478,N_25712);
nor U26099 (N_26099,N_25302,N_25203);
or U26100 (N_26100,N_25616,N_25386);
and U26101 (N_26101,N_25334,N_25411);
or U26102 (N_26102,N_25618,N_25542);
xor U26103 (N_26103,N_25204,N_25718);
or U26104 (N_26104,N_25233,N_25412);
and U26105 (N_26105,N_25310,N_25421);
nor U26106 (N_26106,N_25527,N_25449);
nor U26107 (N_26107,N_25513,N_25489);
or U26108 (N_26108,N_25230,N_25718);
and U26109 (N_26109,N_25506,N_25492);
or U26110 (N_26110,N_25656,N_25226);
and U26111 (N_26111,N_25398,N_25330);
xor U26112 (N_26112,N_25716,N_25574);
and U26113 (N_26113,N_25355,N_25583);
nand U26114 (N_26114,N_25475,N_25730);
or U26115 (N_26115,N_25379,N_25679);
xor U26116 (N_26116,N_25346,N_25502);
and U26117 (N_26117,N_25444,N_25631);
xor U26118 (N_26118,N_25718,N_25736);
or U26119 (N_26119,N_25266,N_25229);
or U26120 (N_26120,N_25515,N_25632);
and U26121 (N_26121,N_25554,N_25235);
and U26122 (N_26122,N_25269,N_25604);
nor U26123 (N_26123,N_25290,N_25560);
nor U26124 (N_26124,N_25276,N_25702);
nand U26125 (N_26125,N_25665,N_25494);
xor U26126 (N_26126,N_25600,N_25395);
nor U26127 (N_26127,N_25677,N_25587);
nand U26128 (N_26128,N_25662,N_25578);
nand U26129 (N_26129,N_25660,N_25757);
nand U26130 (N_26130,N_25479,N_25771);
nor U26131 (N_26131,N_25665,N_25632);
and U26132 (N_26132,N_25697,N_25490);
and U26133 (N_26133,N_25266,N_25430);
and U26134 (N_26134,N_25572,N_25436);
xnor U26135 (N_26135,N_25490,N_25617);
and U26136 (N_26136,N_25327,N_25234);
or U26137 (N_26137,N_25331,N_25221);
or U26138 (N_26138,N_25450,N_25675);
nor U26139 (N_26139,N_25665,N_25776);
xor U26140 (N_26140,N_25404,N_25634);
nor U26141 (N_26141,N_25715,N_25230);
nand U26142 (N_26142,N_25357,N_25284);
nor U26143 (N_26143,N_25637,N_25273);
nand U26144 (N_26144,N_25580,N_25358);
or U26145 (N_26145,N_25682,N_25233);
nor U26146 (N_26146,N_25460,N_25740);
and U26147 (N_26147,N_25733,N_25376);
nor U26148 (N_26148,N_25356,N_25251);
xor U26149 (N_26149,N_25534,N_25750);
and U26150 (N_26150,N_25261,N_25656);
nand U26151 (N_26151,N_25767,N_25470);
nand U26152 (N_26152,N_25711,N_25382);
xor U26153 (N_26153,N_25406,N_25514);
nand U26154 (N_26154,N_25339,N_25279);
nor U26155 (N_26155,N_25371,N_25285);
or U26156 (N_26156,N_25502,N_25770);
or U26157 (N_26157,N_25731,N_25473);
and U26158 (N_26158,N_25272,N_25358);
nand U26159 (N_26159,N_25563,N_25306);
xor U26160 (N_26160,N_25532,N_25480);
or U26161 (N_26161,N_25414,N_25498);
or U26162 (N_26162,N_25627,N_25379);
nand U26163 (N_26163,N_25336,N_25524);
or U26164 (N_26164,N_25667,N_25486);
nor U26165 (N_26165,N_25570,N_25672);
nand U26166 (N_26166,N_25564,N_25704);
nand U26167 (N_26167,N_25242,N_25604);
and U26168 (N_26168,N_25696,N_25504);
and U26169 (N_26169,N_25386,N_25297);
nor U26170 (N_26170,N_25678,N_25286);
xnor U26171 (N_26171,N_25386,N_25612);
and U26172 (N_26172,N_25237,N_25467);
xor U26173 (N_26173,N_25788,N_25577);
nor U26174 (N_26174,N_25753,N_25240);
nand U26175 (N_26175,N_25237,N_25512);
nand U26176 (N_26176,N_25552,N_25644);
nand U26177 (N_26177,N_25458,N_25312);
or U26178 (N_26178,N_25282,N_25626);
nand U26179 (N_26179,N_25546,N_25287);
nor U26180 (N_26180,N_25698,N_25780);
and U26181 (N_26181,N_25618,N_25361);
nand U26182 (N_26182,N_25345,N_25224);
nor U26183 (N_26183,N_25456,N_25403);
nand U26184 (N_26184,N_25652,N_25311);
xor U26185 (N_26185,N_25762,N_25420);
or U26186 (N_26186,N_25625,N_25683);
or U26187 (N_26187,N_25271,N_25332);
xnor U26188 (N_26188,N_25292,N_25344);
and U26189 (N_26189,N_25582,N_25653);
nand U26190 (N_26190,N_25417,N_25642);
xor U26191 (N_26191,N_25284,N_25458);
nor U26192 (N_26192,N_25653,N_25464);
nor U26193 (N_26193,N_25526,N_25272);
xnor U26194 (N_26194,N_25270,N_25486);
and U26195 (N_26195,N_25353,N_25685);
and U26196 (N_26196,N_25293,N_25324);
or U26197 (N_26197,N_25374,N_25600);
nor U26198 (N_26198,N_25614,N_25670);
nand U26199 (N_26199,N_25485,N_25764);
or U26200 (N_26200,N_25281,N_25722);
and U26201 (N_26201,N_25200,N_25371);
nand U26202 (N_26202,N_25701,N_25761);
and U26203 (N_26203,N_25606,N_25635);
nor U26204 (N_26204,N_25430,N_25422);
nand U26205 (N_26205,N_25773,N_25430);
nand U26206 (N_26206,N_25365,N_25499);
or U26207 (N_26207,N_25684,N_25490);
nand U26208 (N_26208,N_25626,N_25794);
xor U26209 (N_26209,N_25741,N_25407);
xor U26210 (N_26210,N_25490,N_25315);
or U26211 (N_26211,N_25475,N_25726);
nor U26212 (N_26212,N_25703,N_25284);
or U26213 (N_26213,N_25724,N_25335);
or U26214 (N_26214,N_25378,N_25423);
nand U26215 (N_26215,N_25779,N_25737);
nor U26216 (N_26216,N_25476,N_25667);
nand U26217 (N_26217,N_25736,N_25399);
or U26218 (N_26218,N_25398,N_25283);
xor U26219 (N_26219,N_25738,N_25462);
nor U26220 (N_26220,N_25304,N_25441);
nand U26221 (N_26221,N_25425,N_25687);
nor U26222 (N_26222,N_25768,N_25624);
xor U26223 (N_26223,N_25551,N_25445);
nand U26224 (N_26224,N_25318,N_25569);
or U26225 (N_26225,N_25502,N_25431);
nand U26226 (N_26226,N_25234,N_25547);
or U26227 (N_26227,N_25233,N_25756);
nand U26228 (N_26228,N_25217,N_25720);
and U26229 (N_26229,N_25376,N_25488);
and U26230 (N_26230,N_25606,N_25751);
nor U26231 (N_26231,N_25578,N_25547);
nor U26232 (N_26232,N_25721,N_25463);
xor U26233 (N_26233,N_25574,N_25409);
xor U26234 (N_26234,N_25537,N_25595);
or U26235 (N_26235,N_25774,N_25345);
or U26236 (N_26236,N_25399,N_25703);
or U26237 (N_26237,N_25615,N_25736);
nor U26238 (N_26238,N_25376,N_25597);
nor U26239 (N_26239,N_25663,N_25318);
and U26240 (N_26240,N_25767,N_25612);
and U26241 (N_26241,N_25228,N_25439);
or U26242 (N_26242,N_25658,N_25782);
and U26243 (N_26243,N_25674,N_25434);
or U26244 (N_26244,N_25783,N_25438);
nor U26245 (N_26245,N_25332,N_25487);
nor U26246 (N_26246,N_25225,N_25785);
or U26247 (N_26247,N_25606,N_25404);
xor U26248 (N_26248,N_25353,N_25383);
xor U26249 (N_26249,N_25770,N_25639);
nor U26250 (N_26250,N_25256,N_25563);
and U26251 (N_26251,N_25360,N_25321);
nor U26252 (N_26252,N_25437,N_25456);
nand U26253 (N_26253,N_25358,N_25273);
nor U26254 (N_26254,N_25721,N_25569);
xor U26255 (N_26255,N_25675,N_25204);
or U26256 (N_26256,N_25341,N_25235);
or U26257 (N_26257,N_25464,N_25788);
xor U26258 (N_26258,N_25596,N_25314);
nand U26259 (N_26259,N_25730,N_25737);
nand U26260 (N_26260,N_25433,N_25478);
or U26261 (N_26261,N_25377,N_25790);
xor U26262 (N_26262,N_25651,N_25367);
nand U26263 (N_26263,N_25617,N_25790);
nand U26264 (N_26264,N_25404,N_25605);
xnor U26265 (N_26265,N_25472,N_25309);
or U26266 (N_26266,N_25634,N_25679);
nor U26267 (N_26267,N_25725,N_25334);
and U26268 (N_26268,N_25494,N_25511);
and U26269 (N_26269,N_25556,N_25451);
nand U26270 (N_26270,N_25305,N_25354);
nand U26271 (N_26271,N_25429,N_25694);
nor U26272 (N_26272,N_25775,N_25623);
xor U26273 (N_26273,N_25511,N_25781);
nor U26274 (N_26274,N_25442,N_25267);
nor U26275 (N_26275,N_25413,N_25663);
nor U26276 (N_26276,N_25789,N_25681);
xor U26277 (N_26277,N_25418,N_25459);
or U26278 (N_26278,N_25767,N_25212);
and U26279 (N_26279,N_25476,N_25313);
or U26280 (N_26280,N_25668,N_25581);
and U26281 (N_26281,N_25615,N_25264);
and U26282 (N_26282,N_25705,N_25748);
xor U26283 (N_26283,N_25740,N_25645);
or U26284 (N_26284,N_25734,N_25305);
and U26285 (N_26285,N_25390,N_25640);
and U26286 (N_26286,N_25746,N_25388);
and U26287 (N_26287,N_25763,N_25309);
xnor U26288 (N_26288,N_25435,N_25753);
xnor U26289 (N_26289,N_25452,N_25498);
and U26290 (N_26290,N_25315,N_25226);
xnor U26291 (N_26291,N_25576,N_25612);
nor U26292 (N_26292,N_25274,N_25408);
or U26293 (N_26293,N_25379,N_25240);
or U26294 (N_26294,N_25675,N_25615);
nand U26295 (N_26295,N_25796,N_25554);
nand U26296 (N_26296,N_25649,N_25312);
or U26297 (N_26297,N_25619,N_25626);
and U26298 (N_26298,N_25600,N_25799);
and U26299 (N_26299,N_25254,N_25465);
or U26300 (N_26300,N_25294,N_25309);
nand U26301 (N_26301,N_25383,N_25709);
and U26302 (N_26302,N_25259,N_25393);
and U26303 (N_26303,N_25509,N_25386);
or U26304 (N_26304,N_25784,N_25385);
nand U26305 (N_26305,N_25431,N_25355);
and U26306 (N_26306,N_25419,N_25402);
xnor U26307 (N_26307,N_25796,N_25397);
xor U26308 (N_26308,N_25755,N_25226);
and U26309 (N_26309,N_25283,N_25235);
nor U26310 (N_26310,N_25241,N_25552);
or U26311 (N_26311,N_25747,N_25464);
nand U26312 (N_26312,N_25699,N_25375);
and U26313 (N_26313,N_25575,N_25739);
and U26314 (N_26314,N_25719,N_25567);
nor U26315 (N_26315,N_25635,N_25753);
or U26316 (N_26316,N_25201,N_25236);
xnor U26317 (N_26317,N_25523,N_25401);
nand U26318 (N_26318,N_25794,N_25247);
and U26319 (N_26319,N_25704,N_25713);
nand U26320 (N_26320,N_25654,N_25312);
nand U26321 (N_26321,N_25550,N_25470);
xnor U26322 (N_26322,N_25634,N_25596);
xor U26323 (N_26323,N_25365,N_25310);
xnor U26324 (N_26324,N_25496,N_25581);
nor U26325 (N_26325,N_25337,N_25300);
xnor U26326 (N_26326,N_25778,N_25366);
and U26327 (N_26327,N_25579,N_25584);
nand U26328 (N_26328,N_25465,N_25544);
or U26329 (N_26329,N_25792,N_25469);
or U26330 (N_26330,N_25625,N_25371);
or U26331 (N_26331,N_25389,N_25516);
nor U26332 (N_26332,N_25695,N_25609);
nor U26333 (N_26333,N_25599,N_25517);
xor U26334 (N_26334,N_25693,N_25233);
xor U26335 (N_26335,N_25558,N_25456);
or U26336 (N_26336,N_25442,N_25666);
xnor U26337 (N_26337,N_25595,N_25527);
and U26338 (N_26338,N_25213,N_25626);
or U26339 (N_26339,N_25593,N_25227);
and U26340 (N_26340,N_25445,N_25701);
nand U26341 (N_26341,N_25742,N_25649);
xnor U26342 (N_26342,N_25460,N_25767);
or U26343 (N_26343,N_25670,N_25643);
and U26344 (N_26344,N_25324,N_25755);
or U26345 (N_26345,N_25293,N_25581);
xnor U26346 (N_26346,N_25532,N_25500);
and U26347 (N_26347,N_25647,N_25710);
and U26348 (N_26348,N_25311,N_25552);
and U26349 (N_26349,N_25273,N_25262);
nand U26350 (N_26350,N_25627,N_25573);
or U26351 (N_26351,N_25400,N_25776);
nand U26352 (N_26352,N_25784,N_25351);
xor U26353 (N_26353,N_25236,N_25372);
nand U26354 (N_26354,N_25579,N_25235);
xnor U26355 (N_26355,N_25696,N_25500);
nand U26356 (N_26356,N_25393,N_25664);
nand U26357 (N_26357,N_25794,N_25769);
nand U26358 (N_26358,N_25328,N_25762);
nand U26359 (N_26359,N_25395,N_25766);
nand U26360 (N_26360,N_25592,N_25540);
nor U26361 (N_26361,N_25719,N_25298);
or U26362 (N_26362,N_25556,N_25440);
nand U26363 (N_26363,N_25734,N_25621);
or U26364 (N_26364,N_25695,N_25224);
or U26365 (N_26365,N_25626,N_25654);
nor U26366 (N_26366,N_25605,N_25755);
and U26367 (N_26367,N_25775,N_25237);
or U26368 (N_26368,N_25414,N_25444);
nand U26369 (N_26369,N_25223,N_25473);
and U26370 (N_26370,N_25207,N_25506);
xor U26371 (N_26371,N_25454,N_25244);
xor U26372 (N_26372,N_25500,N_25216);
and U26373 (N_26373,N_25293,N_25467);
nand U26374 (N_26374,N_25660,N_25797);
and U26375 (N_26375,N_25336,N_25416);
xor U26376 (N_26376,N_25674,N_25520);
or U26377 (N_26377,N_25798,N_25659);
or U26378 (N_26378,N_25706,N_25686);
nand U26379 (N_26379,N_25251,N_25757);
nand U26380 (N_26380,N_25737,N_25666);
nand U26381 (N_26381,N_25265,N_25535);
and U26382 (N_26382,N_25379,N_25749);
nor U26383 (N_26383,N_25733,N_25650);
and U26384 (N_26384,N_25260,N_25596);
and U26385 (N_26385,N_25716,N_25381);
xor U26386 (N_26386,N_25290,N_25365);
nand U26387 (N_26387,N_25511,N_25500);
or U26388 (N_26388,N_25638,N_25344);
nand U26389 (N_26389,N_25334,N_25333);
nor U26390 (N_26390,N_25314,N_25425);
nor U26391 (N_26391,N_25319,N_25562);
or U26392 (N_26392,N_25637,N_25280);
nor U26393 (N_26393,N_25485,N_25600);
nand U26394 (N_26394,N_25549,N_25721);
or U26395 (N_26395,N_25359,N_25685);
and U26396 (N_26396,N_25676,N_25582);
or U26397 (N_26397,N_25789,N_25602);
and U26398 (N_26398,N_25430,N_25699);
nor U26399 (N_26399,N_25567,N_25355);
nor U26400 (N_26400,N_26036,N_26380);
and U26401 (N_26401,N_26110,N_26131);
or U26402 (N_26402,N_26368,N_26136);
nor U26403 (N_26403,N_25808,N_26295);
or U26404 (N_26404,N_25990,N_26203);
nand U26405 (N_26405,N_25982,N_26210);
nand U26406 (N_26406,N_25920,N_25928);
or U26407 (N_26407,N_26090,N_25997);
nor U26408 (N_26408,N_25922,N_26243);
nand U26409 (N_26409,N_25906,N_25848);
nand U26410 (N_26410,N_25913,N_26150);
nand U26411 (N_26411,N_26389,N_26216);
and U26412 (N_26412,N_25855,N_26043);
or U26413 (N_26413,N_25993,N_26335);
or U26414 (N_26414,N_26179,N_25834);
or U26415 (N_26415,N_25974,N_26129);
nor U26416 (N_26416,N_25981,N_26272);
or U26417 (N_26417,N_25950,N_26045);
nand U26418 (N_26418,N_26225,N_26326);
nor U26419 (N_26419,N_25891,N_26311);
and U26420 (N_26420,N_26391,N_26111);
and U26421 (N_26421,N_25843,N_25816);
xor U26422 (N_26422,N_26306,N_26155);
nand U26423 (N_26423,N_26082,N_26357);
nor U26424 (N_26424,N_26120,N_26276);
nor U26425 (N_26425,N_26340,N_26201);
xnor U26426 (N_26426,N_26371,N_26035);
or U26427 (N_26427,N_26133,N_26267);
nor U26428 (N_26428,N_26304,N_25953);
and U26429 (N_26429,N_25998,N_26281);
nand U26430 (N_26430,N_26062,N_26298);
and U26431 (N_26431,N_26399,N_26092);
xor U26432 (N_26432,N_25819,N_26174);
and U26433 (N_26433,N_26382,N_25983);
or U26434 (N_26434,N_26254,N_25870);
nand U26435 (N_26435,N_26152,N_26048);
xnor U26436 (N_26436,N_26183,N_25839);
nand U26437 (N_26437,N_25952,N_26029);
and U26438 (N_26438,N_26051,N_26242);
nor U26439 (N_26439,N_26070,N_25811);
xor U26440 (N_26440,N_25915,N_25844);
and U26441 (N_26441,N_26003,N_25846);
and U26442 (N_26442,N_25988,N_26021);
xnor U26443 (N_26443,N_26031,N_25930);
nor U26444 (N_26444,N_26019,N_26397);
or U26445 (N_26445,N_25987,N_25813);
xor U26446 (N_26446,N_26393,N_26354);
nand U26447 (N_26447,N_25895,N_25858);
nand U26448 (N_26448,N_26080,N_26346);
or U26449 (N_26449,N_25818,N_25901);
and U26450 (N_26450,N_26292,N_26006);
nor U26451 (N_26451,N_26372,N_25944);
nand U26452 (N_26452,N_26213,N_26307);
xnor U26453 (N_26453,N_26094,N_26159);
xor U26454 (N_26454,N_26252,N_26364);
and U26455 (N_26455,N_26379,N_25934);
xor U26456 (N_26456,N_26299,N_26124);
nand U26457 (N_26457,N_25946,N_26227);
or U26458 (N_26458,N_26394,N_26385);
xnor U26459 (N_26459,N_25951,N_25801);
nor U26460 (N_26460,N_26395,N_26322);
and U26461 (N_26461,N_25833,N_26000);
xor U26462 (N_26462,N_25885,N_25905);
and U26463 (N_26463,N_26071,N_26234);
nor U26464 (N_26464,N_26114,N_26205);
nand U26465 (N_26465,N_25931,N_26353);
and U26466 (N_26466,N_26269,N_26245);
xor U26467 (N_26467,N_26121,N_26163);
nor U26468 (N_26468,N_26211,N_26323);
nor U26469 (N_26469,N_25877,N_26332);
or U26470 (N_26470,N_26296,N_26140);
or U26471 (N_26471,N_26233,N_26231);
and U26472 (N_26472,N_26352,N_26009);
nor U26473 (N_26473,N_26343,N_26348);
nand U26474 (N_26474,N_25941,N_26308);
and U26475 (N_26475,N_26142,N_26313);
and U26476 (N_26476,N_26044,N_26146);
nand U26477 (N_26477,N_25856,N_26257);
nand U26478 (N_26478,N_25911,N_26273);
nand U26479 (N_26479,N_26373,N_26190);
nand U26480 (N_26480,N_26042,N_26305);
and U26481 (N_26481,N_25959,N_26162);
or U26482 (N_26482,N_26235,N_26253);
nor U26483 (N_26483,N_26334,N_26219);
nor U26484 (N_26484,N_26109,N_26030);
nand U26485 (N_26485,N_26283,N_26390);
and U26486 (N_26486,N_26108,N_26317);
xor U26487 (N_26487,N_26294,N_25826);
nor U26488 (N_26488,N_26189,N_26087);
or U26489 (N_26489,N_25985,N_25955);
and U26490 (N_26490,N_26293,N_25942);
or U26491 (N_26491,N_26214,N_26081);
and U26492 (N_26492,N_26251,N_25842);
nor U26493 (N_26493,N_26187,N_25845);
or U26494 (N_26494,N_26158,N_26101);
nor U26495 (N_26495,N_26024,N_26270);
or U26496 (N_26496,N_26115,N_25866);
xor U26497 (N_26497,N_26202,N_25824);
nor U26498 (N_26498,N_26383,N_26089);
and U26499 (N_26499,N_26359,N_26369);
nand U26500 (N_26500,N_26025,N_25803);
and U26501 (N_26501,N_25948,N_26139);
nand U26502 (N_26502,N_26229,N_26113);
nand U26503 (N_26503,N_25917,N_25902);
nor U26504 (N_26504,N_26054,N_25840);
xor U26505 (N_26505,N_26010,N_26207);
nor U26506 (N_26506,N_26288,N_26309);
nand U26507 (N_26507,N_26122,N_26100);
xnor U26508 (N_26508,N_26104,N_26318);
and U26509 (N_26509,N_25984,N_26261);
xnor U26510 (N_26510,N_25995,N_26215);
xor U26511 (N_26511,N_26147,N_26223);
xnor U26512 (N_26512,N_25945,N_26191);
xnor U26513 (N_26513,N_25868,N_25936);
nor U26514 (N_26514,N_26208,N_25822);
and U26515 (N_26515,N_26123,N_25933);
nand U26516 (N_26516,N_25859,N_26333);
or U26517 (N_26517,N_26386,N_25832);
nor U26518 (N_26518,N_26017,N_26074);
xnor U26519 (N_26519,N_26388,N_26206);
or U26520 (N_26520,N_26022,N_26028);
or U26521 (N_26521,N_25912,N_25940);
nand U26522 (N_26522,N_25854,N_26173);
xnor U26523 (N_26523,N_26260,N_26002);
and U26524 (N_26524,N_26145,N_25847);
nand U26525 (N_26525,N_26331,N_25973);
nor U26526 (N_26526,N_26095,N_26141);
nor U26527 (N_26527,N_26312,N_25989);
nor U26528 (N_26528,N_26079,N_26169);
and U26529 (N_26529,N_26168,N_26337);
nand U26530 (N_26530,N_26032,N_25888);
nor U26531 (N_26531,N_26197,N_25910);
nand U26532 (N_26532,N_25838,N_26349);
or U26533 (N_26533,N_26297,N_25960);
xor U26534 (N_26534,N_26342,N_25867);
nand U26535 (N_26535,N_26204,N_25850);
nor U26536 (N_26536,N_26078,N_26185);
xnor U26537 (N_26537,N_25865,N_25924);
or U26538 (N_26538,N_26226,N_26246);
or U26539 (N_26539,N_25927,N_26241);
nand U26540 (N_26540,N_25815,N_25863);
xor U26541 (N_26541,N_26020,N_25853);
nand U26542 (N_26542,N_25882,N_25831);
nor U26543 (N_26543,N_26387,N_25925);
nor U26544 (N_26544,N_26135,N_26374);
and U26545 (N_26545,N_26039,N_26012);
xor U26546 (N_26546,N_26336,N_26271);
nand U26547 (N_26547,N_26398,N_26160);
nor U26548 (N_26548,N_25827,N_26344);
and U26549 (N_26549,N_26303,N_26300);
or U26550 (N_26550,N_26023,N_26099);
and U26551 (N_26551,N_25980,N_25809);
or U26552 (N_26552,N_26362,N_26005);
or U26553 (N_26553,N_25898,N_26096);
and U26554 (N_26554,N_26290,N_26107);
and U26555 (N_26555,N_25881,N_25977);
nand U26556 (N_26556,N_25860,N_26118);
and U26557 (N_26557,N_26320,N_26061);
and U26558 (N_26558,N_26265,N_25926);
and U26559 (N_26559,N_25939,N_26329);
nand U26560 (N_26560,N_26112,N_26040);
nand U26561 (N_26561,N_26345,N_25851);
or U26562 (N_26562,N_26171,N_26038);
and U26563 (N_26563,N_26366,N_26076);
xor U26564 (N_26564,N_26165,N_26067);
nand U26565 (N_26565,N_25969,N_26218);
or U26566 (N_26566,N_26161,N_26086);
and U26567 (N_26567,N_26128,N_25810);
nor U26568 (N_26568,N_26148,N_25949);
nor U26569 (N_26569,N_25897,N_26360);
or U26570 (N_26570,N_26105,N_25999);
or U26571 (N_26571,N_26325,N_26355);
nand U26572 (N_26572,N_26011,N_26339);
and U26573 (N_26573,N_25976,N_26262);
nor U26574 (N_26574,N_26209,N_26324);
nor U26575 (N_26575,N_25861,N_26063);
xor U26576 (N_26576,N_26250,N_26268);
nand U26577 (N_26577,N_26199,N_25935);
and U26578 (N_26578,N_25918,N_26278);
xor U26579 (N_26579,N_26164,N_26049);
and U26580 (N_26580,N_25852,N_26098);
or U26581 (N_26581,N_26091,N_26137);
and U26582 (N_26582,N_26068,N_26195);
nor U26583 (N_26583,N_26004,N_26102);
and U26584 (N_26584,N_26230,N_26310);
xnor U26585 (N_26585,N_25879,N_26047);
and U26586 (N_26586,N_25849,N_25943);
and U26587 (N_26587,N_26249,N_25908);
nand U26588 (N_26588,N_25896,N_26351);
xnor U26589 (N_26589,N_26315,N_26154);
or U26590 (N_26590,N_26365,N_25957);
or U26591 (N_26591,N_26277,N_26330);
or U26592 (N_26592,N_25907,N_25805);
nand U26593 (N_26593,N_26378,N_25800);
and U26594 (N_26594,N_26132,N_25975);
xor U26595 (N_26595,N_25894,N_25837);
nand U26596 (N_26596,N_26347,N_25873);
or U26597 (N_26597,N_26376,N_26119);
nand U26598 (N_26598,N_26301,N_25857);
nand U26599 (N_26599,N_25900,N_25884);
xor U26600 (N_26600,N_25874,N_26184);
nor U26601 (N_26601,N_26175,N_26217);
xor U26602 (N_26602,N_26396,N_26319);
nand U26603 (N_26603,N_25992,N_26037);
or U26604 (N_26604,N_26007,N_26274);
and U26605 (N_26605,N_25875,N_26144);
xnor U26606 (N_26606,N_25968,N_25830);
and U26607 (N_26607,N_25864,N_26053);
and U26608 (N_26608,N_26126,N_26259);
nor U26609 (N_26609,N_26156,N_25876);
nor U26610 (N_26610,N_25804,N_26263);
or U26611 (N_26611,N_25823,N_26097);
xor U26612 (N_26612,N_25916,N_26196);
or U26613 (N_26613,N_26279,N_26125);
xnor U26614 (N_26614,N_26224,N_26157);
and U26615 (N_26615,N_25929,N_26255);
xnor U26616 (N_26616,N_26013,N_26280);
and U26617 (N_26617,N_26072,N_26085);
or U26618 (N_26618,N_26327,N_26066);
nor U26619 (N_26619,N_26221,N_26050);
or U26620 (N_26620,N_26064,N_26302);
and U26621 (N_26621,N_25965,N_25956);
nand U26622 (N_26622,N_26055,N_25958);
and U26623 (N_26623,N_25966,N_26392);
nand U26624 (N_26624,N_26170,N_25862);
or U26625 (N_26625,N_26316,N_26338);
nor U26626 (N_26626,N_26266,N_25964);
xor U26627 (N_26627,N_25994,N_25909);
nor U26628 (N_26628,N_26018,N_26033);
nand U26629 (N_26629,N_26172,N_26256);
nor U26630 (N_26630,N_26059,N_26358);
nor U26631 (N_26631,N_25802,N_25872);
xnor U26632 (N_26632,N_26181,N_26321);
and U26633 (N_26633,N_26058,N_26194);
or U26634 (N_26634,N_25841,N_26198);
nor U26635 (N_26635,N_26167,N_26077);
and U26636 (N_26636,N_25821,N_25814);
nor U26637 (N_26637,N_26361,N_26116);
or U26638 (N_26638,N_26093,N_25886);
nand U26639 (N_26639,N_26356,N_25890);
nor U26640 (N_26640,N_25883,N_26248);
and U26641 (N_26641,N_26138,N_26069);
xnor U26642 (N_26642,N_26314,N_25972);
or U26643 (N_26643,N_26177,N_25892);
nor U26644 (N_26644,N_26130,N_26041);
xor U26645 (N_26645,N_25919,N_26240);
xnor U26646 (N_26646,N_25986,N_25967);
nand U26647 (N_26647,N_25835,N_25962);
xor U26648 (N_26648,N_25899,N_26247);
or U26649 (N_26649,N_25947,N_26015);
or U26650 (N_26650,N_25820,N_25807);
xor U26651 (N_26651,N_26117,N_26285);
xnor U26652 (N_26652,N_26151,N_26232);
and U26653 (N_26653,N_26192,N_26381);
and U26654 (N_26654,N_25954,N_26258);
and U26655 (N_26655,N_26212,N_25932);
and U26656 (N_26656,N_26014,N_25812);
xnor U26657 (N_26657,N_26075,N_26088);
nand U26658 (N_26658,N_26244,N_26286);
or U26659 (N_26659,N_26153,N_25829);
nand U26660 (N_26660,N_25938,N_25937);
nand U26661 (N_26661,N_25963,N_25961);
xnor U26662 (N_26662,N_26001,N_26284);
or U26663 (N_26663,N_25978,N_25828);
or U26664 (N_26664,N_26341,N_25970);
nor U26665 (N_26665,N_26220,N_26186);
or U26666 (N_26666,N_26056,N_26375);
or U26667 (N_26667,N_26083,N_25880);
xnor U26668 (N_26668,N_26143,N_25996);
nor U26669 (N_26669,N_26239,N_26060);
nand U26670 (N_26670,N_26134,N_26149);
xnor U26671 (N_26671,N_26188,N_26287);
and U26672 (N_26672,N_25923,N_25979);
xnor U26673 (N_26673,N_25991,N_25904);
xor U26674 (N_26674,N_26282,N_26052);
nand U26675 (N_26675,N_26103,N_26384);
nand U26676 (N_26676,N_26367,N_26289);
nand U26677 (N_26677,N_26237,N_26291);
and U26678 (N_26678,N_25914,N_26034);
nand U26679 (N_26679,N_26057,N_26236);
nand U26680 (N_26680,N_26228,N_26026);
nand U26681 (N_26681,N_25887,N_26073);
or U26682 (N_26682,N_26182,N_26350);
and U26683 (N_26683,N_26027,N_26363);
and U26684 (N_26684,N_25871,N_25806);
or U26685 (N_26685,N_26008,N_25825);
or U26686 (N_26686,N_26238,N_26046);
nand U26687 (N_26687,N_26127,N_26275);
xor U26688 (N_26688,N_26377,N_26016);
nor U26689 (N_26689,N_26065,N_25921);
nor U26690 (N_26690,N_25971,N_26222);
nand U26691 (N_26691,N_26084,N_26200);
xnor U26692 (N_26692,N_26264,N_25869);
nor U26693 (N_26693,N_25903,N_25893);
xor U26694 (N_26694,N_26106,N_26328);
nand U26695 (N_26695,N_26176,N_26178);
xor U26696 (N_26696,N_25817,N_26193);
nor U26697 (N_26697,N_25889,N_25878);
nor U26698 (N_26698,N_26166,N_26370);
nor U26699 (N_26699,N_25836,N_26180);
or U26700 (N_26700,N_25860,N_26281);
and U26701 (N_26701,N_26000,N_25939);
nand U26702 (N_26702,N_26329,N_26240);
and U26703 (N_26703,N_25924,N_25918);
and U26704 (N_26704,N_25823,N_25862);
nor U26705 (N_26705,N_25968,N_26064);
nor U26706 (N_26706,N_25878,N_25990);
nand U26707 (N_26707,N_25982,N_26236);
xnor U26708 (N_26708,N_25968,N_26357);
nor U26709 (N_26709,N_26124,N_26203);
or U26710 (N_26710,N_25887,N_26344);
nand U26711 (N_26711,N_26293,N_26136);
and U26712 (N_26712,N_26380,N_26381);
and U26713 (N_26713,N_26034,N_25927);
xor U26714 (N_26714,N_26156,N_26209);
nor U26715 (N_26715,N_26290,N_26277);
nand U26716 (N_26716,N_26016,N_26181);
or U26717 (N_26717,N_26313,N_25963);
and U26718 (N_26718,N_26281,N_26168);
nand U26719 (N_26719,N_25839,N_26061);
xnor U26720 (N_26720,N_25925,N_25952);
or U26721 (N_26721,N_26047,N_26146);
nor U26722 (N_26722,N_25848,N_25813);
xnor U26723 (N_26723,N_25980,N_25932);
and U26724 (N_26724,N_26339,N_25949);
nand U26725 (N_26725,N_25809,N_26204);
nor U26726 (N_26726,N_25811,N_25947);
and U26727 (N_26727,N_26035,N_26355);
and U26728 (N_26728,N_25885,N_26153);
or U26729 (N_26729,N_25821,N_26012);
xor U26730 (N_26730,N_26067,N_26157);
nor U26731 (N_26731,N_25905,N_26191);
and U26732 (N_26732,N_26300,N_25894);
nand U26733 (N_26733,N_25992,N_25909);
nand U26734 (N_26734,N_26021,N_25883);
xor U26735 (N_26735,N_25881,N_26298);
xor U26736 (N_26736,N_25902,N_25891);
nor U26737 (N_26737,N_26145,N_26349);
nor U26738 (N_26738,N_25944,N_26229);
nor U26739 (N_26739,N_25928,N_26234);
and U26740 (N_26740,N_25905,N_25844);
or U26741 (N_26741,N_26343,N_26378);
xor U26742 (N_26742,N_26055,N_25814);
and U26743 (N_26743,N_25991,N_25876);
nor U26744 (N_26744,N_26073,N_26127);
xor U26745 (N_26745,N_26343,N_26387);
nand U26746 (N_26746,N_26177,N_26032);
and U26747 (N_26747,N_25855,N_25982);
xor U26748 (N_26748,N_25822,N_26343);
nor U26749 (N_26749,N_25894,N_26257);
and U26750 (N_26750,N_26008,N_26010);
or U26751 (N_26751,N_25801,N_26052);
xor U26752 (N_26752,N_25877,N_25861);
or U26753 (N_26753,N_26050,N_26175);
nand U26754 (N_26754,N_26017,N_26029);
nand U26755 (N_26755,N_26067,N_25890);
nor U26756 (N_26756,N_26032,N_26323);
nand U26757 (N_26757,N_25933,N_26022);
xnor U26758 (N_26758,N_25860,N_26367);
or U26759 (N_26759,N_25857,N_25821);
nand U26760 (N_26760,N_26238,N_25942);
xor U26761 (N_26761,N_26144,N_25882);
nand U26762 (N_26762,N_26147,N_26058);
nor U26763 (N_26763,N_25873,N_26037);
and U26764 (N_26764,N_26233,N_26069);
and U26765 (N_26765,N_26111,N_26258);
and U26766 (N_26766,N_26320,N_26335);
and U26767 (N_26767,N_25835,N_25838);
and U26768 (N_26768,N_26319,N_25923);
and U26769 (N_26769,N_26074,N_26376);
nor U26770 (N_26770,N_26196,N_26315);
nand U26771 (N_26771,N_25912,N_25901);
xor U26772 (N_26772,N_25941,N_25988);
nor U26773 (N_26773,N_26034,N_26255);
nand U26774 (N_26774,N_26251,N_26233);
or U26775 (N_26775,N_26110,N_26036);
nand U26776 (N_26776,N_25807,N_25975);
nand U26777 (N_26777,N_26211,N_25924);
and U26778 (N_26778,N_26255,N_25819);
or U26779 (N_26779,N_26150,N_26012);
nand U26780 (N_26780,N_26181,N_26162);
and U26781 (N_26781,N_26142,N_25965);
nor U26782 (N_26782,N_25804,N_26069);
nor U26783 (N_26783,N_26249,N_26043);
or U26784 (N_26784,N_26102,N_26270);
nand U26785 (N_26785,N_25928,N_26155);
xnor U26786 (N_26786,N_26025,N_25941);
and U26787 (N_26787,N_25805,N_26320);
xnor U26788 (N_26788,N_26287,N_26336);
xnor U26789 (N_26789,N_25935,N_26116);
or U26790 (N_26790,N_25943,N_26005);
nor U26791 (N_26791,N_26327,N_26036);
nor U26792 (N_26792,N_26303,N_25942);
xnor U26793 (N_26793,N_26391,N_26192);
nor U26794 (N_26794,N_26358,N_26109);
nor U26795 (N_26795,N_26072,N_26326);
nor U26796 (N_26796,N_26145,N_26061);
xor U26797 (N_26797,N_25916,N_26291);
or U26798 (N_26798,N_25964,N_26330);
or U26799 (N_26799,N_26151,N_26290);
nand U26800 (N_26800,N_25898,N_26226);
nand U26801 (N_26801,N_26033,N_26179);
nor U26802 (N_26802,N_26277,N_26029);
or U26803 (N_26803,N_25946,N_26270);
nand U26804 (N_26804,N_25943,N_25993);
xor U26805 (N_26805,N_26318,N_26371);
nor U26806 (N_26806,N_26187,N_26164);
and U26807 (N_26807,N_26293,N_26244);
nand U26808 (N_26808,N_26083,N_26130);
and U26809 (N_26809,N_25831,N_26275);
xnor U26810 (N_26810,N_25891,N_26372);
nand U26811 (N_26811,N_25871,N_25875);
nor U26812 (N_26812,N_26388,N_26001);
and U26813 (N_26813,N_26315,N_26357);
nor U26814 (N_26814,N_26250,N_25832);
or U26815 (N_26815,N_25943,N_26178);
and U26816 (N_26816,N_26129,N_26218);
and U26817 (N_26817,N_25967,N_26259);
and U26818 (N_26818,N_25846,N_26276);
or U26819 (N_26819,N_25833,N_26378);
or U26820 (N_26820,N_25846,N_26129);
nand U26821 (N_26821,N_26321,N_26024);
or U26822 (N_26822,N_25942,N_26289);
xor U26823 (N_26823,N_26032,N_26110);
nor U26824 (N_26824,N_25832,N_26013);
xor U26825 (N_26825,N_25816,N_26109);
or U26826 (N_26826,N_25883,N_25923);
and U26827 (N_26827,N_25940,N_26212);
xnor U26828 (N_26828,N_26334,N_26343);
and U26829 (N_26829,N_26221,N_25949);
nor U26830 (N_26830,N_26293,N_26108);
nand U26831 (N_26831,N_26009,N_25956);
xnor U26832 (N_26832,N_25832,N_26045);
and U26833 (N_26833,N_26240,N_25947);
or U26834 (N_26834,N_26357,N_25924);
or U26835 (N_26835,N_25891,N_25990);
xor U26836 (N_26836,N_25950,N_25990);
and U26837 (N_26837,N_26271,N_26275);
nand U26838 (N_26838,N_26360,N_25805);
and U26839 (N_26839,N_26360,N_26137);
or U26840 (N_26840,N_26355,N_25996);
or U26841 (N_26841,N_25850,N_26304);
and U26842 (N_26842,N_25978,N_26291);
or U26843 (N_26843,N_25911,N_26011);
nand U26844 (N_26844,N_26218,N_26369);
and U26845 (N_26845,N_25806,N_25980);
xnor U26846 (N_26846,N_25976,N_25812);
nor U26847 (N_26847,N_26141,N_26000);
nor U26848 (N_26848,N_26144,N_26212);
nand U26849 (N_26849,N_26228,N_25813);
xor U26850 (N_26850,N_26227,N_25873);
xor U26851 (N_26851,N_25835,N_26253);
or U26852 (N_26852,N_26129,N_26350);
and U26853 (N_26853,N_26382,N_25985);
and U26854 (N_26854,N_25968,N_26288);
nand U26855 (N_26855,N_25845,N_26255);
xor U26856 (N_26856,N_26138,N_26038);
nand U26857 (N_26857,N_26354,N_26051);
or U26858 (N_26858,N_25961,N_26340);
nor U26859 (N_26859,N_26040,N_26143);
nor U26860 (N_26860,N_26372,N_26325);
nand U26861 (N_26861,N_26287,N_26276);
or U26862 (N_26862,N_26291,N_26163);
nor U26863 (N_26863,N_25948,N_26368);
nand U26864 (N_26864,N_26094,N_26048);
nand U26865 (N_26865,N_26283,N_26071);
or U26866 (N_26866,N_26120,N_26133);
and U26867 (N_26867,N_25821,N_26060);
or U26868 (N_26868,N_25866,N_25881);
nand U26869 (N_26869,N_26109,N_26183);
xor U26870 (N_26870,N_25925,N_26375);
nand U26871 (N_26871,N_26346,N_25983);
and U26872 (N_26872,N_26009,N_26241);
nand U26873 (N_26873,N_26257,N_25940);
or U26874 (N_26874,N_26043,N_25947);
xor U26875 (N_26875,N_26140,N_26242);
nor U26876 (N_26876,N_26131,N_25917);
or U26877 (N_26877,N_26314,N_26391);
nor U26878 (N_26878,N_26347,N_26361);
and U26879 (N_26879,N_25979,N_26011);
or U26880 (N_26880,N_26289,N_26151);
nor U26881 (N_26881,N_25993,N_26103);
nor U26882 (N_26882,N_26220,N_25895);
and U26883 (N_26883,N_26346,N_25857);
xnor U26884 (N_26884,N_26223,N_26315);
xnor U26885 (N_26885,N_26136,N_26323);
and U26886 (N_26886,N_26220,N_26353);
xnor U26887 (N_26887,N_25984,N_26367);
nor U26888 (N_26888,N_26049,N_26036);
xnor U26889 (N_26889,N_26115,N_26225);
or U26890 (N_26890,N_26257,N_26315);
nand U26891 (N_26891,N_26127,N_25887);
and U26892 (N_26892,N_25998,N_25914);
nand U26893 (N_26893,N_25954,N_26357);
and U26894 (N_26894,N_25870,N_26398);
nand U26895 (N_26895,N_25884,N_26109);
or U26896 (N_26896,N_26048,N_26022);
nor U26897 (N_26897,N_26252,N_25837);
nand U26898 (N_26898,N_26099,N_25865);
xor U26899 (N_26899,N_25977,N_26149);
nor U26900 (N_26900,N_26251,N_26383);
and U26901 (N_26901,N_26136,N_26217);
and U26902 (N_26902,N_26116,N_26206);
xor U26903 (N_26903,N_26072,N_26172);
nand U26904 (N_26904,N_26224,N_25916);
or U26905 (N_26905,N_26108,N_25861);
nand U26906 (N_26906,N_26214,N_26321);
or U26907 (N_26907,N_26203,N_26158);
xor U26908 (N_26908,N_26387,N_26018);
or U26909 (N_26909,N_26083,N_26380);
and U26910 (N_26910,N_26096,N_25930);
xnor U26911 (N_26911,N_26046,N_26273);
xnor U26912 (N_26912,N_26145,N_25917);
nor U26913 (N_26913,N_25896,N_26150);
or U26914 (N_26914,N_26251,N_26279);
nand U26915 (N_26915,N_25905,N_25823);
xor U26916 (N_26916,N_26109,N_26334);
nor U26917 (N_26917,N_26093,N_26182);
or U26918 (N_26918,N_26049,N_26290);
nor U26919 (N_26919,N_25927,N_26118);
or U26920 (N_26920,N_26278,N_25850);
xnor U26921 (N_26921,N_25892,N_26355);
nor U26922 (N_26922,N_26097,N_26100);
nand U26923 (N_26923,N_26046,N_26213);
nor U26924 (N_26924,N_26142,N_26012);
and U26925 (N_26925,N_26207,N_25977);
xnor U26926 (N_26926,N_26121,N_26011);
xnor U26927 (N_26927,N_26268,N_26177);
nand U26928 (N_26928,N_25912,N_26041);
xor U26929 (N_26929,N_26000,N_26113);
xnor U26930 (N_26930,N_25987,N_26275);
xor U26931 (N_26931,N_26116,N_26033);
nand U26932 (N_26932,N_26343,N_25962);
and U26933 (N_26933,N_26388,N_26060);
or U26934 (N_26934,N_26308,N_26224);
xnor U26935 (N_26935,N_25908,N_26223);
and U26936 (N_26936,N_26104,N_26226);
or U26937 (N_26937,N_26299,N_26362);
nor U26938 (N_26938,N_26005,N_26239);
and U26939 (N_26939,N_26013,N_26357);
nor U26940 (N_26940,N_25987,N_26065);
nand U26941 (N_26941,N_26134,N_26363);
nand U26942 (N_26942,N_26244,N_25822);
nor U26943 (N_26943,N_26072,N_25890);
and U26944 (N_26944,N_25980,N_26153);
nand U26945 (N_26945,N_26187,N_25959);
or U26946 (N_26946,N_26126,N_26086);
or U26947 (N_26947,N_25850,N_26100);
nand U26948 (N_26948,N_26152,N_26010);
or U26949 (N_26949,N_25990,N_26078);
nand U26950 (N_26950,N_26122,N_25892);
nand U26951 (N_26951,N_26262,N_26251);
and U26952 (N_26952,N_26160,N_26041);
nand U26953 (N_26953,N_26200,N_25947);
nor U26954 (N_26954,N_25887,N_26145);
xnor U26955 (N_26955,N_25960,N_26116);
nand U26956 (N_26956,N_26296,N_26351);
or U26957 (N_26957,N_26132,N_26124);
xnor U26958 (N_26958,N_26010,N_25820);
xnor U26959 (N_26959,N_26329,N_26362);
nor U26960 (N_26960,N_25878,N_25818);
nor U26961 (N_26961,N_25834,N_26161);
xnor U26962 (N_26962,N_25937,N_26174);
nand U26963 (N_26963,N_26366,N_26069);
xnor U26964 (N_26964,N_25883,N_26251);
nor U26965 (N_26965,N_25965,N_26220);
or U26966 (N_26966,N_26182,N_26340);
or U26967 (N_26967,N_26070,N_26119);
xnor U26968 (N_26968,N_25944,N_25907);
xnor U26969 (N_26969,N_26240,N_25998);
or U26970 (N_26970,N_26318,N_26112);
or U26971 (N_26971,N_26218,N_26288);
xnor U26972 (N_26972,N_26394,N_25988);
xnor U26973 (N_26973,N_25897,N_25842);
xnor U26974 (N_26974,N_26124,N_26000);
or U26975 (N_26975,N_25855,N_25803);
and U26976 (N_26976,N_25969,N_25840);
nand U26977 (N_26977,N_26392,N_25887);
nand U26978 (N_26978,N_25919,N_26291);
and U26979 (N_26979,N_26074,N_25897);
or U26980 (N_26980,N_26052,N_26353);
nor U26981 (N_26981,N_25965,N_26081);
or U26982 (N_26982,N_26190,N_26309);
xnor U26983 (N_26983,N_26268,N_25946);
and U26984 (N_26984,N_25881,N_26036);
or U26985 (N_26985,N_26133,N_26308);
and U26986 (N_26986,N_26235,N_26228);
or U26987 (N_26987,N_26070,N_26148);
or U26988 (N_26988,N_26118,N_25911);
nand U26989 (N_26989,N_25937,N_26157);
nor U26990 (N_26990,N_26115,N_25869);
nor U26991 (N_26991,N_25881,N_26299);
or U26992 (N_26992,N_25856,N_26317);
xor U26993 (N_26993,N_26147,N_25879);
xnor U26994 (N_26994,N_26092,N_25888);
nor U26995 (N_26995,N_26172,N_26249);
and U26996 (N_26996,N_25928,N_26196);
nor U26997 (N_26997,N_26117,N_25992);
nor U26998 (N_26998,N_26253,N_26392);
and U26999 (N_26999,N_25980,N_26358);
and U27000 (N_27000,N_26460,N_26809);
nor U27001 (N_27001,N_26626,N_26803);
or U27002 (N_27002,N_26901,N_26814);
xnor U27003 (N_27003,N_26978,N_26605);
nand U27004 (N_27004,N_26417,N_26604);
and U27005 (N_27005,N_26880,N_26671);
and U27006 (N_27006,N_26829,N_26662);
xor U27007 (N_27007,N_26816,N_26543);
and U27008 (N_27008,N_26861,N_26429);
xor U27009 (N_27009,N_26983,N_26697);
nand U27010 (N_27010,N_26629,N_26572);
or U27011 (N_27011,N_26536,N_26775);
nor U27012 (N_27012,N_26591,N_26782);
nor U27013 (N_27013,N_26593,N_26456);
xor U27014 (N_27014,N_26638,N_26815);
and U27015 (N_27015,N_26449,N_26810);
nand U27016 (N_27016,N_26923,N_26461);
nand U27017 (N_27017,N_26806,N_26874);
or U27018 (N_27018,N_26871,N_26989);
nand U27019 (N_27019,N_26661,N_26421);
or U27020 (N_27020,N_26703,N_26792);
nor U27021 (N_27021,N_26659,N_26476);
nand U27022 (N_27022,N_26800,N_26678);
or U27023 (N_27023,N_26700,N_26467);
xnor U27024 (N_27024,N_26845,N_26484);
and U27025 (N_27025,N_26496,N_26439);
nand U27026 (N_27026,N_26905,N_26975);
xor U27027 (N_27027,N_26440,N_26793);
nand U27028 (N_27028,N_26674,N_26633);
or U27029 (N_27029,N_26480,N_26699);
xnor U27030 (N_27030,N_26723,N_26839);
or U27031 (N_27031,N_26881,N_26549);
or U27032 (N_27032,N_26615,N_26527);
nand U27033 (N_27033,N_26813,N_26928);
or U27034 (N_27034,N_26414,N_26955);
nor U27035 (N_27035,N_26812,N_26487);
and U27036 (N_27036,N_26644,N_26654);
and U27037 (N_27037,N_26739,N_26610);
nand U27038 (N_27038,N_26569,N_26450);
or U27039 (N_27039,N_26623,N_26867);
nand U27040 (N_27040,N_26832,N_26885);
and U27041 (N_27041,N_26892,N_26665);
xor U27042 (N_27042,N_26838,N_26943);
or U27043 (N_27043,N_26734,N_26481);
nand U27044 (N_27044,N_26762,N_26941);
and U27045 (N_27045,N_26670,N_26701);
nor U27046 (N_27046,N_26755,N_26620);
xor U27047 (N_27047,N_26986,N_26448);
and U27048 (N_27048,N_26799,N_26691);
or U27049 (N_27049,N_26576,N_26869);
or U27050 (N_27050,N_26916,N_26730);
nand U27051 (N_27051,N_26824,N_26733);
and U27052 (N_27052,N_26817,N_26937);
nor U27053 (N_27053,N_26791,N_26987);
xor U27054 (N_27054,N_26575,N_26835);
nand U27055 (N_27055,N_26447,N_26926);
or U27056 (N_27056,N_26432,N_26742);
nand U27057 (N_27057,N_26876,N_26980);
xor U27058 (N_27058,N_26663,N_26781);
nand U27059 (N_27059,N_26551,N_26680);
and U27060 (N_27060,N_26634,N_26795);
and U27061 (N_27061,N_26667,N_26935);
nor U27062 (N_27062,N_26961,N_26836);
nand U27063 (N_27063,N_26878,N_26993);
xor U27064 (N_27064,N_26495,N_26431);
xor U27065 (N_27065,N_26848,N_26820);
or U27066 (N_27066,N_26519,N_26950);
or U27067 (N_27067,N_26526,N_26681);
nor U27068 (N_27068,N_26466,N_26853);
nor U27069 (N_27069,N_26798,N_26963);
xnor U27070 (N_27070,N_26426,N_26979);
xnor U27071 (N_27071,N_26868,N_26511);
or U27072 (N_27072,N_26607,N_26718);
nor U27073 (N_27073,N_26947,N_26463);
nand U27074 (N_27074,N_26954,N_26532);
xnor U27075 (N_27075,N_26521,N_26689);
and U27076 (N_27076,N_26632,N_26875);
nand U27077 (N_27077,N_26606,N_26584);
nor U27078 (N_27078,N_26690,N_26693);
xnor U27079 (N_27079,N_26722,N_26617);
xor U27080 (N_27080,N_26725,N_26995);
nand U27081 (N_27081,N_26994,N_26927);
or U27082 (N_27082,N_26917,N_26866);
nand U27083 (N_27083,N_26631,N_26929);
and U27084 (N_27084,N_26474,N_26554);
and U27085 (N_27085,N_26915,N_26946);
xor U27086 (N_27086,N_26919,N_26957);
or U27087 (N_27087,N_26992,N_26534);
nor U27088 (N_27088,N_26563,N_26602);
nand U27089 (N_27089,N_26906,N_26523);
xnor U27090 (N_27090,N_26862,N_26828);
nor U27091 (N_27091,N_26408,N_26752);
nor U27092 (N_27092,N_26592,N_26642);
nor U27093 (N_27093,N_26548,N_26647);
nor U27094 (N_27094,N_26415,N_26964);
nor U27095 (N_27095,N_26764,N_26854);
nand U27096 (N_27096,N_26514,N_26518);
nand U27097 (N_27097,N_26985,N_26489);
nand U27098 (N_27098,N_26958,N_26488);
xor U27099 (N_27099,N_26545,N_26404);
and U27100 (N_27100,N_26959,N_26786);
xnor U27101 (N_27101,N_26750,N_26458);
xnor U27102 (N_27102,N_26419,N_26894);
nor U27103 (N_27103,N_26687,N_26745);
nor U27104 (N_27104,N_26729,N_26754);
nand U27105 (N_27105,N_26870,N_26483);
xnor U27106 (N_27106,N_26688,N_26619);
or U27107 (N_27107,N_26973,N_26641);
xnor U27108 (N_27108,N_26589,N_26998);
xnor U27109 (N_27109,N_26865,N_26682);
or U27110 (N_27110,N_26597,N_26857);
nand U27111 (N_27111,N_26457,N_26863);
and U27112 (N_27112,N_26413,N_26897);
and U27113 (N_27113,N_26909,N_26879);
or U27114 (N_27114,N_26451,N_26822);
or U27115 (N_27115,N_26847,N_26564);
xor U27116 (N_27116,N_26706,N_26833);
nand U27117 (N_27117,N_26970,N_26837);
nor U27118 (N_27118,N_26753,N_26741);
nand U27119 (N_27119,N_26748,N_26492);
nor U27120 (N_27120,N_26477,N_26603);
and U27121 (N_27121,N_26738,N_26613);
or U27122 (N_27122,N_26900,N_26911);
xnor U27123 (N_27123,N_26541,N_26473);
or U27124 (N_27124,N_26819,N_26912);
or U27125 (N_27125,N_26506,N_26491);
and U27126 (N_27126,N_26807,N_26988);
xor U27127 (N_27127,N_26616,N_26645);
xor U27128 (N_27128,N_26960,N_26784);
nor U27129 (N_27129,N_26601,N_26965);
and U27130 (N_27130,N_26747,N_26858);
and U27131 (N_27131,N_26756,N_26657);
or U27132 (N_27132,N_26882,N_26403);
and U27133 (N_27133,N_26522,N_26804);
nor U27134 (N_27134,N_26648,N_26560);
and U27135 (N_27135,N_26708,N_26737);
xor U27136 (N_27136,N_26405,N_26702);
nor U27137 (N_27137,N_26427,N_26547);
xnor U27138 (N_27138,N_26772,N_26850);
and U27139 (N_27139,N_26400,N_26505);
nor U27140 (N_27140,N_26893,N_26864);
nor U27141 (N_27141,N_26728,N_26751);
and U27142 (N_27142,N_26410,N_26425);
or U27143 (N_27143,N_26771,N_26468);
nand U27144 (N_27144,N_26778,N_26446);
xnor U27145 (N_27145,N_26889,N_26797);
nor U27146 (N_27146,N_26504,N_26827);
xnor U27147 (N_27147,N_26517,N_26479);
and U27148 (N_27148,N_26673,N_26558);
nand U27149 (N_27149,N_26579,N_26577);
and U27150 (N_27150,N_26774,N_26790);
and U27151 (N_27151,N_26783,N_26769);
and U27152 (N_27152,N_26501,N_26692);
nor U27153 (N_27153,N_26422,N_26945);
nor U27154 (N_27154,N_26891,N_26789);
xor U27155 (N_27155,N_26933,N_26887);
nand U27156 (N_27156,N_26573,N_26849);
nand U27157 (N_27157,N_26788,N_26555);
nor U27158 (N_27158,N_26704,N_26490);
and U27159 (N_27159,N_26493,N_26976);
nor U27160 (N_27160,N_26513,N_26840);
or U27161 (N_27161,N_26581,N_26904);
xnor U27162 (N_27162,N_26903,N_26852);
nand U27163 (N_27163,N_26713,N_26780);
or U27164 (N_27164,N_26842,N_26561);
nand U27165 (N_27165,N_26851,N_26720);
nor U27166 (N_27166,N_26726,N_26990);
xnor U27167 (N_27167,N_26650,N_26643);
nand U27168 (N_27168,N_26808,N_26924);
nand U27169 (N_27169,N_26818,N_26503);
nor U27170 (N_27170,N_26635,N_26760);
nand U27171 (N_27171,N_26719,N_26763);
and U27172 (N_27172,N_26888,N_26707);
xor U27173 (N_27173,N_26710,N_26509);
and U27174 (N_27174,N_26890,N_26658);
nor U27175 (N_27175,N_26464,N_26767);
and U27176 (N_27176,N_26416,N_26672);
or U27177 (N_27177,N_26843,N_26776);
or U27178 (N_27178,N_26434,N_26676);
or U27179 (N_27179,N_26736,N_26420);
xor U27180 (N_27180,N_26469,N_26735);
xor U27181 (N_27181,N_26971,N_26936);
xnor U27182 (N_27182,N_26907,N_26566);
nand U27183 (N_27183,N_26996,N_26991);
and U27184 (N_27184,N_26609,N_26831);
nand U27185 (N_27185,N_26465,N_26587);
and U27186 (N_27186,N_26582,N_26454);
nor U27187 (N_27187,N_26859,N_26442);
and U27188 (N_27188,N_26430,N_26724);
xor U27189 (N_27189,N_26452,N_26721);
nand U27190 (N_27190,N_26540,N_26872);
xor U27191 (N_27191,N_26552,N_26533);
and U27192 (N_27192,N_26627,N_26622);
and U27193 (N_27193,N_26608,N_26500);
xor U27194 (N_27194,N_26712,N_26770);
nor U27195 (N_27195,N_26925,N_26402);
xnor U27196 (N_27196,N_26600,N_26761);
or U27197 (N_27197,N_26482,N_26899);
xnor U27198 (N_27198,N_26588,N_26445);
nand U27199 (N_27199,N_26811,N_26938);
xor U27200 (N_27200,N_26590,N_26636);
nand U27201 (N_27201,N_26982,N_26424);
nand U27202 (N_27202,N_26732,N_26834);
nand U27203 (N_27203,N_26972,N_26966);
and U27204 (N_27204,N_26779,N_26981);
nor U27205 (N_27205,N_26433,N_26902);
and U27206 (N_27206,N_26908,N_26698);
nor U27207 (N_27207,N_26438,N_26746);
and U27208 (N_27208,N_26516,N_26759);
and U27209 (N_27209,N_26614,N_26580);
nand U27210 (N_27210,N_26666,N_26498);
or U27211 (N_27211,N_26727,N_26535);
xor U27212 (N_27212,N_26567,N_26951);
nor U27213 (N_27213,N_26655,N_26565);
or U27214 (N_27214,N_26939,N_26830);
xor U27215 (N_27215,N_26595,N_26715);
and U27216 (N_27216,N_26695,N_26462);
nor U27217 (N_27217,N_26896,N_26962);
nand U27218 (N_27218,N_26537,N_26794);
nand U27219 (N_27219,N_26969,N_26823);
nand U27220 (N_27220,N_26956,N_26883);
xnor U27221 (N_27221,N_26624,N_26967);
and U27222 (N_27222,N_26437,N_26884);
nor U27223 (N_27223,N_26409,N_26436);
xor U27224 (N_27224,N_26596,N_26873);
or U27225 (N_27225,N_26539,N_26570);
nor U27226 (N_27226,N_26546,N_26639);
or U27227 (N_27227,N_26844,N_26948);
and U27228 (N_27228,N_26646,N_26401);
or U27229 (N_27229,N_26583,N_26918);
or U27230 (N_27230,N_26705,N_26997);
and U27231 (N_27231,N_26944,N_26423);
or U27232 (N_27232,N_26675,N_26625);
and U27233 (N_27233,N_26418,N_26621);
xnor U27234 (N_27234,N_26556,N_26685);
nor U27235 (N_27235,N_26709,N_26716);
and U27236 (N_27236,N_26777,N_26796);
xnor U27237 (N_27237,N_26898,N_26411);
nand U27238 (N_27238,N_26571,N_26711);
xor U27239 (N_27239,N_26984,N_26766);
and U27240 (N_27240,N_26512,N_26562);
and U27241 (N_27241,N_26668,N_26550);
xnor U27242 (N_27242,N_26921,N_26508);
nor U27243 (N_27243,N_26441,N_26931);
xnor U27244 (N_27244,N_26686,N_26640);
or U27245 (N_27245,N_26757,N_26826);
and U27246 (N_27246,N_26660,N_26664);
and U27247 (N_27247,N_26805,N_26758);
nor U27248 (N_27248,N_26968,N_26773);
nand U27249 (N_27249,N_26694,N_26598);
and U27250 (N_27250,N_26542,N_26412);
and U27251 (N_27251,N_26740,N_26507);
xor U27252 (N_27252,N_26855,N_26949);
or U27253 (N_27253,N_26649,N_26841);
xor U27254 (N_27254,N_26920,N_26630);
nand U27255 (N_27255,N_26744,N_26628);
nand U27256 (N_27256,N_26435,N_26557);
xnor U27257 (N_27257,N_26914,N_26652);
nand U27258 (N_27258,N_26942,N_26406);
xor U27259 (N_27259,N_26765,N_26787);
nor U27260 (N_27260,N_26599,N_26677);
nor U27261 (N_27261,N_26856,N_26453);
or U27262 (N_27262,N_26821,N_26611);
and U27263 (N_27263,N_26877,N_26802);
nor U27264 (N_27264,N_26651,N_26485);
nand U27265 (N_27265,N_26524,N_26612);
xnor U27266 (N_27266,N_26717,N_26801);
nand U27267 (N_27267,N_26714,N_26679);
and U27268 (N_27268,N_26502,N_26472);
nor U27269 (N_27269,N_26684,N_26768);
or U27270 (N_27270,N_26559,N_26499);
nand U27271 (N_27271,N_26696,N_26578);
nor U27272 (N_27272,N_26913,N_26922);
or U27273 (N_27273,N_26940,N_26637);
and U27274 (N_27274,N_26656,N_26749);
xnor U27275 (N_27275,N_26455,N_26515);
or U27276 (N_27276,N_26618,N_26531);
nand U27277 (N_27277,N_26977,N_26785);
xor U27278 (N_27278,N_26444,N_26910);
and U27279 (N_27279,N_26860,N_26825);
nor U27280 (N_27280,N_26934,N_26528);
xnor U27281 (N_27281,N_26553,N_26594);
nand U27282 (N_27282,N_26475,N_26529);
nand U27283 (N_27283,N_26846,N_26530);
or U27284 (N_27284,N_26653,N_26470);
and U27285 (N_27285,N_26568,N_26525);
xnor U27286 (N_27286,N_26443,N_26520);
nor U27287 (N_27287,N_26974,N_26494);
or U27288 (N_27288,N_26478,N_26731);
and U27289 (N_27289,N_26486,N_26683);
xor U27290 (N_27290,N_26497,N_26471);
or U27291 (N_27291,N_26407,N_26743);
nor U27292 (N_27292,N_26544,N_26538);
or U27293 (N_27293,N_26428,N_26952);
or U27294 (N_27294,N_26999,N_26510);
nand U27295 (N_27295,N_26886,N_26895);
nor U27296 (N_27296,N_26586,N_26930);
nor U27297 (N_27297,N_26932,N_26669);
and U27298 (N_27298,N_26585,N_26953);
nand U27299 (N_27299,N_26459,N_26574);
and U27300 (N_27300,N_26585,N_26996);
nand U27301 (N_27301,N_26714,N_26795);
or U27302 (N_27302,N_26796,N_26846);
xnor U27303 (N_27303,N_26681,N_26705);
xnor U27304 (N_27304,N_26573,N_26806);
xor U27305 (N_27305,N_26869,N_26556);
nand U27306 (N_27306,N_26744,N_26466);
xnor U27307 (N_27307,N_26646,N_26741);
or U27308 (N_27308,N_26805,N_26950);
xnor U27309 (N_27309,N_26842,N_26933);
nor U27310 (N_27310,N_26717,N_26798);
nand U27311 (N_27311,N_26945,N_26409);
xnor U27312 (N_27312,N_26464,N_26695);
nor U27313 (N_27313,N_26626,N_26919);
and U27314 (N_27314,N_26748,N_26563);
nor U27315 (N_27315,N_26868,N_26624);
nand U27316 (N_27316,N_26997,N_26495);
or U27317 (N_27317,N_26825,N_26771);
xnor U27318 (N_27318,N_26799,N_26952);
nor U27319 (N_27319,N_26702,N_26766);
or U27320 (N_27320,N_26495,N_26589);
xnor U27321 (N_27321,N_26921,N_26801);
nand U27322 (N_27322,N_26759,N_26908);
and U27323 (N_27323,N_26831,N_26900);
nor U27324 (N_27324,N_26829,N_26972);
nor U27325 (N_27325,N_26629,N_26947);
and U27326 (N_27326,N_26537,N_26922);
nand U27327 (N_27327,N_26948,N_26487);
nor U27328 (N_27328,N_26962,N_26634);
nor U27329 (N_27329,N_26762,N_26417);
and U27330 (N_27330,N_26940,N_26984);
or U27331 (N_27331,N_26422,N_26589);
or U27332 (N_27332,N_26537,N_26452);
nand U27333 (N_27333,N_26776,N_26548);
and U27334 (N_27334,N_26890,N_26766);
nor U27335 (N_27335,N_26630,N_26742);
nand U27336 (N_27336,N_26404,N_26641);
nor U27337 (N_27337,N_26770,N_26822);
or U27338 (N_27338,N_26495,N_26791);
xnor U27339 (N_27339,N_26648,N_26866);
nor U27340 (N_27340,N_26802,N_26975);
nor U27341 (N_27341,N_26636,N_26977);
xor U27342 (N_27342,N_26664,N_26590);
or U27343 (N_27343,N_26527,N_26439);
or U27344 (N_27344,N_26482,N_26545);
xnor U27345 (N_27345,N_26836,N_26969);
nor U27346 (N_27346,N_26441,N_26540);
or U27347 (N_27347,N_26733,N_26747);
or U27348 (N_27348,N_26991,N_26932);
and U27349 (N_27349,N_26966,N_26629);
nand U27350 (N_27350,N_26533,N_26911);
nor U27351 (N_27351,N_26641,N_26717);
xnor U27352 (N_27352,N_26408,N_26994);
or U27353 (N_27353,N_26449,N_26588);
or U27354 (N_27354,N_26518,N_26555);
and U27355 (N_27355,N_26803,N_26545);
and U27356 (N_27356,N_26759,N_26428);
xor U27357 (N_27357,N_26995,N_26452);
and U27358 (N_27358,N_26579,N_26981);
and U27359 (N_27359,N_26649,N_26755);
nor U27360 (N_27360,N_26668,N_26954);
and U27361 (N_27361,N_26663,N_26437);
nor U27362 (N_27362,N_26489,N_26590);
or U27363 (N_27363,N_26573,N_26435);
or U27364 (N_27364,N_26625,N_26712);
nor U27365 (N_27365,N_26837,N_26666);
xor U27366 (N_27366,N_26408,N_26469);
or U27367 (N_27367,N_26573,N_26954);
nor U27368 (N_27368,N_26412,N_26988);
or U27369 (N_27369,N_26670,N_26536);
or U27370 (N_27370,N_26628,N_26654);
or U27371 (N_27371,N_26604,N_26471);
or U27372 (N_27372,N_26549,N_26695);
or U27373 (N_27373,N_26878,N_26893);
or U27374 (N_27374,N_26644,N_26412);
or U27375 (N_27375,N_26975,N_26484);
xnor U27376 (N_27376,N_26620,N_26659);
or U27377 (N_27377,N_26622,N_26680);
or U27378 (N_27378,N_26510,N_26735);
and U27379 (N_27379,N_26737,N_26437);
and U27380 (N_27380,N_26884,N_26441);
nor U27381 (N_27381,N_26536,N_26852);
and U27382 (N_27382,N_26926,N_26780);
nand U27383 (N_27383,N_26546,N_26448);
nor U27384 (N_27384,N_26930,N_26991);
nor U27385 (N_27385,N_26406,N_26420);
xnor U27386 (N_27386,N_26469,N_26918);
and U27387 (N_27387,N_26623,N_26840);
or U27388 (N_27388,N_26801,N_26813);
and U27389 (N_27389,N_26795,N_26857);
or U27390 (N_27390,N_26992,N_26568);
nand U27391 (N_27391,N_26872,N_26500);
or U27392 (N_27392,N_26547,N_26426);
nor U27393 (N_27393,N_26858,N_26939);
and U27394 (N_27394,N_26924,N_26682);
nand U27395 (N_27395,N_26781,N_26786);
nor U27396 (N_27396,N_26688,N_26589);
nand U27397 (N_27397,N_26542,N_26740);
or U27398 (N_27398,N_26501,N_26871);
nor U27399 (N_27399,N_26492,N_26548);
and U27400 (N_27400,N_26489,N_26677);
xor U27401 (N_27401,N_26523,N_26571);
xnor U27402 (N_27402,N_26444,N_26843);
nor U27403 (N_27403,N_26707,N_26668);
nand U27404 (N_27404,N_26505,N_26670);
or U27405 (N_27405,N_26961,N_26987);
and U27406 (N_27406,N_26896,N_26701);
nand U27407 (N_27407,N_26519,N_26771);
or U27408 (N_27408,N_26794,N_26471);
and U27409 (N_27409,N_26547,N_26430);
xnor U27410 (N_27410,N_26973,N_26954);
xnor U27411 (N_27411,N_26851,N_26955);
xnor U27412 (N_27412,N_26723,N_26943);
xnor U27413 (N_27413,N_26909,N_26439);
and U27414 (N_27414,N_26486,N_26482);
or U27415 (N_27415,N_26775,N_26543);
xnor U27416 (N_27416,N_26646,N_26635);
xor U27417 (N_27417,N_26401,N_26536);
nand U27418 (N_27418,N_26930,N_26488);
nand U27419 (N_27419,N_26725,N_26879);
xor U27420 (N_27420,N_26630,N_26487);
and U27421 (N_27421,N_26900,N_26615);
xnor U27422 (N_27422,N_26410,N_26585);
and U27423 (N_27423,N_26512,N_26819);
or U27424 (N_27424,N_26988,N_26882);
nor U27425 (N_27425,N_26871,N_26862);
nand U27426 (N_27426,N_26598,N_26660);
or U27427 (N_27427,N_26653,N_26648);
and U27428 (N_27428,N_26832,N_26989);
and U27429 (N_27429,N_26778,N_26790);
nand U27430 (N_27430,N_26873,N_26839);
xor U27431 (N_27431,N_26737,N_26593);
nand U27432 (N_27432,N_26440,N_26410);
and U27433 (N_27433,N_26885,N_26530);
xnor U27434 (N_27434,N_26541,N_26905);
xor U27435 (N_27435,N_26676,N_26411);
nand U27436 (N_27436,N_26748,N_26819);
or U27437 (N_27437,N_26481,N_26820);
and U27438 (N_27438,N_26697,N_26543);
and U27439 (N_27439,N_26659,N_26768);
nor U27440 (N_27440,N_26972,N_26438);
or U27441 (N_27441,N_26720,N_26583);
nor U27442 (N_27442,N_26558,N_26676);
or U27443 (N_27443,N_26465,N_26685);
nand U27444 (N_27444,N_26567,N_26418);
xor U27445 (N_27445,N_26706,N_26796);
xnor U27446 (N_27446,N_26970,N_26888);
or U27447 (N_27447,N_26838,N_26420);
or U27448 (N_27448,N_26845,N_26607);
xnor U27449 (N_27449,N_26919,N_26744);
nand U27450 (N_27450,N_26889,N_26660);
nor U27451 (N_27451,N_26523,N_26910);
xnor U27452 (N_27452,N_26883,N_26991);
xnor U27453 (N_27453,N_26785,N_26472);
xnor U27454 (N_27454,N_26828,N_26896);
or U27455 (N_27455,N_26711,N_26883);
and U27456 (N_27456,N_26736,N_26724);
nand U27457 (N_27457,N_26561,N_26931);
or U27458 (N_27458,N_26796,N_26426);
nor U27459 (N_27459,N_26401,N_26884);
xnor U27460 (N_27460,N_26673,N_26481);
xnor U27461 (N_27461,N_26556,N_26432);
xnor U27462 (N_27462,N_26577,N_26978);
nor U27463 (N_27463,N_26482,N_26630);
nor U27464 (N_27464,N_26448,N_26502);
xor U27465 (N_27465,N_26796,N_26862);
and U27466 (N_27466,N_26608,N_26774);
and U27467 (N_27467,N_26868,N_26930);
xnor U27468 (N_27468,N_26753,N_26715);
xnor U27469 (N_27469,N_26602,N_26548);
or U27470 (N_27470,N_26828,N_26560);
nand U27471 (N_27471,N_26673,N_26725);
nor U27472 (N_27472,N_26872,N_26897);
nor U27473 (N_27473,N_26601,N_26853);
xnor U27474 (N_27474,N_26685,N_26686);
or U27475 (N_27475,N_26733,N_26558);
and U27476 (N_27476,N_26846,N_26753);
nor U27477 (N_27477,N_26451,N_26910);
and U27478 (N_27478,N_26431,N_26824);
nand U27479 (N_27479,N_26654,N_26527);
nor U27480 (N_27480,N_26668,N_26702);
and U27481 (N_27481,N_26783,N_26439);
or U27482 (N_27482,N_26455,N_26604);
nand U27483 (N_27483,N_26941,N_26917);
and U27484 (N_27484,N_26831,N_26891);
or U27485 (N_27485,N_26811,N_26997);
or U27486 (N_27486,N_26506,N_26864);
nand U27487 (N_27487,N_26436,N_26558);
or U27488 (N_27488,N_26502,N_26641);
xnor U27489 (N_27489,N_26836,N_26955);
nor U27490 (N_27490,N_26654,N_26499);
xnor U27491 (N_27491,N_26497,N_26704);
xnor U27492 (N_27492,N_26914,N_26723);
and U27493 (N_27493,N_26782,N_26958);
and U27494 (N_27494,N_26684,N_26517);
or U27495 (N_27495,N_26550,N_26884);
xnor U27496 (N_27496,N_26810,N_26930);
or U27497 (N_27497,N_26715,N_26889);
nand U27498 (N_27498,N_26944,N_26629);
and U27499 (N_27499,N_26768,N_26789);
nand U27500 (N_27500,N_26989,N_26533);
nand U27501 (N_27501,N_26675,N_26654);
or U27502 (N_27502,N_26940,N_26948);
and U27503 (N_27503,N_26819,N_26654);
xor U27504 (N_27504,N_26794,N_26688);
nand U27505 (N_27505,N_26960,N_26880);
or U27506 (N_27506,N_26645,N_26988);
or U27507 (N_27507,N_26981,N_26499);
or U27508 (N_27508,N_26860,N_26481);
or U27509 (N_27509,N_26503,N_26738);
xor U27510 (N_27510,N_26467,N_26415);
xnor U27511 (N_27511,N_26796,N_26510);
and U27512 (N_27512,N_26842,N_26975);
xor U27513 (N_27513,N_26854,N_26735);
or U27514 (N_27514,N_26602,N_26516);
nand U27515 (N_27515,N_26854,N_26622);
xor U27516 (N_27516,N_26864,N_26656);
nor U27517 (N_27517,N_26874,N_26575);
nor U27518 (N_27518,N_26451,N_26670);
nor U27519 (N_27519,N_26975,N_26779);
xnor U27520 (N_27520,N_26539,N_26719);
nor U27521 (N_27521,N_26709,N_26552);
nor U27522 (N_27522,N_26883,N_26568);
or U27523 (N_27523,N_26887,N_26897);
and U27524 (N_27524,N_26846,N_26456);
and U27525 (N_27525,N_26479,N_26775);
xor U27526 (N_27526,N_26446,N_26478);
nand U27527 (N_27527,N_26967,N_26990);
nand U27528 (N_27528,N_26605,N_26571);
nor U27529 (N_27529,N_26800,N_26989);
nor U27530 (N_27530,N_26654,N_26930);
nand U27531 (N_27531,N_26712,N_26492);
and U27532 (N_27532,N_26708,N_26746);
nand U27533 (N_27533,N_26975,N_26663);
xor U27534 (N_27534,N_26550,N_26569);
or U27535 (N_27535,N_26546,N_26913);
nand U27536 (N_27536,N_26782,N_26779);
nor U27537 (N_27537,N_26692,N_26935);
xor U27538 (N_27538,N_26606,N_26615);
nand U27539 (N_27539,N_26608,N_26507);
xor U27540 (N_27540,N_26415,N_26400);
nor U27541 (N_27541,N_26409,N_26980);
nand U27542 (N_27542,N_26585,N_26565);
and U27543 (N_27543,N_26765,N_26509);
nor U27544 (N_27544,N_26837,N_26961);
or U27545 (N_27545,N_26535,N_26673);
xor U27546 (N_27546,N_26822,N_26578);
nor U27547 (N_27547,N_26527,N_26636);
and U27548 (N_27548,N_26994,N_26924);
nand U27549 (N_27549,N_26976,N_26984);
nor U27550 (N_27550,N_26688,N_26502);
or U27551 (N_27551,N_26408,N_26589);
or U27552 (N_27552,N_26797,N_26733);
xor U27553 (N_27553,N_26553,N_26763);
and U27554 (N_27554,N_26625,N_26782);
and U27555 (N_27555,N_26811,N_26960);
nand U27556 (N_27556,N_26752,N_26599);
nor U27557 (N_27557,N_26643,N_26985);
or U27558 (N_27558,N_26529,N_26878);
and U27559 (N_27559,N_26964,N_26841);
xnor U27560 (N_27560,N_26684,N_26444);
nand U27561 (N_27561,N_26880,N_26820);
xor U27562 (N_27562,N_26553,N_26417);
xnor U27563 (N_27563,N_26716,N_26851);
nand U27564 (N_27564,N_26436,N_26484);
or U27565 (N_27565,N_26556,N_26471);
nand U27566 (N_27566,N_26911,N_26870);
and U27567 (N_27567,N_26565,N_26966);
and U27568 (N_27568,N_26696,N_26683);
nor U27569 (N_27569,N_26968,N_26722);
and U27570 (N_27570,N_26429,N_26565);
nand U27571 (N_27571,N_26962,N_26945);
nand U27572 (N_27572,N_26847,N_26827);
and U27573 (N_27573,N_26548,N_26926);
and U27574 (N_27574,N_26720,N_26410);
and U27575 (N_27575,N_26675,N_26665);
nand U27576 (N_27576,N_26447,N_26779);
and U27577 (N_27577,N_26534,N_26570);
nand U27578 (N_27578,N_26547,N_26858);
xor U27579 (N_27579,N_26684,N_26767);
nand U27580 (N_27580,N_26592,N_26735);
nand U27581 (N_27581,N_26958,N_26518);
xor U27582 (N_27582,N_26597,N_26895);
or U27583 (N_27583,N_26915,N_26869);
xnor U27584 (N_27584,N_26549,N_26694);
nand U27585 (N_27585,N_26746,N_26794);
nor U27586 (N_27586,N_26508,N_26745);
nor U27587 (N_27587,N_26984,N_26866);
or U27588 (N_27588,N_26596,N_26540);
nor U27589 (N_27589,N_26854,N_26948);
xnor U27590 (N_27590,N_26530,N_26840);
xor U27591 (N_27591,N_26410,N_26855);
xor U27592 (N_27592,N_26986,N_26489);
xnor U27593 (N_27593,N_26432,N_26837);
or U27594 (N_27594,N_26415,N_26619);
nand U27595 (N_27595,N_26415,N_26566);
or U27596 (N_27596,N_26733,N_26664);
and U27597 (N_27597,N_26999,N_26787);
nor U27598 (N_27598,N_26988,N_26639);
nand U27599 (N_27599,N_26746,N_26694);
or U27600 (N_27600,N_27451,N_27272);
or U27601 (N_27601,N_27439,N_27418);
and U27602 (N_27602,N_27155,N_27357);
nor U27603 (N_27603,N_27146,N_27480);
xnor U27604 (N_27604,N_27369,N_27566);
or U27605 (N_27605,N_27364,N_27569);
and U27606 (N_27606,N_27118,N_27564);
nand U27607 (N_27607,N_27406,N_27456);
nor U27608 (N_27608,N_27592,N_27404);
nor U27609 (N_27609,N_27527,N_27265);
or U27610 (N_27610,N_27213,N_27013);
nand U27611 (N_27611,N_27004,N_27572);
or U27612 (N_27612,N_27154,N_27303);
or U27613 (N_27613,N_27542,N_27548);
and U27614 (N_27614,N_27224,N_27356);
and U27615 (N_27615,N_27061,N_27092);
nand U27616 (N_27616,N_27143,N_27546);
xnor U27617 (N_27617,N_27574,N_27120);
nor U27618 (N_27618,N_27207,N_27014);
nand U27619 (N_27619,N_27071,N_27163);
and U27620 (N_27620,N_27295,N_27308);
nor U27621 (N_27621,N_27386,N_27249);
or U27622 (N_27622,N_27210,N_27433);
nand U27623 (N_27623,N_27245,N_27305);
xnor U27624 (N_27624,N_27240,N_27492);
and U27625 (N_27625,N_27286,N_27475);
xor U27626 (N_27626,N_27105,N_27445);
nand U27627 (N_27627,N_27595,N_27549);
nor U27628 (N_27628,N_27132,N_27577);
and U27629 (N_27629,N_27257,N_27522);
nand U27630 (N_27630,N_27221,N_27327);
nand U27631 (N_27631,N_27168,N_27464);
and U27632 (N_27632,N_27270,N_27023);
nor U27633 (N_27633,N_27230,N_27331);
xnor U27634 (N_27634,N_27581,N_27258);
or U27635 (N_27635,N_27485,N_27088);
nand U27636 (N_27636,N_27506,N_27159);
nand U27637 (N_27637,N_27409,N_27179);
xnor U27638 (N_27638,N_27236,N_27205);
and U27639 (N_27639,N_27232,N_27248);
or U27640 (N_27640,N_27174,N_27370);
or U27641 (N_27641,N_27353,N_27568);
nor U27642 (N_27642,N_27276,N_27244);
nand U27643 (N_27643,N_27080,N_27218);
nand U27644 (N_27644,N_27043,N_27314);
nand U27645 (N_27645,N_27556,N_27422);
nor U27646 (N_27646,N_27411,N_27429);
and U27647 (N_27647,N_27032,N_27002);
and U27648 (N_27648,N_27341,N_27339);
nand U27649 (N_27649,N_27321,N_27028);
nor U27650 (N_27650,N_27098,N_27338);
and U27651 (N_27651,N_27350,N_27503);
or U27652 (N_27652,N_27500,N_27366);
and U27653 (N_27653,N_27598,N_27121);
nor U27654 (N_27654,N_27125,N_27173);
or U27655 (N_27655,N_27047,N_27045);
nor U27656 (N_27656,N_27320,N_27130);
and U27657 (N_27657,N_27046,N_27016);
nand U27658 (N_27658,N_27246,N_27507);
nand U27659 (N_27659,N_27058,N_27476);
nand U27660 (N_27660,N_27119,N_27385);
nor U27661 (N_27661,N_27473,N_27442);
nor U27662 (N_27662,N_27192,N_27545);
xnor U27663 (N_27663,N_27031,N_27375);
nand U27664 (N_27664,N_27521,N_27086);
or U27665 (N_27665,N_27127,N_27152);
and U27666 (N_27666,N_27235,N_27565);
nor U27667 (N_27667,N_27465,N_27590);
nand U27668 (N_27668,N_27423,N_27493);
or U27669 (N_27669,N_27233,N_27010);
xor U27670 (N_27670,N_27332,N_27300);
nand U27671 (N_27671,N_27358,N_27291);
xnor U27672 (N_27672,N_27541,N_27172);
and U27673 (N_27673,N_27478,N_27304);
xnor U27674 (N_27674,N_27365,N_27216);
and U27675 (N_27675,N_27191,N_27075);
nand U27676 (N_27676,N_27055,N_27238);
nand U27677 (N_27677,N_27532,N_27381);
nor U27678 (N_27678,N_27591,N_27469);
or U27679 (N_27679,N_27283,N_27355);
or U27680 (N_27680,N_27044,N_27482);
xnor U27681 (N_27681,N_27222,N_27593);
nor U27682 (N_27682,N_27342,N_27042);
xnor U27683 (N_27683,N_27019,N_27229);
xor U27684 (N_27684,N_27368,N_27525);
and U27685 (N_27685,N_27015,N_27535);
nor U27686 (N_27686,N_27101,N_27024);
and U27687 (N_27687,N_27515,N_27250);
nor U27688 (N_27688,N_27307,N_27428);
xnor U27689 (N_27689,N_27150,N_27582);
nand U27690 (N_27690,N_27254,N_27413);
xor U27691 (N_27691,N_27073,N_27274);
nor U27692 (N_27692,N_27519,N_27540);
xor U27693 (N_27693,N_27103,N_27116);
nor U27694 (N_27694,N_27111,N_27193);
nor U27695 (N_27695,N_27051,N_27181);
or U27696 (N_27696,N_27153,N_27264);
and U27697 (N_27697,N_27453,N_27468);
nor U27698 (N_27698,N_27067,N_27074);
or U27699 (N_27699,N_27278,N_27479);
nor U27700 (N_27700,N_27318,N_27234);
and U27701 (N_27701,N_27200,N_27334);
nand U27702 (N_27702,N_27563,N_27544);
and U27703 (N_27703,N_27490,N_27198);
xnor U27704 (N_27704,N_27405,N_27424);
nor U27705 (N_27705,N_27382,N_27460);
and U27706 (N_27706,N_27323,N_27420);
and U27707 (N_27707,N_27017,N_27501);
and U27708 (N_27708,N_27206,N_27547);
nand U27709 (N_27709,N_27580,N_27190);
and U27710 (N_27710,N_27106,N_27378);
xnor U27711 (N_27711,N_27056,N_27310);
or U27712 (N_27712,N_27225,N_27104);
or U27713 (N_27713,N_27062,N_27337);
xor U27714 (N_27714,N_27440,N_27076);
nand U27715 (N_27715,N_27367,N_27066);
nand U27716 (N_27716,N_27054,N_27039);
xnor U27717 (N_27717,N_27037,N_27072);
nor U27718 (N_27718,N_27454,N_27499);
nor U27719 (N_27719,N_27316,N_27114);
nand U27720 (N_27720,N_27538,N_27517);
or U27721 (N_27721,N_27495,N_27040);
nand U27722 (N_27722,N_27313,N_27557);
xor U27723 (N_27723,N_27113,N_27204);
and U27724 (N_27724,N_27554,N_27203);
xor U27725 (N_27725,N_27117,N_27537);
nor U27726 (N_27726,N_27128,N_27164);
nor U27727 (N_27727,N_27183,N_27297);
xnor U27728 (N_27728,N_27397,N_27498);
or U27729 (N_27729,N_27094,N_27349);
xnor U27730 (N_27730,N_27398,N_27448);
nor U27731 (N_27731,N_27534,N_27302);
and U27732 (N_27732,N_27268,N_27588);
nand U27733 (N_27733,N_27166,N_27147);
and U27734 (N_27734,N_27280,N_27059);
and U27735 (N_27735,N_27403,N_27474);
nand U27736 (N_27736,N_27578,N_27135);
xnor U27737 (N_27737,N_27432,N_27005);
nand U27738 (N_27738,N_27371,N_27347);
or U27739 (N_27739,N_27085,N_27387);
xnor U27740 (N_27740,N_27292,N_27211);
or U27741 (N_27741,N_27497,N_27208);
nand U27742 (N_27742,N_27345,N_27596);
and U27743 (N_27743,N_27402,N_27021);
or U27744 (N_27744,N_27057,N_27458);
nand U27745 (N_27745,N_27231,N_27599);
nand U27746 (N_27746,N_27100,N_27443);
xnor U27747 (N_27747,N_27531,N_27570);
or U27748 (N_27748,N_27285,N_27459);
xor U27749 (N_27749,N_27212,N_27144);
or U27750 (N_27750,N_27082,N_27194);
and U27751 (N_27751,N_27068,N_27435);
nand U27752 (N_27752,N_27579,N_27567);
xor U27753 (N_27753,N_27380,N_27145);
xnor U27754 (N_27754,N_27214,N_27396);
or U27755 (N_27755,N_27483,N_27237);
nand U27756 (N_27756,N_27157,N_27457);
or U27757 (N_27757,N_27394,N_27139);
nand U27758 (N_27758,N_27296,N_27512);
or U27759 (N_27759,N_27165,N_27533);
nand U27760 (N_27760,N_27376,N_27555);
or U27761 (N_27761,N_27412,N_27189);
or U27762 (N_27762,N_27575,N_27099);
xor U27763 (N_27763,N_27009,N_27427);
nand U27764 (N_27764,N_27361,N_27414);
or U27765 (N_27765,N_27287,N_27201);
nand U27766 (N_27766,N_27284,N_27187);
and U27767 (N_27767,N_27223,N_27012);
xnor U27768 (N_27768,N_27228,N_27589);
and U27769 (N_27769,N_27518,N_27050);
xor U27770 (N_27770,N_27528,N_27136);
and U27771 (N_27771,N_27444,N_27373);
xnor U27772 (N_27772,N_27426,N_27184);
or U27773 (N_27773,N_27326,N_27354);
xnor U27774 (N_27774,N_27529,N_27097);
or U27775 (N_27775,N_27035,N_27064);
xor U27776 (N_27776,N_27034,N_27573);
nand U27777 (N_27777,N_27176,N_27530);
nor U27778 (N_27778,N_27048,N_27196);
nor U27779 (N_27779,N_27260,N_27550);
xor U27780 (N_27780,N_27175,N_27102);
xor U27781 (N_27781,N_27180,N_27455);
or U27782 (N_27782,N_27077,N_27178);
xor U27783 (N_27783,N_27079,N_27452);
or U27784 (N_27784,N_27470,N_27242);
or U27785 (N_27785,N_27461,N_27388);
and U27786 (N_27786,N_27359,N_27063);
nor U27787 (N_27787,N_27256,N_27571);
or U27788 (N_27788,N_27383,N_27158);
and U27789 (N_27789,N_27131,N_27430);
and U27790 (N_27790,N_27279,N_27003);
or U27791 (N_27791,N_27504,N_27041);
nand U27792 (N_27792,N_27053,N_27195);
nand U27793 (N_27793,N_27025,N_27401);
nor U27794 (N_27794,N_27275,N_27491);
nor U27795 (N_27795,N_27586,N_27161);
and U27796 (N_27796,N_27449,N_27084);
or U27797 (N_27797,N_27309,N_27112);
nand U27798 (N_27798,N_27352,N_27489);
and U27799 (N_27799,N_27516,N_27374);
nand U27800 (N_27800,N_27298,N_27335);
and U27801 (N_27801,N_27049,N_27293);
xnor U27802 (N_27802,N_27438,N_27520);
xor U27803 (N_27803,N_27481,N_27391);
nand U27804 (N_27804,N_27289,N_27407);
nand U27805 (N_27805,N_27149,N_27269);
xnor U27806 (N_27806,N_27227,N_27513);
or U27807 (N_27807,N_27344,N_27502);
and U27808 (N_27808,N_27330,N_27536);
xor U27809 (N_27809,N_27462,N_27087);
nor U27810 (N_27810,N_27301,N_27553);
nand U27811 (N_27811,N_27419,N_27171);
xnor U27812 (N_27812,N_27393,N_27328);
nor U27813 (N_27813,N_27262,N_27510);
and U27814 (N_27814,N_27241,N_27263);
or U27815 (N_27815,N_27038,N_27526);
nor U27816 (N_27816,N_27160,N_27281);
nor U27817 (N_27817,N_27251,N_27362);
xor U27818 (N_27818,N_27141,N_27026);
nand U27819 (N_27819,N_27078,N_27466);
and U27820 (N_27820,N_27255,N_27311);
nor U27821 (N_27821,N_27065,N_27011);
and U27822 (N_27822,N_27346,N_27115);
xnor U27823 (N_27823,N_27007,N_27091);
or U27824 (N_27824,N_27182,N_27089);
and U27825 (N_27825,N_27142,N_27484);
nand U27826 (N_27826,N_27472,N_27093);
nand U27827 (N_27827,N_27508,N_27372);
and U27828 (N_27828,N_27282,N_27496);
nor U27829 (N_27829,N_27299,N_27511);
and U27830 (N_27830,N_27170,N_27239);
and U27831 (N_27831,N_27290,N_27226);
nor U27832 (N_27832,N_27560,N_27273);
nor U27833 (N_27833,N_27390,N_27523);
xor U27834 (N_27834,N_27524,N_27325);
and U27835 (N_27835,N_27266,N_27377);
and U27836 (N_27836,N_27259,N_27199);
xor U27837 (N_27837,N_27509,N_27108);
and U27838 (N_27838,N_27415,N_27018);
nand U27839 (N_27839,N_27329,N_27410);
nand U27840 (N_27840,N_27360,N_27001);
xor U27841 (N_27841,N_27441,N_27417);
or U27842 (N_27842,N_27027,N_27363);
nand U27843 (N_27843,N_27070,N_27122);
nand U27844 (N_27844,N_27243,N_27343);
nor U27845 (N_27845,N_27060,N_27559);
xor U27846 (N_27846,N_27487,N_27436);
nand U27847 (N_27847,N_27551,N_27561);
and U27848 (N_27848,N_27408,N_27202);
nand U27849 (N_27849,N_27215,N_27022);
nand U27850 (N_27850,N_27162,N_27036);
nor U27851 (N_27851,N_27351,N_27583);
xnor U27852 (N_27852,N_27315,N_27425);
or U27853 (N_27853,N_27069,N_27312);
and U27854 (N_27854,N_27514,N_27488);
xnor U27855 (N_27855,N_27123,N_27219);
nor U27856 (N_27856,N_27294,N_27379);
nand U27857 (N_27857,N_27463,N_27124);
xnor U27858 (N_27858,N_27217,N_27095);
and U27859 (N_27859,N_27000,N_27594);
or U27860 (N_27860,N_27340,N_27400);
or U27861 (N_27861,N_27186,N_27169);
or U27862 (N_27862,N_27558,N_27562);
or U27863 (N_27863,N_27185,N_27148);
nand U27864 (N_27864,N_27486,N_27467);
and U27865 (N_27865,N_27395,N_27576);
nand U27866 (N_27866,N_27107,N_27030);
or U27867 (N_27867,N_27322,N_27083);
nor U27868 (N_27868,N_27399,N_27539);
or U27869 (N_27869,N_27505,N_27247);
nor U27870 (N_27870,N_27389,N_27110);
or U27871 (N_27871,N_27450,N_27317);
and U27872 (N_27872,N_27336,N_27177);
nor U27873 (N_27873,N_27288,N_27384);
and U27874 (N_27874,N_27319,N_27434);
or U27875 (N_27875,N_27096,N_27129);
xnor U27876 (N_27876,N_27020,N_27552);
xor U27877 (N_27877,N_27126,N_27008);
and U27878 (N_27878,N_27134,N_27271);
and U27879 (N_27879,N_27156,N_27277);
nor U27880 (N_27880,N_27306,N_27081);
or U27881 (N_27881,N_27584,N_27138);
and U27882 (N_27882,N_27392,N_27140);
xnor U27883 (N_27883,N_27494,N_27197);
nand U27884 (N_27884,N_27133,N_27252);
or U27885 (N_27885,N_27324,N_27090);
or U27886 (N_27886,N_27033,N_27446);
and U27887 (N_27887,N_27437,N_27220);
nand U27888 (N_27888,N_27597,N_27421);
and U27889 (N_27889,N_27006,N_27151);
nand U27890 (N_27890,N_27052,N_27348);
nor U27891 (N_27891,N_27137,N_27431);
nor U27892 (N_27892,N_27471,N_27267);
or U27893 (N_27893,N_27333,N_27029);
nor U27894 (N_27894,N_27587,N_27543);
nand U27895 (N_27895,N_27447,N_27109);
or U27896 (N_27896,N_27416,N_27585);
nor U27897 (N_27897,N_27477,N_27188);
xor U27898 (N_27898,N_27261,N_27167);
or U27899 (N_27899,N_27253,N_27209);
and U27900 (N_27900,N_27330,N_27301);
or U27901 (N_27901,N_27242,N_27436);
or U27902 (N_27902,N_27277,N_27526);
and U27903 (N_27903,N_27522,N_27250);
xor U27904 (N_27904,N_27216,N_27214);
and U27905 (N_27905,N_27284,N_27326);
xor U27906 (N_27906,N_27005,N_27493);
and U27907 (N_27907,N_27311,N_27091);
xor U27908 (N_27908,N_27386,N_27167);
or U27909 (N_27909,N_27430,N_27107);
nand U27910 (N_27910,N_27067,N_27048);
or U27911 (N_27911,N_27288,N_27299);
xnor U27912 (N_27912,N_27477,N_27089);
and U27913 (N_27913,N_27154,N_27328);
nand U27914 (N_27914,N_27368,N_27110);
and U27915 (N_27915,N_27474,N_27021);
nor U27916 (N_27916,N_27519,N_27136);
nor U27917 (N_27917,N_27235,N_27361);
xnor U27918 (N_27918,N_27542,N_27253);
nand U27919 (N_27919,N_27361,N_27102);
xnor U27920 (N_27920,N_27425,N_27359);
and U27921 (N_27921,N_27239,N_27131);
xor U27922 (N_27922,N_27560,N_27137);
and U27923 (N_27923,N_27130,N_27151);
and U27924 (N_27924,N_27397,N_27298);
and U27925 (N_27925,N_27075,N_27133);
nor U27926 (N_27926,N_27215,N_27553);
nand U27927 (N_27927,N_27237,N_27104);
and U27928 (N_27928,N_27425,N_27290);
nor U27929 (N_27929,N_27047,N_27146);
and U27930 (N_27930,N_27541,N_27582);
nand U27931 (N_27931,N_27378,N_27359);
xnor U27932 (N_27932,N_27382,N_27102);
nor U27933 (N_27933,N_27084,N_27265);
nor U27934 (N_27934,N_27390,N_27245);
and U27935 (N_27935,N_27352,N_27321);
nor U27936 (N_27936,N_27168,N_27577);
or U27937 (N_27937,N_27387,N_27462);
nand U27938 (N_27938,N_27295,N_27472);
and U27939 (N_27939,N_27462,N_27012);
nor U27940 (N_27940,N_27387,N_27517);
and U27941 (N_27941,N_27306,N_27111);
xor U27942 (N_27942,N_27338,N_27332);
xnor U27943 (N_27943,N_27379,N_27478);
nor U27944 (N_27944,N_27389,N_27489);
and U27945 (N_27945,N_27096,N_27490);
and U27946 (N_27946,N_27279,N_27004);
xor U27947 (N_27947,N_27446,N_27171);
nand U27948 (N_27948,N_27378,N_27352);
or U27949 (N_27949,N_27304,N_27196);
or U27950 (N_27950,N_27175,N_27496);
nand U27951 (N_27951,N_27486,N_27402);
nor U27952 (N_27952,N_27176,N_27007);
nand U27953 (N_27953,N_27136,N_27035);
or U27954 (N_27954,N_27315,N_27013);
or U27955 (N_27955,N_27048,N_27202);
or U27956 (N_27956,N_27121,N_27166);
nor U27957 (N_27957,N_27337,N_27016);
xor U27958 (N_27958,N_27196,N_27077);
xnor U27959 (N_27959,N_27575,N_27398);
xnor U27960 (N_27960,N_27098,N_27009);
nand U27961 (N_27961,N_27561,N_27553);
nand U27962 (N_27962,N_27519,N_27239);
nand U27963 (N_27963,N_27423,N_27419);
nor U27964 (N_27964,N_27097,N_27202);
or U27965 (N_27965,N_27149,N_27275);
or U27966 (N_27966,N_27303,N_27165);
xor U27967 (N_27967,N_27382,N_27308);
or U27968 (N_27968,N_27349,N_27531);
xor U27969 (N_27969,N_27159,N_27105);
or U27970 (N_27970,N_27119,N_27097);
and U27971 (N_27971,N_27448,N_27561);
nor U27972 (N_27972,N_27333,N_27467);
nor U27973 (N_27973,N_27360,N_27500);
nand U27974 (N_27974,N_27217,N_27532);
and U27975 (N_27975,N_27070,N_27331);
nor U27976 (N_27976,N_27088,N_27131);
nor U27977 (N_27977,N_27312,N_27397);
and U27978 (N_27978,N_27370,N_27474);
nor U27979 (N_27979,N_27040,N_27383);
nor U27980 (N_27980,N_27300,N_27106);
xor U27981 (N_27981,N_27535,N_27541);
nor U27982 (N_27982,N_27240,N_27068);
nor U27983 (N_27983,N_27289,N_27324);
or U27984 (N_27984,N_27481,N_27440);
and U27985 (N_27985,N_27539,N_27203);
nand U27986 (N_27986,N_27573,N_27491);
or U27987 (N_27987,N_27215,N_27087);
xor U27988 (N_27988,N_27282,N_27211);
nor U27989 (N_27989,N_27081,N_27294);
nand U27990 (N_27990,N_27556,N_27401);
nor U27991 (N_27991,N_27251,N_27265);
nand U27992 (N_27992,N_27161,N_27309);
xor U27993 (N_27993,N_27585,N_27592);
xnor U27994 (N_27994,N_27323,N_27100);
nand U27995 (N_27995,N_27074,N_27263);
nand U27996 (N_27996,N_27006,N_27164);
or U27997 (N_27997,N_27292,N_27003);
nand U27998 (N_27998,N_27214,N_27384);
xor U27999 (N_27999,N_27054,N_27375);
nand U28000 (N_28000,N_27401,N_27284);
xor U28001 (N_28001,N_27566,N_27215);
xnor U28002 (N_28002,N_27352,N_27441);
xor U28003 (N_28003,N_27555,N_27254);
xnor U28004 (N_28004,N_27083,N_27434);
or U28005 (N_28005,N_27084,N_27194);
and U28006 (N_28006,N_27401,N_27422);
or U28007 (N_28007,N_27322,N_27484);
or U28008 (N_28008,N_27154,N_27359);
xor U28009 (N_28009,N_27472,N_27053);
xnor U28010 (N_28010,N_27221,N_27389);
nor U28011 (N_28011,N_27328,N_27077);
nor U28012 (N_28012,N_27297,N_27089);
nand U28013 (N_28013,N_27439,N_27006);
nand U28014 (N_28014,N_27449,N_27551);
nor U28015 (N_28015,N_27557,N_27581);
and U28016 (N_28016,N_27414,N_27205);
or U28017 (N_28017,N_27303,N_27110);
nor U28018 (N_28018,N_27031,N_27266);
or U28019 (N_28019,N_27452,N_27211);
xor U28020 (N_28020,N_27180,N_27050);
nand U28021 (N_28021,N_27050,N_27187);
and U28022 (N_28022,N_27143,N_27429);
nand U28023 (N_28023,N_27109,N_27286);
nand U28024 (N_28024,N_27220,N_27010);
or U28025 (N_28025,N_27035,N_27505);
nand U28026 (N_28026,N_27167,N_27226);
xor U28027 (N_28027,N_27417,N_27477);
nand U28028 (N_28028,N_27250,N_27355);
and U28029 (N_28029,N_27506,N_27061);
nor U28030 (N_28030,N_27053,N_27251);
or U28031 (N_28031,N_27173,N_27410);
and U28032 (N_28032,N_27057,N_27108);
or U28033 (N_28033,N_27434,N_27132);
xnor U28034 (N_28034,N_27094,N_27155);
xor U28035 (N_28035,N_27587,N_27391);
nor U28036 (N_28036,N_27243,N_27006);
and U28037 (N_28037,N_27278,N_27521);
nor U28038 (N_28038,N_27033,N_27305);
xnor U28039 (N_28039,N_27521,N_27206);
and U28040 (N_28040,N_27414,N_27463);
and U28041 (N_28041,N_27430,N_27492);
xnor U28042 (N_28042,N_27332,N_27489);
nand U28043 (N_28043,N_27435,N_27387);
nand U28044 (N_28044,N_27364,N_27170);
nand U28045 (N_28045,N_27380,N_27427);
nand U28046 (N_28046,N_27279,N_27083);
or U28047 (N_28047,N_27596,N_27344);
xnor U28048 (N_28048,N_27459,N_27032);
or U28049 (N_28049,N_27197,N_27595);
nor U28050 (N_28050,N_27075,N_27039);
or U28051 (N_28051,N_27520,N_27194);
and U28052 (N_28052,N_27200,N_27330);
xor U28053 (N_28053,N_27338,N_27288);
or U28054 (N_28054,N_27501,N_27285);
nand U28055 (N_28055,N_27306,N_27400);
nor U28056 (N_28056,N_27289,N_27066);
and U28057 (N_28057,N_27506,N_27073);
nor U28058 (N_28058,N_27059,N_27406);
xor U28059 (N_28059,N_27319,N_27332);
and U28060 (N_28060,N_27334,N_27182);
nand U28061 (N_28061,N_27307,N_27246);
or U28062 (N_28062,N_27366,N_27068);
xor U28063 (N_28063,N_27066,N_27292);
nor U28064 (N_28064,N_27572,N_27063);
xnor U28065 (N_28065,N_27050,N_27366);
nand U28066 (N_28066,N_27269,N_27234);
or U28067 (N_28067,N_27337,N_27597);
nor U28068 (N_28068,N_27269,N_27226);
or U28069 (N_28069,N_27297,N_27327);
nand U28070 (N_28070,N_27321,N_27582);
or U28071 (N_28071,N_27462,N_27453);
nand U28072 (N_28072,N_27455,N_27161);
and U28073 (N_28073,N_27219,N_27335);
nor U28074 (N_28074,N_27382,N_27152);
nor U28075 (N_28075,N_27310,N_27383);
nand U28076 (N_28076,N_27138,N_27151);
or U28077 (N_28077,N_27318,N_27511);
nand U28078 (N_28078,N_27489,N_27483);
nor U28079 (N_28079,N_27310,N_27389);
nor U28080 (N_28080,N_27354,N_27415);
nand U28081 (N_28081,N_27494,N_27373);
xnor U28082 (N_28082,N_27251,N_27559);
and U28083 (N_28083,N_27482,N_27070);
xnor U28084 (N_28084,N_27452,N_27297);
nand U28085 (N_28085,N_27445,N_27436);
xor U28086 (N_28086,N_27378,N_27291);
or U28087 (N_28087,N_27011,N_27241);
and U28088 (N_28088,N_27113,N_27366);
and U28089 (N_28089,N_27542,N_27545);
nor U28090 (N_28090,N_27062,N_27262);
and U28091 (N_28091,N_27564,N_27397);
or U28092 (N_28092,N_27027,N_27231);
nor U28093 (N_28093,N_27069,N_27032);
or U28094 (N_28094,N_27586,N_27324);
xnor U28095 (N_28095,N_27433,N_27322);
nand U28096 (N_28096,N_27423,N_27411);
nor U28097 (N_28097,N_27295,N_27085);
or U28098 (N_28098,N_27051,N_27305);
nand U28099 (N_28099,N_27044,N_27029);
or U28100 (N_28100,N_27352,N_27366);
and U28101 (N_28101,N_27384,N_27539);
xor U28102 (N_28102,N_27470,N_27096);
and U28103 (N_28103,N_27226,N_27362);
or U28104 (N_28104,N_27444,N_27462);
nand U28105 (N_28105,N_27265,N_27340);
or U28106 (N_28106,N_27166,N_27235);
nor U28107 (N_28107,N_27457,N_27019);
xnor U28108 (N_28108,N_27008,N_27409);
nand U28109 (N_28109,N_27059,N_27020);
nor U28110 (N_28110,N_27486,N_27555);
xor U28111 (N_28111,N_27557,N_27249);
xnor U28112 (N_28112,N_27064,N_27478);
xor U28113 (N_28113,N_27163,N_27092);
nor U28114 (N_28114,N_27332,N_27078);
and U28115 (N_28115,N_27489,N_27383);
nor U28116 (N_28116,N_27498,N_27451);
and U28117 (N_28117,N_27140,N_27581);
and U28118 (N_28118,N_27182,N_27062);
nor U28119 (N_28119,N_27340,N_27194);
or U28120 (N_28120,N_27244,N_27544);
nand U28121 (N_28121,N_27124,N_27178);
and U28122 (N_28122,N_27521,N_27165);
nor U28123 (N_28123,N_27368,N_27391);
nand U28124 (N_28124,N_27280,N_27029);
nand U28125 (N_28125,N_27301,N_27394);
nand U28126 (N_28126,N_27426,N_27016);
nor U28127 (N_28127,N_27453,N_27562);
and U28128 (N_28128,N_27390,N_27262);
and U28129 (N_28129,N_27146,N_27261);
and U28130 (N_28130,N_27554,N_27407);
and U28131 (N_28131,N_27534,N_27579);
and U28132 (N_28132,N_27024,N_27243);
nand U28133 (N_28133,N_27439,N_27453);
and U28134 (N_28134,N_27336,N_27003);
or U28135 (N_28135,N_27215,N_27491);
or U28136 (N_28136,N_27066,N_27240);
xor U28137 (N_28137,N_27573,N_27440);
or U28138 (N_28138,N_27525,N_27309);
xnor U28139 (N_28139,N_27229,N_27294);
nand U28140 (N_28140,N_27246,N_27516);
nand U28141 (N_28141,N_27001,N_27132);
nand U28142 (N_28142,N_27022,N_27371);
xnor U28143 (N_28143,N_27024,N_27047);
and U28144 (N_28144,N_27399,N_27472);
nor U28145 (N_28145,N_27465,N_27134);
xnor U28146 (N_28146,N_27496,N_27427);
or U28147 (N_28147,N_27244,N_27400);
and U28148 (N_28148,N_27057,N_27460);
nand U28149 (N_28149,N_27083,N_27259);
or U28150 (N_28150,N_27035,N_27121);
xnor U28151 (N_28151,N_27095,N_27365);
and U28152 (N_28152,N_27496,N_27420);
and U28153 (N_28153,N_27419,N_27008);
or U28154 (N_28154,N_27182,N_27257);
or U28155 (N_28155,N_27365,N_27570);
and U28156 (N_28156,N_27452,N_27002);
xor U28157 (N_28157,N_27392,N_27479);
xnor U28158 (N_28158,N_27454,N_27001);
or U28159 (N_28159,N_27266,N_27591);
nand U28160 (N_28160,N_27518,N_27147);
nand U28161 (N_28161,N_27197,N_27279);
or U28162 (N_28162,N_27533,N_27578);
nand U28163 (N_28163,N_27222,N_27523);
xor U28164 (N_28164,N_27187,N_27005);
nand U28165 (N_28165,N_27113,N_27005);
and U28166 (N_28166,N_27397,N_27238);
xnor U28167 (N_28167,N_27096,N_27340);
nor U28168 (N_28168,N_27415,N_27444);
and U28169 (N_28169,N_27057,N_27050);
xnor U28170 (N_28170,N_27086,N_27507);
and U28171 (N_28171,N_27237,N_27572);
nand U28172 (N_28172,N_27295,N_27491);
xor U28173 (N_28173,N_27160,N_27034);
xor U28174 (N_28174,N_27117,N_27466);
or U28175 (N_28175,N_27034,N_27495);
nand U28176 (N_28176,N_27148,N_27453);
or U28177 (N_28177,N_27184,N_27500);
nor U28178 (N_28178,N_27251,N_27106);
and U28179 (N_28179,N_27584,N_27489);
and U28180 (N_28180,N_27126,N_27374);
nor U28181 (N_28181,N_27369,N_27312);
nor U28182 (N_28182,N_27114,N_27325);
and U28183 (N_28183,N_27002,N_27503);
and U28184 (N_28184,N_27385,N_27317);
nor U28185 (N_28185,N_27221,N_27120);
or U28186 (N_28186,N_27036,N_27014);
nor U28187 (N_28187,N_27160,N_27586);
nand U28188 (N_28188,N_27029,N_27522);
nand U28189 (N_28189,N_27422,N_27272);
and U28190 (N_28190,N_27581,N_27560);
and U28191 (N_28191,N_27059,N_27506);
or U28192 (N_28192,N_27465,N_27434);
and U28193 (N_28193,N_27389,N_27448);
and U28194 (N_28194,N_27388,N_27152);
or U28195 (N_28195,N_27408,N_27467);
nand U28196 (N_28196,N_27425,N_27208);
or U28197 (N_28197,N_27563,N_27035);
nor U28198 (N_28198,N_27211,N_27062);
or U28199 (N_28199,N_27250,N_27203);
nor U28200 (N_28200,N_27679,N_27800);
nor U28201 (N_28201,N_27916,N_27904);
and U28202 (N_28202,N_28070,N_27753);
or U28203 (N_28203,N_27759,N_27912);
nor U28204 (N_28204,N_28192,N_27752);
xnor U28205 (N_28205,N_27937,N_28137);
or U28206 (N_28206,N_27844,N_27953);
nor U28207 (N_28207,N_28186,N_27863);
nor U28208 (N_28208,N_27721,N_28102);
or U28209 (N_28209,N_27809,N_27660);
xor U28210 (N_28210,N_28030,N_27890);
or U28211 (N_28211,N_27667,N_27996);
xnor U28212 (N_28212,N_27949,N_27730);
and U28213 (N_28213,N_27606,N_27669);
nor U28214 (N_28214,N_28129,N_27799);
nand U28215 (N_28215,N_28150,N_28028);
nor U28216 (N_28216,N_27817,N_27784);
and U28217 (N_28217,N_28121,N_27713);
or U28218 (N_28218,N_28040,N_27968);
nand U28219 (N_28219,N_28105,N_27615);
xnor U28220 (N_28220,N_28057,N_27936);
nand U28221 (N_28221,N_27607,N_27914);
nor U28222 (N_28222,N_27899,N_27655);
nor U28223 (N_28223,N_27847,N_27820);
nand U28224 (N_28224,N_27872,N_28094);
nor U28225 (N_28225,N_28145,N_28130);
xnor U28226 (N_28226,N_27742,N_28103);
nand U28227 (N_28227,N_27991,N_28037);
nand U28228 (N_28228,N_27868,N_27958);
and U28229 (N_28229,N_27616,N_27771);
xnor U28230 (N_28230,N_28166,N_27774);
nand U28231 (N_28231,N_28020,N_27952);
nor U28232 (N_28232,N_28060,N_28193);
and U28233 (N_28233,N_28104,N_27964);
and U28234 (N_28234,N_28163,N_28144);
nand U28235 (N_28235,N_27941,N_28189);
nand U28236 (N_28236,N_28119,N_28046);
or U28237 (N_28237,N_27959,N_27779);
and U28238 (N_28238,N_27884,N_27642);
nor U28239 (N_28239,N_28076,N_27950);
and U28240 (N_28240,N_27707,N_27861);
nand U28241 (N_28241,N_27609,N_27775);
nor U28242 (N_28242,N_27989,N_28125);
or U28243 (N_28243,N_28009,N_28045);
or U28244 (N_28244,N_27954,N_28048);
nor U28245 (N_28245,N_27836,N_27645);
nor U28246 (N_28246,N_27757,N_27696);
nand U28247 (N_28247,N_27641,N_28098);
and U28248 (N_28248,N_28069,N_27824);
or U28249 (N_28249,N_27691,N_27782);
nand U28250 (N_28250,N_27961,N_27746);
nand U28251 (N_28251,N_27903,N_27876);
and U28252 (N_28252,N_28126,N_27613);
or U28253 (N_28253,N_28086,N_27789);
or U28254 (N_28254,N_28199,N_28197);
nand U28255 (N_28255,N_27705,N_27732);
xor U28256 (N_28256,N_28047,N_27990);
or U28257 (N_28257,N_27726,N_27710);
xnor U28258 (N_28258,N_27638,N_27818);
or U28259 (N_28259,N_27913,N_27687);
nor U28260 (N_28260,N_27815,N_27915);
xor U28261 (N_28261,N_27689,N_27973);
or U28262 (N_28262,N_28007,N_28136);
or U28263 (N_28263,N_28117,N_27835);
nand U28264 (N_28264,N_28053,N_28061);
nand U28265 (N_28265,N_28169,N_27640);
or U28266 (N_28266,N_28156,N_28001);
nand U28267 (N_28267,N_27804,N_27881);
xnor U28268 (N_28268,N_27825,N_28074);
and U28269 (N_28269,N_27887,N_27860);
xnor U28270 (N_28270,N_27834,N_27602);
or U28271 (N_28271,N_28008,N_27933);
nand U28272 (N_28272,N_27902,N_27802);
and U28273 (N_28273,N_27711,N_28078);
xor U28274 (N_28274,N_27853,N_27988);
xnor U28275 (N_28275,N_27859,N_27893);
and U28276 (N_28276,N_27764,N_27692);
and U28277 (N_28277,N_27895,N_28172);
or U28278 (N_28278,N_27808,N_28187);
and U28279 (N_28279,N_27866,N_27729);
nor U28280 (N_28280,N_27967,N_28112);
nand U28281 (N_28281,N_28088,N_28158);
and U28282 (N_28282,N_27788,N_27674);
nand U28283 (N_28283,N_27886,N_27891);
or U28284 (N_28284,N_27747,N_27908);
xnor U28285 (N_28285,N_28021,N_27944);
and U28286 (N_28286,N_28149,N_28182);
or U28287 (N_28287,N_27928,N_27971);
and U28288 (N_28288,N_27617,N_28143);
nand U28289 (N_28289,N_27931,N_27661);
xor U28290 (N_28290,N_27748,N_28023);
nor U28291 (N_28291,N_27624,N_27813);
or U28292 (N_28292,N_27977,N_28153);
or U28293 (N_28293,N_27731,N_27702);
nor U28294 (N_28294,N_27735,N_27997);
nand U28295 (N_28295,N_28183,N_28075);
and U28296 (N_28296,N_27805,N_27681);
nand U28297 (N_28297,N_28000,N_27811);
or U28298 (N_28298,N_27797,N_28190);
xor U28299 (N_28299,N_28185,N_28024);
and U28300 (N_28300,N_27871,N_28132);
xnor U28301 (N_28301,N_27637,N_28004);
nor U28302 (N_28302,N_27634,N_28106);
xor U28303 (N_28303,N_27827,N_27942);
xor U28304 (N_28304,N_27984,N_27776);
or U28305 (N_28305,N_27858,N_27882);
xnor U28306 (N_28306,N_27810,N_28177);
and U28307 (N_28307,N_28174,N_27668);
xnor U28308 (N_28308,N_27749,N_27956);
nor U28309 (N_28309,N_28133,N_28015);
xnor U28310 (N_28310,N_28109,N_28176);
xor U28311 (N_28311,N_27750,N_27676);
and U28312 (N_28312,N_28180,N_27673);
or U28313 (N_28313,N_28139,N_27926);
xor U28314 (N_28314,N_27756,N_27986);
and U28315 (N_28315,N_27940,N_27694);
nor U28316 (N_28316,N_28017,N_27932);
nor U28317 (N_28317,N_27662,N_27626);
and U28318 (N_28318,N_27970,N_27966);
nor U28319 (N_28319,N_27650,N_27639);
or U28320 (N_28320,N_27683,N_27651);
and U28321 (N_28321,N_27727,N_27722);
and U28322 (N_28322,N_27690,N_27869);
and U28323 (N_28323,N_27695,N_27923);
nand U28324 (N_28324,N_28033,N_27981);
nand U28325 (N_28325,N_27894,N_27843);
or U28326 (N_28326,N_27832,N_27955);
nor U28327 (N_28327,N_27604,N_28099);
nor U28328 (N_28328,N_27803,N_28170);
nor U28329 (N_28329,N_27874,N_27880);
xnor U28330 (N_28330,N_28111,N_28128);
or U28331 (N_28331,N_28101,N_27801);
nor U28332 (N_28332,N_27737,N_27885);
nand U28333 (N_28333,N_27744,N_27920);
or U28334 (N_28334,N_27649,N_27703);
xor U28335 (N_28335,N_27814,N_27889);
or U28336 (N_28336,N_28115,N_27905);
nand U28337 (N_28337,N_27733,N_27699);
xor U28338 (N_28338,N_27630,N_27939);
or U28339 (N_28339,N_28113,N_27957);
nand U28340 (N_28340,N_27706,N_27664);
nor U28341 (N_28341,N_28097,N_27963);
xor U28342 (N_28342,N_27773,N_27704);
nand U28343 (N_28343,N_27930,N_27678);
nor U28344 (N_28344,N_28054,N_28173);
or U28345 (N_28345,N_27601,N_28087);
xnor U28346 (N_28346,N_28071,N_27877);
xnor U28347 (N_28347,N_27765,N_27998);
nand U28348 (N_28348,N_28077,N_28140);
xnor U28349 (N_28349,N_27845,N_27736);
or U28350 (N_28350,N_27646,N_28151);
nand U28351 (N_28351,N_27921,N_27793);
nand U28352 (N_28352,N_28014,N_28161);
and U28353 (N_28353,N_28036,N_27812);
nor U28354 (N_28354,N_27697,N_27723);
or U28355 (N_28355,N_28191,N_28067);
xor U28356 (N_28356,N_27900,N_27778);
or U28357 (N_28357,N_28083,N_27943);
nand U28358 (N_28358,N_27842,N_27741);
nand U28359 (N_28359,N_27856,N_27982);
nand U28360 (N_28360,N_27851,N_27978);
nand U28361 (N_28361,N_28059,N_28168);
and U28362 (N_28362,N_27918,N_27648);
xor U28363 (N_28363,N_27924,N_27854);
nor U28364 (N_28364,N_27850,N_27717);
xnor U28365 (N_28365,N_27897,N_27794);
nor U28366 (N_28366,N_27701,N_27635);
or U28367 (N_28367,N_27795,N_27770);
xor U28368 (N_28368,N_27724,N_28082);
or U28369 (N_28369,N_27969,N_27734);
nor U28370 (N_28370,N_27980,N_27829);
xor U28371 (N_28371,N_27992,N_28039);
and U28372 (N_28372,N_27680,N_28035);
nand U28373 (N_28373,N_27629,N_28164);
nor U28374 (N_28374,N_27623,N_27838);
xnor U28375 (N_28375,N_27875,N_28012);
and U28376 (N_28376,N_27987,N_27917);
nand U28377 (N_28377,N_27700,N_28114);
nor U28378 (N_28378,N_28044,N_27947);
and U28379 (N_28379,N_27614,N_28019);
and U28380 (N_28380,N_27766,N_27828);
xor U28381 (N_28381,N_28162,N_28108);
and U28382 (N_28382,N_27663,N_27960);
or U28383 (N_28383,N_28134,N_28127);
xor U28384 (N_28384,N_28049,N_28065);
xnor U28385 (N_28385,N_28051,N_28124);
nor U28386 (N_28386,N_27677,N_27754);
nand U28387 (N_28387,N_28079,N_27688);
xor U28388 (N_28388,N_27929,N_28095);
nor U28389 (N_28389,N_27995,N_27792);
or U28390 (N_28390,N_27656,N_27619);
and U28391 (N_28391,N_27781,N_27823);
nor U28392 (N_28392,N_27934,N_28135);
or U28393 (N_28393,N_27807,N_28026);
or U28394 (N_28394,N_27919,N_27994);
and U28395 (N_28395,N_27666,N_27708);
or U28396 (N_28396,N_27867,N_27892);
and U28397 (N_28397,N_28123,N_27848);
and U28398 (N_28398,N_27870,N_27879);
or U28399 (N_28399,N_27948,N_27974);
and U28400 (N_28400,N_28159,N_28052);
nor U28401 (N_28401,N_27654,N_27927);
or U28402 (N_28402,N_28118,N_28038);
nor U28403 (N_28403,N_28043,N_27719);
xor U28404 (N_28404,N_28062,N_28160);
xnor U28405 (N_28405,N_27993,N_28181);
nor U28406 (N_28406,N_28034,N_27612);
and U28407 (N_28407,N_28155,N_27883);
xnor U28408 (N_28408,N_27740,N_27611);
nand U28409 (N_28409,N_28116,N_28188);
xnor U28410 (N_28410,N_27846,N_28096);
or U28411 (N_28411,N_27849,N_28018);
xor U28412 (N_28412,N_27653,N_28050);
and U28413 (N_28413,N_28157,N_27657);
and U28414 (N_28414,N_27772,N_27620);
and U28415 (N_28415,N_28002,N_27841);
and U28416 (N_28416,N_27743,N_27643);
nand U28417 (N_28417,N_28147,N_27714);
and U28418 (N_28418,N_27983,N_27762);
nand U28419 (N_28419,N_28016,N_27855);
and U28420 (N_28420,N_28178,N_27672);
and U28421 (N_28421,N_28175,N_27786);
or U28422 (N_28422,N_28165,N_28184);
and U28423 (N_28423,N_28022,N_27685);
or U28424 (N_28424,N_27783,N_27852);
nand U28425 (N_28425,N_27684,N_27985);
nand U28426 (N_28426,N_28089,N_28032);
and U28427 (N_28427,N_27659,N_28056);
or U28428 (N_28428,N_28092,N_27922);
nor U28429 (N_28429,N_27715,N_27682);
and U28430 (N_28430,N_28010,N_28003);
nor U28431 (N_28431,N_27608,N_28058);
and U28432 (N_28432,N_27901,N_27888);
or U28433 (N_28433,N_28063,N_27864);
or U28434 (N_28434,N_27755,N_28091);
nor U28435 (N_28435,N_27898,N_27739);
xnor U28436 (N_28436,N_27600,N_27972);
and U28437 (N_28437,N_27796,N_27911);
nor U28438 (N_28438,N_27720,N_28085);
nor U28439 (N_28439,N_27605,N_28171);
nor U28440 (N_28440,N_28005,N_27925);
nor U28441 (N_28441,N_28041,N_27761);
nand U28442 (N_28442,N_27821,N_28068);
or U28443 (N_28443,N_28011,N_27806);
or U28444 (N_28444,N_27857,N_27831);
nand U28445 (N_28445,N_27822,N_28081);
xor U28446 (N_28446,N_28110,N_27633);
xnor U28447 (N_28447,N_28122,N_27618);
or U28448 (N_28448,N_27709,N_28029);
nand U28449 (N_28449,N_27878,N_27693);
nor U28450 (N_28450,N_27862,N_28179);
xnor U28451 (N_28451,N_27790,N_28093);
and U28452 (N_28452,N_27946,N_28138);
and U28453 (N_28453,N_28055,N_27671);
or U28454 (N_28454,N_27760,N_27839);
nor U28455 (N_28455,N_28080,N_27816);
nor U28456 (N_28456,N_27837,N_28031);
xnor U28457 (N_28457,N_28141,N_27769);
xnor U28458 (N_28458,N_27798,N_28064);
nand U28459 (N_28459,N_27725,N_27819);
nor U28460 (N_28460,N_27979,N_27826);
xnor U28461 (N_28461,N_28142,N_27658);
nor U28462 (N_28462,N_27698,N_27647);
nor U28463 (N_28463,N_27945,N_28198);
or U28464 (N_28464,N_27665,N_27787);
nand U28465 (N_28465,N_27716,N_27909);
or U28466 (N_28466,N_27627,N_27830);
and U28467 (N_28467,N_27728,N_28148);
nor U28468 (N_28468,N_28152,N_27628);
xor U28469 (N_28469,N_27670,N_28196);
and U28470 (N_28470,N_27951,N_27751);
nor U28471 (N_28471,N_27718,N_27652);
or U28472 (N_28472,N_27632,N_28167);
nor U28473 (N_28473,N_27910,N_27610);
nand U28474 (N_28474,N_27865,N_28195);
nor U28475 (N_28475,N_27785,N_27935);
nand U28476 (N_28476,N_27768,N_28027);
nand U28477 (N_28477,N_27621,N_27631);
and U28478 (N_28478,N_27777,N_28107);
nand U28479 (N_28479,N_28090,N_27636);
or U28480 (N_28480,N_27962,N_28042);
or U28481 (N_28481,N_27833,N_27675);
xnor U28482 (N_28482,N_27603,N_27791);
nand U28483 (N_28483,N_27745,N_27738);
or U28484 (N_28484,N_28072,N_27873);
and U28485 (N_28485,N_27644,N_28146);
xnor U28486 (N_28486,N_28073,N_27840);
and U28487 (N_28487,N_28006,N_28013);
and U28488 (N_28488,N_27758,N_28025);
and U28489 (N_28489,N_27896,N_28084);
or U28490 (N_28490,N_28120,N_27906);
or U28491 (N_28491,N_27975,N_27938);
nor U28492 (N_28492,N_27686,N_27625);
or U28493 (N_28493,N_28154,N_27622);
nor U28494 (N_28494,N_27763,N_27907);
or U28495 (N_28495,N_28100,N_27780);
nor U28496 (N_28496,N_27965,N_27999);
nand U28497 (N_28497,N_28066,N_28131);
nand U28498 (N_28498,N_27976,N_27767);
nor U28499 (N_28499,N_28194,N_27712);
nand U28500 (N_28500,N_27930,N_27884);
and U28501 (N_28501,N_27772,N_27926);
and U28502 (N_28502,N_27632,N_27821);
nor U28503 (N_28503,N_28078,N_28143);
and U28504 (N_28504,N_28093,N_27607);
or U28505 (N_28505,N_27803,N_27715);
nor U28506 (N_28506,N_27778,N_27636);
nor U28507 (N_28507,N_27935,N_27879);
xor U28508 (N_28508,N_27728,N_28048);
xnor U28509 (N_28509,N_28139,N_27736);
or U28510 (N_28510,N_27998,N_28068);
and U28511 (N_28511,N_27715,N_27784);
xnor U28512 (N_28512,N_27670,N_27960);
and U28513 (N_28513,N_27685,N_27755);
nand U28514 (N_28514,N_27724,N_28168);
nand U28515 (N_28515,N_28129,N_27737);
and U28516 (N_28516,N_27753,N_28055);
nor U28517 (N_28517,N_28088,N_27838);
or U28518 (N_28518,N_28027,N_27686);
nor U28519 (N_28519,N_27986,N_28172);
xnor U28520 (N_28520,N_27657,N_28176);
and U28521 (N_28521,N_27900,N_27961);
and U28522 (N_28522,N_27628,N_27823);
xnor U28523 (N_28523,N_28112,N_28016);
xnor U28524 (N_28524,N_27648,N_27707);
or U28525 (N_28525,N_28114,N_27674);
and U28526 (N_28526,N_28121,N_27973);
xor U28527 (N_28527,N_27744,N_28169);
xor U28528 (N_28528,N_28026,N_27761);
nand U28529 (N_28529,N_27657,N_27872);
or U28530 (N_28530,N_28162,N_27906);
nor U28531 (N_28531,N_27915,N_28165);
xnor U28532 (N_28532,N_28046,N_27756);
nand U28533 (N_28533,N_27868,N_28140);
nor U28534 (N_28534,N_27683,N_27848);
or U28535 (N_28535,N_27861,N_27748);
and U28536 (N_28536,N_27682,N_27849);
nand U28537 (N_28537,N_27784,N_27761);
nand U28538 (N_28538,N_27885,N_28087);
and U28539 (N_28539,N_28048,N_27920);
xnor U28540 (N_28540,N_27911,N_28024);
xor U28541 (N_28541,N_27928,N_27606);
xnor U28542 (N_28542,N_27650,N_27833);
xor U28543 (N_28543,N_28183,N_27603);
xor U28544 (N_28544,N_27870,N_27820);
xnor U28545 (N_28545,N_27959,N_28066);
and U28546 (N_28546,N_28130,N_27692);
and U28547 (N_28547,N_28010,N_27940);
nor U28548 (N_28548,N_28018,N_27789);
or U28549 (N_28549,N_27649,N_27617);
xnor U28550 (N_28550,N_27897,N_27836);
or U28551 (N_28551,N_28129,N_27782);
nand U28552 (N_28552,N_28120,N_27930);
and U28553 (N_28553,N_27639,N_27757);
or U28554 (N_28554,N_27714,N_28008);
or U28555 (N_28555,N_28027,N_28082);
or U28556 (N_28556,N_28190,N_27622);
or U28557 (N_28557,N_27634,N_27977);
nor U28558 (N_28558,N_27771,N_27682);
nand U28559 (N_28559,N_27737,N_27887);
or U28560 (N_28560,N_28013,N_27711);
nor U28561 (N_28561,N_27765,N_28016);
or U28562 (N_28562,N_27728,N_28088);
nand U28563 (N_28563,N_27944,N_27940);
xnor U28564 (N_28564,N_27654,N_28180);
nor U28565 (N_28565,N_27617,N_28044);
or U28566 (N_28566,N_28160,N_27618);
and U28567 (N_28567,N_27838,N_27629);
or U28568 (N_28568,N_27914,N_28012);
or U28569 (N_28569,N_28112,N_27754);
xnor U28570 (N_28570,N_27691,N_27784);
and U28571 (N_28571,N_27711,N_27938);
xor U28572 (N_28572,N_28139,N_28158);
xor U28573 (N_28573,N_27669,N_27737);
or U28574 (N_28574,N_28074,N_28070);
nor U28575 (N_28575,N_27833,N_28145);
xnor U28576 (N_28576,N_27934,N_27803);
nor U28577 (N_28577,N_27733,N_27973);
nor U28578 (N_28578,N_28034,N_28059);
nand U28579 (N_28579,N_27951,N_28006);
xnor U28580 (N_28580,N_27862,N_28063);
nor U28581 (N_28581,N_28037,N_28036);
nor U28582 (N_28582,N_28026,N_27869);
and U28583 (N_28583,N_28163,N_27702);
nor U28584 (N_28584,N_27838,N_28050);
and U28585 (N_28585,N_27830,N_28096);
xor U28586 (N_28586,N_28101,N_27854);
or U28587 (N_28587,N_27743,N_27722);
xnor U28588 (N_28588,N_28136,N_27623);
or U28589 (N_28589,N_27622,N_27646);
or U28590 (N_28590,N_27871,N_27652);
and U28591 (N_28591,N_28046,N_27618);
or U28592 (N_28592,N_27970,N_28162);
nor U28593 (N_28593,N_27912,N_28134);
or U28594 (N_28594,N_27995,N_27945);
xnor U28595 (N_28595,N_27900,N_28077);
nor U28596 (N_28596,N_28160,N_27787);
nand U28597 (N_28597,N_28151,N_27749);
nor U28598 (N_28598,N_28156,N_27992);
nand U28599 (N_28599,N_28174,N_28006);
nand U28600 (N_28600,N_28148,N_27829);
xor U28601 (N_28601,N_28175,N_27921);
xnor U28602 (N_28602,N_27865,N_27908);
nand U28603 (N_28603,N_27765,N_28096);
and U28604 (N_28604,N_27883,N_27798);
nor U28605 (N_28605,N_27903,N_27931);
xor U28606 (N_28606,N_27960,N_27659);
and U28607 (N_28607,N_28108,N_28098);
xor U28608 (N_28608,N_27644,N_27646);
nor U28609 (N_28609,N_27621,N_27817);
or U28610 (N_28610,N_28177,N_28037);
nand U28611 (N_28611,N_28140,N_28164);
or U28612 (N_28612,N_28099,N_27631);
nand U28613 (N_28613,N_28191,N_27995);
nand U28614 (N_28614,N_27924,N_28037);
xnor U28615 (N_28615,N_28176,N_27902);
or U28616 (N_28616,N_27873,N_28166);
and U28617 (N_28617,N_27772,N_28102);
nor U28618 (N_28618,N_27926,N_27976);
nand U28619 (N_28619,N_27725,N_27864);
nor U28620 (N_28620,N_27901,N_27777);
nor U28621 (N_28621,N_28082,N_27966);
nor U28622 (N_28622,N_28039,N_27971);
nand U28623 (N_28623,N_28099,N_27871);
nor U28624 (N_28624,N_28113,N_27894);
nand U28625 (N_28625,N_28086,N_27854);
xnor U28626 (N_28626,N_27843,N_28078);
xnor U28627 (N_28627,N_27738,N_27789);
and U28628 (N_28628,N_28042,N_27995);
nand U28629 (N_28629,N_28138,N_28022);
nor U28630 (N_28630,N_28021,N_27764);
or U28631 (N_28631,N_28036,N_27811);
or U28632 (N_28632,N_27946,N_27660);
xor U28633 (N_28633,N_28130,N_27608);
nor U28634 (N_28634,N_28112,N_28160);
nor U28635 (N_28635,N_28154,N_27650);
and U28636 (N_28636,N_28046,N_28017);
xnor U28637 (N_28637,N_27919,N_27740);
nand U28638 (N_28638,N_27939,N_28030);
and U28639 (N_28639,N_27636,N_28101);
nor U28640 (N_28640,N_27955,N_28042);
nor U28641 (N_28641,N_27706,N_27654);
xor U28642 (N_28642,N_27898,N_28043);
and U28643 (N_28643,N_28058,N_27807);
nand U28644 (N_28644,N_28053,N_27852);
xnor U28645 (N_28645,N_28038,N_27965);
nand U28646 (N_28646,N_27816,N_27749);
nand U28647 (N_28647,N_27713,N_27943);
xor U28648 (N_28648,N_27943,N_27938);
or U28649 (N_28649,N_27808,N_27803);
nor U28650 (N_28650,N_28193,N_28108);
or U28651 (N_28651,N_27986,N_27650);
or U28652 (N_28652,N_27743,N_27676);
nand U28653 (N_28653,N_28164,N_27915);
and U28654 (N_28654,N_28142,N_27708);
nor U28655 (N_28655,N_27674,N_27770);
nand U28656 (N_28656,N_27786,N_27633);
nand U28657 (N_28657,N_28067,N_27824);
and U28658 (N_28658,N_27881,N_27819);
xnor U28659 (N_28659,N_27959,N_27682);
nand U28660 (N_28660,N_27775,N_27604);
nor U28661 (N_28661,N_28152,N_27713);
and U28662 (N_28662,N_27835,N_27845);
xnor U28663 (N_28663,N_27792,N_28083);
or U28664 (N_28664,N_27683,N_28109);
nor U28665 (N_28665,N_27798,N_28168);
nand U28666 (N_28666,N_27772,N_27865);
or U28667 (N_28667,N_27844,N_27739);
or U28668 (N_28668,N_27942,N_27653);
nor U28669 (N_28669,N_27616,N_27912);
or U28670 (N_28670,N_27848,N_27807);
xnor U28671 (N_28671,N_27974,N_27872);
nor U28672 (N_28672,N_28158,N_27976);
and U28673 (N_28673,N_27651,N_28093);
and U28674 (N_28674,N_27664,N_27704);
nor U28675 (N_28675,N_28180,N_27629);
xor U28676 (N_28676,N_27729,N_27742);
xnor U28677 (N_28677,N_27847,N_27609);
xor U28678 (N_28678,N_27639,N_27600);
or U28679 (N_28679,N_28015,N_28176);
xnor U28680 (N_28680,N_28005,N_28130);
xnor U28681 (N_28681,N_27803,N_28072);
nor U28682 (N_28682,N_27724,N_27747);
nor U28683 (N_28683,N_28024,N_28105);
xnor U28684 (N_28684,N_28072,N_28121);
and U28685 (N_28685,N_27947,N_27924);
xor U28686 (N_28686,N_28106,N_27708);
and U28687 (N_28687,N_27853,N_27983);
xor U28688 (N_28688,N_28170,N_27630);
nor U28689 (N_28689,N_28198,N_27743);
xnor U28690 (N_28690,N_27780,N_27615);
nand U28691 (N_28691,N_28067,N_28072);
nor U28692 (N_28692,N_27846,N_27653);
or U28693 (N_28693,N_28139,N_27808);
and U28694 (N_28694,N_27960,N_27884);
xor U28695 (N_28695,N_27696,N_27862);
nor U28696 (N_28696,N_28147,N_28125);
xnor U28697 (N_28697,N_28185,N_27879);
xnor U28698 (N_28698,N_27914,N_28060);
or U28699 (N_28699,N_27981,N_27820);
xor U28700 (N_28700,N_27999,N_28143);
and U28701 (N_28701,N_27845,N_27763);
or U28702 (N_28702,N_28118,N_27976);
xnor U28703 (N_28703,N_28093,N_28160);
and U28704 (N_28704,N_27721,N_27603);
or U28705 (N_28705,N_27854,N_27871);
and U28706 (N_28706,N_27821,N_28143);
nor U28707 (N_28707,N_28001,N_27885);
nand U28708 (N_28708,N_27631,N_27616);
or U28709 (N_28709,N_27833,N_28025);
nand U28710 (N_28710,N_28082,N_27642);
and U28711 (N_28711,N_28027,N_27943);
nand U28712 (N_28712,N_27657,N_27859);
nor U28713 (N_28713,N_27640,N_27848);
and U28714 (N_28714,N_27955,N_27890);
xnor U28715 (N_28715,N_27739,N_27967);
xnor U28716 (N_28716,N_28022,N_27728);
nor U28717 (N_28717,N_27656,N_27943);
or U28718 (N_28718,N_27657,N_27841);
and U28719 (N_28719,N_27702,N_27788);
nand U28720 (N_28720,N_27670,N_27836);
nand U28721 (N_28721,N_27698,N_27877);
and U28722 (N_28722,N_27765,N_27798);
nor U28723 (N_28723,N_28016,N_27821);
xnor U28724 (N_28724,N_27740,N_27660);
xor U28725 (N_28725,N_27779,N_27967);
nand U28726 (N_28726,N_27874,N_27891);
nor U28727 (N_28727,N_28085,N_27667);
or U28728 (N_28728,N_27948,N_27740);
nor U28729 (N_28729,N_27742,N_27941);
nand U28730 (N_28730,N_27805,N_27917);
nor U28731 (N_28731,N_27996,N_27812);
or U28732 (N_28732,N_27863,N_28074);
nor U28733 (N_28733,N_27831,N_27674);
xor U28734 (N_28734,N_27879,N_28017);
and U28735 (N_28735,N_27823,N_27858);
or U28736 (N_28736,N_28063,N_27690);
or U28737 (N_28737,N_27997,N_28019);
nor U28738 (N_28738,N_27982,N_27906);
nand U28739 (N_28739,N_27735,N_27762);
xnor U28740 (N_28740,N_27709,N_27886);
nand U28741 (N_28741,N_27687,N_28034);
and U28742 (N_28742,N_27803,N_27840);
or U28743 (N_28743,N_28190,N_28084);
and U28744 (N_28744,N_27770,N_28041);
and U28745 (N_28745,N_28192,N_27823);
nand U28746 (N_28746,N_28125,N_28154);
nor U28747 (N_28747,N_28056,N_27712);
and U28748 (N_28748,N_27982,N_27650);
or U28749 (N_28749,N_27691,N_28133);
nor U28750 (N_28750,N_28175,N_27875);
and U28751 (N_28751,N_27819,N_28054);
and U28752 (N_28752,N_27899,N_27644);
or U28753 (N_28753,N_27729,N_27677);
and U28754 (N_28754,N_27876,N_28010);
nor U28755 (N_28755,N_28010,N_27760);
xnor U28756 (N_28756,N_28153,N_27714);
nand U28757 (N_28757,N_27825,N_27717);
and U28758 (N_28758,N_27727,N_27992);
nor U28759 (N_28759,N_27647,N_27776);
or U28760 (N_28760,N_28160,N_27881);
and U28761 (N_28761,N_27964,N_27847);
xor U28762 (N_28762,N_27940,N_27791);
nand U28763 (N_28763,N_27767,N_27601);
nand U28764 (N_28764,N_27798,N_27952);
nor U28765 (N_28765,N_28104,N_28168);
and U28766 (N_28766,N_28175,N_27989);
and U28767 (N_28767,N_27900,N_28047);
and U28768 (N_28768,N_27743,N_27789);
or U28769 (N_28769,N_27648,N_27840);
nand U28770 (N_28770,N_27877,N_28153);
nand U28771 (N_28771,N_27891,N_27753);
nand U28772 (N_28772,N_28199,N_27613);
nand U28773 (N_28773,N_27986,N_27828);
xor U28774 (N_28774,N_28012,N_27988);
nand U28775 (N_28775,N_27771,N_28174);
and U28776 (N_28776,N_27850,N_27682);
xor U28777 (N_28777,N_27611,N_27836);
or U28778 (N_28778,N_28156,N_27636);
xnor U28779 (N_28779,N_27696,N_28061);
xor U28780 (N_28780,N_28166,N_27686);
nor U28781 (N_28781,N_28171,N_27662);
nand U28782 (N_28782,N_27633,N_27821);
and U28783 (N_28783,N_27617,N_27819);
nand U28784 (N_28784,N_27913,N_28142);
or U28785 (N_28785,N_27668,N_27935);
xor U28786 (N_28786,N_27776,N_28186);
and U28787 (N_28787,N_28183,N_27902);
nand U28788 (N_28788,N_28063,N_27961);
xor U28789 (N_28789,N_27889,N_28062);
nor U28790 (N_28790,N_28056,N_27679);
nor U28791 (N_28791,N_28146,N_28108);
or U28792 (N_28792,N_27719,N_27722);
nor U28793 (N_28793,N_27990,N_27985);
or U28794 (N_28794,N_27790,N_28098);
nand U28795 (N_28795,N_27716,N_28199);
or U28796 (N_28796,N_28051,N_27823);
and U28797 (N_28797,N_27748,N_27738);
nor U28798 (N_28798,N_27766,N_27854);
and U28799 (N_28799,N_28014,N_28001);
nand U28800 (N_28800,N_28261,N_28344);
nand U28801 (N_28801,N_28770,N_28517);
xnor U28802 (N_28802,N_28444,N_28438);
nor U28803 (N_28803,N_28667,N_28233);
nand U28804 (N_28804,N_28270,N_28217);
nand U28805 (N_28805,N_28677,N_28469);
xor U28806 (N_28806,N_28293,N_28290);
and U28807 (N_28807,N_28616,N_28523);
xor U28808 (N_28808,N_28708,N_28568);
xnor U28809 (N_28809,N_28787,N_28447);
nor U28810 (N_28810,N_28572,N_28535);
and U28811 (N_28811,N_28487,N_28796);
or U28812 (N_28812,N_28686,N_28559);
or U28813 (N_28813,N_28727,N_28521);
nand U28814 (N_28814,N_28285,N_28624);
xnor U28815 (N_28815,N_28751,N_28382);
nand U28816 (N_28816,N_28211,N_28370);
nand U28817 (N_28817,N_28338,N_28530);
nand U28818 (N_28818,N_28248,N_28458);
nand U28819 (N_28819,N_28761,N_28341);
and U28820 (N_28820,N_28762,N_28273);
nand U28821 (N_28821,N_28281,N_28703);
nand U28822 (N_28822,N_28631,N_28561);
xor U28823 (N_28823,N_28556,N_28260);
and U28824 (N_28824,N_28660,N_28543);
nand U28825 (N_28825,N_28700,N_28665);
or U28826 (N_28826,N_28429,N_28691);
and U28827 (N_28827,N_28606,N_28736);
nand U28828 (N_28828,N_28268,N_28671);
or U28829 (N_28829,N_28701,N_28308);
or U28830 (N_28830,N_28760,N_28638);
and U28831 (N_28831,N_28764,N_28239);
and U28832 (N_28832,N_28777,N_28299);
nor U28833 (N_28833,N_28611,N_28791);
nor U28834 (N_28834,N_28790,N_28361);
xor U28835 (N_28835,N_28250,N_28694);
nor U28836 (N_28836,N_28367,N_28402);
xor U28837 (N_28837,N_28567,N_28702);
or U28838 (N_28838,N_28358,N_28291);
xor U28839 (N_28839,N_28496,N_28489);
xnor U28840 (N_28840,N_28715,N_28235);
xnor U28841 (N_28841,N_28420,N_28735);
nor U28842 (N_28842,N_28615,N_28357);
xor U28843 (N_28843,N_28733,N_28728);
xnor U28844 (N_28844,N_28442,N_28599);
xor U28845 (N_28845,N_28410,N_28474);
or U28846 (N_28846,N_28448,N_28778);
xor U28847 (N_28847,N_28334,N_28242);
or U28848 (N_28848,N_28670,N_28780);
nor U28849 (N_28849,N_28666,N_28722);
nand U28850 (N_28850,N_28411,N_28688);
xnor U28851 (N_28851,N_28204,N_28656);
nand U28852 (N_28852,N_28680,N_28397);
nand U28853 (N_28853,N_28594,N_28513);
or U28854 (N_28854,N_28505,N_28768);
nand U28855 (N_28855,N_28466,N_28421);
xnor U28856 (N_28856,N_28414,N_28560);
nor U28857 (N_28857,N_28277,N_28541);
or U28858 (N_28858,N_28462,N_28351);
nand U28859 (N_28859,N_28659,N_28732);
nand U28860 (N_28860,N_28743,N_28303);
or U28861 (N_28861,N_28409,N_28550);
nand U28862 (N_28862,N_28475,N_28203);
xor U28863 (N_28863,N_28707,N_28704);
and U28864 (N_28864,N_28753,N_28600);
nand U28865 (N_28865,N_28269,N_28364);
nand U28866 (N_28866,N_28349,N_28288);
xnor U28867 (N_28867,N_28548,N_28545);
or U28868 (N_28868,N_28336,N_28380);
or U28869 (N_28869,N_28573,N_28365);
and U28870 (N_28870,N_28637,N_28734);
xor U28871 (N_28871,N_28276,N_28223);
xor U28872 (N_28872,N_28330,N_28418);
xnor U28873 (N_28873,N_28481,N_28316);
and U28874 (N_28874,N_28394,N_28679);
or U28875 (N_28875,N_28328,N_28640);
or U28876 (N_28876,N_28699,N_28214);
xnor U28877 (N_28877,N_28566,N_28354);
nand U28878 (N_28878,N_28746,N_28473);
or U28879 (N_28879,N_28675,N_28588);
or U28880 (N_28880,N_28398,N_28754);
nand U28881 (N_28881,N_28205,N_28445);
nor U28882 (N_28882,N_28546,N_28633);
nor U28883 (N_28883,N_28710,N_28564);
nand U28884 (N_28884,N_28267,N_28283);
or U28885 (N_28885,N_28230,N_28663);
nand U28886 (N_28886,N_28511,N_28292);
and U28887 (N_28887,N_28298,N_28297);
nor U28888 (N_28888,N_28635,N_28578);
xor U28889 (N_28889,N_28782,N_28323);
xor U28890 (N_28890,N_28634,N_28678);
or U28891 (N_28891,N_28621,N_28306);
xor U28892 (N_28892,N_28213,N_28519);
nor U28893 (N_28893,N_28725,N_28717);
or U28894 (N_28894,N_28779,N_28209);
nor U28895 (N_28895,N_28377,N_28212);
and U28896 (N_28896,N_28492,N_28741);
or U28897 (N_28897,N_28747,N_28504);
or U28898 (N_28898,N_28789,N_28221);
nand U28899 (N_28899,N_28372,N_28730);
nand U28900 (N_28900,N_28799,N_28472);
or U28901 (N_28901,N_28431,N_28480);
nand U28902 (N_28902,N_28527,N_28363);
and U28903 (N_28903,N_28580,N_28681);
or U28904 (N_28904,N_28262,N_28646);
and U28905 (N_28905,N_28396,N_28713);
and U28906 (N_28906,N_28430,N_28459);
or U28907 (N_28907,N_28254,N_28247);
and U28908 (N_28908,N_28463,N_28720);
and U28909 (N_28909,N_28416,N_28243);
nor U28910 (N_28910,N_28272,N_28571);
nor U28911 (N_28911,N_28724,N_28238);
and U28912 (N_28912,N_28698,N_28625);
nor U28913 (N_28913,N_28767,N_28661);
or U28914 (N_28914,N_28723,N_28554);
nand U28915 (N_28915,N_28674,N_28352);
xor U28916 (N_28916,N_28765,N_28643);
nor U28917 (N_28917,N_28256,N_28552);
or U28918 (N_28918,N_28692,N_28461);
nor U28919 (N_28919,N_28296,N_28636);
xor U28920 (N_28920,N_28534,N_28451);
xnor U28921 (N_28921,N_28274,N_28423);
xnor U28922 (N_28922,N_28404,N_28426);
and U28923 (N_28923,N_28331,N_28343);
nor U28924 (N_28924,N_28300,N_28479);
and U28925 (N_28925,N_28729,N_28249);
nand U28926 (N_28926,N_28207,N_28391);
xor U28927 (N_28927,N_28798,N_28537);
and U28928 (N_28928,N_28226,N_28584);
xnor U28929 (N_28929,N_28575,N_28645);
nand U28930 (N_28930,N_28648,N_28608);
or U28931 (N_28931,N_28651,N_28266);
or U28932 (N_28932,N_28501,N_28201);
nor U28933 (N_28933,N_28403,N_28325);
nand U28934 (N_28934,N_28289,N_28630);
nand U28935 (N_28935,N_28520,N_28719);
or U28936 (N_28936,N_28539,N_28776);
nor U28937 (N_28937,N_28326,N_28465);
nor U28938 (N_28938,N_28373,N_28607);
nor U28939 (N_28939,N_28467,N_28378);
nor U28940 (N_28940,N_28553,N_28353);
xor U28941 (N_28941,N_28536,N_28622);
nor U28942 (N_28942,N_28485,N_28718);
or U28943 (N_28943,N_28345,N_28440);
and U28944 (N_28944,N_28310,N_28314);
nor U28945 (N_28945,N_28641,N_28533);
nand U28946 (N_28946,N_28785,N_28346);
xnor U28947 (N_28947,N_28200,N_28449);
nor U28948 (N_28948,N_28569,N_28726);
xnor U28949 (N_28949,N_28202,N_28794);
nand U28950 (N_28950,N_28731,N_28781);
or U28951 (N_28951,N_28639,N_28547);
or U28952 (N_28952,N_28453,N_28524);
and U28953 (N_28953,N_28738,N_28225);
xor U28954 (N_28954,N_28313,N_28216);
or U28955 (N_28955,N_28662,N_28763);
or U28956 (N_28956,N_28294,N_28590);
and U28957 (N_28957,N_28356,N_28401);
nand U28958 (N_28958,N_28407,N_28493);
nand U28959 (N_28959,N_28716,N_28251);
or U28960 (N_28960,N_28234,N_28497);
nor U28961 (N_28961,N_28457,N_28450);
and U28962 (N_28962,N_28525,N_28602);
nand U28963 (N_28963,N_28476,N_28333);
nor U28964 (N_28964,N_28437,N_28605);
nand U28965 (N_28965,N_28766,N_28752);
or U28966 (N_28966,N_28478,N_28522);
xor U28967 (N_28967,N_28593,N_28684);
or U28968 (N_28968,N_28379,N_28604);
and U28969 (N_28969,N_28742,N_28603);
nor U28970 (N_28970,N_28287,N_28695);
or U28971 (N_28971,N_28263,N_28388);
xnor U28972 (N_28972,N_28585,N_28755);
nor U28973 (N_28973,N_28312,N_28240);
xnor U28974 (N_28974,N_28516,N_28337);
nor U28975 (N_28975,N_28264,N_28494);
or U28976 (N_28976,N_28750,N_28619);
nand U28977 (N_28977,N_28280,N_28632);
nand U28978 (N_28978,N_28653,N_28406);
and U28979 (N_28979,N_28424,N_28227);
or U28980 (N_28980,N_28508,N_28232);
or U28981 (N_28981,N_28598,N_28446);
nand U28982 (N_28982,N_28721,N_28419);
xor U28983 (N_28983,N_28339,N_28400);
nand U28984 (N_28984,N_28757,N_28460);
nor U28985 (N_28985,N_28540,N_28528);
and U28986 (N_28986,N_28538,N_28577);
or U28987 (N_28987,N_28311,N_28609);
xnor U28988 (N_28988,N_28745,N_28515);
and U28989 (N_28989,N_28626,N_28302);
nor U28990 (N_28990,N_28390,N_28712);
or U28991 (N_28991,N_28512,N_28792);
and U28992 (N_28992,N_28514,N_28434);
and U28993 (N_28993,N_28231,N_28574);
and U28994 (N_28994,N_28284,N_28301);
or U28995 (N_28995,N_28456,N_28687);
nand U28996 (N_28996,N_28652,N_28386);
nor U28997 (N_28997,N_28529,N_28581);
or U28998 (N_28998,N_28773,N_28237);
and U28999 (N_28999,N_28455,N_28384);
xor U29000 (N_29000,N_28433,N_28376);
and U29001 (N_29001,N_28749,N_28595);
or U29002 (N_29002,N_28714,N_28374);
nor U29003 (N_29003,N_28706,N_28241);
nand U29004 (N_29004,N_28244,N_28592);
xor U29005 (N_29005,N_28286,N_28644);
nor U29006 (N_29006,N_28617,N_28558);
nand U29007 (N_29007,N_28542,N_28775);
nand U29008 (N_29008,N_28389,N_28623);
nand U29009 (N_29009,N_28565,N_28486);
nand U29010 (N_29010,N_28642,N_28413);
or U29011 (N_29011,N_28591,N_28618);
xnor U29012 (N_29012,N_28507,N_28464);
nor U29013 (N_29013,N_28366,N_28612);
nor U29014 (N_29014,N_28484,N_28348);
or U29015 (N_29015,N_28555,N_28582);
or U29016 (N_29016,N_28218,N_28347);
or U29017 (N_29017,N_28499,N_28305);
xnor U29018 (N_29018,N_28696,N_28628);
nor U29019 (N_29019,N_28482,N_28549);
xnor U29020 (N_29020,N_28428,N_28422);
xor U29021 (N_29021,N_28509,N_28206);
nand U29022 (N_29022,N_28408,N_28412);
and U29023 (N_29023,N_28253,N_28664);
nand U29024 (N_29024,N_28786,N_28210);
nand U29025 (N_29025,N_28557,N_28693);
and U29026 (N_29026,N_28470,N_28257);
or U29027 (N_29027,N_28208,N_28669);
nand U29028 (N_29028,N_28689,N_28387);
nand U29029 (N_29029,N_28614,N_28375);
xor U29030 (N_29030,N_28368,N_28676);
and U29031 (N_29031,N_28685,N_28335);
or U29032 (N_29032,N_28647,N_28759);
or U29033 (N_29033,N_28705,N_28282);
nor U29034 (N_29034,N_28405,N_28756);
xnor U29035 (N_29035,N_28562,N_28295);
or U29036 (N_29036,N_28246,N_28392);
or U29037 (N_29037,N_28583,N_28435);
xor U29038 (N_29038,N_28551,N_28627);
and U29039 (N_29039,N_28629,N_28769);
nor U29040 (N_29040,N_28531,N_28395);
nand U29041 (N_29041,N_28327,N_28359);
nand U29042 (N_29042,N_28417,N_28672);
nand U29043 (N_29043,N_28441,N_28383);
or U29044 (N_29044,N_28432,N_28252);
or U29045 (N_29045,N_28668,N_28321);
nand U29046 (N_29046,N_28613,N_28657);
xor U29047 (N_29047,N_28381,N_28744);
nand U29048 (N_29048,N_28393,N_28436);
or U29049 (N_29049,N_28362,N_28222);
and U29050 (N_29050,N_28518,N_28307);
nand U29051 (N_29051,N_28255,N_28783);
nand U29052 (N_29052,N_28570,N_28793);
and U29053 (N_29053,N_28771,N_28774);
or U29054 (N_29054,N_28772,N_28697);
nor U29055 (N_29055,N_28491,N_28610);
or U29056 (N_29056,N_28683,N_28526);
or U29057 (N_29057,N_28490,N_28506);
and U29058 (N_29058,N_28690,N_28332);
xnor U29059 (N_29059,N_28737,N_28329);
nand U29060 (N_29060,N_28258,N_28399);
nand U29061 (N_29061,N_28502,N_28318);
nor U29062 (N_29062,N_28649,N_28655);
or U29063 (N_29063,N_28454,N_28620);
or U29064 (N_29064,N_28275,N_28265);
nor U29065 (N_29065,N_28587,N_28650);
xnor U29066 (N_29066,N_28579,N_28215);
and U29067 (N_29067,N_28415,N_28340);
nand U29068 (N_29068,N_28317,N_28740);
nor U29069 (N_29069,N_28360,N_28477);
and U29070 (N_29070,N_28452,N_28350);
nor U29071 (N_29071,N_28425,N_28788);
nand U29072 (N_29072,N_28219,N_28320);
xnor U29073 (N_29073,N_28309,N_28278);
nand U29074 (N_29074,N_28711,N_28601);
or U29075 (N_29075,N_28279,N_28544);
nor U29076 (N_29076,N_28503,N_28224);
and U29077 (N_29077,N_28589,N_28498);
or U29078 (N_29078,N_28563,N_28271);
nor U29079 (N_29079,N_28709,N_28228);
nand U29080 (N_29080,N_28483,N_28532);
nor U29081 (N_29081,N_28784,N_28324);
nor U29082 (N_29082,N_28654,N_28427);
xnor U29083 (N_29083,N_28342,N_28500);
nand U29084 (N_29084,N_28795,N_28658);
nor U29085 (N_29085,N_28385,N_28797);
and U29086 (N_29086,N_28510,N_28229);
nand U29087 (N_29087,N_28748,N_28322);
and U29088 (N_29088,N_28471,N_28586);
or U29089 (N_29089,N_28673,N_28355);
xnor U29090 (N_29090,N_28495,N_28220);
nand U29091 (N_29091,N_28443,N_28369);
xnor U29092 (N_29092,N_28596,N_28468);
nor U29093 (N_29093,N_28245,N_28259);
nand U29094 (N_29094,N_28488,N_28597);
xnor U29095 (N_29095,N_28739,N_28371);
or U29096 (N_29096,N_28439,N_28758);
and U29097 (N_29097,N_28315,N_28304);
nand U29098 (N_29098,N_28236,N_28319);
nand U29099 (N_29099,N_28682,N_28576);
or U29100 (N_29100,N_28530,N_28739);
nand U29101 (N_29101,N_28231,N_28350);
or U29102 (N_29102,N_28522,N_28774);
nor U29103 (N_29103,N_28597,N_28276);
and U29104 (N_29104,N_28492,N_28592);
xor U29105 (N_29105,N_28542,N_28235);
or U29106 (N_29106,N_28468,N_28470);
and U29107 (N_29107,N_28230,N_28432);
xor U29108 (N_29108,N_28765,N_28319);
nor U29109 (N_29109,N_28598,N_28443);
nand U29110 (N_29110,N_28401,N_28224);
or U29111 (N_29111,N_28526,N_28608);
nand U29112 (N_29112,N_28758,N_28633);
xor U29113 (N_29113,N_28202,N_28420);
nor U29114 (N_29114,N_28596,N_28387);
nand U29115 (N_29115,N_28564,N_28345);
nand U29116 (N_29116,N_28713,N_28637);
and U29117 (N_29117,N_28254,N_28424);
and U29118 (N_29118,N_28373,N_28317);
or U29119 (N_29119,N_28212,N_28581);
nor U29120 (N_29120,N_28444,N_28436);
nand U29121 (N_29121,N_28711,N_28481);
nand U29122 (N_29122,N_28358,N_28286);
and U29123 (N_29123,N_28517,N_28738);
nand U29124 (N_29124,N_28566,N_28548);
xor U29125 (N_29125,N_28725,N_28443);
nand U29126 (N_29126,N_28571,N_28768);
or U29127 (N_29127,N_28319,N_28288);
nor U29128 (N_29128,N_28262,N_28548);
or U29129 (N_29129,N_28722,N_28232);
nand U29130 (N_29130,N_28668,N_28566);
or U29131 (N_29131,N_28328,N_28451);
and U29132 (N_29132,N_28265,N_28727);
xnor U29133 (N_29133,N_28652,N_28352);
or U29134 (N_29134,N_28457,N_28399);
xor U29135 (N_29135,N_28375,N_28621);
nand U29136 (N_29136,N_28765,N_28744);
or U29137 (N_29137,N_28717,N_28531);
and U29138 (N_29138,N_28796,N_28477);
nand U29139 (N_29139,N_28486,N_28737);
or U29140 (N_29140,N_28367,N_28527);
xor U29141 (N_29141,N_28601,N_28262);
nand U29142 (N_29142,N_28441,N_28273);
or U29143 (N_29143,N_28494,N_28203);
nand U29144 (N_29144,N_28435,N_28219);
or U29145 (N_29145,N_28644,N_28262);
xnor U29146 (N_29146,N_28796,N_28598);
xor U29147 (N_29147,N_28226,N_28689);
and U29148 (N_29148,N_28315,N_28647);
and U29149 (N_29149,N_28694,N_28541);
nand U29150 (N_29150,N_28636,N_28431);
nand U29151 (N_29151,N_28594,N_28325);
or U29152 (N_29152,N_28586,N_28254);
and U29153 (N_29153,N_28706,N_28625);
nand U29154 (N_29154,N_28798,N_28426);
and U29155 (N_29155,N_28465,N_28565);
or U29156 (N_29156,N_28680,N_28311);
or U29157 (N_29157,N_28255,N_28727);
and U29158 (N_29158,N_28634,N_28433);
nor U29159 (N_29159,N_28427,N_28411);
xnor U29160 (N_29160,N_28756,N_28573);
xor U29161 (N_29161,N_28768,N_28775);
nor U29162 (N_29162,N_28201,N_28526);
and U29163 (N_29163,N_28448,N_28281);
or U29164 (N_29164,N_28586,N_28218);
or U29165 (N_29165,N_28385,N_28764);
xor U29166 (N_29166,N_28703,N_28279);
or U29167 (N_29167,N_28210,N_28585);
nand U29168 (N_29168,N_28217,N_28480);
xor U29169 (N_29169,N_28617,N_28760);
and U29170 (N_29170,N_28346,N_28429);
or U29171 (N_29171,N_28351,N_28204);
nor U29172 (N_29172,N_28434,N_28272);
nor U29173 (N_29173,N_28466,N_28378);
xnor U29174 (N_29174,N_28556,N_28508);
and U29175 (N_29175,N_28488,N_28683);
xor U29176 (N_29176,N_28212,N_28742);
xnor U29177 (N_29177,N_28231,N_28284);
or U29178 (N_29178,N_28369,N_28326);
nor U29179 (N_29179,N_28286,N_28643);
and U29180 (N_29180,N_28765,N_28478);
xnor U29181 (N_29181,N_28348,N_28504);
and U29182 (N_29182,N_28498,N_28627);
or U29183 (N_29183,N_28274,N_28797);
xnor U29184 (N_29184,N_28564,N_28765);
nand U29185 (N_29185,N_28315,N_28214);
nor U29186 (N_29186,N_28280,N_28235);
and U29187 (N_29187,N_28472,N_28263);
nand U29188 (N_29188,N_28672,N_28273);
nand U29189 (N_29189,N_28418,N_28214);
nor U29190 (N_29190,N_28319,N_28272);
and U29191 (N_29191,N_28638,N_28784);
nand U29192 (N_29192,N_28769,N_28666);
and U29193 (N_29193,N_28472,N_28520);
or U29194 (N_29194,N_28669,N_28723);
xor U29195 (N_29195,N_28265,N_28321);
xnor U29196 (N_29196,N_28330,N_28494);
xor U29197 (N_29197,N_28367,N_28641);
nor U29198 (N_29198,N_28617,N_28702);
or U29199 (N_29199,N_28271,N_28403);
xnor U29200 (N_29200,N_28280,N_28606);
and U29201 (N_29201,N_28413,N_28211);
or U29202 (N_29202,N_28418,N_28435);
and U29203 (N_29203,N_28778,N_28232);
nand U29204 (N_29204,N_28579,N_28304);
nor U29205 (N_29205,N_28357,N_28435);
nor U29206 (N_29206,N_28664,N_28784);
or U29207 (N_29207,N_28322,N_28377);
or U29208 (N_29208,N_28697,N_28339);
nand U29209 (N_29209,N_28324,N_28573);
nor U29210 (N_29210,N_28333,N_28393);
and U29211 (N_29211,N_28329,N_28724);
nand U29212 (N_29212,N_28419,N_28630);
and U29213 (N_29213,N_28747,N_28535);
and U29214 (N_29214,N_28580,N_28672);
nand U29215 (N_29215,N_28775,N_28407);
or U29216 (N_29216,N_28477,N_28344);
and U29217 (N_29217,N_28722,N_28314);
nor U29218 (N_29218,N_28687,N_28631);
xor U29219 (N_29219,N_28429,N_28222);
or U29220 (N_29220,N_28573,N_28304);
or U29221 (N_29221,N_28485,N_28620);
nor U29222 (N_29222,N_28280,N_28502);
and U29223 (N_29223,N_28725,N_28538);
nand U29224 (N_29224,N_28595,N_28729);
xor U29225 (N_29225,N_28656,N_28738);
and U29226 (N_29226,N_28440,N_28557);
or U29227 (N_29227,N_28229,N_28237);
xnor U29228 (N_29228,N_28457,N_28537);
nor U29229 (N_29229,N_28466,N_28484);
and U29230 (N_29230,N_28390,N_28210);
xor U29231 (N_29231,N_28599,N_28788);
or U29232 (N_29232,N_28772,N_28738);
xor U29233 (N_29233,N_28628,N_28672);
xnor U29234 (N_29234,N_28624,N_28720);
and U29235 (N_29235,N_28426,N_28594);
or U29236 (N_29236,N_28446,N_28516);
or U29237 (N_29237,N_28707,N_28523);
xnor U29238 (N_29238,N_28457,N_28434);
nor U29239 (N_29239,N_28365,N_28771);
or U29240 (N_29240,N_28494,N_28377);
or U29241 (N_29241,N_28551,N_28263);
nor U29242 (N_29242,N_28706,N_28661);
or U29243 (N_29243,N_28684,N_28202);
or U29244 (N_29244,N_28732,N_28427);
or U29245 (N_29245,N_28680,N_28508);
and U29246 (N_29246,N_28413,N_28551);
nor U29247 (N_29247,N_28533,N_28534);
or U29248 (N_29248,N_28416,N_28468);
xnor U29249 (N_29249,N_28222,N_28252);
or U29250 (N_29250,N_28445,N_28232);
or U29251 (N_29251,N_28492,N_28515);
and U29252 (N_29252,N_28726,N_28214);
xor U29253 (N_29253,N_28624,N_28704);
nor U29254 (N_29254,N_28728,N_28281);
nand U29255 (N_29255,N_28664,N_28498);
nor U29256 (N_29256,N_28294,N_28688);
or U29257 (N_29257,N_28506,N_28647);
xor U29258 (N_29258,N_28661,N_28791);
xor U29259 (N_29259,N_28489,N_28692);
nand U29260 (N_29260,N_28692,N_28293);
or U29261 (N_29261,N_28401,N_28675);
and U29262 (N_29262,N_28224,N_28609);
xor U29263 (N_29263,N_28734,N_28248);
nand U29264 (N_29264,N_28258,N_28642);
nor U29265 (N_29265,N_28689,N_28708);
nand U29266 (N_29266,N_28294,N_28346);
nand U29267 (N_29267,N_28452,N_28620);
xnor U29268 (N_29268,N_28681,N_28686);
and U29269 (N_29269,N_28798,N_28271);
nor U29270 (N_29270,N_28684,N_28524);
nor U29271 (N_29271,N_28752,N_28331);
or U29272 (N_29272,N_28222,N_28258);
and U29273 (N_29273,N_28390,N_28640);
nand U29274 (N_29274,N_28334,N_28617);
and U29275 (N_29275,N_28621,N_28258);
or U29276 (N_29276,N_28779,N_28756);
and U29277 (N_29277,N_28569,N_28580);
and U29278 (N_29278,N_28419,N_28542);
and U29279 (N_29279,N_28667,N_28540);
xnor U29280 (N_29280,N_28374,N_28543);
and U29281 (N_29281,N_28617,N_28389);
or U29282 (N_29282,N_28506,N_28788);
nand U29283 (N_29283,N_28291,N_28616);
nand U29284 (N_29284,N_28381,N_28261);
and U29285 (N_29285,N_28219,N_28781);
xnor U29286 (N_29286,N_28631,N_28265);
nand U29287 (N_29287,N_28788,N_28547);
nand U29288 (N_29288,N_28289,N_28746);
and U29289 (N_29289,N_28388,N_28402);
or U29290 (N_29290,N_28239,N_28760);
nor U29291 (N_29291,N_28718,N_28346);
nor U29292 (N_29292,N_28445,N_28428);
nor U29293 (N_29293,N_28303,N_28607);
and U29294 (N_29294,N_28772,N_28308);
nand U29295 (N_29295,N_28339,N_28630);
and U29296 (N_29296,N_28657,N_28543);
xnor U29297 (N_29297,N_28210,N_28705);
nor U29298 (N_29298,N_28598,N_28678);
xnor U29299 (N_29299,N_28361,N_28678);
nand U29300 (N_29300,N_28303,N_28660);
nor U29301 (N_29301,N_28781,N_28347);
and U29302 (N_29302,N_28578,N_28365);
xor U29303 (N_29303,N_28408,N_28607);
xor U29304 (N_29304,N_28612,N_28686);
nand U29305 (N_29305,N_28349,N_28201);
or U29306 (N_29306,N_28579,N_28517);
nand U29307 (N_29307,N_28452,N_28527);
or U29308 (N_29308,N_28377,N_28532);
nand U29309 (N_29309,N_28237,N_28531);
and U29310 (N_29310,N_28764,N_28673);
and U29311 (N_29311,N_28555,N_28276);
nor U29312 (N_29312,N_28777,N_28379);
nand U29313 (N_29313,N_28649,N_28499);
nor U29314 (N_29314,N_28213,N_28399);
xnor U29315 (N_29315,N_28487,N_28481);
and U29316 (N_29316,N_28379,N_28582);
xnor U29317 (N_29317,N_28730,N_28256);
nand U29318 (N_29318,N_28721,N_28376);
and U29319 (N_29319,N_28468,N_28523);
and U29320 (N_29320,N_28581,N_28315);
and U29321 (N_29321,N_28643,N_28248);
xnor U29322 (N_29322,N_28641,N_28483);
nand U29323 (N_29323,N_28702,N_28459);
nand U29324 (N_29324,N_28501,N_28513);
nor U29325 (N_29325,N_28255,N_28781);
and U29326 (N_29326,N_28455,N_28311);
nor U29327 (N_29327,N_28340,N_28782);
and U29328 (N_29328,N_28265,N_28566);
and U29329 (N_29329,N_28425,N_28289);
and U29330 (N_29330,N_28533,N_28509);
nor U29331 (N_29331,N_28548,N_28522);
nor U29332 (N_29332,N_28738,N_28309);
nand U29333 (N_29333,N_28692,N_28294);
nand U29334 (N_29334,N_28580,N_28728);
and U29335 (N_29335,N_28783,N_28768);
xnor U29336 (N_29336,N_28262,N_28590);
nand U29337 (N_29337,N_28483,N_28679);
or U29338 (N_29338,N_28610,N_28425);
or U29339 (N_29339,N_28619,N_28675);
nand U29340 (N_29340,N_28781,N_28298);
or U29341 (N_29341,N_28594,N_28634);
nor U29342 (N_29342,N_28243,N_28608);
xor U29343 (N_29343,N_28262,N_28459);
or U29344 (N_29344,N_28712,N_28416);
or U29345 (N_29345,N_28623,N_28789);
nor U29346 (N_29346,N_28740,N_28302);
and U29347 (N_29347,N_28786,N_28325);
nor U29348 (N_29348,N_28781,N_28367);
xnor U29349 (N_29349,N_28477,N_28519);
xor U29350 (N_29350,N_28568,N_28466);
or U29351 (N_29351,N_28536,N_28772);
or U29352 (N_29352,N_28402,N_28561);
nor U29353 (N_29353,N_28316,N_28309);
nand U29354 (N_29354,N_28478,N_28378);
and U29355 (N_29355,N_28604,N_28698);
xnor U29356 (N_29356,N_28675,N_28643);
xor U29357 (N_29357,N_28578,N_28567);
nand U29358 (N_29358,N_28210,N_28665);
nand U29359 (N_29359,N_28460,N_28476);
and U29360 (N_29360,N_28642,N_28767);
nand U29361 (N_29361,N_28576,N_28262);
nand U29362 (N_29362,N_28333,N_28574);
xor U29363 (N_29363,N_28388,N_28363);
nand U29364 (N_29364,N_28554,N_28213);
or U29365 (N_29365,N_28739,N_28794);
nand U29366 (N_29366,N_28642,N_28752);
xor U29367 (N_29367,N_28267,N_28336);
and U29368 (N_29368,N_28270,N_28223);
xnor U29369 (N_29369,N_28753,N_28616);
nor U29370 (N_29370,N_28433,N_28638);
or U29371 (N_29371,N_28231,N_28566);
nand U29372 (N_29372,N_28391,N_28428);
xnor U29373 (N_29373,N_28678,N_28566);
nand U29374 (N_29374,N_28606,N_28313);
and U29375 (N_29375,N_28716,N_28371);
or U29376 (N_29376,N_28749,N_28239);
or U29377 (N_29377,N_28476,N_28264);
xnor U29378 (N_29378,N_28560,N_28411);
and U29379 (N_29379,N_28241,N_28710);
xnor U29380 (N_29380,N_28504,N_28655);
xor U29381 (N_29381,N_28770,N_28231);
nor U29382 (N_29382,N_28224,N_28561);
nand U29383 (N_29383,N_28212,N_28369);
or U29384 (N_29384,N_28373,N_28695);
nand U29385 (N_29385,N_28640,N_28609);
nand U29386 (N_29386,N_28299,N_28706);
nor U29387 (N_29387,N_28339,N_28763);
nor U29388 (N_29388,N_28403,N_28328);
nor U29389 (N_29389,N_28636,N_28790);
or U29390 (N_29390,N_28695,N_28311);
and U29391 (N_29391,N_28469,N_28770);
or U29392 (N_29392,N_28252,N_28319);
nor U29393 (N_29393,N_28449,N_28495);
xor U29394 (N_29394,N_28503,N_28612);
nand U29395 (N_29395,N_28474,N_28370);
nor U29396 (N_29396,N_28487,N_28751);
and U29397 (N_29397,N_28758,N_28722);
and U29398 (N_29398,N_28441,N_28735);
xnor U29399 (N_29399,N_28277,N_28662);
and U29400 (N_29400,N_29222,N_29362);
nor U29401 (N_29401,N_29034,N_29159);
xor U29402 (N_29402,N_28913,N_28886);
and U29403 (N_29403,N_29345,N_29020);
or U29404 (N_29404,N_28853,N_28863);
nor U29405 (N_29405,N_28993,N_28815);
or U29406 (N_29406,N_29316,N_29381);
nand U29407 (N_29407,N_28986,N_29385);
nor U29408 (N_29408,N_29231,N_28874);
nand U29409 (N_29409,N_29165,N_28946);
xor U29410 (N_29410,N_28884,N_28980);
xnor U29411 (N_29411,N_29321,N_29080);
nor U29412 (N_29412,N_29185,N_29326);
and U29413 (N_29413,N_28995,N_28933);
xnor U29414 (N_29414,N_28904,N_29086);
or U29415 (N_29415,N_28911,N_29047);
nand U29416 (N_29416,N_28826,N_29073);
xnor U29417 (N_29417,N_29288,N_29143);
xnor U29418 (N_29418,N_29351,N_29352);
nand U29419 (N_29419,N_29277,N_28875);
nand U29420 (N_29420,N_29271,N_28991);
nor U29421 (N_29421,N_28846,N_28998);
and U29422 (N_29422,N_29037,N_28961);
nand U29423 (N_29423,N_29105,N_29010);
or U29424 (N_29424,N_28811,N_29066);
and U29425 (N_29425,N_29386,N_29198);
and U29426 (N_29426,N_29358,N_29071);
xnor U29427 (N_29427,N_29097,N_29171);
or U29428 (N_29428,N_29084,N_29077);
nand U29429 (N_29429,N_29335,N_28832);
xor U29430 (N_29430,N_29221,N_28951);
nor U29431 (N_29431,N_28974,N_28966);
or U29432 (N_29432,N_28841,N_29090);
or U29433 (N_29433,N_28836,N_29272);
xnor U29434 (N_29434,N_29180,N_28804);
nor U29435 (N_29435,N_29327,N_29085);
xnor U29436 (N_29436,N_29233,N_28945);
and U29437 (N_29437,N_29348,N_28947);
nand U29438 (N_29438,N_28979,N_28950);
and U29439 (N_29439,N_28916,N_29065);
nand U29440 (N_29440,N_29078,N_29319);
nand U29441 (N_29441,N_28935,N_29164);
nor U29442 (N_29442,N_29199,N_29259);
and U29443 (N_29443,N_29098,N_29058);
or U29444 (N_29444,N_28909,N_28956);
nor U29445 (N_29445,N_29242,N_29330);
and U29446 (N_29446,N_29117,N_29152);
xor U29447 (N_29447,N_29081,N_29336);
and U29448 (N_29448,N_28807,N_29009);
xnor U29449 (N_29449,N_29234,N_29297);
nor U29450 (N_29450,N_29060,N_29119);
or U29451 (N_29451,N_29120,N_29217);
nand U29452 (N_29452,N_29295,N_29053);
nand U29453 (N_29453,N_28900,N_29001);
nor U29454 (N_29454,N_29167,N_29377);
or U29455 (N_29455,N_29156,N_29162);
nor U29456 (N_29456,N_29170,N_29032);
nor U29457 (N_29457,N_29296,N_29359);
xor U29458 (N_29458,N_29372,N_29396);
nor U29459 (N_29459,N_29252,N_29107);
xnor U29460 (N_29460,N_29339,N_29289);
xnor U29461 (N_29461,N_29276,N_29137);
nand U29462 (N_29462,N_28849,N_28948);
nand U29463 (N_29463,N_28862,N_29063);
nand U29464 (N_29464,N_29203,N_29240);
or U29465 (N_29465,N_28924,N_29184);
nand U29466 (N_29466,N_29226,N_29031);
and U29467 (N_29467,N_29318,N_28859);
nand U29468 (N_29468,N_28960,N_28883);
or U29469 (N_29469,N_29310,N_29245);
and U29470 (N_29470,N_28972,N_29347);
or U29471 (N_29471,N_29102,N_29390);
nor U29472 (N_29472,N_29267,N_28871);
xnor U29473 (N_29473,N_29148,N_28968);
and U29474 (N_29474,N_29087,N_29304);
or U29475 (N_29475,N_29215,N_29206);
and U29476 (N_29476,N_28821,N_29363);
or U29477 (N_29477,N_29298,N_29354);
nor U29478 (N_29478,N_29302,N_29290);
and U29479 (N_29479,N_29204,N_29263);
nand U29480 (N_29480,N_29168,N_28930);
xor U29481 (N_29481,N_29025,N_29052);
or U29482 (N_29482,N_29370,N_29173);
nand U29483 (N_29483,N_28828,N_29187);
and U29484 (N_29484,N_28982,N_29264);
nor U29485 (N_29485,N_29213,N_28850);
xor U29486 (N_29486,N_29244,N_29067);
and U29487 (N_29487,N_29256,N_29192);
and U29488 (N_29488,N_29306,N_28905);
and U29489 (N_29489,N_28941,N_29328);
and U29490 (N_29490,N_28997,N_29398);
nand U29491 (N_29491,N_29301,N_28842);
nand U29492 (N_29492,N_29103,N_28838);
or U29493 (N_29493,N_28805,N_28897);
and U29494 (N_29494,N_29388,N_29254);
or U29495 (N_29495,N_28877,N_29135);
nor U29496 (N_29496,N_29273,N_29161);
nor U29497 (N_29497,N_28989,N_29142);
nor U29498 (N_29498,N_28919,N_29323);
nor U29499 (N_29499,N_28891,N_28880);
or U29500 (N_29500,N_29341,N_28819);
nand U29501 (N_29501,N_29279,N_28810);
nor U29502 (N_29502,N_29131,N_28867);
xor U29503 (N_29503,N_28834,N_29208);
xor U29504 (N_29504,N_29228,N_28845);
or U29505 (N_29505,N_29325,N_29030);
nand U29506 (N_29506,N_29041,N_29366);
xnor U29507 (N_29507,N_29261,N_28872);
nor U29508 (N_29508,N_29044,N_29106);
nor U29509 (N_29509,N_29183,N_29286);
nor U29510 (N_29510,N_29280,N_28975);
xnor U29511 (N_29511,N_29145,N_29054);
nor U29512 (N_29512,N_29068,N_29178);
nor U29513 (N_29513,N_29257,N_29153);
nand U29514 (N_29514,N_29196,N_28990);
and U29515 (N_29515,N_29380,N_29337);
xor U29516 (N_29516,N_29344,N_29223);
xnor U29517 (N_29517,N_29013,N_29056);
nand U29518 (N_29518,N_29284,N_29094);
nor U29519 (N_29519,N_29309,N_28940);
nor U29520 (N_29520,N_28813,N_29003);
nand U29521 (N_29521,N_29104,N_28976);
and U29522 (N_29522,N_29093,N_29195);
nand U29523 (N_29523,N_29146,N_28868);
or U29524 (N_29524,N_28923,N_28823);
nand U29525 (N_29525,N_28920,N_29389);
and U29526 (N_29526,N_28939,N_29250);
nand U29527 (N_29527,N_29128,N_29384);
nor U29528 (N_29528,N_28906,N_29134);
nand U29529 (N_29529,N_29189,N_28914);
nor U29530 (N_29530,N_29191,N_29157);
nand U29531 (N_29531,N_29091,N_28866);
or U29532 (N_29532,N_29059,N_29110);
xor U29533 (N_29533,N_29202,N_29308);
nand U29534 (N_29534,N_29227,N_29055);
or U29535 (N_29535,N_29114,N_29023);
nand U29536 (N_29536,N_29334,N_29311);
nor U29537 (N_29537,N_29040,N_28944);
xor U29538 (N_29538,N_28921,N_29082);
nand U29539 (N_29539,N_29194,N_28889);
or U29540 (N_29540,N_28912,N_28808);
and U29541 (N_29541,N_28926,N_29241);
or U29542 (N_29542,N_29147,N_29004);
xnor U29543 (N_29543,N_29355,N_29265);
and U29544 (N_29544,N_29207,N_28977);
nand U29545 (N_29545,N_28869,N_29266);
nand U29546 (N_29546,N_28927,N_29230);
xnor U29547 (N_29547,N_29375,N_28844);
and U29548 (N_29548,N_28999,N_29211);
nor U29549 (N_29549,N_29190,N_28931);
nand U29550 (N_29550,N_29038,N_29101);
and U29551 (N_29551,N_28822,N_28988);
nor U29552 (N_29552,N_29006,N_29281);
nor U29553 (N_29553,N_28981,N_29033);
and U29554 (N_29554,N_28802,N_28858);
or U29555 (N_29555,N_29070,N_29018);
and U29556 (N_29556,N_29155,N_29229);
or U29557 (N_29557,N_29210,N_29099);
and U29558 (N_29558,N_28922,N_29039);
nor U29559 (N_29559,N_29140,N_29092);
or U29560 (N_29560,N_29019,N_29393);
and U29561 (N_29561,N_28907,N_29166);
nand U29562 (N_29562,N_29248,N_29305);
or U29563 (N_29563,N_29343,N_29239);
nand U29564 (N_29564,N_29181,N_28820);
xor U29565 (N_29565,N_29219,N_29200);
and U29566 (N_29566,N_29176,N_29216);
nor U29567 (N_29567,N_29232,N_28952);
or U29568 (N_29568,N_28861,N_28894);
and U29569 (N_29569,N_29111,N_29121);
xor U29570 (N_29570,N_28840,N_29046);
or U29571 (N_29571,N_29365,N_29075);
nand U29572 (N_29572,N_28817,N_29303);
nand U29573 (N_29573,N_29236,N_28984);
xor U29574 (N_29574,N_29291,N_29247);
nand U29575 (N_29575,N_29154,N_29238);
xor U29576 (N_29576,N_29048,N_28896);
or U29577 (N_29577,N_29011,N_29374);
nor U29578 (N_29578,N_28812,N_29074);
and U29579 (N_29579,N_29262,N_29283);
nand U29580 (N_29580,N_29095,N_29397);
and U29581 (N_29581,N_29144,N_29324);
or U29582 (N_29582,N_28870,N_28954);
nor U29583 (N_29583,N_29116,N_29367);
xnor U29584 (N_29584,N_29069,N_29005);
xor U29585 (N_29585,N_28852,N_28965);
or U29586 (N_29586,N_29149,N_28854);
or U29587 (N_29587,N_29287,N_28942);
or U29588 (N_29588,N_28903,N_29130);
nor U29589 (N_29589,N_28809,N_28806);
nand U29590 (N_29590,N_29050,N_29051);
xor U29591 (N_29591,N_28899,N_29282);
xor U29592 (N_29592,N_28892,N_29182);
and U29593 (N_29593,N_29392,N_29373);
xnor U29594 (N_29594,N_28833,N_29399);
xor U29595 (N_29595,N_29395,N_29057);
nor U29596 (N_29596,N_28978,N_29260);
nor U29597 (N_29597,N_29109,N_28901);
nand U29598 (N_29598,N_29076,N_29123);
xnor U29599 (N_29599,N_29061,N_29017);
nor U29600 (N_29600,N_29320,N_28938);
nor U29601 (N_29601,N_29079,N_29322);
and U29602 (N_29602,N_29249,N_29338);
and U29603 (N_29603,N_29193,N_28888);
nand U29604 (N_29604,N_29258,N_29350);
and U29605 (N_29605,N_28800,N_28918);
and U29606 (N_29606,N_29112,N_28837);
xor U29607 (N_29607,N_29064,N_29382);
or U29608 (N_29608,N_29270,N_28992);
nor U29609 (N_29609,N_29138,N_29314);
nand U29610 (N_29610,N_29133,N_29225);
xor U29611 (N_29611,N_29361,N_28856);
xnor U29612 (N_29612,N_29042,N_29124);
and U29613 (N_29613,N_29356,N_28855);
nand U29614 (N_29614,N_29237,N_29049);
nor U29615 (N_29615,N_29235,N_29293);
xor U29616 (N_29616,N_29294,N_29022);
or U29617 (N_29617,N_28835,N_28898);
or U29618 (N_29618,N_28973,N_28848);
nor U29619 (N_29619,N_29072,N_29368);
nand U29620 (N_29620,N_28873,N_29333);
nor U29621 (N_29621,N_29197,N_29088);
or U29622 (N_29622,N_28893,N_29122);
nand U29623 (N_29623,N_28937,N_29150);
or U29624 (N_29624,N_29172,N_29364);
and U29625 (N_29625,N_28879,N_29186);
nor U29626 (N_29626,N_29127,N_29315);
nand U29627 (N_29627,N_29027,N_29205);
nand U29628 (N_29628,N_29371,N_29201);
nor U29629 (N_29629,N_29243,N_28949);
nand U29630 (N_29630,N_28887,N_28851);
and U29631 (N_29631,N_29307,N_28908);
and U29632 (N_29632,N_28929,N_29118);
xor U29633 (N_29633,N_29224,N_28890);
xnor U29634 (N_29634,N_29214,N_28818);
nand U29635 (N_29635,N_28928,N_28843);
nor U29636 (N_29636,N_29342,N_29021);
or U29637 (N_29637,N_29340,N_28934);
nor U29638 (N_29638,N_29285,N_28994);
xnor U29639 (N_29639,N_29028,N_29132);
or U29640 (N_29640,N_28983,N_28996);
nand U29641 (N_29641,N_29312,N_29353);
nor U29642 (N_29642,N_28957,N_29062);
xnor U29643 (N_29643,N_29126,N_28970);
nand U29644 (N_29644,N_29043,N_28953);
or U29645 (N_29645,N_29188,N_29125);
or U29646 (N_29646,N_29002,N_29169);
and U29647 (N_29647,N_29349,N_29100);
xor U29648 (N_29648,N_29163,N_29151);
and U29649 (N_29649,N_29139,N_29275);
and U29650 (N_29650,N_29383,N_29278);
nor U29651 (N_29651,N_28881,N_29220);
xor U29652 (N_29652,N_28829,N_28865);
xor U29653 (N_29653,N_29015,N_29357);
nor U29654 (N_29654,N_28932,N_28878);
xnor U29655 (N_29655,N_28839,N_29141);
nor U29656 (N_29656,N_29036,N_28876);
or U29657 (N_29657,N_29269,N_28803);
nand U29658 (N_29658,N_29376,N_28827);
xor U29659 (N_29659,N_29212,N_29083);
xor U29660 (N_29660,N_29299,N_29113);
and U29661 (N_29661,N_28964,N_29007);
nor U29662 (N_29662,N_28985,N_29012);
or U29663 (N_29663,N_28831,N_29253);
nor U29664 (N_29664,N_29332,N_28971);
and U29665 (N_29665,N_29158,N_28857);
and U29666 (N_29666,N_29174,N_29251);
and U29667 (N_29667,N_28816,N_28943);
xnor U29668 (N_29668,N_28814,N_29292);
and U29669 (N_29669,N_29014,N_28801);
nand U29670 (N_29670,N_29089,N_29029);
and U29671 (N_29671,N_29209,N_28962);
nor U29672 (N_29672,N_29313,N_29331);
or U29673 (N_29673,N_28967,N_29160);
nand U29674 (N_29674,N_28955,N_28825);
nor U29675 (N_29675,N_29394,N_28969);
or U29676 (N_29676,N_29179,N_29115);
nor U29677 (N_29677,N_29379,N_29026);
nand U29678 (N_29678,N_29391,N_29255);
nand U29679 (N_29679,N_28910,N_29175);
or U29680 (N_29680,N_28987,N_28830);
xnor U29681 (N_29681,N_28959,N_28958);
or U29682 (N_29682,N_29024,N_28915);
and U29683 (N_29683,N_28925,N_28847);
nor U29684 (N_29684,N_28885,N_29360);
nor U29685 (N_29685,N_29008,N_29000);
and U29686 (N_29686,N_29016,N_28824);
and U29687 (N_29687,N_29136,N_28895);
nor U29688 (N_29688,N_29096,N_29378);
nor U29689 (N_29689,N_29246,N_28902);
or U29690 (N_29690,N_29317,N_28936);
nor U29691 (N_29691,N_29369,N_28917);
nand U29692 (N_29692,N_29108,N_28864);
nand U29693 (N_29693,N_29329,N_29177);
xnor U29694 (N_29694,N_29268,N_28860);
or U29695 (N_29695,N_29346,N_29035);
xnor U29696 (N_29696,N_28963,N_29274);
xor U29697 (N_29697,N_29129,N_28882);
and U29698 (N_29698,N_29387,N_29045);
nor U29699 (N_29699,N_29218,N_29300);
nor U29700 (N_29700,N_29073,N_29035);
and U29701 (N_29701,N_29283,N_29347);
xnor U29702 (N_29702,N_28993,N_29321);
and U29703 (N_29703,N_29357,N_28926);
nor U29704 (N_29704,N_28963,N_29001);
or U29705 (N_29705,N_29209,N_29239);
nand U29706 (N_29706,N_29390,N_29356);
or U29707 (N_29707,N_28992,N_28829);
nand U29708 (N_29708,N_29257,N_29118);
or U29709 (N_29709,N_29298,N_29262);
xnor U29710 (N_29710,N_29324,N_29385);
or U29711 (N_29711,N_29375,N_29102);
xor U29712 (N_29712,N_29362,N_28901);
and U29713 (N_29713,N_29175,N_28830);
nand U29714 (N_29714,N_29146,N_29300);
or U29715 (N_29715,N_29098,N_28850);
or U29716 (N_29716,N_29349,N_29377);
xor U29717 (N_29717,N_29195,N_28946);
nand U29718 (N_29718,N_28989,N_29354);
nand U29719 (N_29719,N_28804,N_28950);
xnor U29720 (N_29720,N_29246,N_28923);
xor U29721 (N_29721,N_29394,N_29072);
and U29722 (N_29722,N_29017,N_29072);
nor U29723 (N_29723,N_29181,N_28866);
xor U29724 (N_29724,N_28939,N_29044);
xnor U29725 (N_29725,N_29396,N_29235);
xor U29726 (N_29726,N_29192,N_29200);
and U29727 (N_29727,N_28924,N_29101);
nand U29728 (N_29728,N_28985,N_29321);
and U29729 (N_29729,N_28929,N_29053);
nand U29730 (N_29730,N_29041,N_29376);
nor U29731 (N_29731,N_29322,N_29281);
xnor U29732 (N_29732,N_29098,N_29164);
nor U29733 (N_29733,N_29357,N_28867);
or U29734 (N_29734,N_29292,N_29229);
nand U29735 (N_29735,N_29141,N_28880);
or U29736 (N_29736,N_29304,N_28963);
or U29737 (N_29737,N_29001,N_29119);
and U29738 (N_29738,N_28868,N_29166);
or U29739 (N_29739,N_29378,N_29310);
xnor U29740 (N_29740,N_29374,N_28991);
nor U29741 (N_29741,N_29012,N_28839);
xor U29742 (N_29742,N_29276,N_28818);
nand U29743 (N_29743,N_29038,N_28920);
or U29744 (N_29744,N_29086,N_29023);
nand U29745 (N_29745,N_28836,N_29061);
nand U29746 (N_29746,N_28892,N_28808);
nand U29747 (N_29747,N_29002,N_29036);
nor U29748 (N_29748,N_29341,N_28824);
nor U29749 (N_29749,N_29241,N_28947);
nor U29750 (N_29750,N_29305,N_29188);
nor U29751 (N_29751,N_28984,N_29015);
and U29752 (N_29752,N_29156,N_28856);
xnor U29753 (N_29753,N_29183,N_28876);
or U29754 (N_29754,N_29174,N_28919);
or U29755 (N_29755,N_29151,N_29327);
nor U29756 (N_29756,N_28989,N_29323);
nor U29757 (N_29757,N_29245,N_28810);
xnor U29758 (N_29758,N_28899,N_29009);
xor U29759 (N_29759,N_29374,N_29063);
and U29760 (N_29760,N_29017,N_29242);
xor U29761 (N_29761,N_29093,N_29143);
or U29762 (N_29762,N_29369,N_29129);
and U29763 (N_29763,N_28995,N_29030);
and U29764 (N_29764,N_29155,N_29352);
or U29765 (N_29765,N_29269,N_28811);
nand U29766 (N_29766,N_29299,N_28838);
nand U29767 (N_29767,N_29066,N_28814);
nand U29768 (N_29768,N_28801,N_28930);
xnor U29769 (N_29769,N_29219,N_29268);
nand U29770 (N_29770,N_29307,N_28991);
nand U29771 (N_29771,N_29363,N_29328);
xor U29772 (N_29772,N_29187,N_28843);
xor U29773 (N_29773,N_29076,N_29063);
and U29774 (N_29774,N_28815,N_29319);
nor U29775 (N_29775,N_29151,N_29186);
nand U29776 (N_29776,N_29222,N_28822);
and U29777 (N_29777,N_28805,N_29249);
nor U29778 (N_29778,N_28906,N_29344);
nand U29779 (N_29779,N_29111,N_28886);
nor U29780 (N_29780,N_29055,N_28914);
xor U29781 (N_29781,N_29036,N_29129);
or U29782 (N_29782,N_29282,N_28986);
nor U29783 (N_29783,N_29036,N_28973);
nor U29784 (N_29784,N_29358,N_29231);
nor U29785 (N_29785,N_29308,N_28857);
or U29786 (N_29786,N_29326,N_28960);
xnor U29787 (N_29787,N_29030,N_29312);
and U29788 (N_29788,N_29341,N_29027);
and U29789 (N_29789,N_29185,N_29288);
xor U29790 (N_29790,N_29386,N_29263);
and U29791 (N_29791,N_29314,N_29000);
nor U29792 (N_29792,N_29001,N_28843);
or U29793 (N_29793,N_29263,N_28935);
and U29794 (N_29794,N_28858,N_29245);
or U29795 (N_29795,N_28849,N_29147);
and U29796 (N_29796,N_29335,N_29124);
xnor U29797 (N_29797,N_29350,N_29216);
nand U29798 (N_29798,N_28891,N_29382);
nor U29799 (N_29799,N_29145,N_29045);
and U29800 (N_29800,N_29311,N_29120);
nand U29801 (N_29801,N_29118,N_28848);
nand U29802 (N_29802,N_29227,N_29203);
nand U29803 (N_29803,N_28996,N_28989);
or U29804 (N_29804,N_28842,N_29221);
nor U29805 (N_29805,N_28908,N_29291);
xnor U29806 (N_29806,N_29256,N_28985);
or U29807 (N_29807,N_29028,N_29074);
xor U29808 (N_29808,N_29155,N_29234);
xor U29809 (N_29809,N_29317,N_29081);
nand U29810 (N_29810,N_29169,N_28993);
nor U29811 (N_29811,N_28848,N_29314);
and U29812 (N_29812,N_29014,N_28985);
xor U29813 (N_29813,N_29083,N_29214);
or U29814 (N_29814,N_28997,N_29334);
or U29815 (N_29815,N_29213,N_28949);
or U29816 (N_29816,N_29064,N_29239);
or U29817 (N_29817,N_29252,N_29291);
or U29818 (N_29818,N_29372,N_28975);
nand U29819 (N_29819,N_29218,N_28840);
nand U29820 (N_29820,N_29171,N_28903);
or U29821 (N_29821,N_28851,N_28800);
and U29822 (N_29822,N_29109,N_28836);
nor U29823 (N_29823,N_29104,N_29278);
xor U29824 (N_29824,N_29149,N_29177);
nor U29825 (N_29825,N_29201,N_29146);
or U29826 (N_29826,N_29346,N_29293);
and U29827 (N_29827,N_29235,N_29284);
xnor U29828 (N_29828,N_28847,N_29322);
nor U29829 (N_29829,N_29017,N_29370);
and U29830 (N_29830,N_29170,N_29334);
xor U29831 (N_29831,N_29252,N_29138);
xor U29832 (N_29832,N_28897,N_28981);
nor U29833 (N_29833,N_28879,N_28850);
nand U29834 (N_29834,N_29274,N_29190);
xor U29835 (N_29835,N_28827,N_28961);
or U29836 (N_29836,N_28942,N_29143);
and U29837 (N_29837,N_29243,N_29159);
and U29838 (N_29838,N_29321,N_29156);
or U29839 (N_29839,N_28935,N_28951);
nand U29840 (N_29840,N_28956,N_28882);
xnor U29841 (N_29841,N_29384,N_28949);
or U29842 (N_29842,N_29285,N_29225);
nor U29843 (N_29843,N_29196,N_28932);
and U29844 (N_29844,N_29025,N_29387);
or U29845 (N_29845,N_29144,N_29161);
or U29846 (N_29846,N_29048,N_29314);
or U29847 (N_29847,N_29340,N_29016);
nand U29848 (N_29848,N_28919,N_29282);
nand U29849 (N_29849,N_28819,N_29191);
nor U29850 (N_29850,N_29128,N_29131);
nor U29851 (N_29851,N_28951,N_28862);
nor U29852 (N_29852,N_29299,N_29168);
xnor U29853 (N_29853,N_28901,N_29004);
nor U29854 (N_29854,N_29136,N_29188);
or U29855 (N_29855,N_29065,N_29131);
nor U29856 (N_29856,N_29142,N_28915);
nand U29857 (N_29857,N_29010,N_28875);
xnor U29858 (N_29858,N_29042,N_29102);
and U29859 (N_29859,N_28951,N_29223);
and U29860 (N_29860,N_29197,N_29191);
or U29861 (N_29861,N_29279,N_28954);
and U29862 (N_29862,N_28957,N_28814);
and U29863 (N_29863,N_29092,N_29330);
and U29864 (N_29864,N_29128,N_29119);
xnor U29865 (N_29865,N_28963,N_29082);
or U29866 (N_29866,N_29362,N_29230);
xnor U29867 (N_29867,N_29313,N_28869);
nand U29868 (N_29868,N_29019,N_29027);
nor U29869 (N_29869,N_28902,N_29055);
xor U29870 (N_29870,N_29191,N_29070);
nand U29871 (N_29871,N_29158,N_29113);
or U29872 (N_29872,N_29208,N_29253);
nand U29873 (N_29873,N_29311,N_29034);
nand U29874 (N_29874,N_29277,N_28901);
xor U29875 (N_29875,N_28832,N_28872);
nand U29876 (N_29876,N_29215,N_29111);
or U29877 (N_29877,N_29244,N_28993);
nor U29878 (N_29878,N_29043,N_29316);
xnor U29879 (N_29879,N_29046,N_29184);
nor U29880 (N_29880,N_29203,N_29122);
or U29881 (N_29881,N_29136,N_29156);
nor U29882 (N_29882,N_28849,N_28959);
xor U29883 (N_29883,N_29093,N_29259);
nor U29884 (N_29884,N_29386,N_29356);
and U29885 (N_29885,N_29109,N_29390);
nand U29886 (N_29886,N_29323,N_29344);
and U29887 (N_29887,N_28829,N_29307);
or U29888 (N_29888,N_29109,N_29238);
nor U29889 (N_29889,N_28854,N_29345);
nand U29890 (N_29890,N_29302,N_29080);
nand U29891 (N_29891,N_28868,N_29091);
xor U29892 (N_29892,N_28828,N_29343);
and U29893 (N_29893,N_29241,N_29201);
and U29894 (N_29894,N_29201,N_28982);
or U29895 (N_29895,N_29364,N_28993);
nand U29896 (N_29896,N_29219,N_29281);
nor U29897 (N_29897,N_28808,N_29103);
or U29898 (N_29898,N_28986,N_29322);
nand U29899 (N_29899,N_29013,N_29344);
xnor U29900 (N_29900,N_29041,N_29019);
nand U29901 (N_29901,N_29042,N_28943);
and U29902 (N_29902,N_29117,N_29098);
and U29903 (N_29903,N_29284,N_28802);
xnor U29904 (N_29904,N_29003,N_29358);
and U29905 (N_29905,N_29042,N_29315);
nand U29906 (N_29906,N_28903,N_29124);
nand U29907 (N_29907,N_29395,N_29099);
or U29908 (N_29908,N_29287,N_29110);
xor U29909 (N_29909,N_29153,N_29040);
and U29910 (N_29910,N_28873,N_29187);
xnor U29911 (N_29911,N_29287,N_29399);
nor U29912 (N_29912,N_29220,N_28911);
nand U29913 (N_29913,N_29198,N_28849);
or U29914 (N_29914,N_28930,N_29357);
xnor U29915 (N_29915,N_28868,N_29199);
and U29916 (N_29916,N_28928,N_29245);
nor U29917 (N_29917,N_29064,N_29062);
or U29918 (N_29918,N_28972,N_28884);
nand U29919 (N_29919,N_28845,N_29350);
xor U29920 (N_29920,N_29120,N_28965);
or U29921 (N_29921,N_28904,N_28995);
nand U29922 (N_29922,N_29162,N_29119);
xor U29923 (N_29923,N_29049,N_28879);
nor U29924 (N_29924,N_29267,N_28935);
and U29925 (N_29925,N_29223,N_28849);
nor U29926 (N_29926,N_29332,N_29042);
nor U29927 (N_29927,N_29009,N_29360);
and U29928 (N_29928,N_28854,N_29293);
or U29929 (N_29929,N_29042,N_29006);
nor U29930 (N_29930,N_29123,N_29030);
nand U29931 (N_29931,N_28984,N_29073);
and U29932 (N_29932,N_28951,N_28903);
nor U29933 (N_29933,N_28996,N_29318);
nor U29934 (N_29934,N_29087,N_29141);
xnor U29935 (N_29935,N_29209,N_29010);
nand U29936 (N_29936,N_29356,N_29157);
and U29937 (N_29937,N_29270,N_29257);
and U29938 (N_29938,N_29154,N_29068);
and U29939 (N_29939,N_29377,N_29302);
or U29940 (N_29940,N_28834,N_29135);
xnor U29941 (N_29941,N_29074,N_29281);
nand U29942 (N_29942,N_29032,N_29079);
or U29943 (N_29943,N_28910,N_29188);
nor U29944 (N_29944,N_29300,N_28886);
nand U29945 (N_29945,N_29135,N_29380);
nand U29946 (N_29946,N_28835,N_29167);
nand U29947 (N_29947,N_29161,N_29138);
nand U29948 (N_29948,N_29012,N_29385);
nor U29949 (N_29949,N_29356,N_29130);
or U29950 (N_29950,N_28982,N_29159);
nor U29951 (N_29951,N_29101,N_29041);
and U29952 (N_29952,N_28800,N_29186);
or U29953 (N_29953,N_28958,N_28870);
nand U29954 (N_29954,N_28987,N_29212);
and U29955 (N_29955,N_28886,N_29060);
nor U29956 (N_29956,N_29243,N_29204);
nand U29957 (N_29957,N_29305,N_29007);
nor U29958 (N_29958,N_29121,N_29125);
nor U29959 (N_29959,N_28849,N_28955);
xor U29960 (N_29960,N_29372,N_29063);
and U29961 (N_29961,N_29315,N_28984);
nand U29962 (N_29962,N_28951,N_29290);
nand U29963 (N_29963,N_29309,N_28960);
and U29964 (N_29964,N_29227,N_28923);
nor U29965 (N_29965,N_29318,N_28989);
nor U29966 (N_29966,N_29219,N_28825);
nand U29967 (N_29967,N_29147,N_29025);
xnor U29968 (N_29968,N_29158,N_29267);
or U29969 (N_29969,N_29272,N_28804);
and U29970 (N_29970,N_29125,N_29089);
nand U29971 (N_29971,N_28943,N_29089);
nand U29972 (N_29972,N_29031,N_29121);
or U29973 (N_29973,N_29172,N_29197);
and U29974 (N_29974,N_28821,N_29326);
and U29975 (N_29975,N_29284,N_29333);
and U29976 (N_29976,N_28823,N_29282);
and U29977 (N_29977,N_29131,N_28845);
nor U29978 (N_29978,N_29258,N_29382);
xnor U29979 (N_29979,N_28952,N_28939);
and U29980 (N_29980,N_29073,N_28820);
and U29981 (N_29981,N_29139,N_29171);
and U29982 (N_29982,N_28973,N_29365);
and U29983 (N_29983,N_29305,N_28914);
or U29984 (N_29984,N_28908,N_29195);
or U29985 (N_29985,N_28889,N_29264);
xnor U29986 (N_29986,N_29238,N_29355);
nor U29987 (N_29987,N_28935,N_29018);
and U29988 (N_29988,N_29232,N_29183);
nor U29989 (N_29989,N_29157,N_29014);
nand U29990 (N_29990,N_29127,N_29294);
xnor U29991 (N_29991,N_29340,N_29048);
or U29992 (N_29992,N_28882,N_29028);
xor U29993 (N_29993,N_28930,N_28838);
nand U29994 (N_29994,N_29381,N_29036);
and U29995 (N_29995,N_29140,N_28949);
or U29996 (N_29996,N_29305,N_28839);
and U29997 (N_29997,N_29328,N_29033);
xor U29998 (N_29998,N_28802,N_29007);
or U29999 (N_29999,N_29055,N_28874);
xnor UO_0 (O_0,N_29418,N_29803);
nand UO_1 (O_1,N_29914,N_29404);
and UO_2 (O_2,N_29848,N_29641);
and UO_3 (O_3,N_29956,N_29950);
and UO_4 (O_4,N_29713,N_29810);
and UO_5 (O_5,N_29596,N_29629);
xor UO_6 (O_6,N_29603,N_29465);
nand UO_7 (O_7,N_29422,N_29822);
or UO_8 (O_8,N_29577,N_29482);
and UO_9 (O_9,N_29421,N_29484);
xnor UO_10 (O_10,N_29543,N_29586);
and UO_11 (O_11,N_29698,N_29488);
xnor UO_12 (O_12,N_29636,N_29718);
and UO_13 (O_13,N_29682,N_29521);
nand UO_14 (O_14,N_29964,N_29783);
nand UO_15 (O_15,N_29533,N_29683);
and UO_16 (O_16,N_29691,N_29758);
xnor UO_17 (O_17,N_29562,N_29568);
nand UO_18 (O_18,N_29487,N_29694);
xnor UO_19 (O_19,N_29760,N_29880);
and UO_20 (O_20,N_29643,N_29445);
and UO_21 (O_21,N_29440,N_29670);
or UO_22 (O_22,N_29687,N_29967);
or UO_23 (O_23,N_29419,N_29846);
nand UO_24 (O_24,N_29744,N_29504);
or UO_25 (O_25,N_29785,N_29613);
nor UO_26 (O_26,N_29998,N_29917);
xnor UO_27 (O_27,N_29429,N_29566);
nor UO_28 (O_28,N_29497,N_29700);
or UO_29 (O_29,N_29711,N_29767);
and UO_30 (O_30,N_29721,N_29431);
or UO_31 (O_31,N_29551,N_29692);
or UO_32 (O_32,N_29823,N_29420);
nand UO_33 (O_33,N_29769,N_29768);
xnor UO_34 (O_34,N_29411,N_29836);
or UO_35 (O_35,N_29853,N_29689);
xnor UO_36 (O_36,N_29983,N_29978);
nand UO_37 (O_37,N_29786,N_29696);
nand UO_38 (O_38,N_29802,N_29776);
or UO_39 (O_39,N_29732,N_29885);
and UO_40 (O_40,N_29623,N_29847);
nand UO_41 (O_41,N_29915,N_29944);
nand UO_42 (O_42,N_29717,N_29437);
and UO_43 (O_43,N_29932,N_29993);
or UO_44 (O_44,N_29473,N_29526);
or UO_45 (O_45,N_29883,N_29478);
nor UO_46 (O_46,N_29812,N_29742);
and UO_47 (O_47,N_29708,N_29879);
nand UO_48 (O_48,N_29626,N_29483);
nor UO_49 (O_49,N_29984,N_29576);
and UO_50 (O_50,N_29875,N_29740);
nand UO_51 (O_51,N_29726,N_29624);
nand UO_52 (O_52,N_29664,N_29505);
or UO_53 (O_53,N_29756,N_29597);
xnor UO_54 (O_54,N_29741,N_29720);
nor UO_55 (O_55,N_29549,N_29731);
xor UO_56 (O_56,N_29674,N_29757);
or UO_57 (O_57,N_29637,N_29793);
nand UO_58 (O_58,N_29922,N_29938);
and UO_59 (O_59,N_29840,N_29554);
nor UO_60 (O_60,N_29842,N_29787);
nor UO_61 (O_61,N_29936,N_29555);
or UO_62 (O_62,N_29680,N_29456);
nor UO_63 (O_63,N_29621,N_29648);
and UO_64 (O_64,N_29738,N_29426);
and UO_65 (O_65,N_29489,N_29889);
and UO_66 (O_66,N_29759,N_29415);
nand UO_67 (O_67,N_29729,N_29963);
and UO_68 (O_68,N_29750,N_29662);
nand UO_69 (O_69,N_29408,N_29468);
nand UO_70 (O_70,N_29684,N_29477);
and UO_71 (O_71,N_29450,N_29941);
xor UO_72 (O_72,N_29806,N_29512);
nand UO_73 (O_73,N_29818,N_29471);
and UO_74 (O_74,N_29706,N_29977);
nor UO_75 (O_75,N_29658,N_29645);
or UO_76 (O_76,N_29704,N_29650);
nor UO_77 (O_77,N_29646,N_29898);
xor UO_78 (O_78,N_29816,N_29417);
or UO_79 (O_79,N_29778,N_29858);
and UO_80 (O_80,N_29985,N_29438);
and UO_81 (O_81,N_29605,N_29868);
nor UO_82 (O_82,N_29693,N_29739);
xor UO_83 (O_83,N_29509,N_29407);
or UO_84 (O_84,N_29588,N_29951);
xor UO_85 (O_85,N_29994,N_29954);
nor UO_86 (O_86,N_29957,N_29801);
and UO_87 (O_87,N_29814,N_29892);
xnor UO_88 (O_88,N_29463,N_29519);
or UO_89 (O_89,N_29556,N_29890);
or UO_90 (O_90,N_29530,N_29867);
xor UO_91 (O_91,N_29598,N_29775);
nand UO_92 (O_92,N_29929,N_29628);
xor UO_93 (O_93,N_29886,N_29714);
or UO_94 (O_94,N_29707,N_29686);
and UO_95 (O_95,N_29608,N_29607);
nand UO_96 (O_96,N_29668,N_29515);
or UO_97 (O_97,N_29773,N_29746);
nand UO_98 (O_98,N_29869,N_29534);
or UO_99 (O_99,N_29745,N_29548);
nor UO_100 (O_100,N_29499,N_29833);
xor UO_101 (O_101,N_29472,N_29953);
xnor UO_102 (O_102,N_29653,N_29884);
or UO_103 (O_103,N_29736,N_29486);
xnor UO_104 (O_104,N_29545,N_29552);
nor UO_105 (O_105,N_29513,N_29894);
nand UO_106 (O_106,N_29843,N_29563);
and UO_107 (O_107,N_29986,N_29857);
nand UO_108 (O_108,N_29452,N_29480);
or UO_109 (O_109,N_29930,N_29595);
nor UO_110 (O_110,N_29864,N_29719);
nand UO_111 (O_111,N_29651,N_29981);
nor UO_112 (O_112,N_29474,N_29454);
nand UO_113 (O_113,N_29874,N_29616);
and UO_114 (O_114,N_29856,N_29400);
xor UO_115 (O_115,N_29850,N_29677);
xnor UO_116 (O_116,N_29784,N_29667);
nor UO_117 (O_117,N_29798,N_29860);
and UO_118 (O_118,N_29462,N_29966);
or UO_119 (O_119,N_29699,N_29679);
xnor UO_120 (O_120,N_29432,N_29444);
and UO_121 (O_121,N_29439,N_29755);
nand UO_122 (O_122,N_29678,N_29730);
nand UO_123 (O_123,N_29428,N_29647);
nor UO_124 (O_124,N_29792,N_29446);
nor UO_125 (O_125,N_29579,N_29459);
or UO_126 (O_126,N_29457,N_29561);
xnor UO_127 (O_127,N_29939,N_29441);
and UO_128 (O_128,N_29476,N_29491);
and UO_129 (O_129,N_29433,N_29617);
or UO_130 (O_130,N_29600,N_29945);
or UO_131 (O_131,N_29522,N_29751);
xor UO_132 (O_132,N_29878,N_29615);
nor UO_133 (O_133,N_29413,N_29649);
and UO_134 (O_134,N_29982,N_29817);
xnor UO_135 (O_135,N_29839,N_29734);
and UO_136 (O_136,N_29702,N_29834);
xnor UO_137 (O_137,N_29451,N_29537);
or UO_138 (O_138,N_29992,N_29779);
nand UO_139 (O_139,N_29761,N_29927);
nand UO_140 (O_140,N_29791,N_29952);
or UO_141 (O_141,N_29747,N_29763);
nand UO_142 (O_142,N_29771,N_29573);
nand UO_143 (O_143,N_29508,N_29820);
and UO_144 (O_144,N_29788,N_29835);
nor UO_145 (O_145,N_29908,N_29520);
xnor UO_146 (O_146,N_29965,N_29620);
xnor UO_147 (O_147,N_29777,N_29976);
nand UO_148 (O_148,N_29479,N_29523);
xor UO_149 (O_149,N_29910,N_29673);
and UO_150 (O_150,N_29987,N_29961);
nor UO_151 (O_151,N_29581,N_29940);
and UO_152 (O_152,N_29642,N_29701);
or UO_153 (O_153,N_29709,N_29622);
xor UO_154 (O_154,N_29988,N_29435);
xor UO_155 (O_155,N_29436,N_29676);
nand UO_156 (O_156,N_29838,N_29547);
xnor UO_157 (O_157,N_29453,N_29602);
nand UO_158 (O_158,N_29580,N_29527);
nor UO_159 (O_159,N_29873,N_29830);
and UO_160 (O_160,N_29490,N_29989);
nand UO_161 (O_161,N_29690,N_29943);
xor UO_162 (O_162,N_29980,N_29837);
xor UO_163 (O_163,N_29583,N_29485);
nand UO_164 (O_164,N_29449,N_29780);
nor UO_165 (O_165,N_29852,N_29671);
nor UO_166 (O_166,N_29423,N_29410);
nand UO_167 (O_167,N_29971,N_29772);
nand UO_168 (O_168,N_29824,N_29665);
or UO_169 (O_169,N_29619,N_29614);
nor UO_170 (O_170,N_29593,N_29753);
and UO_171 (O_171,N_29639,N_29968);
and UO_172 (O_172,N_29946,N_29916);
nand UO_173 (O_173,N_29913,N_29789);
nor UO_174 (O_174,N_29909,N_29416);
and UO_175 (O_175,N_29825,N_29924);
and UO_176 (O_176,N_29669,N_29849);
or UO_177 (O_177,N_29974,N_29712);
nor UO_178 (O_178,N_29895,N_29805);
or UO_179 (O_179,N_29722,N_29795);
and UO_180 (O_180,N_29782,N_29409);
nor UO_181 (O_181,N_29401,N_29501);
nor UO_182 (O_182,N_29752,N_29900);
and UO_183 (O_183,N_29770,N_29705);
and UO_184 (O_184,N_29827,N_29995);
nor UO_185 (O_185,N_29506,N_29625);
and UO_186 (O_186,N_29854,N_29743);
xnor UO_187 (O_187,N_29790,N_29609);
and UO_188 (O_188,N_29675,N_29498);
nand UO_189 (O_189,N_29443,N_29990);
or UO_190 (O_190,N_29447,N_29905);
and UO_191 (O_191,N_29996,N_29507);
nand UO_192 (O_192,N_29610,N_29774);
and UO_193 (O_193,N_29503,N_29962);
nand UO_194 (O_194,N_29832,N_29887);
nor UO_195 (O_195,N_29861,N_29800);
nand UO_196 (O_196,N_29466,N_29592);
xnor UO_197 (O_197,N_29765,N_29872);
and UO_198 (O_198,N_29553,N_29564);
and UO_199 (O_199,N_29425,N_29975);
and UO_200 (O_200,N_29899,N_29542);
xnor UO_201 (O_201,N_29928,N_29796);
nand UO_202 (O_202,N_29599,N_29627);
xor UO_203 (O_203,N_29862,N_29538);
nand UO_204 (O_204,N_29403,N_29871);
xor UO_205 (O_205,N_29728,N_29589);
nand UO_206 (O_206,N_29469,N_29574);
and UO_207 (O_207,N_29402,N_29819);
nand UO_208 (O_208,N_29808,N_29826);
nand UO_209 (O_209,N_29582,N_29470);
xor UO_210 (O_210,N_29630,N_29933);
or UO_211 (O_211,N_29460,N_29781);
xor UO_212 (O_212,N_29524,N_29934);
or UO_213 (O_213,N_29494,N_29813);
and UO_214 (O_214,N_29727,N_29412);
nor UO_215 (O_215,N_29536,N_29518);
or UO_216 (O_216,N_29570,N_29749);
and UO_217 (O_217,N_29735,N_29937);
xnor UO_218 (O_218,N_29517,N_29902);
and UO_219 (O_219,N_29427,N_29635);
and UO_220 (O_220,N_29764,N_29859);
xnor UO_221 (O_221,N_29912,N_29666);
and UO_222 (O_222,N_29529,N_29558);
and UO_223 (O_223,N_29970,N_29888);
or UO_224 (O_224,N_29559,N_29882);
nor UO_225 (O_225,N_29661,N_29601);
or UO_226 (O_226,N_29541,N_29514);
or UO_227 (O_227,N_29973,N_29644);
and UO_228 (O_228,N_29502,N_29672);
xor UO_229 (O_229,N_29587,N_29811);
or UO_230 (O_230,N_29851,N_29931);
or UO_231 (O_231,N_29455,N_29475);
nor UO_232 (O_232,N_29815,N_29531);
and UO_233 (O_233,N_29560,N_29493);
xor UO_234 (O_234,N_29461,N_29863);
nand UO_235 (O_235,N_29578,N_29640);
xor UO_236 (O_236,N_29896,N_29500);
and UO_237 (O_237,N_29845,N_29585);
nor UO_238 (O_238,N_29958,N_29652);
and UO_239 (O_239,N_29540,N_29414);
nor UO_240 (O_240,N_29604,N_29997);
nand UO_241 (O_241,N_29688,N_29565);
nor UO_242 (O_242,N_29959,N_29999);
xnor UO_243 (O_243,N_29525,N_29663);
nand UO_244 (O_244,N_29893,N_29881);
xnor UO_245 (O_245,N_29804,N_29550);
nand UO_246 (O_246,N_29492,N_29901);
or UO_247 (O_247,N_29424,N_29631);
and UO_248 (O_248,N_29511,N_29703);
nand UO_249 (O_249,N_29737,N_29877);
and UO_250 (O_250,N_29430,N_29972);
or UO_251 (O_251,N_29481,N_29546);
nor UO_252 (O_252,N_29535,N_29891);
nand UO_253 (O_253,N_29733,N_29590);
xor UO_254 (O_254,N_29935,N_29904);
or UO_255 (O_255,N_29442,N_29496);
xnor UO_256 (O_256,N_29657,N_29841);
nor UO_257 (O_257,N_29544,N_29633);
xor UO_258 (O_258,N_29870,N_29611);
xor UO_259 (O_259,N_29528,N_29942);
xnor UO_260 (O_260,N_29710,N_29748);
or UO_261 (O_261,N_29448,N_29794);
nand UO_262 (O_262,N_29612,N_29809);
nand UO_263 (O_263,N_29495,N_29865);
and UO_264 (O_264,N_29571,N_29911);
or UO_265 (O_265,N_29539,N_29716);
and UO_266 (O_266,N_29949,N_29557);
xor UO_267 (O_267,N_29926,N_29697);
xor UO_268 (O_268,N_29960,N_29855);
nand UO_269 (O_269,N_29406,N_29632);
and UO_270 (O_270,N_29659,N_29569);
and UO_271 (O_271,N_29516,N_29762);
nor UO_272 (O_272,N_29458,N_29921);
nor UO_273 (O_273,N_29844,N_29828);
or UO_274 (O_274,N_29799,N_29923);
xor UO_275 (O_275,N_29634,N_29723);
xor UO_276 (O_276,N_29754,N_29695);
and UO_277 (O_277,N_29979,N_29715);
nand UO_278 (O_278,N_29681,N_29532);
xnor UO_279 (O_279,N_29991,N_29906);
or UO_280 (O_280,N_29925,N_29405);
nand UO_281 (O_281,N_29907,N_29903);
and UO_282 (O_282,N_29591,N_29866);
and UO_283 (O_283,N_29725,N_29969);
and UO_284 (O_284,N_29918,N_29685);
nand UO_285 (O_285,N_29920,N_29947);
xnor UO_286 (O_286,N_29955,N_29821);
nand UO_287 (O_287,N_29594,N_29897);
or UO_288 (O_288,N_29606,N_29948);
nand UO_289 (O_289,N_29797,N_29655);
and UO_290 (O_290,N_29572,N_29575);
and UO_291 (O_291,N_29766,N_29567);
nor UO_292 (O_292,N_29876,N_29831);
xnor UO_293 (O_293,N_29584,N_29638);
or UO_294 (O_294,N_29618,N_29654);
or UO_295 (O_295,N_29919,N_29510);
xor UO_296 (O_296,N_29434,N_29807);
nand UO_297 (O_297,N_29656,N_29464);
nor UO_298 (O_298,N_29724,N_29467);
nand UO_299 (O_299,N_29660,N_29829);
xnor UO_300 (O_300,N_29659,N_29670);
or UO_301 (O_301,N_29864,N_29612);
xor UO_302 (O_302,N_29564,N_29457);
nand UO_303 (O_303,N_29707,N_29984);
xnor UO_304 (O_304,N_29720,N_29681);
and UO_305 (O_305,N_29590,N_29504);
nand UO_306 (O_306,N_29658,N_29656);
xnor UO_307 (O_307,N_29674,N_29640);
and UO_308 (O_308,N_29498,N_29924);
or UO_309 (O_309,N_29414,N_29411);
and UO_310 (O_310,N_29914,N_29988);
nor UO_311 (O_311,N_29508,N_29813);
xnor UO_312 (O_312,N_29728,N_29534);
or UO_313 (O_313,N_29429,N_29798);
xnor UO_314 (O_314,N_29935,N_29758);
and UO_315 (O_315,N_29922,N_29691);
nor UO_316 (O_316,N_29632,N_29967);
nor UO_317 (O_317,N_29406,N_29971);
or UO_318 (O_318,N_29829,N_29573);
nor UO_319 (O_319,N_29980,N_29732);
nand UO_320 (O_320,N_29764,N_29822);
xor UO_321 (O_321,N_29931,N_29412);
and UO_322 (O_322,N_29474,N_29849);
nor UO_323 (O_323,N_29839,N_29708);
and UO_324 (O_324,N_29977,N_29575);
xnor UO_325 (O_325,N_29551,N_29962);
or UO_326 (O_326,N_29848,N_29688);
nand UO_327 (O_327,N_29797,N_29709);
nand UO_328 (O_328,N_29806,N_29624);
nor UO_329 (O_329,N_29788,N_29930);
nand UO_330 (O_330,N_29519,N_29810);
and UO_331 (O_331,N_29993,N_29726);
nand UO_332 (O_332,N_29573,N_29538);
nor UO_333 (O_333,N_29800,N_29497);
xor UO_334 (O_334,N_29981,N_29805);
or UO_335 (O_335,N_29810,N_29993);
nand UO_336 (O_336,N_29969,N_29483);
xor UO_337 (O_337,N_29625,N_29698);
xor UO_338 (O_338,N_29739,N_29980);
or UO_339 (O_339,N_29764,N_29865);
or UO_340 (O_340,N_29714,N_29951);
or UO_341 (O_341,N_29760,N_29976);
or UO_342 (O_342,N_29608,N_29428);
nand UO_343 (O_343,N_29486,N_29617);
nand UO_344 (O_344,N_29664,N_29774);
or UO_345 (O_345,N_29823,N_29809);
nor UO_346 (O_346,N_29726,N_29563);
nand UO_347 (O_347,N_29701,N_29937);
xnor UO_348 (O_348,N_29864,N_29433);
or UO_349 (O_349,N_29727,N_29969);
xor UO_350 (O_350,N_29921,N_29880);
xor UO_351 (O_351,N_29741,N_29494);
or UO_352 (O_352,N_29625,N_29462);
xnor UO_353 (O_353,N_29861,N_29529);
nor UO_354 (O_354,N_29473,N_29795);
or UO_355 (O_355,N_29869,N_29922);
or UO_356 (O_356,N_29648,N_29701);
nor UO_357 (O_357,N_29757,N_29625);
xnor UO_358 (O_358,N_29617,N_29764);
or UO_359 (O_359,N_29844,N_29489);
nand UO_360 (O_360,N_29868,N_29405);
xor UO_361 (O_361,N_29521,N_29846);
nor UO_362 (O_362,N_29989,N_29700);
nand UO_363 (O_363,N_29901,N_29955);
nor UO_364 (O_364,N_29725,N_29709);
nand UO_365 (O_365,N_29493,N_29834);
xnor UO_366 (O_366,N_29771,N_29463);
and UO_367 (O_367,N_29434,N_29671);
nor UO_368 (O_368,N_29550,N_29497);
or UO_369 (O_369,N_29977,N_29774);
nand UO_370 (O_370,N_29929,N_29851);
nor UO_371 (O_371,N_29553,N_29725);
nor UO_372 (O_372,N_29956,N_29640);
xnor UO_373 (O_373,N_29809,N_29745);
nand UO_374 (O_374,N_29930,N_29862);
xor UO_375 (O_375,N_29812,N_29660);
and UO_376 (O_376,N_29718,N_29835);
nand UO_377 (O_377,N_29595,N_29618);
or UO_378 (O_378,N_29493,N_29454);
nand UO_379 (O_379,N_29941,N_29510);
nor UO_380 (O_380,N_29703,N_29705);
and UO_381 (O_381,N_29571,N_29775);
nand UO_382 (O_382,N_29965,N_29724);
or UO_383 (O_383,N_29982,N_29862);
and UO_384 (O_384,N_29680,N_29902);
xnor UO_385 (O_385,N_29845,N_29536);
nor UO_386 (O_386,N_29507,N_29984);
xnor UO_387 (O_387,N_29964,N_29989);
or UO_388 (O_388,N_29764,N_29867);
nor UO_389 (O_389,N_29921,N_29581);
nor UO_390 (O_390,N_29812,N_29409);
nor UO_391 (O_391,N_29821,N_29692);
xor UO_392 (O_392,N_29706,N_29884);
and UO_393 (O_393,N_29734,N_29837);
nor UO_394 (O_394,N_29899,N_29681);
and UO_395 (O_395,N_29644,N_29995);
xnor UO_396 (O_396,N_29513,N_29989);
xor UO_397 (O_397,N_29810,N_29736);
xnor UO_398 (O_398,N_29494,N_29730);
xor UO_399 (O_399,N_29936,N_29583);
or UO_400 (O_400,N_29997,N_29660);
xnor UO_401 (O_401,N_29981,N_29707);
and UO_402 (O_402,N_29529,N_29591);
nand UO_403 (O_403,N_29465,N_29900);
nor UO_404 (O_404,N_29612,N_29710);
nand UO_405 (O_405,N_29671,N_29773);
nand UO_406 (O_406,N_29443,N_29493);
or UO_407 (O_407,N_29972,N_29734);
xnor UO_408 (O_408,N_29421,N_29548);
or UO_409 (O_409,N_29431,N_29656);
xnor UO_410 (O_410,N_29929,N_29777);
nand UO_411 (O_411,N_29758,N_29623);
nand UO_412 (O_412,N_29663,N_29880);
or UO_413 (O_413,N_29549,N_29473);
nand UO_414 (O_414,N_29934,N_29881);
and UO_415 (O_415,N_29865,N_29807);
and UO_416 (O_416,N_29618,N_29740);
nor UO_417 (O_417,N_29417,N_29488);
xor UO_418 (O_418,N_29463,N_29682);
or UO_419 (O_419,N_29694,N_29554);
nand UO_420 (O_420,N_29552,N_29553);
nand UO_421 (O_421,N_29967,N_29507);
or UO_422 (O_422,N_29877,N_29427);
and UO_423 (O_423,N_29562,N_29942);
nor UO_424 (O_424,N_29485,N_29729);
and UO_425 (O_425,N_29458,N_29766);
nor UO_426 (O_426,N_29783,N_29595);
or UO_427 (O_427,N_29985,N_29601);
nor UO_428 (O_428,N_29447,N_29550);
and UO_429 (O_429,N_29964,N_29548);
and UO_430 (O_430,N_29596,N_29702);
nand UO_431 (O_431,N_29414,N_29536);
nand UO_432 (O_432,N_29863,N_29802);
nand UO_433 (O_433,N_29627,N_29899);
and UO_434 (O_434,N_29503,N_29739);
nand UO_435 (O_435,N_29944,N_29523);
nand UO_436 (O_436,N_29598,N_29876);
or UO_437 (O_437,N_29978,N_29546);
xor UO_438 (O_438,N_29985,N_29953);
nand UO_439 (O_439,N_29457,N_29623);
xor UO_440 (O_440,N_29786,N_29928);
nor UO_441 (O_441,N_29531,N_29575);
xor UO_442 (O_442,N_29458,N_29676);
or UO_443 (O_443,N_29527,N_29455);
xor UO_444 (O_444,N_29932,N_29981);
nor UO_445 (O_445,N_29899,N_29631);
or UO_446 (O_446,N_29681,N_29993);
nand UO_447 (O_447,N_29745,N_29931);
xnor UO_448 (O_448,N_29521,N_29796);
nor UO_449 (O_449,N_29870,N_29624);
or UO_450 (O_450,N_29521,N_29947);
or UO_451 (O_451,N_29738,N_29513);
and UO_452 (O_452,N_29642,N_29908);
or UO_453 (O_453,N_29560,N_29767);
or UO_454 (O_454,N_29737,N_29590);
or UO_455 (O_455,N_29774,N_29952);
or UO_456 (O_456,N_29969,N_29518);
or UO_457 (O_457,N_29931,N_29743);
or UO_458 (O_458,N_29908,N_29545);
or UO_459 (O_459,N_29812,N_29907);
or UO_460 (O_460,N_29695,N_29820);
or UO_461 (O_461,N_29692,N_29970);
xor UO_462 (O_462,N_29587,N_29719);
xnor UO_463 (O_463,N_29525,N_29480);
nand UO_464 (O_464,N_29626,N_29607);
xnor UO_465 (O_465,N_29788,N_29637);
or UO_466 (O_466,N_29403,N_29921);
or UO_467 (O_467,N_29430,N_29991);
or UO_468 (O_468,N_29490,N_29521);
and UO_469 (O_469,N_29415,N_29869);
nand UO_470 (O_470,N_29402,N_29513);
nor UO_471 (O_471,N_29715,N_29977);
xnor UO_472 (O_472,N_29950,N_29878);
nor UO_473 (O_473,N_29851,N_29705);
xor UO_474 (O_474,N_29677,N_29548);
or UO_475 (O_475,N_29439,N_29719);
nand UO_476 (O_476,N_29644,N_29741);
or UO_477 (O_477,N_29637,N_29827);
or UO_478 (O_478,N_29714,N_29510);
and UO_479 (O_479,N_29521,N_29750);
nand UO_480 (O_480,N_29822,N_29734);
or UO_481 (O_481,N_29824,N_29980);
nand UO_482 (O_482,N_29583,N_29860);
or UO_483 (O_483,N_29456,N_29889);
nand UO_484 (O_484,N_29404,N_29463);
nand UO_485 (O_485,N_29796,N_29829);
nor UO_486 (O_486,N_29685,N_29526);
and UO_487 (O_487,N_29763,N_29500);
or UO_488 (O_488,N_29482,N_29506);
nand UO_489 (O_489,N_29697,N_29786);
xnor UO_490 (O_490,N_29512,N_29604);
xnor UO_491 (O_491,N_29839,N_29725);
or UO_492 (O_492,N_29727,N_29829);
and UO_493 (O_493,N_29975,N_29754);
xor UO_494 (O_494,N_29948,N_29805);
or UO_495 (O_495,N_29642,N_29470);
nand UO_496 (O_496,N_29862,N_29458);
or UO_497 (O_497,N_29957,N_29640);
nand UO_498 (O_498,N_29725,N_29454);
xnor UO_499 (O_499,N_29980,N_29469);
and UO_500 (O_500,N_29503,N_29702);
and UO_501 (O_501,N_29915,N_29802);
xnor UO_502 (O_502,N_29431,N_29760);
nor UO_503 (O_503,N_29630,N_29842);
nand UO_504 (O_504,N_29880,N_29901);
and UO_505 (O_505,N_29889,N_29515);
or UO_506 (O_506,N_29661,N_29783);
xor UO_507 (O_507,N_29920,N_29956);
or UO_508 (O_508,N_29750,N_29536);
or UO_509 (O_509,N_29477,N_29529);
and UO_510 (O_510,N_29470,N_29602);
nand UO_511 (O_511,N_29780,N_29616);
and UO_512 (O_512,N_29405,N_29793);
xnor UO_513 (O_513,N_29618,N_29919);
xor UO_514 (O_514,N_29651,N_29832);
or UO_515 (O_515,N_29729,N_29922);
and UO_516 (O_516,N_29995,N_29922);
nand UO_517 (O_517,N_29891,N_29757);
or UO_518 (O_518,N_29529,N_29626);
xor UO_519 (O_519,N_29427,N_29957);
xnor UO_520 (O_520,N_29779,N_29669);
xor UO_521 (O_521,N_29432,N_29694);
nand UO_522 (O_522,N_29949,N_29728);
nor UO_523 (O_523,N_29576,N_29961);
or UO_524 (O_524,N_29691,N_29532);
nand UO_525 (O_525,N_29536,N_29723);
nand UO_526 (O_526,N_29615,N_29770);
nor UO_527 (O_527,N_29935,N_29676);
xnor UO_528 (O_528,N_29727,N_29404);
or UO_529 (O_529,N_29513,N_29996);
and UO_530 (O_530,N_29552,N_29767);
or UO_531 (O_531,N_29695,N_29825);
and UO_532 (O_532,N_29512,N_29969);
xnor UO_533 (O_533,N_29747,N_29762);
xnor UO_534 (O_534,N_29639,N_29641);
or UO_535 (O_535,N_29670,N_29560);
xnor UO_536 (O_536,N_29564,N_29972);
xor UO_537 (O_537,N_29530,N_29850);
and UO_538 (O_538,N_29462,N_29596);
nand UO_539 (O_539,N_29904,N_29424);
and UO_540 (O_540,N_29460,N_29576);
and UO_541 (O_541,N_29716,N_29407);
or UO_542 (O_542,N_29619,N_29973);
nand UO_543 (O_543,N_29520,N_29401);
xnor UO_544 (O_544,N_29526,N_29641);
nor UO_545 (O_545,N_29977,N_29796);
nor UO_546 (O_546,N_29539,N_29508);
and UO_547 (O_547,N_29726,N_29845);
xnor UO_548 (O_548,N_29913,N_29756);
xor UO_549 (O_549,N_29841,N_29442);
nand UO_550 (O_550,N_29552,N_29713);
xnor UO_551 (O_551,N_29668,N_29698);
or UO_552 (O_552,N_29848,N_29710);
and UO_553 (O_553,N_29428,N_29636);
nor UO_554 (O_554,N_29666,N_29623);
or UO_555 (O_555,N_29710,N_29838);
and UO_556 (O_556,N_29525,N_29572);
and UO_557 (O_557,N_29812,N_29807);
nor UO_558 (O_558,N_29866,N_29409);
or UO_559 (O_559,N_29961,N_29728);
xor UO_560 (O_560,N_29885,N_29595);
xor UO_561 (O_561,N_29469,N_29544);
or UO_562 (O_562,N_29400,N_29653);
nor UO_563 (O_563,N_29604,N_29930);
nand UO_564 (O_564,N_29433,N_29600);
xnor UO_565 (O_565,N_29798,N_29864);
nor UO_566 (O_566,N_29757,N_29729);
or UO_567 (O_567,N_29683,N_29404);
nand UO_568 (O_568,N_29633,N_29840);
and UO_569 (O_569,N_29776,N_29525);
xor UO_570 (O_570,N_29749,N_29943);
or UO_571 (O_571,N_29595,N_29757);
or UO_572 (O_572,N_29806,N_29728);
nand UO_573 (O_573,N_29518,N_29443);
or UO_574 (O_574,N_29724,N_29877);
xnor UO_575 (O_575,N_29597,N_29760);
xnor UO_576 (O_576,N_29567,N_29620);
and UO_577 (O_577,N_29513,N_29951);
xnor UO_578 (O_578,N_29736,N_29456);
nand UO_579 (O_579,N_29731,N_29625);
or UO_580 (O_580,N_29867,N_29487);
nand UO_581 (O_581,N_29952,N_29794);
and UO_582 (O_582,N_29842,N_29458);
nor UO_583 (O_583,N_29681,N_29844);
or UO_584 (O_584,N_29938,N_29567);
nor UO_585 (O_585,N_29812,N_29473);
nor UO_586 (O_586,N_29913,N_29855);
nor UO_587 (O_587,N_29833,N_29737);
nand UO_588 (O_588,N_29692,N_29746);
nor UO_589 (O_589,N_29545,N_29820);
xor UO_590 (O_590,N_29763,N_29728);
nor UO_591 (O_591,N_29779,N_29847);
and UO_592 (O_592,N_29539,N_29575);
and UO_593 (O_593,N_29969,N_29820);
nor UO_594 (O_594,N_29571,N_29617);
nand UO_595 (O_595,N_29904,N_29776);
and UO_596 (O_596,N_29480,N_29703);
nor UO_597 (O_597,N_29860,N_29760);
and UO_598 (O_598,N_29564,N_29443);
or UO_599 (O_599,N_29973,N_29549);
or UO_600 (O_600,N_29950,N_29929);
and UO_601 (O_601,N_29906,N_29934);
nand UO_602 (O_602,N_29711,N_29564);
nand UO_603 (O_603,N_29607,N_29699);
or UO_604 (O_604,N_29876,N_29666);
xor UO_605 (O_605,N_29527,N_29784);
xnor UO_606 (O_606,N_29412,N_29780);
xor UO_607 (O_607,N_29773,N_29649);
and UO_608 (O_608,N_29478,N_29945);
or UO_609 (O_609,N_29482,N_29887);
or UO_610 (O_610,N_29840,N_29600);
or UO_611 (O_611,N_29548,N_29524);
xnor UO_612 (O_612,N_29574,N_29526);
nand UO_613 (O_613,N_29597,N_29959);
or UO_614 (O_614,N_29995,N_29765);
xor UO_615 (O_615,N_29460,N_29699);
xnor UO_616 (O_616,N_29797,N_29913);
and UO_617 (O_617,N_29974,N_29598);
or UO_618 (O_618,N_29744,N_29635);
nand UO_619 (O_619,N_29782,N_29959);
and UO_620 (O_620,N_29502,N_29791);
xor UO_621 (O_621,N_29997,N_29814);
or UO_622 (O_622,N_29438,N_29973);
nand UO_623 (O_623,N_29703,N_29536);
or UO_624 (O_624,N_29706,N_29961);
xnor UO_625 (O_625,N_29833,N_29482);
nor UO_626 (O_626,N_29539,N_29519);
or UO_627 (O_627,N_29435,N_29823);
and UO_628 (O_628,N_29804,N_29486);
xnor UO_629 (O_629,N_29737,N_29957);
xnor UO_630 (O_630,N_29526,N_29451);
and UO_631 (O_631,N_29493,N_29781);
nor UO_632 (O_632,N_29524,N_29586);
nand UO_633 (O_633,N_29514,N_29922);
xor UO_634 (O_634,N_29513,N_29589);
and UO_635 (O_635,N_29686,N_29886);
and UO_636 (O_636,N_29987,N_29504);
xor UO_637 (O_637,N_29648,N_29603);
xor UO_638 (O_638,N_29848,N_29624);
nor UO_639 (O_639,N_29840,N_29863);
and UO_640 (O_640,N_29455,N_29864);
nor UO_641 (O_641,N_29614,N_29988);
and UO_642 (O_642,N_29724,N_29994);
and UO_643 (O_643,N_29556,N_29855);
xnor UO_644 (O_644,N_29574,N_29583);
xnor UO_645 (O_645,N_29537,N_29715);
nor UO_646 (O_646,N_29999,N_29952);
nand UO_647 (O_647,N_29726,N_29461);
nor UO_648 (O_648,N_29400,N_29444);
nand UO_649 (O_649,N_29909,N_29796);
nand UO_650 (O_650,N_29929,N_29925);
nand UO_651 (O_651,N_29656,N_29830);
nor UO_652 (O_652,N_29607,N_29417);
and UO_653 (O_653,N_29740,N_29835);
xnor UO_654 (O_654,N_29896,N_29736);
nor UO_655 (O_655,N_29605,N_29793);
or UO_656 (O_656,N_29871,N_29822);
nand UO_657 (O_657,N_29558,N_29942);
xor UO_658 (O_658,N_29483,N_29632);
xnor UO_659 (O_659,N_29760,N_29444);
xnor UO_660 (O_660,N_29560,N_29648);
nor UO_661 (O_661,N_29539,N_29442);
nand UO_662 (O_662,N_29434,N_29633);
nor UO_663 (O_663,N_29621,N_29433);
or UO_664 (O_664,N_29874,N_29947);
nand UO_665 (O_665,N_29624,N_29925);
and UO_666 (O_666,N_29988,N_29742);
xnor UO_667 (O_667,N_29742,N_29740);
or UO_668 (O_668,N_29648,N_29993);
nor UO_669 (O_669,N_29855,N_29753);
nor UO_670 (O_670,N_29626,N_29959);
or UO_671 (O_671,N_29679,N_29455);
and UO_672 (O_672,N_29629,N_29420);
nand UO_673 (O_673,N_29618,N_29836);
or UO_674 (O_674,N_29926,N_29998);
nand UO_675 (O_675,N_29765,N_29517);
xnor UO_676 (O_676,N_29747,N_29897);
or UO_677 (O_677,N_29916,N_29721);
or UO_678 (O_678,N_29417,N_29504);
nor UO_679 (O_679,N_29403,N_29554);
and UO_680 (O_680,N_29836,N_29950);
or UO_681 (O_681,N_29580,N_29845);
or UO_682 (O_682,N_29543,N_29815);
nor UO_683 (O_683,N_29442,N_29678);
xor UO_684 (O_684,N_29437,N_29695);
xor UO_685 (O_685,N_29667,N_29578);
or UO_686 (O_686,N_29879,N_29965);
nor UO_687 (O_687,N_29840,N_29620);
nand UO_688 (O_688,N_29977,N_29570);
nand UO_689 (O_689,N_29406,N_29458);
xor UO_690 (O_690,N_29927,N_29870);
or UO_691 (O_691,N_29417,N_29847);
and UO_692 (O_692,N_29984,N_29699);
and UO_693 (O_693,N_29439,N_29722);
xnor UO_694 (O_694,N_29568,N_29993);
xnor UO_695 (O_695,N_29798,N_29650);
nand UO_696 (O_696,N_29974,N_29744);
nor UO_697 (O_697,N_29658,N_29663);
and UO_698 (O_698,N_29812,N_29628);
xnor UO_699 (O_699,N_29814,N_29659);
or UO_700 (O_700,N_29951,N_29577);
nand UO_701 (O_701,N_29540,N_29519);
nor UO_702 (O_702,N_29735,N_29923);
or UO_703 (O_703,N_29608,N_29551);
nor UO_704 (O_704,N_29565,N_29902);
and UO_705 (O_705,N_29580,N_29883);
xnor UO_706 (O_706,N_29870,N_29859);
nand UO_707 (O_707,N_29468,N_29579);
xor UO_708 (O_708,N_29570,N_29696);
or UO_709 (O_709,N_29586,N_29721);
xor UO_710 (O_710,N_29841,N_29423);
xnor UO_711 (O_711,N_29955,N_29683);
and UO_712 (O_712,N_29608,N_29981);
xor UO_713 (O_713,N_29663,N_29967);
nand UO_714 (O_714,N_29494,N_29905);
xor UO_715 (O_715,N_29572,N_29507);
nor UO_716 (O_716,N_29971,N_29662);
or UO_717 (O_717,N_29759,N_29779);
and UO_718 (O_718,N_29424,N_29491);
and UO_719 (O_719,N_29730,N_29465);
xnor UO_720 (O_720,N_29740,N_29854);
and UO_721 (O_721,N_29540,N_29927);
xnor UO_722 (O_722,N_29937,N_29844);
and UO_723 (O_723,N_29607,N_29454);
nor UO_724 (O_724,N_29493,N_29815);
nand UO_725 (O_725,N_29995,N_29837);
nor UO_726 (O_726,N_29758,N_29835);
or UO_727 (O_727,N_29736,N_29619);
nor UO_728 (O_728,N_29779,N_29437);
xor UO_729 (O_729,N_29418,N_29922);
nor UO_730 (O_730,N_29523,N_29619);
and UO_731 (O_731,N_29756,N_29834);
nor UO_732 (O_732,N_29862,N_29837);
and UO_733 (O_733,N_29424,N_29487);
xor UO_734 (O_734,N_29722,N_29827);
nor UO_735 (O_735,N_29438,N_29488);
nor UO_736 (O_736,N_29450,N_29560);
and UO_737 (O_737,N_29992,N_29463);
and UO_738 (O_738,N_29462,N_29642);
nand UO_739 (O_739,N_29567,N_29690);
and UO_740 (O_740,N_29982,N_29443);
and UO_741 (O_741,N_29980,N_29468);
or UO_742 (O_742,N_29433,N_29927);
nand UO_743 (O_743,N_29405,N_29548);
nor UO_744 (O_744,N_29883,N_29494);
and UO_745 (O_745,N_29699,N_29574);
xor UO_746 (O_746,N_29427,N_29521);
and UO_747 (O_747,N_29642,N_29958);
and UO_748 (O_748,N_29971,N_29427);
or UO_749 (O_749,N_29846,N_29737);
xnor UO_750 (O_750,N_29454,N_29827);
nand UO_751 (O_751,N_29733,N_29936);
or UO_752 (O_752,N_29559,N_29500);
xnor UO_753 (O_753,N_29708,N_29540);
and UO_754 (O_754,N_29886,N_29606);
nand UO_755 (O_755,N_29480,N_29751);
xnor UO_756 (O_756,N_29575,N_29821);
or UO_757 (O_757,N_29661,N_29714);
or UO_758 (O_758,N_29913,N_29818);
or UO_759 (O_759,N_29933,N_29878);
nand UO_760 (O_760,N_29880,N_29762);
and UO_761 (O_761,N_29444,N_29479);
or UO_762 (O_762,N_29840,N_29672);
and UO_763 (O_763,N_29915,N_29951);
xor UO_764 (O_764,N_29442,N_29703);
or UO_765 (O_765,N_29736,N_29936);
nor UO_766 (O_766,N_29962,N_29766);
and UO_767 (O_767,N_29712,N_29708);
nor UO_768 (O_768,N_29416,N_29897);
nor UO_769 (O_769,N_29423,N_29906);
or UO_770 (O_770,N_29501,N_29690);
and UO_771 (O_771,N_29434,N_29468);
nor UO_772 (O_772,N_29997,N_29536);
or UO_773 (O_773,N_29651,N_29810);
nor UO_774 (O_774,N_29442,N_29468);
nand UO_775 (O_775,N_29924,N_29575);
nand UO_776 (O_776,N_29933,N_29702);
nand UO_777 (O_777,N_29556,N_29455);
xor UO_778 (O_778,N_29738,N_29485);
nor UO_779 (O_779,N_29456,N_29686);
and UO_780 (O_780,N_29813,N_29886);
nor UO_781 (O_781,N_29833,N_29757);
nand UO_782 (O_782,N_29591,N_29887);
nand UO_783 (O_783,N_29936,N_29865);
or UO_784 (O_784,N_29729,N_29904);
and UO_785 (O_785,N_29495,N_29815);
and UO_786 (O_786,N_29982,N_29634);
and UO_787 (O_787,N_29425,N_29956);
xor UO_788 (O_788,N_29815,N_29501);
xor UO_789 (O_789,N_29627,N_29788);
or UO_790 (O_790,N_29996,N_29405);
or UO_791 (O_791,N_29877,N_29483);
nand UO_792 (O_792,N_29957,N_29700);
nand UO_793 (O_793,N_29958,N_29874);
or UO_794 (O_794,N_29555,N_29443);
or UO_795 (O_795,N_29723,N_29454);
xor UO_796 (O_796,N_29698,N_29528);
nor UO_797 (O_797,N_29446,N_29541);
or UO_798 (O_798,N_29546,N_29638);
xnor UO_799 (O_799,N_29634,N_29623);
xnor UO_800 (O_800,N_29460,N_29484);
nand UO_801 (O_801,N_29911,N_29802);
nor UO_802 (O_802,N_29519,N_29816);
nand UO_803 (O_803,N_29448,N_29817);
or UO_804 (O_804,N_29647,N_29549);
nor UO_805 (O_805,N_29462,N_29913);
nand UO_806 (O_806,N_29770,N_29742);
nand UO_807 (O_807,N_29672,N_29433);
or UO_808 (O_808,N_29510,N_29452);
xor UO_809 (O_809,N_29522,N_29428);
and UO_810 (O_810,N_29861,N_29702);
or UO_811 (O_811,N_29671,N_29618);
or UO_812 (O_812,N_29873,N_29609);
and UO_813 (O_813,N_29745,N_29471);
nand UO_814 (O_814,N_29775,N_29549);
xnor UO_815 (O_815,N_29496,N_29574);
or UO_816 (O_816,N_29617,N_29933);
or UO_817 (O_817,N_29772,N_29927);
and UO_818 (O_818,N_29988,N_29590);
and UO_819 (O_819,N_29454,N_29844);
nor UO_820 (O_820,N_29744,N_29540);
xnor UO_821 (O_821,N_29457,N_29802);
and UO_822 (O_822,N_29486,N_29862);
xnor UO_823 (O_823,N_29878,N_29785);
nor UO_824 (O_824,N_29826,N_29973);
xnor UO_825 (O_825,N_29624,N_29798);
and UO_826 (O_826,N_29601,N_29725);
nand UO_827 (O_827,N_29906,N_29584);
nand UO_828 (O_828,N_29766,N_29673);
nor UO_829 (O_829,N_29949,N_29438);
nor UO_830 (O_830,N_29941,N_29405);
or UO_831 (O_831,N_29576,N_29432);
nand UO_832 (O_832,N_29494,N_29824);
nand UO_833 (O_833,N_29519,N_29733);
nand UO_834 (O_834,N_29912,N_29423);
nor UO_835 (O_835,N_29524,N_29563);
nor UO_836 (O_836,N_29796,N_29596);
nor UO_837 (O_837,N_29664,N_29963);
xnor UO_838 (O_838,N_29947,N_29626);
nand UO_839 (O_839,N_29533,N_29715);
nor UO_840 (O_840,N_29800,N_29773);
xor UO_841 (O_841,N_29464,N_29984);
or UO_842 (O_842,N_29541,N_29402);
or UO_843 (O_843,N_29879,N_29992);
xnor UO_844 (O_844,N_29649,N_29740);
and UO_845 (O_845,N_29891,N_29444);
and UO_846 (O_846,N_29575,N_29868);
or UO_847 (O_847,N_29467,N_29703);
nand UO_848 (O_848,N_29563,N_29819);
xnor UO_849 (O_849,N_29484,N_29406);
nand UO_850 (O_850,N_29477,N_29681);
and UO_851 (O_851,N_29592,N_29418);
nand UO_852 (O_852,N_29667,N_29661);
and UO_853 (O_853,N_29791,N_29441);
nor UO_854 (O_854,N_29415,N_29638);
nand UO_855 (O_855,N_29986,N_29401);
xnor UO_856 (O_856,N_29992,N_29769);
or UO_857 (O_857,N_29995,N_29735);
xnor UO_858 (O_858,N_29998,N_29761);
or UO_859 (O_859,N_29963,N_29894);
and UO_860 (O_860,N_29896,N_29715);
or UO_861 (O_861,N_29758,N_29946);
nor UO_862 (O_862,N_29757,N_29402);
nor UO_863 (O_863,N_29794,N_29677);
and UO_864 (O_864,N_29639,N_29772);
xor UO_865 (O_865,N_29694,N_29677);
nor UO_866 (O_866,N_29995,N_29676);
and UO_867 (O_867,N_29680,N_29849);
or UO_868 (O_868,N_29999,N_29637);
and UO_869 (O_869,N_29788,N_29572);
xnor UO_870 (O_870,N_29719,N_29804);
and UO_871 (O_871,N_29844,N_29973);
nand UO_872 (O_872,N_29777,N_29819);
nor UO_873 (O_873,N_29856,N_29911);
nand UO_874 (O_874,N_29600,N_29961);
xor UO_875 (O_875,N_29642,N_29843);
or UO_876 (O_876,N_29533,N_29703);
nor UO_877 (O_877,N_29827,N_29892);
nor UO_878 (O_878,N_29842,N_29965);
nor UO_879 (O_879,N_29680,N_29833);
nand UO_880 (O_880,N_29709,N_29488);
nand UO_881 (O_881,N_29824,N_29591);
and UO_882 (O_882,N_29845,N_29840);
and UO_883 (O_883,N_29452,N_29772);
xnor UO_884 (O_884,N_29917,N_29619);
or UO_885 (O_885,N_29923,N_29685);
xor UO_886 (O_886,N_29506,N_29961);
or UO_887 (O_887,N_29925,N_29489);
and UO_888 (O_888,N_29919,N_29595);
or UO_889 (O_889,N_29432,N_29459);
nand UO_890 (O_890,N_29937,N_29917);
nand UO_891 (O_891,N_29585,N_29943);
nand UO_892 (O_892,N_29842,N_29427);
and UO_893 (O_893,N_29650,N_29898);
and UO_894 (O_894,N_29949,N_29872);
xor UO_895 (O_895,N_29632,N_29589);
nand UO_896 (O_896,N_29826,N_29497);
or UO_897 (O_897,N_29965,N_29583);
xnor UO_898 (O_898,N_29811,N_29857);
or UO_899 (O_899,N_29531,N_29600);
nor UO_900 (O_900,N_29552,N_29524);
xnor UO_901 (O_901,N_29931,N_29987);
and UO_902 (O_902,N_29416,N_29479);
nor UO_903 (O_903,N_29462,N_29417);
xnor UO_904 (O_904,N_29752,N_29858);
and UO_905 (O_905,N_29919,N_29945);
or UO_906 (O_906,N_29516,N_29562);
nor UO_907 (O_907,N_29905,N_29844);
and UO_908 (O_908,N_29561,N_29943);
or UO_909 (O_909,N_29423,N_29649);
nand UO_910 (O_910,N_29893,N_29599);
nand UO_911 (O_911,N_29473,N_29710);
xor UO_912 (O_912,N_29906,N_29548);
xnor UO_913 (O_913,N_29655,N_29605);
nor UO_914 (O_914,N_29638,N_29431);
nand UO_915 (O_915,N_29624,N_29830);
xnor UO_916 (O_916,N_29898,N_29419);
nor UO_917 (O_917,N_29724,N_29460);
and UO_918 (O_918,N_29472,N_29687);
or UO_919 (O_919,N_29689,N_29649);
nand UO_920 (O_920,N_29823,N_29661);
and UO_921 (O_921,N_29957,N_29678);
nor UO_922 (O_922,N_29670,N_29488);
or UO_923 (O_923,N_29957,N_29635);
nor UO_924 (O_924,N_29602,N_29462);
or UO_925 (O_925,N_29919,N_29785);
nand UO_926 (O_926,N_29628,N_29862);
nor UO_927 (O_927,N_29489,N_29486);
or UO_928 (O_928,N_29789,N_29505);
or UO_929 (O_929,N_29555,N_29788);
nand UO_930 (O_930,N_29792,N_29885);
nor UO_931 (O_931,N_29763,N_29773);
nand UO_932 (O_932,N_29482,N_29773);
xor UO_933 (O_933,N_29592,N_29787);
xnor UO_934 (O_934,N_29533,N_29633);
and UO_935 (O_935,N_29408,N_29466);
or UO_936 (O_936,N_29984,N_29582);
and UO_937 (O_937,N_29900,N_29979);
nor UO_938 (O_938,N_29461,N_29566);
and UO_939 (O_939,N_29719,N_29445);
nand UO_940 (O_940,N_29947,N_29952);
nor UO_941 (O_941,N_29745,N_29893);
and UO_942 (O_942,N_29789,N_29943);
xor UO_943 (O_943,N_29993,N_29754);
and UO_944 (O_944,N_29619,N_29618);
nand UO_945 (O_945,N_29562,N_29574);
nor UO_946 (O_946,N_29752,N_29966);
and UO_947 (O_947,N_29413,N_29960);
nand UO_948 (O_948,N_29479,N_29403);
nor UO_949 (O_949,N_29595,N_29442);
nand UO_950 (O_950,N_29575,N_29522);
or UO_951 (O_951,N_29864,N_29944);
nand UO_952 (O_952,N_29733,N_29981);
and UO_953 (O_953,N_29805,N_29677);
xnor UO_954 (O_954,N_29430,N_29830);
xnor UO_955 (O_955,N_29492,N_29853);
and UO_956 (O_956,N_29468,N_29676);
nor UO_957 (O_957,N_29753,N_29989);
nor UO_958 (O_958,N_29856,N_29971);
or UO_959 (O_959,N_29871,N_29981);
and UO_960 (O_960,N_29613,N_29734);
nor UO_961 (O_961,N_29995,N_29436);
nor UO_962 (O_962,N_29862,N_29640);
nand UO_963 (O_963,N_29493,N_29510);
nor UO_964 (O_964,N_29492,N_29929);
xnor UO_965 (O_965,N_29612,N_29912);
nor UO_966 (O_966,N_29994,N_29440);
nor UO_967 (O_967,N_29819,N_29957);
xnor UO_968 (O_968,N_29863,N_29715);
xor UO_969 (O_969,N_29814,N_29729);
nand UO_970 (O_970,N_29511,N_29461);
or UO_971 (O_971,N_29676,N_29924);
and UO_972 (O_972,N_29913,N_29415);
nand UO_973 (O_973,N_29403,N_29714);
and UO_974 (O_974,N_29556,N_29765);
and UO_975 (O_975,N_29569,N_29732);
and UO_976 (O_976,N_29433,N_29629);
or UO_977 (O_977,N_29585,N_29770);
xnor UO_978 (O_978,N_29564,N_29677);
or UO_979 (O_979,N_29730,N_29933);
nor UO_980 (O_980,N_29963,N_29472);
or UO_981 (O_981,N_29897,N_29473);
or UO_982 (O_982,N_29562,N_29603);
nor UO_983 (O_983,N_29636,N_29522);
nor UO_984 (O_984,N_29627,N_29947);
or UO_985 (O_985,N_29492,N_29410);
xnor UO_986 (O_986,N_29762,N_29951);
nand UO_987 (O_987,N_29482,N_29466);
xnor UO_988 (O_988,N_29414,N_29730);
nor UO_989 (O_989,N_29494,N_29839);
nand UO_990 (O_990,N_29903,N_29894);
nor UO_991 (O_991,N_29935,N_29669);
or UO_992 (O_992,N_29612,N_29552);
and UO_993 (O_993,N_29764,N_29543);
xnor UO_994 (O_994,N_29680,N_29451);
or UO_995 (O_995,N_29750,N_29886);
or UO_996 (O_996,N_29852,N_29572);
and UO_997 (O_997,N_29520,N_29922);
or UO_998 (O_998,N_29701,N_29471);
xor UO_999 (O_999,N_29898,N_29785);
or UO_1000 (O_1000,N_29560,N_29745);
xor UO_1001 (O_1001,N_29583,N_29474);
nand UO_1002 (O_1002,N_29560,N_29624);
and UO_1003 (O_1003,N_29871,N_29573);
xnor UO_1004 (O_1004,N_29804,N_29928);
and UO_1005 (O_1005,N_29664,N_29466);
and UO_1006 (O_1006,N_29994,N_29572);
and UO_1007 (O_1007,N_29698,N_29629);
xnor UO_1008 (O_1008,N_29527,N_29631);
xnor UO_1009 (O_1009,N_29457,N_29723);
nand UO_1010 (O_1010,N_29818,N_29753);
nand UO_1011 (O_1011,N_29530,N_29794);
xor UO_1012 (O_1012,N_29507,N_29408);
or UO_1013 (O_1013,N_29642,N_29823);
and UO_1014 (O_1014,N_29749,N_29624);
or UO_1015 (O_1015,N_29639,N_29406);
and UO_1016 (O_1016,N_29712,N_29835);
and UO_1017 (O_1017,N_29942,N_29706);
nor UO_1018 (O_1018,N_29983,N_29445);
or UO_1019 (O_1019,N_29567,N_29644);
and UO_1020 (O_1020,N_29874,N_29684);
xor UO_1021 (O_1021,N_29459,N_29858);
nor UO_1022 (O_1022,N_29908,N_29728);
xnor UO_1023 (O_1023,N_29798,N_29965);
xnor UO_1024 (O_1024,N_29820,N_29498);
nor UO_1025 (O_1025,N_29473,N_29933);
xor UO_1026 (O_1026,N_29686,N_29621);
nand UO_1027 (O_1027,N_29406,N_29833);
nor UO_1028 (O_1028,N_29853,N_29871);
nor UO_1029 (O_1029,N_29853,N_29731);
and UO_1030 (O_1030,N_29959,N_29711);
xor UO_1031 (O_1031,N_29960,N_29507);
or UO_1032 (O_1032,N_29471,N_29918);
or UO_1033 (O_1033,N_29739,N_29790);
xor UO_1034 (O_1034,N_29685,N_29475);
nor UO_1035 (O_1035,N_29833,N_29928);
xor UO_1036 (O_1036,N_29863,N_29520);
and UO_1037 (O_1037,N_29661,N_29754);
xor UO_1038 (O_1038,N_29691,N_29746);
xnor UO_1039 (O_1039,N_29520,N_29495);
or UO_1040 (O_1040,N_29511,N_29809);
and UO_1041 (O_1041,N_29715,N_29619);
nor UO_1042 (O_1042,N_29898,N_29686);
xnor UO_1043 (O_1043,N_29434,N_29539);
and UO_1044 (O_1044,N_29813,N_29976);
xnor UO_1045 (O_1045,N_29531,N_29591);
xnor UO_1046 (O_1046,N_29820,N_29798);
or UO_1047 (O_1047,N_29557,N_29919);
and UO_1048 (O_1048,N_29953,N_29733);
and UO_1049 (O_1049,N_29718,N_29678);
and UO_1050 (O_1050,N_29926,N_29649);
xor UO_1051 (O_1051,N_29892,N_29558);
nor UO_1052 (O_1052,N_29745,N_29629);
nand UO_1053 (O_1053,N_29437,N_29450);
nor UO_1054 (O_1054,N_29946,N_29784);
nand UO_1055 (O_1055,N_29911,N_29916);
and UO_1056 (O_1056,N_29943,N_29727);
or UO_1057 (O_1057,N_29828,N_29665);
nand UO_1058 (O_1058,N_29454,N_29728);
and UO_1059 (O_1059,N_29792,N_29905);
or UO_1060 (O_1060,N_29533,N_29595);
or UO_1061 (O_1061,N_29859,N_29681);
xor UO_1062 (O_1062,N_29938,N_29402);
and UO_1063 (O_1063,N_29968,N_29553);
nor UO_1064 (O_1064,N_29559,N_29730);
and UO_1065 (O_1065,N_29447,N_29601);
and UO_1066 (O_1066,N_29726,N_29736);
xor UO_1067 (O_1067,N_29544,N_29814);
or UO_1068 (O_1068,N_29807,N_29512);
or UO_1069 (O_1069,N_29802,N_29588);
xnor UO_1070 (O_1070,N_29840,N_29510);
and UO_1071 (O_1071,N_29817,N_29810);
or UO_1072 (O_1072,N_29973,N_29897);
and UO_1073 (O_1073,N_29511,N_29636);
and UO_1074 (O_1074,N_29671,N_29984);
or UO_1075 (O_1075,N_29503,N_29444);
and UO_1076 (O_1076,N_29855,N_29631);
xor UO_1077 (O_1077,N_29970,N_29997);
nor UO_1078 (O_1078,N_29974,N_29495);
nand UO_1079 (O_1079,N_29763,N_29482);
xor UO_1080 (O_1080,N_29633,N_29784);
nand UO_1081 (O_1081,N_29657,N_29714);
nor UO_1082 (O_1082,N_29645,N_29728);
and UO_1083 (O_1083,N_29948,N_29683);
or UO_1084 (O_1084,N_29768,N_29582);
xnor UO_1085 (O_1085,N_29714,N_29976);
xor UO_1086 (O_1086,N_29529,N_29556);
and UO_1087 (O_1087,N_29666,N_29629);
xnor UO_1088 (O_1088,N_29470,N_29825);
nor UO_1089 (O_1089,N_29748,N_29879);
nor UO_1090 (O_1090,N_29808,N_29843);
nand UO_1091 (O_1091,N_29564,N_29802);
or UO_1092 (O_1092,N_29616,N_29531);
nand UO_1093 (O_1093,N_29709,N_29546);
or UO_1094 (O_1094,N_29419,N_29767);
xnor UO_1095 (O_1095,N_29803,N_29633);
or UO_1096 (O_1096,N_29573,N_29692);
nand UO_1097 (O_1097,N_29604,N_29607);
nand UO_1098 (O_1098,N_29679,N_29438);
nand UO_1099 (O_1099,N_29572,N_29939);
or UO_1100 (O_1100,N_29786,N_29757);
nand UO_1101 (O_1101,N_29429,N_29576);
xnor UO_1102 (O_1102,N_29863,N_29687);
and UO_1103 (O_1103,N_29636,N_29777);
or UO_1104 (O_1104,N_29946,N_29703);
nor UO_1105 (O_1105,N_29618,N_29693);
nand UO_1106 (O_1106,N_29754,N_29755);
and UO_1107 (O_1107,N_29769,N_29861);
nand UO_1108 (O_1108,N_29710,N_29443);
nand UO_1109 (O_1109,N_29753,N_29738);
and UO_1110 (O_1110,N_29912,N_29433);
and UO_1111 (O_1111,N_29978,N_29792);
or UO_1112 (O_1112,N_29753,N_29660);
xor UO_1113 (O_1113,N_29884,N_29757);
xor UO_1114 (O_1114,N_29686,N_29869);
or UO_1115 (O_1115,N_29880,N_29836);
nor UO_1116 (O_1116,N_29868,N_29612);
or UO_1117 (O_1117,N_29720,N_29837);
nor UO_1118 (O_1118,N_29631,N_29500);
or UO_1119 (O_1119,N_29604,N_29537);
nor UO_1120 (O_1120,N_29653,N_29454);
or UO_1121 (O_1121,N_29986,N_29465);
or UO_1122 (O_1122,N_29656,N_29838);
or UO_1123 (O_1123,N_29770,N_29994);
xor UO_1124 (O_1124,N_29468,N_29796);
and UO_1125 (O_1125,N_29580,N_29654);
and UO_1126 (O_1126,N_29898,N_29971);
or UO_1127 (O_1127,N_29901,N_29520);
xnor UO_1128 (O_1128,N_29740,N_29883);
nand UO_1129 (O_1129,N_29778,N_29543);
and UO_1130 (O_1130,N_29753,N_29590);
nor UO_1131 (O_1131,N_29703,N_29813);
or UO_1132 (O_1132,N_29731,N_29590);
and UO_1133 (O_1133,N_29421,N_29865);
nand UO_1134 (O_1134,N_29586,N_29991);
xor UO_1135 (O_1135,N_29813,N_29778);
and UO_1136 (O_1136,N_29742,N_29501);
xor UO_1137 (O_1137,N_29676,N_29634);
nor UO_1138 (O_1138,N_29739,N_29592);
and UO_1139 (O_1139,N_29790,N_29430);
and UO_1140 (O_1140,N_29836,N_29688);
and UO_1141 (O_1141,N_29999,N_29890);
or UO_1142 (O_1142,N_29929,N_29890);
or UO_1143 (O_1143,N_29559,N_29844);
and UO_1144 (O_1144,N_29546,N_29542);
nor UO_1145 (O_1145,N_29941,N_29504);
and UO_1146 (O_1146,N_29468,N_29959);
nor UO_1147 (O_1147,N_29435,N_29778);
or UO_1148 (O_1148,N_29689,N_29828);
and UO_1149 (O_1149,N_29903,N_29748);
nand UO_1150 (O_1150,N_29739,N_29736);
nor UO_1151 (O_1151,N_29719,N_29458);
xor UO_1152 (O_1152,N_29891,N_29567);
or UO_1153 (O_1153,N_29430,N_29839);
or UO_1154 (O_1154,N_29901,N_29720);
and UO_1155 (O_1155,N_29933,N_29503);
nand UO_1156 (O_1156,N_29956,N_29597);
nor UO_1157 (O_1157,N_29558,N_29752);
or UO_1158 (O_1158,N_29737,N_29744);
nor UO_1159 (O_1159,N_29905,N_29582);
xor UO_1160 (O_1160,N_29712,N_29553);
or UO_1161 (O_1161,N_29538,N_29837);
nand UO_1162 (O_1162,N_29870,N_29851);
and UO_1163 (O_1163,N_29610,N_29860);
xnor UO_1164 (O_1164,N_29980,N_29807);
or UO_1165 (O_1165,N_29977,N_29832);
nor UO_1166 (O_1166,N_29413,N_29831);
and UO_1167 (O_1167,N_29832,N_29706);
or UO_1168 (O_1168,N_29646,N_29763);
nand UO_1169 (O_1169,N_29727,N_29703);
nand UO_1170 (O_1170,N_29548,N_29594);
and UO_1171 (O_1171,N_29970,N_29543);
nor UO_1172 (O_1172,N_29684,N_29946);
nand UO_1173 (O_1173,N_29653,N_29453);
or UO_1174 (O_1174,N_29873,N_29591);
nor UO_1175 (O_1175,N_29542,N_29442);
and UO_1176 (O_1176,N_29482,N_29844);
nand UO_1177 (O_1177,N_29508,N_29677);
nand UO_1178 (O_1178,N_29671,N_29666);
or UO_1179 (O_1179,N_29547,N_29572);
or UO_1180 (O_1180,N_29729,N_29977);
xnor UO_1181 (O_1181,N_29964,N_29464);
xnor UO_1182 (O_1182,N_29465,N_29959);
and UO_1183 (O_1183,N_29558,N_29585);
nand UO_1184 (O_1184,N_29636,N_29434);
and UO_1185 (O_1185,N_29407,N_29433);
nor UO_1186 (O_1186,N_29989,N_29730);
nor UO_1187 (O_1187,N_29931,N_29643);
xnor UO_1188 (O_1188,N_29579,N_29788);
nand UO_1189 (O_1189,N_29582,N_29955);
xor UO_1190 (O_1190,N_29929,N_29733);
xnor UO_1191 (O_1191,N_29883,N_29670);
nand UO_1192 (O_1192,N_29433,N_29984);
nor UO_1193 (O_1193,N_29746,N_29652);
or UO_1194 (O_1194,N_29520,N_29778);
xnor UO_1195 (O_1195,N_29645,N_29442);
xnor UO_1196 (O_1196,N_29546,N_29550);
xnor UO_1197 (O_1197,N_29936,N_29574);
or UO_1198 (O_1198,N_29563,N_29827);
and UO_1199 (O_1199,N_29908,N_29930);
or UO_1200 (O_1200,N_29637,N_29975);
nor UO_1201 (O_1201,N_29408,N_29605);
xnor UO_1202 (O_1202,N_29478,N_29728);
xor UO_1203 (O_1203,N_29923,N_29888);
or UO_1204 (O_1204,N_29765,N_29607);
or UO_1205 (O_1205,N_29438,N_29456);
nand UO_1206 (O_1206,N_29952,N_29666);
or UO_1207 (O_1207,N_29542,N_29744);
nor UO_1208 (O_1208,N_29799,N_29410);
xor UO_1209 (O_1209,N_29970,N_29584);
nor UO_1210 (O_1210,N_29620,N_29465);
xnor UO_1211 (O_1211,N_29688,N_29468);
or UO_1212 (O_1212,N_29736,N_29966);
nor UO_1213 (O_1213,N_29669,N_29498);
nand UO_1214 (O_1214,N_29602,N_29618);
or UO_1215 (O_1215,N_29439,N_29409);
and UO_1216 (O_1216,N_29547,N_29909);
and UO_1217 (O_1217,N_29772,N_29517);
or UO_1218 (O_1218,N_29782,N_29843);
or UO_1219 (O_1219,N_29465,N_29439);
nor UO_1220 (O_1220,N_29896,N_29636);
and UO_1221 (O_1221,N_29464,N_29504);
xor UO_1222 (O_1222,N_29407,N_29986);
and UO_1223 (O_1223,N_29734,N_29401);
nand UO_1224 (O_1224,N_29552,N_29847);
nand UO_1225 (O_1225,N_29635,N_29625);
nand UO_1226 (O_1226,N_29585,N_29427);
xnor UO_1227 (O_1227,N_29624,N_29525);
or UO_1228 (O_1228,N_29757,N_29970);
and UO_1229 (O_1229,N_29947,N_29925);
nor UO_1230 (O_1230,N_29572,N_29881);
nor UO_1231 (O_1231,N_29656,N_29903);
nor UO_1232 (O_1232,N_29483,N_29591);
or UO_1233 (O_1233,N_29483,N_29903);
nor UO_1234 (O_1234,N_29977,N_29410);
or UO_1235 (O_1235,N_29774,N_29754);
and UO_1236 (O_1236,N_29480,N_29405);
or UO_1237 (O_1237,N_29551,N_29462);
xnor UO_1238 (O_1238,N_29405,N_29707);
and UO_1239 (O_1239,N_29656,N_29519);
and UO_1240 (O_1240,N_29844,N_29757);
and UO_1241 (O_1241,N_29739,N_29713);
or UO_1242 (O_1242,N_29831,N_29525);
nor UO_1243 (O_1243,N_29857,N_29911);
xnor UO_1244 (O_1244,N_29534,N_29872);
xnor UO_1245 (O_1245,N_29470,N_29952);
nor UO_1246 (O_1246,N_29887,N_29562);
nor UO_1247 (O_1247,N_29541,N_29876);
nor UO_1248 (O_1248,N_29945,N_29770);
nor UO_1249 (O_1249,N_29936,N_29822);
or UO_1250 (O_1250,N_29554,N_29911);
xor UO_1251 (O_1251,N_29830,N_29768);
or UO_1252 (O_1252,N_29415,N_29647);
and UO_1253 (O_1253,N_29495,N_29483);
nor UO_1254 (O_1254,N_29711,N_29946);
xor UO_1255 (O_1255,N_29668,N_29823);
or UO_1256 (O_1256,N_29663,N_29934);
nor UO_1257 (O_1257,N_29508,N_29906);
xnor UO_1258 (O_1258,N_29617,N_29763);
nand UO_1259 (O_1259,N_29480,N_29735);
or UO_1260 (O_1260,N_29838,N_29890);
nor UO_1261 (O_1261,N_29455,N_29871);
nand UO_1262 (O_1262,N_29941,N_29808);
nand UO_1263 (O_1263,N_29481,N_29827);
or UO_1264 (O_1264,N_29428,N_29873);
or UO_1265 (O_1265,N_29955,N_29779);
nor UO_1266 (O_1266,N_29466,N_29572);
xor UO_1267 (O_1267,N_29590,N_29478);
nor UO_1268 (O_1268,N_29617,N_29892);
xor UO_1269 (O_1269,N_29766,N_29703);
or UO_1270 (O_1270,N_29562,N_29661);
xor UO_1271 (O_1271,N_29919,N_29654);
xnor UO_1272 (O_1272,N_29666,N_29752);
nand UO_1273 (O_1273,N_29914,N_29712);
or UO_1274 (O_1274,N_29930,N_29496);
nor UO_1275 (O_1275,N_29656,N_29507);
xor UO_1276 (O_1276,N_29738,N_29663);
nor UO_1277 (O_1277,N_29709,N_29799);
nor UO_1278 (O_1278,N_29565,N_29443);
or UO_1279 (O_1279,N_29682,N_29774);
xnor UO_1280 (O_1280,N_29948,N_29945);
and UO_1281 (O_1281,N_29471,N_29878);
or UO_1282 (O_1282,N_29420,N_29434);
or UO_1283 (O_1283,N_29509,N_29480);
or UO_1284 (O_1284,N_29411,N_29758);
xor UO_1285 (O_1285,N_29425,N_29450);
and UO_1286 (O_1286,N_29602,N_29793);
nor UO_1287 (O_1287,N_29915,N_29451);
nand UO_1288 (O_1288,N_29743,N_29815);
or UO_1289 (O_1289,N_29913,N_29435);
and UO_1290 (O_1290,N_29518,N_29729);
or UO_1291 (O_1291,N_29653,N_29994);
nand UO_1292 (O_1292,N_29927,N_29905);
nand UO_1293 (O_1293,N_29517,N_29690);
xnor UO_1294 (O_1294,N_29645,N_29754);
nor UO_1295 (O_1295,N_29522,N_29865);
xor UO_1296 (O_1296,N_29539,N_29544);
nor UO_1297 (O_1297,N_29687,N_29826);
nor UO_1298 (O_1298,N_29954,N_29804);
xnor UO_1299 (O_1299,N_29612,N_29501);
or UO_1300 (O_1300,N_29538,N_29633);
nor UO_1301 (O_1301,N_29714,N_29414);
or UO_1302 (O_1302,N_29539,N_29549);
and UO_1303 (O_1303,N_29922,N_29584);
nor UO_1304 (O_1304,N_29566,N_29832);
and UO_1305 (O_1305,N_29649,N_29418);
or UO_1306 (O_1306,N_29577,N_29643);
or UO_1307 (O_1307,N_29609,N_29483);
xor UO_1308 (O_1308,N_29719,N_29452);
and UO_1309 (O_1309,N_29738,N_29545);
nand UO_1310 (O_1310,N_29930,N_29906);
xor UO_1311 (O_1311,N_29566,N_29750);
xnor UO_1312 (O_1312,N_29503,N_29504);
or UO_1313 (O_1313,N_29764,N_29752);
xor UO_1314 (O_1314,N_29468,N_29940);
nor UO_1315 (O_1315,N_29724,N_29755);
nand UO_1316 (O_1316,N_29903,N_29671);
nor UO_1317 (O_1317,N_29580,N_29775);
nand UO_1318 (O_1318,N_29852,N_29505);
or UO_1319 (O_1319,N_29719,N_29473);
or UO_1320 (O_1320,N_29888,N_29554);
or UO_1321 (O_1321,N_29780,N_29494);
and UO_1322 (O_1322,N_29417,N_29651);
and UO_1323 (O_1323,N_29682,N_29926);
nand UO_1324 (O_1324,N_29970,N_29871);
or UO_1325 (O_1325,N_29559,N_29995);
xnor UO_1326 (O_1326,N_29433,N_29951);
and UO_1327 (O_1327,N_29595,N_29990);
or UO_1328 (O_1328,N_29952,N_29480);
or UO_1329 (O_1329,N_29518,N_29893);
and UO_1330 (O_1330,N_29631,N_29539);
nor UO_1331 (O_1331,N_29518,N_29858);
and UO_1332 (O_1332,N_29800,N_29852);
nand UO_1333 (O_1333,N_29702,N_29808);
nand UO_1334 (O_1334,N_29535,N_29716);
nor UO_1335 (O_1335,N_29812,N_29723);
or UO_1336 (O_1336,N_29618,N_29449);
nand UO_1337 (O_1337,N_29729,N_29647);
nand UO_1338 (O_1338,N_29405,N_29654);
nor UO_1339 (O_1339,N_29639,N_29798);
and UO_1340 (O_1340,N_29665,N_29571);
or UO_1341 (O_1341,N_29521,N_29446);
or UO_1342 (O_1342,N_29782,N_29757);
nor UO_1343 (O_1343,N_29882,N_29968);
nand UO_1344 (O_1344,N_29686,N_29496);
xor UO_1345 (O_1345,N_29682,N_29515);
or UO_1346 (O_1346,N_29576,N_29452);
nand UO_1347 (O_1347,N_29762,N_29633);
or UO_1348 (O_1348,N_29770,N_29904);
or UO_1349 (O_1349,N_29533,N_29596);
and UO_1350 (O_1350,N_29733,N_29749);
xor UO_1351 (O_1351,N_29551,N_29414);
nor UO_1352 (O_1352,N_29645,N_29673);
and UO_1353 (O_1353,N_29847,N_29698);
nand UO_1354 (O_1354,N_29993,N_29854);
or UO_1355 (O_1355,N_29913,N_29900);
xor UO_1356 (O_1356,N_29519,N_29941);
and UO_1357 (O_1357,N_29908,N_29707);
nor UO_1358 (O_1358,N_29548,N_29793);
nand UO_1359 (O_1359,N_29976,N_29524);
and UO_1360 (O_1360,N_29993,N_29443);
or UO_1361 (O_1361,N_29877,N_29489);
and UO_1362 (O_1362,N_29657,N_29861);
or UO_1363 (O_1363,N_29681,N_29893);
or UO_1364 (O_1364,N_29441,N_29457);
xor UO_1365 (O_1365,N_29962,N_29713);
xnor UO_1366 (O_1366,N_29786,N_29846);
xnor UO_1367 (O_1367,N_29813,N_29523);
nor UO_1368 (O_1368,N_29964,N_29522);
xor UO_1369 (O_1369,N_29636,N_29568);
and UO_1370 (O_1370,N_29835,N_29901);
nor UO_1371 (O_1371,N_29799,N_29897);
nand UO_1372 (O_1372,N_29519,N_29606);
or UO_1373 (O_1373,N_29863,N_29410);
or UO_1374 (O_1374,N_29920,N_29759);
or UO_1375 (O_1375,N_29496,N_29972);
nand UO_1376 (O_1376,N_29898,N_29746);
or UO_1377 (O_1377,N_29647,N_29621);
nand UO_1378 (O_1378,N_29939,N_29597);
nand UO_1379 (O_1379,N_29911,N_29689);
nor UO_1380 (O_1380,N_29552,N_29956);
nor UO_1381 (O_1381,N_29719,N_29495);
xnor UO_1382 (O_1382,N_29995,N_29536);
and UO_1383 (O_1383,N_29576,N_29894);
or UO_1384 (O_1384,N_29556,N_29829);
xor UO_1385 (O_1385,N_29558,N_29691);
or UO_1386 (O_1386,N_29912,N_29491);
and UO_1387 (O_1387,N_29646,N_29604);
or UO_1388 (O_1388,N_29507,N_29665);
nor UO_1389 (O_1389,N_29576,N_29953);
nand UO_1390 (O_1390,N_29943,N_29760);
nand UO_1391 (O_1391,N_29602,N_29785);
xnor UO_1392 (O_1392,N_29748,N_29934);
nand UO_1393 (O_1393,N_29590,N_29845);
nand UO_1394 (O_1394,N_29992,N_29826);
nor UO_1395 (O_1395,N_29880,N_29852);
nand UO_1396 (O_1396,N_29605,N_29607);
nand UO_1397 (O_1397,N_29938,N_29855);
nand UO_1398 (O_1398,N_29836,N_29615);
and UO_1399 (O_1399,N_29602,N_29983);
xnor UO_1400 (O_1400,N_29690,N_29811);
nand UO_1401 (O_1401,N_29848,N_29804);
and UO_1402 (O_1402,N_29654,N_29569);
nand UO_1403 (O_1403,N_29935,N_29643);
or UO_1404 (O_1404,N_29794,N_29566);
and UO_1405 (O_1405,N_29650,N_29894);
and UO_1406 (O_1406,N_29742,N_29999);
and UO_1407 (O_1407,N_29505,N_29518);
and UO_1408 (O_1408,N_29447,N_29918);
or UO_1409 (O_1409,N_29544,N_29463);
nand UO_1410 (O_1410,N_29620,N_29484);
or UO_1411 (O_1411,N_29595,N_29865);
xor UO_1412 (O_1412,N_29594,N_29665);
or UO_1413 (O_1413,N_29809,N_29835);
nand UO_1414 (O_1414,N_29551,N_29965);
or UO_1415 (O_1415,N_29695,N_29694);
or UO_1416 (O_1416,N_29765,N_29976);
and UO_1417 (O_1417,N_29655,N_29854);
xor UO_1418 (O_1418,N_29672,N_29656);
or UO_1419 (O_1419,N_29415,N_29964);
and UO_1420 (O_1420,N_29730,N_29757);
nor UO_1421 (O_1421,N_29676,N_29786);
nor UO_1422 (O_1422,N_29966,N_29420);
nor UO_1423 (O_1423,N_29508,N_29453);
or UO_1424 (O_1424,N_29773,N_29663);
xor UO_1425 (O_1425,N_29837,N_29444);
nand UO_1426 (O_1426,N_29593,N_29611);
nand UO_1427 (O_1427,N_29420,N_29662);
and UO_1428 (O_1428,N_29475,N_29447);
nand UO_1429 (O_1429,N_29561,N_29618);
and UO_1430 (O_1430,N_29689,N_29940);
nand UO_1431 (O_1431,N_29561,N_29658);
or UO_1432 (O_1432,N_29774,N_29446);
xnor UO_1433 (O_1433,N_29788,N_29781);
nand UO_1434 (O_1434,N_29455,N_29920);
xnor UO_1435 (O_1435,N_29722,N_29873);
or UO_1436 (O_1436,N_29932,N_29955);
and UO_1437 (O_1437,N_29824,N_29614);
or UO_1438 (O_1438,N_29863,N_29803);
xnor UO_1439 (O_1439,N_29699,N_29936);
and UO_1440 (O_1440,N_29901,N_29488);
nand UO_1441 (O_1441,N_29769,N_29845);
or UO_1442 (O_1442,N_29744,N_29557);
nor UO_1443 (O_1443,N_29619,N_29572);
nor UO_1444 (O_1444,N_29903,N_29957);
nor UO_1445 (O_1445,N_29774,N_29715);
nor UO_1446 (O_1446,N_29526,N_29632);
nor UO_1447 (O_1447,N_29462,N_29963);
nor UO_1448 (O_1448,N_29446,N_29821);
nor UO_1449 (O_1449,N_29753,N_29782);
and UO_1450 (O_1450,N_29515,N_29553);
or UO_1451 (O_1451,N_29693,N_29463);
or UO_1452 (O_1452,N_29974,N_29664);
nand UO_1453 (O_1453,N_29463,N_29986);
or UO_1454 (O_1454,N_29584,N_29473);
and UO_1455 (O_1455,N_29887,N_29693);
xnor UO_1456 (O_1456,N_29409,N_29597);
xor UO_1457 (O_1457,N_29730,N_29934);
and UO_1458 (O_1458,N_29547,N_29403);
nor UO_1459 (O_1459,N_29921,N_29702);
or UO_1460 (O_1460,N_29894,N_29552);
nor UO_1461 (O_1461,N_29593,N_29444);
nor UO_1462 (O_1462,N_29557,N_29582);
xnor UO_1463 (O_1463,N_29417,N_29802);
nor UO_1464 (O_1464,N_29651,N_29968);
nand UO_1465 (O_1465,N_29901,N_29597);
xnor UO_1466 (O_1466,N_29547,N_29759);
xnor UO_1467 (O_1467,N_29739,N_29494);
nand UO_1468 (O_1468,N_29606,N_29662);
nor UO_1469 (O_1469,N_29596,N_29781);
nand UO_1470 (O_1470,N_29804,N_29509);
nand UO_1471 (O_1471,N_29581,N_29490);
nand UO_1472 (O_1472,N_29835,N_29510);
xnor UO_1473 (O_1473,N_29810,N_29774);
nand UO_1474 (O_1474,N_29723,N_29491);
xnor UO_1475 (O_1475,N_29566,N_29721);
nor UO_1476 (O_1476,N_29693,N_29866);
xnor UO_1477 (O_1477,N_29903,N_29496);
nor UO_1478 (O_1478,N_29826,N_29422);
or UO_1479 (O_1479,N_29681,N_29647);
nor UO_1480 (O_1480,N_29510,N_29508);
nand UO_1481 (O_1481,N_29422,N_29449);
nor UO_1482 (O_1482,N_29683,N_29791);
or UO_1483 (O_1483,N_29495,N_29904);
or UO_1484 (O_1484,N_29838,N_29934);
or UO_1485 (O_1485,N_29652,N_29563);
nor UO_1486 (O_1486,N_29688,N_29938);
xnor UO_1487 (O_1487,N_29796,N_29423);
or UO_1488 (O_1488,N_29621,N_29551);
and UO_1489 (O_1489,N_29614,N_29782);
or UO_1490 (O_1490,N_29684,N_29905);
nor UO_1491 (O_1491,N_29517,N_29854);
xor UO_1492 (O_1492,N_29937,N_29506);
nand UO_1493 (O_1493,N_29540,N_29626);
nand UO_1494 (O_1494,N_29600,N_29694);
or UO_1495 (O_1495,N_29452,N_29501);
nor UO_1496 (O_1496,N_29847,N_29452);
or UO_1497 (O_1497,N_29690,N_29475);
and UO_1498 (O_1498,N_29867,N_29533);
xnor UO_1499 (O_1499,N_29668,N_29405);
xnor UO_1500 (O_1500,N_29978,N_29896);
or UO_1501 (O_1501,N_29876,N_29578);
nor UO_1502 (O_1502,N_29672,N_29539);
nand UO_1503 (O_1503,N_29646,N_29525);
nor UO_1504 (O_1504,N_29497,N_29929);
or UO_1505 (O_1505,N_29792,N_29846);
nand UO_1506 (O_1506,N_29570,N_29564);
or UO_1507 (O_1507,N_29967,N_29866);
nor UO_1508 (O_1508,N_29638,N_29879);
nand UO_1509 (O_1509,N_29483,N_29942);
nor UO_1510 (O_1510,N_29734,N_29473);
nand UO_1511 (O_1511,N_29620,N_29518);
and UO_1512 (O_1512,N_29804,N_29401);
xnor UO_1513 (O_1513,N_29712,N_29718);
and UO_1514 (O_1514,N_29498,N_29932);
or UO_1515 (O_1515,N_29814,N_29601);
nand UO_1516 (O_1516,N_29824,N_29573);
and UO_1517 (O_1517,N_29659,N_29470);
nor UO_1518 (O_1518,N_29401,N_29732);
nand UO_1519 (O_1519,N_29431,N_29477);
and UO_1520 (O_1520,N_29851,N_29708);
or UO_1521 (O_1521,N_29806,N_29740);
nor UO_1522 (O_1522,N_29529,N_29584);
nor UO_1523 (O_1523,N_29886,N_29640);
nor UO_1524 (O_1524,N_29959,N_29430);
nor UO_1525 (O_1525,N_29858,N_29714);
nor UO_1526 (O_1526,N_29644,N_29591);
nor UO_1527 (O_1527,N_29556,N_29998);
and UO_1528 (O_1528,N_29496,N_29671);
and UO_1529 (O_1529,N_29999,N_29757);
xor UO_1530 (O_1530,N_29587,N_29595);
or UO_1531 (O_1531,N_29549,N_29733);
and UO_1532 (O_1532,N_29861,N_29544);
nand UO_1533 (O_1533,N_29948,N_29443);
or UO_1534 (O_1534,N_29895,N_29888);
nor UO_1535 (O_1535,N_29626,N_29636);
xor UO_1536 (O_1536,N_29800,N_29644);
nor UO_1537 (O_1537,N_29593,N_29605);
nand UO_1538 (O_1538,N_29615,N_29448);
and UO_1539 (O_1539,N_29425,N_29714);
or UO_1540 (O_1540,N_29648,N_29960);
nor UO_1541 (O_1541,N_29546,N_29953);
and UO_1542 (O_1542,N_29979,N_29532);
nor UO_1543 (O_1543,N_29623,N_29699);
and UO_1544 (O_1544,N_29445,N_29834);
or UO_1545 (O_1545,N_29688,N_29840);
and UO_1546 (O_1546,N_29796,N_29592);
xnor UO_1547 (O_1547,N_29494,N_29722);
nor UO_1548 (O_1548,N_29948,N_29844);
or UO_1549 (O_1549,N_29489,N_29480);
or UO_1550 (O_1550,N_29773,N_29957);
and UO_1551 (O_1551,N_29468,N_29459);
xor UO_1552 (O_1552,N_29618,N_29423);
or UO_1553 (O_1553,N_29866,N_29926);
xor UO_1554 (O_1554,N_29408,N_29902);
or UO_1555 (O_1555,N_29935,N_29675);
xor UO_1556 (O_1556,N_29718,N_29660);
nand UO_1557 (O_1557,N_29800,N_29556);
or UO_1558 (O_1558,N_29910,N_29912);
nand UO_1559 (O_1559,N_29453,N_29560);
or UO_1560 (O_1560,N_29576,N_29948);
or UO_1561 (O_1561,N_29488,N_29494);
and UO_1562 (O_1562,N_29607,N_29813);
and UO_1563 (O_1563,N_29911,N_29943);
and UO_1564 (O_1564,N_29498,N_29526);
xor UO_1565 (O_1565,N_29984,N_29411);
nand UO_1566 (O_1566,N_29901,N_29749);
xnor UO_1567 (O_1567,N_29907,N_29569);
or UO_1568 (O_1568,N_29985,N_29688);
nand UO_1569 (O_1569,N_29425,N_29742);
or UO_1570 (O_1570,N_29886,N_29803);
nor UO_1571 (O_1571,N_29766,N_29818);
nand UO_1572 (O_1572,N_29435,N_29605);
or UO_1573 (O_1573,N_29612,N_29746);
and UO_1574 (O_1574,N_29786,N_29443);
or UO_1575 (O_1575,N_29466,N_29598);
nor UO_1576 (O_1576,N_29745,N_29545);
nand UO_1577 (O_1577,N_29643,N_29635);
nand UO_1578 (O_1578,N_29817,N_29834);
and UO_1579 (O_1579,N_29802,N_29771);
xor UO_1580 (O_1580,N_29525,N_29777);
nand UO_1581 (O_1581,N_29761,N_29508);
nor UO_1582 (O_1582,N_29454,N_29753);
or UO_1583 (O_1583,N_29588,N_29753);
nor UO_1584 (O_1584,N_29800,N_29928);
or UO_1585 (O_1585,N_29663,N_29406);
xor UO_1586 (O_1586,N_29927,N_29835);
nand UO_1587 (O_1587,N_29784,N_29894);
nand UO_1588 (O_1588,N_29663,N_29820);
xnor UO_1589 (O_1589,N_29912,N_29817);
nand UO_1590 (O_1590,N_29924,N_29896);
and UO_1591 (O_1591,N_29782,N_29906);
xor UO_1592 (O_1592,N_29407,N_29482);
nor UO_1593 (O_1593,N_29865,N_29757);
nor UO_1594 (O_1594,N_29694,N_29667);
or UO_1595 (O_1595,N_29773,N_29768);
or UO_1596 (O_1596,N_29755,N_29952);
nand UO_1597 (O_1597,N_29500,N_29731);
nand UO_1598 (O_1598,N_29655,N_29645);
or UO_1599 (O_1599,N_29932,N_29711);
nand UO_1600 (O_1600,N_29806,N_29996);
or UO_1601 (O_1601,N_29787,N_29510);
or UO_1602 (O_1602,N_29682,N_29679);
nand UO_1603 (O_1603,N_29678,N_29811);
xor UO_1604 (O_1604,N_29456,N_29417);
nor UO_1605 (O_1605,N_29926,N_29933);
and UO_1606 (O_1606,N_29993,N_29633);
and UO_1607 (O_1607,N_29900,N_29978);
nand UO_1608 (O_1608,N_29822,N_29938);
nor UO_1609 (O_1609,N_29980,N_29777);
or UO_1610 (O_1610,N_29427,N_29493);
or UO_1611 (O_1611,N_29522,N_29568);
xnor UO_1612 (O_1612,N_29582,N_29805);
and UO_1613 (O_1613,N_29901,N_29613);
and UO_1614 (O_1614,N_29956,N_29507);
xor UO_1615 (O_1615,N_29443,N_29680);
and UO_1616 (O_1616,N_29408,N_29942);
nand UO_1617 (O_1617,N_29675,N_29788);
nand UO_1618 (O_1618,N_29451,N_29656);
nand UO_1619 (O_1619,N_29934,N_29595);
nand UO_1620 (O_1620,N_29816,N_29683);
nand UO_1621 (O_1621,N_29585,N_29779);
xor UO_1622 (O_1622,N_29482,N_29882);
nor UO_1623 (O_1623,N_29400,N_29534);
or UO_1624 (O_1624,N_29744,N_29534);
xor UO_1625 (O_1625,N_29912,N_29963);
or UO_1626 (O_1626,N_29963,N_29842);
nor UO_1627 (O_1627,N_29572,N_29993);
nor UO_1628 (O_1628,N_29936,N_29970);
or UO_1629 (O_1629,N_29963,N_29837);
nor UO_1630 (O_1630,N_29882,N_29468);
nor UO_1631 (O_1631,N_29918,N_29937);
nand UO_1632 (O_1632,N_29505,N_29897);
nand UO_1633 (O_1633,N_29522,N_29778);
nor UO_1634 (O_1634,N_29823,N_29854);
nand UO_1635 (O_1635,N_29535,N_29547);
nand UO_1636 (O_1636,N_29985,N_29827);
and UO_1637 (O_1637,N_29829,N_29598);
nor UO_1638 (O_1638,N_29899,N_29585);
xor UO_1639 (O_1639,N_29403,N_29826);
xor UO_1640 (O_1640,N_29519,N_29643);
and UO_1641 (O_1641,N_29427,N_29442);
and UO_1642 (O_1642,N_29791,N_29800);
nand UO_1643 (O_1643,N_29652,N_29601);
or UO_1644 (O_1644,N_29978,N_29838);
nor UO_1645 (O_1645,N_29403,N_29546);
and UO_1646 (O_1646,N_29886,N_29699);
and UO_1647 (O_1647,N_29825,N_29821);
nand UO_1648 (O_1648,N_29673,N_29662);
xor UO_1649 (O_1649,N_29445,N_29644);
nor UO_1650 (O_1650,N_29872,N_29809);
and UO_1651 (O_1651,N_29904,N_29742);
nand UO_1652 (O_1652,N_29870,N_29619);
nor UO_1653 (O_1653,N_29819,N_29460);
or UO_1654 (O_1654,N_29438,N_29667);
or UO_1655 (O_1655,N_29971,N_29773);
or UO_1656 (O_1656,N_29708,N_29985);
and UO_1657 (O_1657,N_29872,N_29821);
or UO_1658 (O_1658,N_29579,N_29473);
nor UO_1659 (O_1659,N_29459,N_29466);
xnor UO_1660 (O_1660,N_29741,N_29735);
or UO_1661 (O_1661,N_29852,N_29820);
nor UO_1662 (O_1662,N_29425,N_29939);
or UO_1663 (O_1663,N_29857,N_29657);
and UO_1664 (O_1664,N_29933,N_29745);
and UO_1665 (O_1665,N_29825,N_29418);
nand UO_1666 (O_1666,N_29844,N_29543);
nand UO_1667 (O_1667,N_29838,N_29917);
or UO_1668 (O_1668,N_29489,N_29700);
and UO_1669 (O_1669,N_29469,N_29669);
xnor UO_1670 (O_1670,N_29443,N_29791);
and UO_1671 (O_1671,N_29808,N_29536);
xor UO_1672 (O_1672,N_29798,N_29630);
nor UO_1673 (O_1673,N_29950,N_29665);
nand UO_1674 (O_1674,N_29680,N_29612);
or UO_1675 (O_1675,N_29553,N_29789);
xnor UO_1676 (O_1676,N_29493,N_29513);
nand UO_1677 (O_1677,N_29801,N_29441);
nor UO_1678 (O_1678,N_29921,N_29881);
and UO_1679 (O_1679,N_29743,N_29572);
xor UO_1680 (O_1680,N_29532,N_29641);
nand UO_1681 (O_1681,N_29959,N_29873);
nor UO_1682 (O_1682,N_29465,N_29763);
nor UO_1683 (O_1683,N_29719,N_29465);
and UO_1684 (O_1684,N_29659,N_29428);
or UO_1685 (O_1685,N_29410,N_29814);
nor UO_1686 (O_1686,N_29815,N_29598);
or UO_1687 (O_1687,N_29865,N_29968);
xor UO_1688 (O_1688,N_29599,N_29819);
nand UO_1689 (O_1689,N_29510,N_29666);
nand UO_1690 (O_1690,N_29813,N_29896);
xor UO_1691 (O_1691,N_29922,N_29500);
nor UO_1692 (O_1692,N_29467,N_29862);
or UO_1693 (O_1693,N_29667,N_29805);
nor UO_1694 (O_1694,N_29755,N_29646);
xor UO_1695 (O_1695,N_29992,N_29480);
or UO_1696 (O_1696,N_29692,N_29886);
xnor UO_1697 (O_1697,N_29776,N_29627);
or UO_1698 (O_1698,N_29494,N_29609);
or UO_1699 (O_1699,N_29778,N_29576);
or UO_1700 (O_1700,N_29816,N_29707);
or UO_1701 (O_1701,N_29794,N_29432);
and UO_1702 (O_1702,N_29459,N_29469);
xor UO_1703 (O_1703,N_29710,N_29517);
xor UO_1704 (O_1704,N_29878,N_29627);
and UO_1705 (O_1705,N_29916,N_29875);
and UO_1706 (O_1706,N_29726,N_29678);
xnor UO_1707 (O_1707,N_29888,N_29740);
or UO_1708 (O_1708,N_29917,N_29665);
and UO_1709 (O_1709,N_29859,N_29413);
and UO_1710 (O_1710,N_29827,N_29671);
nor UO_1711 (O_1711,N_29734,N_29447);
nor UO_1712 (O_1712,N_29528,N_29715);
xnor UO_1713 (O_1713,N_29912,N_29585);
nor UO_1714 (O_1714,N_29625,N_29714);
or UO_1715 (O_1715,N_29589,N_29526);
nor UO_1716 (O_1716,N_29735,N_29912);
nor UO_1717 (O_1717,N_29717,N_29920);
xnor UO_1718 (O_1718,N_29488,N_29776);
and UO_1719 (O_1719,N_29741,N_29836);
nor UO_1720 (O_1720,N_29713,N_29933);
and UO_1721 (O_1721,N_29945,N_29608);
xor UO_1722 (O_1722,N_29455,N_29528);
and UO_1723 (O_1723,N_29886,N_29846);
nand UO_1724 (O_1724,N_29770,N_29407);
xor UO_1725 (O_1725,N_29607,N_29672);
and UO_1726 (O_1726,N_29587,N_29708);
xnor UO_1727 (O_1727,N_29432,N_29851);
nor UO_1728 (O_1728,N_29660,N_29983);
and UO_1729 (O_1729,N_29734,N_29652);
nor UO_1730 (O_1730,N_29641,N_29902);
xor UO_1731 (O_1731,N_29908,N_29712);
and UO_1732 (O_1732,N_29489,N_29880);
xor UO_1733 (O_1733,N_29746,N_29666);
or UO_1734 (O_1734,N_29597,N_29648);
nand UO_1735 (O_1735,N_29515,N_29468);
and UO_1736 (O_1736,N_29402,N_29872);
and UO_1737 (O_1737,N_29952,N_29493);
xor UO_1738 (O_1738,N_29620,N_29705);
nor UO_1739 (O_1739,N_29676,N_29432);
nand UO_1740 (O_1740,N_29541,N_29695);
xor UO_1741 (O_1741,N_29926,N_29617);
xor UO_1742 (O_1742,N_29565,N_29897);
nand UO_1743 (O_1743,N_29542,N_29637);
nand UO_1744 (O_1744,N_29809,N_29790);
and UO_1745 (O_1745,N_29618,N_29556);
xor UO_1746 (O_1746,N_29647,N_29911);
and UO_1747 (O_1747,N_29786,N_29762);
nor UO_1748 (O_1748,N_29640,N_29689);
xor UO_1749 (O_1749,N_29678,N_29907);
xnor UO_1750 (O_1750,N_29431,N_29514);
nand UO_1751 (O_1751,N_29870,N_29882);
nand UO_1752 (O_1752,N_29492,N_29541);
and UO_1753 (O_1753,N_29758,N_29574);
or UO_1754 (O_1754,N_29968,N_29810);
nor UO_1755 (O_1755,N_29909,N_29998);
nand UO_1756 (O_1756,N_29576,N_29855);
nor UO_1757 (O_1757,N_29422,N_29818);
xor UO_1758 (O_1758,N_29938,N_29961);
nand UO_1759 (O_1759,N_29444,N_29409);
xor UO_1760 (O_1760,N_29516,N_29755);
and UO_1761 (O_1761,N_29525,N_29655);
or UO_1762 (O_1762,N_29729,N_29955);
or UO_1763 (O_1763,N_29795,N_29733);
nand UO_1764 (O_1764,N_29929,N_29480);
xnor UO_1765 (O_1765,N_29782,N_29657);
or UO_1766 (O_1766,N_29861,N_29605);
and UO_1767 (O_1767,N_29523,N_29907);
or UO_1768 (O_1768,N_29416,N_29892);
nor UO_1769 (O_1769,N_29702,N_29501);
xnor UO_1770 (O_1770,N_29723,N_29735);
or UO_1771 (O_1771,N_29584,N_29417);
or UO_1772 (O_1772,N_29985,N_29626);
xnor UO_1773 (O_1773,N_29757,N_29995);
nor UO_1774 (O_1774,N_29921,N_29988);
nor UO_1775 (O_1775,N_29472,N_29877);
or UO_1776 (O_1776,N_29807,N_29568);
xnor UO_1777 (O_1777,N_29644,N_29923);
and UO_1778 (O_1778,N_29562,N_29951);
and UO_1779 (O_1779,N_29497,N_29973);
xor UO_1780 (O_1780,N_29427,N_29451);
and UO_1781 (O_1781,N_29515,N_29904);
nor UO_1782 (O_1782,N_29703,N_29835);
xor UO_1783 (O_1783,N_29682,N_29914);
xor UO_1784 (O_1784,N_29763,N_29524);
or UO_1785 (O_1785,N_29762,N_29528);
or UO_1786 (O_1786,N_29459,N_29738);
nor UO_1787 (O_1787,N_29823,N_29719);
or UO_1788 (O_1788,N_29668,N_29974);
nand UO_1789 (O_1789,N_29969,N_29933);
or UO_1790 (O_1790,N_29801,N_29992);
nor UO_1791 (O_1791,N_29987,N_29990);
nor UO_1792 (O_1792,N_29705,N_29449);
xnor UO_1793 (O_1793,N_29649,N_29439);
and UO_1794 (O_1794,N_29476,N_29767);
nand UO_1795 (O_1795,N_29417,N_29963);
and UO_1796 (O_1796,N_29418,N_29439);
xor UO_1797 (O_1797,N_29965,N_29994);
nor UO_1798 (O_1798,N_29706,N_29416);
xnor UO_1799 (O_1799,N_29935,N_29922);
or UO_1800 (O_1800,N_29896,N_29881);
and UO_1801 (O_1801,N_29914,N_29476);
nor UO_1802 (O_1802,N_29492,N_29756);
xor UO_1803 (O_1803,N_29476,N_29986);
or UO_1804 (O_1804,N_29821,N_29627);
xnor UO_1805 (O_1805,N_29712,N_29450);
xor UO_1806 (O_1806,N_29884,N_29938);
and UO_1807 (O_1807,N_29461,N_29902);
nor UO_1808 (O_1808,N_29541,N_29410);
xnor UO_1809 (O_1809,N_29641,N_29733);
nor UO_1810 (O_1810,N_29436,N_29640);
or UO_1811 (O_1811,N_29552,N_29962);
nand UO_1812 (O_1812,N_29862,N_29663);
nand UO_1813 (O_1813,N_29765,N_29554);
xor UO_1814 (O_1814,N_29514,N_29814);
and UO_1815 (O_1815,N_29878,N_29691);
nand UO_1816 (O_1816,N_29590,N_29451);
nand UO_1817 (O_1817,N_29544,N_29462);
nor UO_1818 (O_1818,N_29650,N_29445);
nand UO_1819 (O_1819,N_29617,N_29586);
or UO_1820 (O_1820,N_29987,N_29410);
and UO_1821 (O_1821,N_29755,N_29601);
or UO_1822 (O_1822,N_29830,N_29856);
nor UO_1823 (O_1823,N_29678,N_29855);
nor UO_1824 (O_1824,N_29638,N_29440);
nand UO_1825 (O_1825,N_29697,N_29520);
nor UO_1826 (O_1826,N_29838,N_29644);
or UO_1827 (O_1827,N_29873,N_29409);
or UO_1828 (O_1828,N_29612,N_29910);
and UO_1829 (O_1829,N_29956,N_29611);
nand UO_1830 (O_1830,N_29936,N_29826);
nand UO_1831 (O_1831,N_29838,N_29470);
nand UO_1832 (O_1832,N_29871,N_29923);
xnor UO_1833 (O_1833,N_29933,N_29984);
nor UO_1834 (O_1834,N_29446,N_29713);
nor UO_1835 (O_1835,N_29476,N_29993);
and UO_1836 (O_1836,N_29571,N_29722);
or UO_1837 (O_1837,N_29785,N_29870);
xnor UO_1838 (O_1838,N_29900,N_29680);
nand UO_1839 (O_1839,N_29595,N_29766);
and UO_1840 (O_1840,N_29412,N_29874);
or UO_1841 (O_1841,N_29861,N_29878);
nand UO_1842 (O_1842,N_29813,N_29783);
nor UO_1843 (O_1843,N_29957,N_29949);
xnor UO_1844 (O_1844,N_29529,N_29446);
nor UO_1845 (O_1845,N_29860,N_29607);
nor UO_1846 (O_1846,N_29789,N_29674);
xor UO_1847 (O_1847,N_29668,N_29757);
and UO_1848 (O_1848,N_29784,N_29464);
xnor UO_1849 (O_1849,N_29870,N_29647);
nor UO_1850 (O_1850,N_29453,N_29638);
nand UO_1851 (O_1851,N_29933,N_29605);
and UO_1852 (O_1852,N_29584,N_29937);
and UO_1853 (O_1853,N_29902,N_29867);
or UO_1854 (O_1854,N_29629,N_29798);
or UO_1855 (O_1855,N_29676,N_29823);
xnor UO_1856 (O_1856,N_29988,N_29412);
nand UO_1857 (O_1857,N_29821,N_29411);
or UO_1858 (O_1858,N_29929,N_29940);
nor UO_1859 (O_1859,N_29691,N_29612);
nand UO_1860 (O_1860,N_29665,N_29956);
xnor UO_1861 (O_1861,N_29782,N_29760);
nand UO_1862 (O_1862,N_29759,N_29819);
nand UO_1863 (O_1863,N_29935,N_29455);
nor UO_1864 (O_1864,N_29897,N_29603);
nand UO_1865 (O_1865,N_29942,N_29448);
xnor UO_1866 (O_1866,N_29552,N_29933);
or UO_1867 (O_1867,N_29810,N_29860);
xnor UO_1868 (O_1868,N_29907,N_29931);
nand UO_1869 (O_1869,N_29704,N_29627);
xnor UO_1870 (O_1870,N_29985,N_29872);
and UO_1871 (O_1871,N_29674,N_29898);
xor UO_1872 (O_1872,N_29939,N_29650);
and UO_1873 (O_1873,N_29919,N_29578);
or UO_1874 (O_1874,N_29413,N_29758);
nand UO_1875 (O_1875,N_29860,N_29925);
nand UO_1876 (O_1876,N_29581,N_29726);
or UO_1877 (O_1877,N_29619,N_29510);
nand UO_1878 (O_1878,N_29544,N_29433);
nor UO_1879 (O_1879,N_29447,N_29454);
nand UO_1880 (O_1880,N_29792,N_29588);
xor UO_1881 (O_1881,N_29933,N_29491);
or UO_1882 (O_1882,N_29620,N_29897);
or UO_1883 (O_1883,N_29897,N_29854);
and UO_1884 (O_1884,N_29587,N_29803);
or UO_1885 (O_1885,N_29410,N_29698);
nand UO_1886 (O_1886,N_29898,N_29500);
nor UO_1887 (O_1887,N_29966,N_29619);
nand UO_1888 (O_1888,N_29890,N_29974);
nand UO_1889 (O_1889,N_29715,N_29975);
xnor UO_1890 (O_1890,N_29970,N_29873);
nor UO_1891 (O_1891,N_29658,N_29897);
or UO_1892 (O_1892,N_29883,N_29571);
nand UO_1893 (O_1893,N_29966,N_29611);
or UO_1894 (O_1894,N_29461,N_29939);
nand UO_1895 (O_1895,N_29531,N_29813);
and UO_1896 (O_1896,N_29512,N_29666);
nor UO_1897 (O_1897,N_29532,N_29442);
or UO_1898 (O_1898,N_29458,N_29799);
nor UO_1899 (O_1899,N_29567,N_29797);
xor UO_1900 (O_1900,N_29909,N_29924);
xnor UO_1901 (O_1901,N_29493,N_29697);
nand UO_1902 (O_1902,N_29488,N_29472);
nand UO_1903 (O_1903,N_29513,N_29566);
or UO_1904 (O_1904,N_29793,N_29747);
xor UO_1905 (O_1905,N_29822,N_29713);
xnor UO_1906 (O_1906,N_29978,N_29588);
nand UO_1907 (O_1907,N_29885,N_29870);
nand UO_1908 (O_1908,N_29513,N_29975);
or UO_1909 (O_1909,N_29480,N_29953);
nand UO_1910 (O_1910,N_29954,N_29933);
and UO_1911 (O_1911,N_29766,N_29739);
xnor UO_1912 (O_1912,N_29867,N_29478);
or UO_1913 (O_1913,N_29867,N_29594);
or UO_1914 (O_1914,N_29713,N_29487);
or UO_1915 (O_1915,N_29536,N_29731);
or UO_1916 (O_1916,N_29540,N_29848);
nand UO_1917 (O_1917,N_29423,N_29817);
nor UO_1918 (O_1918,N_29461,N_29759);
nand UO_1919 (O_1919,N_29675,N_29571);
xor UO_1920 (O_1920,N_29863,N_29705);
or UO_1921 (O_1921,N_29465,N_29643);
nor UO_1922 (O_1922,N_29969,N_29605);
nand UO_1923 (O_1923,N_29712,N_29673);
nand UO_1924 (O_1924,N_29909,N_29969);
or UO_1925 (O_1925,N_29408,N_29727);
nor UO_1926 (O_1926,N_29561,N_29911);
or UO_1927 (O_1927,N_29879,N_29440);
nand UO_1928 (O_1928,N_29909,N_29627);
or UO_1929 (O_1929,N_29890,N_29846);
nand UO_1930 (O_1930,N_29866,N_29569);
nand UO_1931 (O_1931,N_29632,N_29778);
xnor UO_1932 (O_1932,N_29622,N_29460);
nand UO_1933 (O_1933,N_29966,N_29836);
nand UO_1934 (O_1934,N_29810,N_29820);
and UO_1935 (O_1935,N_29665,N_29942);
and UO_1936 (O_1936,N_29509,N_29549);
and UO_1937 (O_1937,N_29886,N_29440);
nor UO_1938 (O_1938,N_29878,N_29414);
xor UO_1939 (O_1939,N_29439,N_29700);
xor UO_1940 (O_1940,N_29604,N_29868);
xor UO_1941 (O_1941,N_29910,N_29922);
nor UO_1942 (O_1942,N_29913,N_29606);
xor UO_1943 (O_1943,N_29852,N_29575);
xnor UO_1944 (O_1944,N_29832,N_29422);
and UO_1945 (O_1945,N_29758,N_29916);
xor UO_1946 (O_1946,N_29624,N_29861);
and UO_1947 (O_1947,N_29429,N_29423);
xnor UO_1948 (O_1948,N_29613,N_29565);
nand UO_1949 (O_1949,N_29400,N_29845);
and UO_1950 (O_1950,N_29553,N_29418);
nand UO_1951 (O_1951,N_29608,N_29647);
and UO_1952 (O_1952,N_29990,N_29956);
nand UO_1953 (O_1953,N_29491,N_29410);
and UO_1954 (O_1954,N_29524,N_29651);
nand UO_1955 (O_1955,N_29839,N_29953);
or UO_1956 (O_1956,N_29947,N_29636);
xor UO_1957 (O_1957,N_29910,N_29672);
and UO_1958 (O_1958,N_29443,N_29886);
nand UO_1959 (O_1959,N_29900,N_29862);
nor UO_1960 (O_1960,N_29682,N_29851);
or UO_1961 (O_1961,N_29841,N_29732);
and UO_1962 (O_1962,N_29797,N_29802);
xnor UO_1963 (O_1963,N_29882,N_29532);
and UO_1964 (O_1964,N_29666,N_29788);
nor UO_1965 (O_1965,N_29754,N_29512);
nand UO_1966 (O_1966,N_29620,N_29434);
nand UO_1967 (O_1967,N_29852,N_29838);
nand UO_1968 (O_1968,N_29431,N_29425);
or UO_1969 (O_1969,N_29679,N_29788);
or UO_1970 (O_1970,N_29485,N_29447);
and UO_1971 (O_1971,N_29543,N_29993);
or UO_1972 (O_1972,N_29873,N_29407);
or UO_1973 (O_1973,N_29520,N_29582);
and UO_1974 (O_1974,N_29838,N_29630);
and UO_1975 (O_1975,N_29530,N_29691);
nor UO_1976 (O_1976,N_29836,N_29697);
or UO_1977 (O_1977,N_29720,N_29948);
nor UO_1978 (O_1978,N_29788,N_29951);
xor UO_1979 (O_1979,N_29627,N_29810);
nor UO_1980 (O_1980,N_29431,N_29814);
and UO_1981 (O_1981,N_29547,N_29498);
and UO_1982 (O_1982,N_29979,N_29448);
xor UO_1983 (O_1983,N_29985,N_29705);
or UO_1984 (O_1984,N_29639,N_29922);
nor UO_1985 (O_1985,N_29911,N_29691);
xnor UO_1986 (O_1986,N_29729,N_29920);
nor UO_1987 (O_1987,N_29706,N_29599);
or UO_1988 (O_1988,N_29786,N_29916);
and UO_1989 (O_1989,N_29599,N_29924);
xor UO_1990 (O_1990,N_29873,N_29908);
xor UO_1991 (O_1991,N_29458,N_29693);
nand UO_1992 (O_1992,N_29660,N_29452);
and UO_1993 (O_1993,N_29757,N_29955);
nor UO_1994 (O_1994,N_29955,N_29745);
nand UO_1995 (O_1995,N_29937,N_29749);
or UO_1996 (O_1996,N_29855,N_29914);
nor UO_1997 (O_1997,N_29529,N_29560);
or UO_1998 (O_1998,N_29741,N_29918);
nand UO_1999 (O_1999,N_29705,N_29658);
nand UO_2000 (O_2000,N_29733,N_29660);
nand UO_2001 (O_2001,N_29434,N_29751);
xnor UO_2002 (O_2002,N_29582,N_29810);
nor UO_2003 (O_2003,N_29466,N_29456);
nor UO_2004 (O_2004,N_29569,N_29814);
nand UO_2005 (O_2005,N_29537,N_29714);
xnor UO_2006 (O_2006,N_29781,N_29625);
nand UO_2007 (O_2007,N_29587,N_29941);
xor UO_2008 (O_2008,N_29708,N_29647);
nor UO_2009 (O_2009,N_29978,N_29744);
xnor UO_2010 (O_2010,N_29901,N_29617);
nor UO_2011 (O_2011,N_29982,N_29776);
xor UO_2012 (O_2012,N_29421,N_29969);
and UO_2013 (O_2013,N_29778,N_29630);
nand UO_2014 (O_2014,N_29800,N_29687);
xnor UO_2015 (O_2015,N_29422,N_29649);
and UO_2016 (O_2016,N_29787,N_29718);
xnor UO_2017 (O_2017,N_29487,N_29705);
or UO_2018 (O_2018,N_29446,N_29565);
or UO_2019 (O_2019,N_29910,N_29739);
nand UO_2020 (O_2020,N_29745,N_29587);
xor UO_2021 (O_2021,N_29843,N_29670);
nand UO_2022 (O_2022,N_29515,N_29877);
xnor UO_2023 (O_2023,N_29685,N_29891);
or UO_2024 (O_2024,N_29934,N_29401);
or UO_2025 (O_2025,N_29543,N_29823);
nand UO_2026 (O_2026,N_29414,N_29692);
and UO_2027 (O_2027,N_29645,N_29763);
nor UO_2028 (O_2028,N_29873,N_29901);
or UO_2029 (O_2029,N_29550,N_29417);
nor UO_2030 (O_2030,N_29677,N_29523);
and UO_2031 (O_2031,N_29418,N_29440);
nor UO_2032 (O_2032,N_29641,N_29486);
and UO_2033 (O_2033,N_29993,N_29657);
and UO_2034 (O_2034,N_29559,N_29745);
nand UO_2035 (O_2035,N_29408,N_29904);
nand UO_2036 (O_2036,N_29774,N_29419);
or UO_2037 (O_2037,N_29858,N_29465);
xnor UO_2038 (O_2038,N_29898,N_29633);
or UO_2039 (O_2039,N_29563,N_29433);
and UO_2040 (O_2040,N_29795,N_29447);
xnor UO_2041 (O_2041,N_29573,N_29681);
or UO_2042 (O_2042,N_29461,N_29830);
xor UO_2043 (O_2043,N_29687,N_29700);
or UO_2044 (O_2044,N_29474,N_29637);
nor UO_2045 (O_2045,N_29510,N_29809);
nand UO_2046 (O_2046,N_29666,N_29400);
nor UO_2047 (O_2047,N_29833,N_29653);
and UO_2048 (O_2048,N_29696,N_29740);
nand UO_2049 (O_2049,N_29482,N_29868);
xnor UO_2050 (O_2050,N_29876,N_29976);
nor UO_2051 (O_2051,N_29488,N_29700);
or UO_2052 (O_2052,N_29576,N_29463);
xor UO_2053 (O_2053,N_29597,N_29580);
and UO_2054 (O_2054,N_29591,N_29658);
or UO_2055 (O_2055,N_29535,N_29679);
or UO_2056 (O_2056,N_29542,N_29488);
or UO_2057 (O_2057,N_29936,N_29560);
and UO_2058 (O_2058,N_29590,N_29901);
nor UO_2059 (O_2059,N_29549,N_29914);
nand UO_2060 (O_2060,N_29493,N_29634);
and UO_2061 (O_2061,N_29647,N_29625);
xor UO_2062 (O_2062,N_29526,N_29841);
or UO_2063 (O_2063,N_29511,N_29535);
or UO_2064 (O_2064,N_29849,N_29642);
nor UO_2065 (O_2065,N_29620,N_29995);
and UO_2066 (O_2066,N_29888,N_29818);
xor UO_2067 (O_2067,N_29780,N_29785);
or UO_2068 (O_2068,N_29809,N_29656);
nand UO_2069 (O_2069,N_29889,N_29425);
xnor UO_2070 (O_2070,N_29971,N_29446);
nor UO_2071 (O_2071,N_29648,N_29421);
nor UO_2072 (O_2072,N_29520,N_29719);
nand UO_2073 (O_2073,N_29927,N_29509);
nand UO_2074 (O_2074,N_29735,N_29561);
nand UO_2075 (O_2075,N_29588,N_29694);
nor UO_2076 (O_2076,N_29799,N_29801);
and UO_2077 (O_2077,N_29789,N_29988);
or UO_2078 (O_2078,N_29568,N_29711);
or UO_2079 (O_2079,N_29560,N_29600);
nand UO_2080 (O_2080,N_29561,N_29775);
nand UO_2081 (O_2081,N_29857,N_29821);
or UO_2082 (O_2082,N_29596,N_29985);
xor UO_2083 (O_2083,N_29784,N_29858);
xnor UO_2084 (O_2084,N_29422,N_29770);
xnor UO_2085 (O_2085,N_29691,N_29517);
and UO_2086 (O_2086,N_29963,N_29823);
and UO_2087 (O_2087,N_29584,N_29766);
and UO_2088 (O_2088,N_29418,N_29517);
nand UO_2089 (O_2089,N_29514,N_29998);
xnor UO_2090 (O_2090,N_29632,N_29575);
or UO_2091 (O_2091,N_29457,N_29704);
xnor UO_2092 (O_2092,N_29933,N_29736);
nand UO_2093 (O_2093,N_29822,N_29483);
nor UO_2094 (O_2094,N_29556,N_29934);
and UO_2095 (O_2095,N_29889,N_29980);
or UO_2096 (O_2096,N_29450,N_29404);
and UO_2097 (O_2097,N_29639,N_29417);
nand UO_2098 (O_2098,N_29874,N_29877);
nand UO_2099 (O_2099,N_29604,N_29797);
or UO_2100 (O_2100,N_29937,N_29700);
xnor UO_2101 (O_2101,N_29463,N_29457);
nand UO_2102 (O_2102,N_29928,N_29463);
nor UO_2103 (O_2103,N_29595,N_29844);
nor UO_2104 (O_2104,N_29464,N_29818);
xor UO_2105 (O_2105,N_29771,N_29645);
nand UO_2106 (O_2106,N_29670,N_29471);
nor UO_2107 (O_2107,N_29679,N_29638);
xor UO_2108 (O_2108,N_29601,N_29669);
and UO_2109 (O_2109,N_29641,N_29625);
and UO_2110 (O_2110,N_29798,N_29719);
nand UO_2111 (O_2111,N_29891,N_29734);
nand UO_2112 (O_2112,N_29631,N_29738);
nand UO_2113 (O_2113,N_29726,N_29536);
nand UO_2114 (O_2114,N_29988,N_29554);
nand UO_2115 (O_2115,N_29721,N_29627);
or UO_2116 (O_2116,N_29744,N_29820);
or UO_2117 (O_2117,N_29403,N_29661);
nor UO_2118 (O_2118,N_29560,N_29588);
nand UO_2119 (O_2119,N_29969,N_29902);
and UO_2120 (O_2120,N_29947,N_29492);
or UO_2121 (O_2121,N_29999,N_29708);
xnor UO_2122 (O_2122,N_29720,N_29878);
or UO_2123 (O_2123,N_29677,N_29753);
and UO_2124 (O_2124,N_29557,N_29745);
nand UO_2125 (O_2125,N_29641,N_29934);
nand UO_2126 (O_2126,N_29716,N_29700);
and UO_2127 (O_2127,N_29869,N_29672);
xor UO_2128 (O_2128,N_29400,N_29435);
nor UO_2129 (O_2129,N_29515,N_29597);
or UO_2130 (O_2130,N_29975,N_29697);
or UO_2131 (O_2131,N_29627,N_29797);
xnor UO_2132 (O_2132,N_29663,N_29547);
or UO_2133 (O_2133,N_29653,N_29646);
or UO_2134 (O_2134,N_29407,N_29631);
or UO_2135 (O_2135,N_29799,N_29645);
nand UO_2136 (O_2136,N_29478,N_29499);
xnor UO_2137 (O_2137,N_29631,N_29869);
xnor UO_2138 (O_2138,N_29495,N_29884);
or UO_2139 (O_2139,N_29751,N_29629);
nand UO_2140 (O_2140,N_29471,N_29795);
xnor UO_2141 (O_2141,N_29541,N_29758);
xor UO_2142 (O_2142,N_29559,N_29681);
or UO_2143 (O_2143,N_29676,N_29478);
and UO_2144 (O_2144,N_29523,N_29899);
xnor UO_2145 (O_2145,N_29459,N_29608);
or UO_2146 (O_2146,N_29877,N_29726);
xor UO_2147 (O_2147,N_29969,N_29643);
nor UO_2148 (O_2148,N_29592,N_29851);
xor UO_2149 (O_2149,N_29971,N_29984);
nor UO_2150 (O_2150,N_29595,N_29760);
nor UO_2151 (O_2151,N_29461,N_29464);
nor UO_2152 (O_2152,N_29896,N_29613);
or UO_2153 (O_2153,N_29677,N_29557);
nor UO_2154 (O_2154,N_29451,N_29931);
or UO_2155 (O_2155,N_29455,N_29721);
nand UO_2156 (O_2156,N_29905,N_29633);
nand UO_2157 (O_2157,N_29952,N_29441);
nand UO_2158 (O_2158,N_29617,N_29967);
xor UO_2159 (O_2159,N_29626,N_29700);
nand UO_2160 (O_2160,N_29679,N_29706);
nor UO_2161 (O_2161,N_29503,N_29512);
xor UO_2162 (O_2162,N_29509,N_29767);
xnor UO_2163 (O_2163,N_29702,N_29679);
and UO_2164 (O_2164,N_29976,N_29897);
nor UO_2165 (O_2165,N_29725,N_29885);
xnor UO_2166 (O_2166,N_29451,N_29547);
and UO_2167 (O_2167,N_29743,N_29677);
nand UO_2168 (O_2168,N_29915,N_29513);
or UO_2169 (O_2169,N_29483,N_29554);
xor UO_2170 (O_2170,N_29890,N_29487);
xor UO_2171 (O_2171,N_29684,N_29897);
nand UO_2172 (O_2172,N_29544,N_29710);
or UO_2173 (O_2173,N_29929,N_29693);
and UO_2174 (O_2174,N_29655,N_29572);
nand UO_2175 (O_2175,N_29572,N_29576);
or UO_2176 (O_2176,N_29516,N_29812);
nor UO_2177 (O_2177,N_29939,N_29486);
or UO_2178 (O_2178,N_29976,N_29960);
nor UO_2179 (O_2179,N_29521,N_29814);
and UO_2180 (O_2180,N_29497,N_29716);
and UO_2181 (O_2181,N_29714,N_29782);
or UO_2182 (O_2182,N_29620,N_29976);
and UO_2183 (O_2183,N_29884,N_29693);
xnor UO_2184 (O_2184,N_29847,N_29983);
nand UO_2185 (O_2185,N_29660,N_29746);
nor UO_2186 (O_2186,N_29593,N_29704);
and UO_2187 (O_2187,N_29628,N_29615);
nor UO_2188 (O_2188,N_29674,N_29669);
xor UO_2189 (O_2189,N_29743,N_29759);
nand UO_2190 (O_2190,N_29665,N_29521);
xnor UO_2191 (O_2191,N_29667,N_29556);
nand UO_2192 (O_2192,N_29898,N_29904);
xor UO_2193 (O_2193,N_29997,N_29945);
xnor UO_2194 (O_2194,N_29786,N_29918);
nor UO_2195 (O_2195,N_29470,N_29789);
or UO_2196 (O_2196,N_29806,N_29655);
and UO_2197 (O_2197,N_29409,N_29472);
or UO_2198 (O_2198,N_29550,N_29924);
and UO_2199 (O_2199,N_29816,N_29837);
nand UO_2200 (O_2200,N_29688,N_29577);
and UO_2201 (O_2201,N_29643,N_29893);
or UO_2202 (O_2202,N_29478,N_29943);
nand UO_2203 (O_2203,N_29628,N_29569);
and UO_2204 (O_2204,N_29541,N_29588);
nor UO_2205 (O_2205,N_29673,N_29550);
and UO_2206 (O_2206,N_29452,N_29622);
or UO_2207 (O_2207,N_29690,N_29435);
nor UO_2208 (O_2208,N_29717,N_29843);
and UO_2209 (O_2209,N_29731,N_29771);
xnor UO_2210 (O_2210,N_29403,N_29708);
xnor UO_2211 (O_2211,N_29442,N_29481);
nor UO_2212 (O_2212,N_29947,N_29408);
nor UO_2213 (O_2213,N_29593,N_29980);
and UO_2214 (O_2214,N_29861,N_29687);
nand UO_2215 (O_2215,N_29689,N_29782);
and UO_2216 (O_2216,N_29841,N_29842);
nor UO_2217 (O_2217,N_29658,N_29503);
nor UO_2218 (O_2218,N_29758,N_29594);
nand UO_2219 (O_2219,N_29598,N_29799);
nor UO_2220 (O_2220,N_29521,N_29799);
and UO_2221 (O_2221,N_29699,N_29869);
nor UO_2222 (O_2222,N_29802,N_29962);
or UO_2223 (O_2223,N_29841,N_29998);
or UO_2224 (O_2224,N_29597,N_29728);
xor UO_2225 (O_2225,N_29420,N_29786);
and UO_2226 (O_2226,N_29837,N_29582);
nand UO_2227 (O_2227,N_29970,N_29699);
nand UO_2228 (O_2228,N_29788,N_29590);
nand UO_2229 (O_2229,N_29956,N_29520);
and UO_2230 (O_2230,N_29650,N_29461);
nor UO_2231 (O_2231,N_29629,N_29607);
nand UO_2232 (O_2232,N_29601,N_29589);
and UO_2233 (O_2233,N_29441,N_29970);
nor UO_2234 (O_2234,N_29495,N_29455);
nor UO_2235 (O_2235,N_29965,N_29547);
nor UO_2236 (O_2236,N_29485,N_29784);
nand UO_2237 (O_2237,N_29527,N_29468);
xnor UO_2238 (O_2238,N_29724,N_29997);
or UO_2239 (O_2239,N_29838,N_29646);
xnor UO_2240 (O_2240,N_29976,N_29482);
xor UO_2241 (O_2241,N_29407,N_29627);
xnor UO_2242 (O_2242,N_29548,N_29552);
and UO_2243 (O_2243,N_29818,N_29627);
or UO_2244 (O_2244,N_29831,N_29710);
xnor UO_2245 (O_2245,N_29992,N_29429);
xnor UO_2246 (O_2246,N_29569,N_29994);
and UO_2247 (O_2247,N_29841,N_29420);
and UO_2248 (O_2248,N_29675,N_29676);
and UO_2249 (O_2249,N_29658,N_29796);
nor UO_2250 (O_2250,N_29753,N_29800);
or UO_2251 (O_2251,N_29992,N_29780);
nor UO_2252 (O_2252,N_29586,N_29433);
nand UO_2253 (O_2253,N_29874,N_29640);
nand UO_2254 (O_2254,N_29518,N_29855);
nor UO_2255 (O_2255,N_29593,N_29410);
xor UO_2256 (O_2256,N_29634,N_29815);
nand UO_2257 (O_2257,N_29426,N_29994);
xor UO_2258 (O_2258,N_29745,N_29549);
xor UO_2259 (O_2259,N_29903,N_29826);
nand UO_2260 (O_2260,N_29491,N_29885);
or UO_2261 (O_2261,N_29487,N_29931);
and UO_2262 (O_2262,N_29917,N_29578);
and UO_2263 (O_2263,N_29408,N_29937);
xor UO_2264 (O_2264,N_29604,N_29738);
nor UO_2265 (O_2265,N_29898,N_29678);
nor UO_2266 (O_2266,N_29688,N_29524);
xor UO_2267 (O_2267,N_29585,N_29549);
or UO_2268 (O_2268,N_29478,N_29528);
nand UO_2269 (O_2269,N_29757,N_29658);
xor UO_2270 (O_2270,N_29528,N_29436);
or UO_2271 (O_2271,N_29725,N_29908);
nand UO_2272 (O_2272,N_29971,N_29677);
or UO_2273 (O_2273,N_29536,N_29550);
nand UO_2274 (O_2274,N_29970,N_29773);
xor UO_2275 (O_2275,N_29674,N_29762);
nand UO_2276 (O_2276,N_29675,N_29450);
or UO_2277 (O_2277,N_29943,N_29798);
or UO_2278 (O_2278,N_29931,N_29923);
xnor UO_2279 (O_2279,N_29500,N_29762);
nand UO_2280 (O_2280,N_29589,N_29844);
nand UO_2281 (O_2281,N_29622,N_29786);
xnor UO_2282 (O_2282,N_29757,N_29787);
or UO_2283 (O_2283,N_29693,N_29474);
xor UO_2284 (O_2284,N_29779,N_29565);
and UO_2285 (O_2285,N_29514,N_29408);
and UO_2286 (O_2286,N_29407,N_29892);
xor UO_2287 (O_2287,N_29858,N_29416);
and UO_2288 (O_2288,N_29530,N_29470);
nor UO_2289 (O_2289,N_29434,N_29441);
and UO_2290 (O_2290,N_29568,N_29962);
nand UO_2291 (O_2291,N_29426,N_29476);
xnor UO_2292 (O_2292,N_29628,N_29681);
or UO_2293 (O_2293,N_29580,N_29593);
xnor UO_2294 (O_2294,N_29605,N_29815);
xnor UO_2295 (O_2295,N_29604,N_29908);
and UO_2296 (O_2296,N_29824,N_29891);
nor UO_2297 (O_2297,N_29752,N_29960);
and UO_2298 (O_2298,N_29863,N_29953);
nand UO_2299 (O_2299,N_29958,N_29770);
and UO_2300 (O_2300,N_29567,N_29457);
or UO_2301 (O_2301,N_29632,N_29987);
or UO_2302 (O_2302,N_29590,N_29467);
or UO_2303 (O_2303,N_29935,N_29587);
or UO_2304 (O_2304,N_29508,N_29502);
or UO_2305 (O_2305,N_29405,N_29857);
xor UO_2306 (O_2306,N_29568,N_29961);
xnor UO_2307 (O_2307,N_29969,N_29670);
xor UO_2308 (O_2308,N_29930,N_29892);
or UO_2309 (O_2309,N_29467,N_29769);
xor UO_2310 (O_2310,N_29610,N_29683);
nand UO_2311 (O_2311,N_29448,N_29841);
xnor UO_2312 (O_2312,N_29605,N_29720);
nor UO_2313 (O_2313,N_29555,N_29722);
and UO_2314 (O_2314,N_29827,N_29924);
xnor UO_2315 (O_2315,N_29539,N_29593);
or UO_2316 (O_2316,N_29986,N_29791);
or UO_2317 (O_2317,N_29415,N_29410);
nor UO_2318 (O_2318,N_29881,N_29474);
and UO_2319 (O_2319,N_29998,N_29945);
nand UO_2320 (O_2320,N_29757,N_29547);
nand UO_2321 (O_2321,N_29732,N_29549);
or UO_2322 (O_2322,N_29602,N_29920);
nand UO_2323 (O_2323,N_29839,N_29861);
xor UO_2324 (O_2324,N_29619,N_29733);
xnor UO_2325 (O_2325,N_29779,N_29851);
and UO_2326 (O_2326,N_29942,N_29687);
and UO_2327 (O_2327,N_29614,N_29913);
and UO_2328 (O_2328,N_29810,N_29475);
or UO_2329 (O_2329,N_29636,N_29583);
xnor UO_2330 (O_2330,N_29886,N_29974);
or UO_2331 (O_2331,N_29834,N_29844);
nand UO_2332 (O_2332,N_29457,N_29937);
xor UO_2333 (O_2333,N_29616,N_29405);
nor UO_2334 (O_2334,N_29440,N_29475);
and UO_2335 (O_2335,N_29722,N_29502);
nand UO_2336 (O_2336,N_29506,N_29915);
nor UO_2337 (O_2337,N_29897,N_29847);
xor UO_2338 (O_2338,N_29811,N_29826);
nor UO_2339 (O_2339,N_29521,N_29612);
or UO_2340 (O_2340,N_29489,N_29586);
xnor UO_2341 (O_2341,N_29945,N_29488);
and UO_2342 (O_2342,N_29651,N_29976);
nand UO_2343 (O_2343,N_29793,N_29638);
and UO_2344 (O_2344,N_29695,N_29683);
or UO_2345 (O_2345,N_29645,N_29811);
xnor UO_2346 (O_2346,N_29691,N_29881);
or UO_2347 (O_2347,N_29463,N_29529);
nor UO_2348 (O_2348,N_29432,N_29438);
nand UO_2349 (O_2349,N_29896,N_29423);
nand UO_2350 (O_2350,N_29568,N_29645);
xnor UO_2351 (O_2351,N_29871,N_29810);
or UO_2352 (O_2352,N_29641,N_29913);
and UO_2353 (O_2353,N_29483,N_29400);
nor UO_2354 (O_2354,N_29970,N_29453);
or UO_2355 (O_2355,N_29887,N_29981);
xnor UO_2356 (O_2356,N_29892,N_29532);
xor UO_2357 (O_2357,N_29618,N_29878);
xor UO_2358 (O_2358,N_29736,N_29568);
xnor UO_2359 (O_2359,N_29638,N_29438);
or UO_2360 (O_2360,N_29972,N_29977);
nor UO_2361 (O_2361,N_29541,N_29565);
xor UO_2362 (O_2362,N_29609,N_29639);
xnor UO_2363 (O_2363,N_29639,N_29833);
nand UO_2364 (O_2364,N_29486,N_29703);
xnor UO_2365 (O_2365,N_29771,N_29759);
nor UO_2366 (O_2366,N_29610,N_29613);
and UO_2367 (O_2367,N_29543,N_29687);
or UO_2368 (O_2368,N_29925,N_29724);
nor UO_2369 (O_2369,N_29405,N_29975);
and UO_2370 (O_2370,N_29734,N_29631);
xor UO_2371 (O_2371,N_29711,N_29887);
nand UO_2372 (O_2372,N_29537,N_29587);
xor UO_2373 (O_2373,N_29749,N_29547);
nor UO_2374 (O_2374,N_29811,N_29951);
or UO_2375 (O_2375,N_29453,N_29460);
nand UO_2376 (O_2376,N_29739,N_29612);
xor UO_2377 (O_2377,N_29975,N_29732);
and UO_2378 (O_2378,N_29693,N_29967);
and UO_2379 (O_2379,N_29929,N_29894);
and UO_2380 (O_2380,N_29524,N_29783);
xor UO_2381 (O_2381,N_29476,N_29960);
nand UO_2382 (O_2382,N_29981,N_29697);
or UO_2383 (O_2383,N_29991,N_29587);
and UO_2384 (O_2384,N_29983,N_29720);
or UO_2385 (O_2385,N_29614,N_29584);
and UO_2386 (O_2386,N_29622,N_29428);
nand UO_2387 (O_2387,N_29642,N_29775);
nand UO_2388 (O_2388,N_29587,N_29809);
and UO_2389 (O_2389,N_29845,N_29593);
xor UO_2390 (O_2390,N_29406,N_29461);
nor UO_2391 (O_2391,N_29674,N_29455);
and UO_2392 (O_2392,N_29848,N_29946);
nor UO_2393 (O_2393,N_29724,N_29538);
nor UO_2394 (O_2394,N_29449,N_29567);
or UO_2395 (O_2395,N_29854,N_29678);
and UO_2396 (O_2396,N_29446,N_29856);
nor UO_2397 (O_2397,N_29836,N_29575);
nand UO_2398 (O_2398,N_29664,N_29852);
xor UO_2399 (O_2399,N_29792,N_29491);
or UO_2400 (O_2400,N_29577,N_29906);
or UO_2401 (O_2401,N_29985,N_29741);
xnor UO_2402 (O_2402,N_29849,N_29788);
xnor UO_2403 (O_2403,N_29932,N_29915);
nor UO_2404 (O_2404,N_29956,N_29696);
xnor UO_2405 (O_2405,N_29579,N_29760);
nand UO_2406 (O_2406,N_29757,N_29979);
and UO_2407 (O_2407,N_29601,N_29865);
and UO_2408 (O_2408,N_29787,N_29465);
or UO_2409 (O_2409,N_29755,N_29756);
nor UO_2410 (O_2410,N_29789,N_29415);
xor UO_2411 (O_2411,N_29468,N_29954);
nor UO_2412 (O_2412,N_29633,N_29516);
and UO_2413 (O_2413,N_29811,N_29721);
or UO_2414 (O_2414,N_29568,N_29407);
or UO_2415 (O_2415,N_29756,N_29414);
nand UO_2416 (O_2416,N_29467,N_29582);
or UO_2417 (O_2417,N_29674,N_29900);
nand UO_2418 (O_2418,N_29418,N_29678);
xor UO_2419 (O_2419,N_29656,N_29684);
nand UO_2420 (O_2420,N_29898,N_29947);
nor UO_2421 (O_2421,N_29997,N_29904);
or UO_2422 (O_2422,N_29925,N_29499);
xor UO_2423 (O_2423,N_29583,N_29422);
nor UO_2424 (O_2424,N_29814,N_29861);
nand UO_2425 (O_2425,N_29516,N_29885);
and UO_2426 (O_2426,N_29665,N_29697);
nand UO_2427 (O_2427,N_29472,N_29751);
nor UO_2428 (O_2428,N_29791,N_29489);
and UO_2429 (O_2429,N_29637,N_29708);
and UO_2430 (O_2430,N_29839,N_29503);
or UO_2431 (O_2431,N_29885,N_29609);
xor UO_2432 (O_2432,N_29797,N_29839);
nand UO_2433 (O_2433,N_29428,N_29607);
xnor UO_2434 (O_2434,N_29646,N_29883);
nand UO_2435 (O_2435,N_29605,N_29489);
xor UO_2436 (O_2436,N_29671,N_29540);
or UO_2437 (O_2437,N_29744,N_29794);
nand UO_2438 (O_2438,N_29493,N_29703);
xnor UO_2439 (O_2439,N_29495,N_29832);
nand UO_2440 (O_2440,N_29487,N_29446);
xor UO_2441 (O_2441,N_29447,N_29677);
and UO_2442 (O_2442,N_29557,N_29959);
nor UO_2443 (O_2443,N_29863,N_29591);
and UO_2444 (O_2444,N_29847,N_29544);
or UO_2445 (O_2445,N_29873,N_29953);
or UO_2446 (O_2446,N_29962,N_29837);
xor UO_2447 (O_2447,N_29502,N_29963);
xor UO_2448 (O_2448,N_29479,N_29569);
nor UO_2449 (O_2449,N_29481,N_29889);
nor UO_2450 (O_2450,N_29972,N_29746);
xnor UO_2451 (O_2451,N_29627,N_29520);
nor UO_2452 (O_2452,N_29421,N_29667);
and UO_2453 (O_2453,N_29798,N_29757);
or UO_2454 (O_2454,N_29907,N_29930);
xnor UO_2455 (O_2455,N_29787,N_29845);
nand UO_2456 (O_2456,N_29963,N_29704);
xnor UO_2457 (O_2457,N_29782,N_29641);
nor UO_2458 (O_2458,N_29863,N_29534);
nand UO_2459 (O_2459,N_29809,N_29450);
xor UO_2460 (O_2460,N_29995,N_29692);
and UO_2461 (O_2461,N_29979,N_29903);
xnor UO_2462 (O_2462,N_29473,N_29639);
xnor UO_2463 (O_2463,N_29907,N_29776);
nand UO_2464 (O_2464,N_29787,N_29527);
nor UO_2465 (O_2465,N_29879,N_29579);
xnor UO_2466 (O_2466,N_29773,N_29676);
xnor UO_2467 (O_2467,N_29835,N_29728);
nor UO_2468 (O_2468,N_29542,N_29980);
xnor UO_2469 (O_2469,N_29917,N_29511);
nand UO_2470 (O_2470,N_29995,N_29463);
nor UO_2471 (O_2471,N_29765,N_29875);
nand UO_2472 (O_2472,N_29422,N_29980);
nor UO_2473 (O_2473,N_29782,N_29982);
nand UO_2474 (O_2474,N_29440,N_29460);
nand UO_2475 (O_2475,N_29918,N_29718);
xor UO_2476 (O_2476,N_29458,N_29461);
or UO_2477 (O_2477,N_29462,N_29449);
nor UO_2478 (O_2478,N_29921,N_29535);
nor UO_2479 (O_2479,N_29576,N_29919);
nand UO_2480 (O_2480,N_29965,N_29731);
nand UO_2481 (O_2481,N_29740,N_29439);
and UO_2482 (O_2482,N_29942,N_29843);
nor UO_2483 (O_2483,N_29596,N_29983);
xor UO_2484 (O_2484,N_29757,N_29506);
and UO_2485 (O_2485,N_29820,N_29993);
nor UO_2486 (O_2486,N_29497,N_29958);
nand UO_2487 (O_2487,N_29616,N_29988);
nor UO_2488 (O_2488,N_29677,N_29513);
and UO_2489 (O_2489,N_29989,N_29517);
nor UO_2490 (O_2490,N_29783,N_29625);
xnor UO_2491 (O_2491,N_29450,N_29457);
nand UO_2492 (O_2492,N_29747,N_29501);
nor UO_2493 (O_2493,N_29847,N_29576);
and UO_2494 (O_2494,N_29940,N_29583);
nand UO_2495 (O_2495,N_29459,N_29936);
nand UO_2496 (O_2496,N_29780,N_29513);
nor UO_2497 (O_2497,N_29502,N_29576);
and UO_2498 (O_2498,N_29935,N_29583);
xnor UO_2499 (O_2499,N_29834,N_29951);
or UO_2500 (O_2500,N_29744,N_29659);
nand UO_2501 (O_2501,N_29788,N_29615);
nand UO_2502 (O_2502,N_29694,N_29603);
or UO_2503 (O_2503,N_29612,N_29761);
nand UO_2504 (O_2504,N_29551,N_29426);
nand UO_2505 (O_2505,N_29841,N_29533);
nand UO_2506 (O_2506,N_29983,N_29850);
and UO_2507 (O_2507,N_29583,N_29430);
nand UO_2508 (O_2508,N_29657,N_29970);
and UO_2509 (O_2509,N_29824,N_29904);
and UO_2510 (O_2510,N_29842,N_29462);
xor UO_2511 (O_2511,N_29623,N_29865);
xnor UO_2512 (O_2512,N_29416,N_29795);
xor UO_2513 (O_2513,N_29941,N_29729);
or UO_2514 (O_2514,N_29799,N_29584);
or UO_2515 (O_2515,N_29840,N_29481);
or UO_2516 (O_2516,N_29884,N_29915);
or UO_2517 (O_2517,N_29898,N_29864);
and UO_2518 (O_2518,N_29546,N_29404);
or UO_2519 (O_2519,N_29578,N_29864);
xor UO_2520 (O_2520,N_29695,N_29454);
and UO_2521 (O_2521,N_29617,N_29468);
nor UO_2522 (O_2522,N_29726,N_29415);
nor UO_2523 (O_2523,N_29684,N_29530);
xor UO_2524 (O_2524,N_29932,N_29525);
or UO_2525 (O_2525,N_29517,N_29912);
and UO_2526 (O_2526,N_29763,N_29916);
xnor UO_2527 (O_2527,N_29519,N_29501);
xnor UO_2528 (O_2528,N_29868,N_29740);
nand UO_2529 (O_2529,N_29491,N_29700);
nor UO_2530 (O_2530,N_29550,N_29674);
xor UO_2531 (O_2531,N_29868,N_29825);
nand UO_2532 (O_2532,N_29549,N_29608);
nor UO_2533 (O_2533,N_29492,N_29862);
and UO_2534 (O_2534,N_29422,N_29735);
and UO_2535 (O_2535,N_29806,N_29744);
nor UO_2536 (O_2536,N_29924,N_29687);
or UO_2537 (O_2537,N_29804,N_29478);
or UO_2538 (O_2538,N_29517,N_29472);
nor UO_2539 (O_2539,N_29845,N_29776);
and UO_2540 (O_2540,N_29734,N_29851);
nor UO_2541 (O_2541,N_29654,N_29530);
and UO_2542 (O_2542,N_29428,N_29834);
and UO_2543 (O_2543,N_29968,N_29530);
nand UO_2544 (O_2544,N_29667,N_29617);
or UO_2545 (O_2545,N_29893,N_29612);
xor UO_2546 (O_2546,N_29942,N_29436);
xnor UO_2547 (O_2547,N_29927,N_29997);
xor UO_2548 (O_2548,N_29744,N_29998);
xnor UO_2549 (O_2549,N_29730,N_29423);
nand UO_2550 (O_2550,N_29693,N_29706);
xor UO_2551 (O_2551,N_29930,N_29877);
and UO_2552 (O_2552,N_29476,N_29626);
and UO_2553 (O_2553,N_29473,N_29741);
or UO_2554 (O_2554,N_29401,N_29906);
nor UO_2555 (O_2555,N_29411,N_29885);
and UO_2556 (O_2556,N_29559,N_29717);
nor UO_2557 (O_2557,N_29515,N_29496);
nor UO_2558 (O_2558,N_29401,N_29554);
and UO_2559 (O_2559,N_29433,N_29973);
nor UO_2560 (O_2560,N_29465,N_29764);
nand UO_2561 (O_2561,N_29701,N_29723);
nand UO_2562 (O_2562,N_29507,N_29774);
and UO_2563 (O_2563,N_29865,N_29409);
and UO_2564 (O_2564,N_29692,N_29888);
nand UO_2565 (O_2565,N_29522,N_29565);
nor UO_2566 (O_2566,N_29583,N_29593);
and UO_2567 (O_2567,N_29542,N_29513);
or UO_2568 (O_2568,N_29569,N_29851);
or UO_2569 (O_2569,N_29534,N_29836);
and UO_2570 (O_2570,N_29766,N_29785);
nand UO_2571 (O_2571,N_29964,N_29489);
or UO_2572 (O_2572,N_29800,N_29608);
nand UO_2573 (O_2573,N_29968,N_29933);
and UO_2574 (O_2574,N_29607,N_29850);
and UO_2575 (O_2575,N_29612,N_29471);
nand UO_2576 (O_2576,N_29680,N_29500);
and UO_2577 (O_2577,N_29514,N_29674);
xnor UO_2578 (O_2578,N_29920,N_29986);
or UO_2579 (O_2579,N_29565,N_29505);
nor UO_2580 (O_2580,N_29481,N_29579);
nor UO_2581 (O_2581,N_29468,N_29911);
nand UO_2582 (O_2582,N_29743,N_29739);
nor UO_2583 (O_2583,N_29952,N_29579);
and UO_2584 (O_2584,N_29734,N_29527);
nor UO_2585 (O_2585,N_29413,N_29966);
nand UO_2586 (O_2586,N_29509,N_29556);
or UO_2587 (O_2587,N_29526,N_29818);
nor UO_2588 (O_2588,N_29553,N_29777);
nand UO_2589 (O_2589,N_29610,N_29828);
nor UO_2590 (O_2590,N_29850,N_29935);
and UO_2591 (O_2591,N_29501,N_29887);
xnor UO_2592 (O_2592,N_29586,N_29957);
and UO_2593 (O_2593,N_29463,N_29518);
xnor UO_2594 (O_2594,N_29711,N_29646);
or UO_2595 (O_2595,N_29648,N_29469);
xnor UO_2596 (O_2596,N_29855,N_29893);
xnor UO_2597 (O_2597,N_29548,N_29998);
nand UO_2598 (O_2598,N_29801,N_29710);
nand UO_2599 (O_2599,N_29450,N_29624);
nor UO_2600 (O_2600,N_29480,N_29564);
or UO_2601 (O_2601,N_29890,N_29485);
and UO_2602 (O_2602,N_29478,N_29544);
xnor UO_2603 (O_2603,N_29953,N_29753);
nand UO_2604 (O_2604,N_29734,N_29896);
and UO_2605 (O_2605,N_29627,N_29981);
nor UO_2606 (O_2606,N_29441,N_29889);
xor UO_2607 (O_2607,N_29796,N_29499);
or UO_2608 (O_2608,N_29612,N_29958);
and UO_2609 (O_2609,N_29894,N_29861);
and UO_2610 (O_2610,N_29621,N_29426);
xor UO_2611 (O_2611,N_29955,N_29879);
nand UO_2612 (O_2612,N_29413,N_29777);
and UO_2613 (O_2613,N_29417,N_29777);
or UO_2614 (O_2614,N_29538,N_29577);
or UO_2615 (O_2615,N_29976,N_29851);
xnor UO_2616 (O_2616,N_29962,N_29569);
nor UO_2617 (O_2617,N_29614,N_29768);
nor UO_2618 (O_2618,N_29400,N_29733);
nor UO_2619 (O_2619,N_29845,N_29445);
and UO_2620 (O_2620,N_29491,N_29816);
nor UO_2621 (O_2621,N_29660,N_29888);
or UO_2622 (O_2622,N_29878,N_29732);
or UO_2623 (O_2623,N_29940,N_29802);
nor UO_2624 (O_2624,N_29801,N_29432);
and UO_2625 (O_2625,N_29530,N_29504);
or UO_2626 (O_2626,N_29497,N_29426);
and UO_2627 (O_2627,N_29977,N_29425);
and UO_2628 (O_2628,N_29417,N_29764);
or UO_2629 (O_2629,N_29899,N_29476);
nor UO_2630 (O_2630,N_29687,N_29899);
nor UO_2631 (O_2631,N_29477,N_29977);
nand UO_2632 (O_2632,N_29599,N_29968);
xnor UO_2633 (O_2633,N_29857,N_29879);
and UO_2634 (O_2634,N_29625,N_29996);
and UO_2635 (O_2635,N_29428,N_29616);
nand UO_2636 (O_2636,N_29882,N_29457);
and UO_2637 (O_2637,N_29873,N_29627);
or UO_2638 (O_2638,N_29632,N_29877);
xor UO_2639 (O_2639,N_29707,N_29676);
nand UO_2640 (O_2640,N_29751,N_29451);
or UO_2641 (O_2641,N_29455,N_29886);
nor UO_2642 (O_2642,N_29578,N_29461);
and UO_2643 (O_2643,N_29559,N_29560);
xor UO_2644 (O_2644,N_29450,N_29643);
xnor UO_2645 (O_2645,N_29550,N_29983);
xor UO_2646 (O_2646,N_29914,N_29445);
xnor UO_2647 (O_2647,N_29591,N_29712);
or UO_2648 (O_2648,N_29437,N_29710);
nand UO_2649 (O_2649,N_29919,N_29824);
and UO_2650 (O_2650,N_29450,N_29902);
nand UO_2651 (O_2651,N_29663,N_29724);
xor UO_2652 (O_2652,N_29467,N_29461);
nor UO_2653 (O_2653,N_29803,N_29671);
nand UO_2654 (O_2654,N_29854,N_29676);
nand UO_2655 (O_2655,N_29754,N_29689);
xnor UO_2656 (O_2656,N_29985,N_29968);
and UO_2657 (O_2657,N_29776,N_29902);
or UO_2658 (O_2658,N_29923,N_29790);
nand UO_2659 (O_2659,N_29951,N_29890);
nor UO_2660 (O_2660,N_29962,N_29605);
or UO_2661 (O_2661,N_29663,N_29950);
or UO_2662 (O_2662,N_29888,N_29518);
xor UO_2663 (O_2663,N_29714,N_29424);
nand UO_2664 (O_2664,N_29659,N_29573);
nand UO_2665 (O_2665,N_29472,N_29761);
nand UO_2666 (O_2666,N_29901,N_29849);
and UO_2667 (O_2667,N_29980,N_29559);
and UO_2668 (O_2668,N_29867,N_29820);
or UO_2669 (O_2669,N_29617,N_29881);
and UO_2670 (O_2670,N_29924,N_29811);
nand UO_2671 (O_2671,N_29653,N_29615);
nand UO_2672 (O_2672,N_29622,N_29869);
and UO_2673 (O_2673,N_29422,N_29839);
and UO_2674 (O_2674,N_29790,N_29961);
and UO_2675 (O_2675,N_29776,N_29617);
nand UO_2676 (O_2676,N_29703,N_29852);
xnor UO_2677 (O_2677,N_29890,N_29852);
nor UO_2678 (O_2678,N_29894,N_29548);
xor UO_2679 (O_2679,N_29930,N_29453);
nand UO_2680 (O_2680,N_29582,N_29733);
nor UO_2681 (O_2681,N_29870,N_29456);
xor UO_2682 (O_2682,N_29404,N_29735);
or UO_2683 (O_2683,N_29872,N_29425);
nor UO_2684 (O_2684,N_29790,N_29778);
or UO_2685 (O_2685,N_29921,N_29677);
or UO_2686 (O_2686,N_29852,N_29484);
nor UO_2687 (O_2687,N_29988,N_29543);
xor UO_2688 (O_2688,N_29568,N_29502);
nor UO_2689 (O_2689,N_29569,N_29754);
or UO_2690 (O_2690,N_29975,N_29872);
nor UO_2691 (O_2691,N_29748,N_29878);
and UO_2692 (O_2692,N_29409,N_29708);
nand UO_2693 (O_2693,N_29581,N_29888);
and UO_2694 (O_2694,N_29866,N_29550);
and UO_2695 (O_2695,N_29497,N_29768);
and UO_2696 (O_2696,N_29781,N_29758);
xnor UO_2697 (O_2697,N_29588,N_29467);
or UO_2698 (O_2698,N_29874,N_29464);
and UO_2699 (O_2699,N_29421,N_29438);
nor UO_2700 (O_2700,N_29488,N_29978);
or UO_2701 (O_2701,N_29731,N_29610);
or UO_2702 (O_2702,N_29447,N_29458);
and UO_2703 (O_2703,N_29454,N_29726);
nor UO_2704 (O_2704,N_29707,N_29789);
xor UO_2705 (O_2705,N_29553,N_29445);
and UO_2706 (O_2706,N_29842,N_29926);
xor UO_2707 (O_2707,N_29813,N_29894);
and UO_2708 (O_2708,N_29658,N_29776);
and UO_2709 (O_2709,N_29488,N_29882);
nand UO_2710 (O_2710,N_29741,N_29414);
nor UO_2711 (O_2711,N_29694,N_29800);
nor UO_2712 (O_2712,N_29730,N_29750);
or UO_2713 (O_2713,N_29662,N_29939);
nor UO_2714 (O_2714,N_29710,N_29424);
xor UO_2715 (O_2715,N_29535,N_29915);
or UO_2716 (O_2716,N_29556,N_29944);
nor UO_2717 (O_2717,N_29661,N_29481);
nand UO_2718 (O_2718,N_29589,N_29507);
and UO_2719 (O_2719,N_29629,N_29862);
nor UO_2720 (O_2720,N_29472,N_29590);
nand UO_2721 (O_2721,N_29978,N_29894);
xnor UO_2722 (O_2722,N_29564,N_29958);
and UO_2723 (O_2723,N_29476,N_29716);
or UO_2724 (O_2724,N_29444,N_29543);
nor UO_2725 (O_2725,N_29459,N_29583);
nand UO_2726 (O_2726,N_29799,N_29407);
xor UO_2727 (O_2727,N_29762,N_29739);
or UO_2728 (O_2728,N_29585,N_29741);
nand UO_2729 (O_2729,N_29563,N_29547);
nand UO_2730 (O_2730,N_29420,N_29895);
xor UO_2731 (O_2731,N_29494,N_29611);
or UO_2732 (O_2732,N_29745,N_29837);
and UO_2733 (O_2733,N_29788,N_29497);
nand UO_2734 (O_2734,N_29549,N_29429);
nand UO_2735 (O_2735,N_29429,N_29422);
xnor UO_2736 (O_2736,N_29766,N_29707);
nor UO_2737 (O_2737,N_29680,N_29547);
or UO_2738 (O_2738,N_29633,N_29563);
or UO_2739 (O_2739,N_29963,N_29486);
and UO_2740 (O_2740,N_29642,N_29950);
nand UO_2741 (O_2741,N_29920,N_29466);
nand UO_2742 (O_2742,N_29945,N_29416);
nand UO_2743 (O_2743,N_29480,N_29719);
and UO_2744 (O_2744,N_29554,N_29608);
nor UO_2745 (O_2745,N_29802,N_29695);
or UO_2746 (O_2746,N_29955,N_29841);
nor UO_2747 (O_2747,N_29925,N_29445);
nor UO_2748 (O_2748,N_29567,N_29883);
xor UO_2749 (O_2749,N_29651,N_29686);
xnor UO_2750 (O_2750,N_29508,N_29922);
and UO_2751 (O_2751,N_29554,N_29849);
and UO_2752 (O_2752,N_29427,N_29717);
nor UO_2753 (O_2753,N_29940,N_29580);
or UO_2754 (O_2754,N_29773,N_29960);
xnor UO_2755 (O_2755,N_29784,N_29811);
and UO_2756 (O_2756,N_29687,N_29425);
or UO_2757 (O_2757,N_29439,N_29970);
xnor UO_2758 (O_2758,N_29586,N_29682);
nand UO_2759 (O_2759,N_29772,N_29507);
xnor UO_2760 (O_2760,N_29677,N_29825);
or UO_2761 (O_2761,N_29510,N_29562);
nand UO_2762 (O_2762,N_29654,N_29719);
or UO_2763 (O_2763,N_29981,N_29997);
nor UO_2764 (O_2764,N_29868,N_29483);
or UO_2765 (O_2765,N_29875,N_29524);
or UO_2766 (O_2766,N_29825,N_29831);
and UO_2767 (O_2767,N_29794,N_29923);
xnor UO_2768 (O_2768,N_29799,N_29993);
and UO_2769 (O_2769,N_29807,N_29569);
or UO_2770 (O_2770,N_29475,N_29555);
or UO_2771 (O_2771,N_29405,N_29859);
or UO_2772 (O_2772,N_29588,N_29440);
nand UO_2773 (O_2773,N_29515,N_29747);
nor UO_2774 (O_2774,N_29701,N_29661);
nand UO_2775 (O_2775,N_29812,N_29721);
or UO_2776 (O_2776,N_29605,N_29896);
or UO_2777 (O_2777,N_29718,N_29856);
and UO_2778 (O_2778,N_29911,N_29651);
and UO_2779 (O_2779,N_29647,N_29823);
nand UO_2780 (O_2780,N_29823,N_29501);
or UO_2781 (O_2781,N_29978,N_29771);
and UO_2782 (O_2782,N_29816,N_29704);
xnor UO_2783 (O_2783,N_29525,N_29988);
xor UO_2784 (O_2784,N_29758,N_29673);
or UO_2785 (O_2785,N_29599,N_29538);
nor UO_2786 (O_2786,N_29508,N_29624);
or UO_2787 (O_2787,N_29847,N_29539);
xnor UO_2788 (O_2788,N_29940,N_29697);
xnor UO_2789 (O_2789,N_29798,N_29440);
nand UO_2790 (O_2790,N_29616,N_29467);
xor UO_2791 (O_2791,N_29632,N_29405);
xor UO_2792 (O_2792,N_29427,N_29736);
xor UO_2793 (O_2793,N_29908,N_29925);
nand UO_2794 (O_2794,N_29673,N_29467);
nand UO_2795 (O_2795,N_29619,N_29892);
nand UO_2796 (O_2796,N_29851,N_29481);
nand UO_2797 (O_2797,N_29434,N_29733);
and UO_2798 (O_2798,N_29525,N_29873);
or UO_2799 (O_2799,N_29854,N_29644);
nor UO_2800 (O_2800,N_29979,N_29964);
nand UO_2801 (O_2801,N_29571,N_29869);
and UO_2802 (O_2802,N_29469,N_29770);
and UO_2803 (O_2803,N_29575,N_29810);
or UO_2804 (O_2804,N_29831,N_29669);
nor UO_2805 (O_2805,N_29950,N_29763);
and UO_2806 (O_2806,N_29562,N_29695);
nand UO_2807 (O_2807,N_29804,N_29602);
nor UO_2808 (O_2808,N_29652,N_29811);
nand UO_2809 (O_2809,N_29448,N_29522);
or UO_2810 (O_2810,N_29740,N_29648);
or UO_2811 (O_2811,N_29966,N_29978);
or UO_2812 (O_2812,N_29993,N_29757);
xnor UO_2813 (O_2813,N_29655,N_29457);
or UO_2814 (O_2814,N_29563,N_29811);
and UO_2815 (O_2815,N_29881,N_29883);
xnor UO_2816 (O_2816,N_29939,N_29727);
nor UO_2817 (O_2817,N_29630,N_29544);
nor UO_2818 (O_2818,N_29813,N_29752);
nand UO_2819 (O_2819,N_29843,N_29680);
nor UO_2820 (O_2820,N_29924,N_29793);
and UO_2821 (O_2821,N_29493,N_29676);
and UO_2822 (O_2822,N_29770,N_29896);
xnor UO_2823 (O_2823,N_29842,N_29647);
nand UO_2824 (O_2824,N_29941,N_29950);
nand UO_2825 (O_2825,N_29505,N_29727);
nand UO_2826 (O_2826,N_29480,N_29411);
nand UO_2827 (O_2827,N_29833,N_29924);
nor UO_2828 (O_2828,N_29494,N_29783);
nor UO_2829 (O_2829,N_29973,N_29543);
xor UO_2830 (O_2830,N_29623,N_29760);
and UO_2831 (O_2831,N_29846,N_29769);
nand UO_2832 (O_2832,N_29744,N_29450);
and UO_2833 (O_2833,N_29491,N_29457);
xor UO_2834 (O_2834,N_29724,N_29715);
and UO_2835 (O_2835,N_29822,N_29861);
xnor UO_2836 (O_2836,N_29528,N_29659);
and UO_2837 (O_2837,N_29952,N_29507);
nand UO_2838 (O_2838,N_29551,N_29654);
or UO_2839 (O_2839,N_29439,N_29888);
xnor UO_2840 (O_2840,N_29651,N_29698);
nand UO_2841 (O_2841,N_29959,N_29755);
or UO_2842 (O_2842,N_29808,N_29861);
or UO_2843 (O_2843,N_29515,N_29488);
nand UO_2844 (O_2844,N_29819,N_29937);
nand UO_2845 (O_2845,N_29699,N_29701);
xnor UO_2846 (O_2846,N_29688,N_29903);
nor UO_2847 (O_2847,N_29707,N_29836);
or UO_2848 (O_2848,N_29787,N_29966);
nor UO_2849 (O_2849,N_29918,N_29802);
nor UO_2850 (O_2850,N_29733,N_29573);
and UO_2851 (O_2851,N_29579,N_29457);
or UO_2852 (O_2852,N_29921,N_29757);
nor UO_2853 (O_2853,N_29558,N_29447);
nor UO_2854 (O_2854,N_29667,N_29901);
xnor UO_2855 (O_2855,N_29719,N_29562);
nand UO_2856 (O_2856,N_29837,N_29998);
xor UO_2857 (O_2857,N_29904,N_29466);
nor UO_2858 (O_2858,N_29774,N_29407);
xnor UO_2859 (O_2859,N_29997,N_29863);
or UO_2860 (O_2860,N_29440,N_29402);
nand UO_2861 (O_2861,N_29546,N_29919);
and UO_2862 (O_2862,N_29589,N_29474);
xnor UO_2863 (O_2863,N_29651,N_29496);
nor UO_2864 (O_2864,N_29846,N_29734);
xnor UO_2865 (O_2865,N_29959,N_29837);
nand UO_2866 (O_2866,N_29452,N_29959);
nand UO_2867 (O_2867,N_29413,N_29891);
and UO_2868 (O_2868,N_29954,N_29756);
xor UO_2869 (O_2869,N_29446,N_29998);
nor UO_2870 (O_2870,N_29826,N_29914);
and UO_2871 (O_2871,N_29929,N_29714);
or UO_2872 (O_2872,N_29462,N_29601);
and UO_2873 (O_2873,N_29430,N_29704);
nand UO_2874 (O_2874,N_29547,N_29842);
or UO_2875 (O_2875,N_29877,N_29947);
xnor UO_2876 (O_2876,N_29536,N_29802);
and UO_2877 (O_2877,N_29503,N_29587);
xnor UO_2878 (O_2878,N_29750,N_29863);
and UO_2879 (O_2879,N_29667,N_29994);
xor UO_2880 (O_2880,N_29587,N_29621);
and UO_2881 (O_2881,N_29881,N_29407);
or UO_2882 (O_2882,N_29877,N_29915);
nor UO_2883 (O_2883,N_29950,N_29938);
xor UO_2884 (O_2884,N_29760,N_29939);
or UO_2885 (O_2885,N_29598,N_29759);
and UO_2886 (O_2886,N_29437,N_29582);
or UO_2887 (O_2887,N_29632,N_29932);
or UO_2888 (O_2888,N_29919,N_29764);
or UO_2889 (O_2889,N_29723,N_29713);
or UO_2890 (O_2890,N_29898,N_29730);
xnor UO_2891 (O_2891,N_29819,N_29737);
or UO_2892 (O_2892,N_29864,N_29536);
nor UO_2893 (O_2893,N_29527,N_29711);
nor UO_2894 (O_2894,N_29557,N_29401);
or UO_2895 (O_2895,N_29735,N_29839);
xnor UO_2896 (O_2896,N_29559,N_29992);
xnor UO_2897 (O_2897,N_29480,N_29776);
and UO_2898 (O_2898,N_29641,N_29833);
nand UO_2899 (O_2899,N_29562,N_29866);
nor UO_2900 (O_2900,N_29435,N_29980);
or UO_2901 (O_2901,N_29629,N_29837);
or UO_2902 (O_2902,N_29497,N_29654);
nor UO_2903 (O_2903,N_29422,N_29495);
nand UO_2904 (O_2904,N_29804,N_29979);
nor UO_2905 (O_2905,N_29729,N_29524);
nand UO_2906 (O_2906,N_29842,N_29953);
nand UO_2907 (O_2907,N_29748,N_29728);
and UO_2908 (O_2908,N_29832,N_29719);
or UO_2909 (O_2909,N_29609,N_29856);
or UO_2910 (O_2910,N_29607,N_29684);
nor UO_2911 (O_2911,N_29978,N_29979);
nor UO_2912 (O_2912,N_29888,N_29460);
or UO_2913 (O_2913,N_29597,N_29684);
nand UO_2914 (O_2914,N_29907,N_29507);
and UO_2915 (O_2915,N_29524,N_29843);
nand UO_2916 (O_2916,N_29698,N_29626);
nor UO_2917 (O_2917,N_29443,N_29975);
or UO_2918 (O_2918,N_29653,N_29504);
nor UO_2919 (O_2919,N_29758,N_29617);
and UO_2920 (O_2920,N_29553,N_29426);
xnor UO_2921 (O_2921,N_29895,N_29609);
xnor UO_2922 (O_2922,N_29525,N_29606);
xor UO_2923 (O_2923,N_29839,N_29563);
and UO_2924 (O_2924,N_29692,N_29820);
or UO_2925 (O_2925,N_29985,N_29754);
xor UO_2926 (O_2926,N_29888,N_29723);
nor UO_2927 (O_2927,N_29761,N_29490);
xnor UO_2928 (O_2928,N_29510,N_29616);
nand UO_2929 (O_2929,N_29513,N_29635);
xor UO_2930 (O_2930,N_29943,N_29445);
nand UO_2931 (O_2931,N_29853,N_29696);
nand UO_2932 (O_2932,N_29616,N_29431);
and UO_2933 (O_2933,N_29816,N_29761);
and UO_2934 (O_2934,N_29998,N_29422);
nand UO_2935 (O_2935,N_29799,N_29968);
and UO_2936 (O_2936,N_29873,N_29993);
nor UO_2937 (O_2937,N_29939,N_29973);
nor UO_2938 (O_2938,N_29582,N_29961);
xnor UO_2939 (O_2939,N_29899,N_29401);
or UO_2940 (O_2940,N_29460,N_29966);
nor UO_2941 (O_2941,N_29934,N_29942);
xnor UO_2942 (O_2942,N_29854,N_29597);
nand UO_2943 (O_2943,N_29810,N_29704);
nand UO_2944 (O_2944,N_29801,N_29736);
nand UO_2945 (O_2945,N_29479,N_29917);
or UO_2946 (O_2946,N_29971,N_29558);
and UO_2947 (O_2947,N_29407,N_29593);
or UO_2948 (O_2948,N_29704,N_29458);
nand UO_2949 (O_2949,N_29977,N_29521);
or UO_2950 (O_2950,N_29550,N_29442);
nand UO_2951 (O_2951,N_29578,N_29899);
nor UO_2952 (O_2952,N_29657,N_29847);
xnor UO_2953 (O_2953,N_29814,N_29494);
or UO_2954 (O_2954,N_29969,N_29453);
nor UO_2955 (O_2955,N_29493,N_29673);
nand UO_2956 (O_2956,N_29957,N_29634);
nor UO_2957 (O_2957,N_29938,N_29715);
nor UO_2958 (O_2958,N_29966,N_29490);
and UO_2959 (O_2959,N_29562,N_29842);
and UO_2960 (O_2960,N_29422,N_29602);
nand UO_2961 (O_2961,N_29837,N_29642);
xor UO_2962 (O_2962,N_29778,N_29703);
or UO_2963 (O_2963,N_29896,N_29665);
xor UO_2964 (O_2964,N_29971,N_29836);
nor UO_2965 (O_2965,N_29732,N_29851);
and UO_2966 (O_2966,N_29576,N_29659);
xnor UO_2967 (O_2967,N_29583,N_29873);
nor UO_2968 (O_2968,N_29449,N_29639);
nand UO_2969 (O_2969,N_29950,N_29930);
nand UO_2970 (O_2970,N_29734,N_29569);
or UO_2971 (O_2971,N_29655,N_29848);
nor UO_2972 (O_2972,N_29470,N_29703);
nand UO_2973 (O_2973,N_29629,N_29993);
xor UO_2974 (O_2974,N_29768,N_29793);
and UO_2975 (O_2975,N_29872,N_29817);
or UO_2976 (O_2976,N_29822,N_29957);
or UO_2977 (O_2977,N_29476,N_29777);
and UO_2978 (O_2978,N_29920,N_29499);
and UO_2979 (O_2979,N_29754,N_29936);
xor UO_2980 (O_2980,N_29811,N_29706);
or UO_2981 (O_2981,N_29444,N_29601);
nand UO_2982 (O_2982,N_29799,N_29798);
nor UO_2983 (O_2983,N_29932,N_29974);
and UO_2984 (O_2984,N_29753,N_29701);
or UO_2985 (O_2985,N_29881,N_29603);
or UO_2986 (O_2986,N_29655,N_29811);
xor UO_2987 (O_2987,N_29537,N_29626);
and UO_2988 (O_2988,N_29601,N_29980);
or UO_2989 (O_2989,N_29403,N_29822);
and UO_2990 (O_2990,N_29746,N_29996);
xnor UO_2991 (O_2991,N_29798,N_29880);
or UO_2992 (O_2992,N_29427,N_29522);
and UO_2993 (O_2993,N_29761,N_29566);
xor UO_2994 (O_2994,N_29661,N_29936);
nor UO_2995 (O_2995,N_29821,N_29817);
and UO_2996 (O_2996,N_29906,N_29883);
nand UO_2997 (O_2997,N_29418,N_29444);
xor UO_2998 (O_2998,N_29545,N_29968);
nand UO_2999 (O_2999,N_29726,N_29456);
and UO_3000 (O_3000,N_29687,N_29876);
and UO_3001 (O_3001,N_29446,N_29563);
nor UO_3002 (O_3002,N_29773,N_29893);
or UO_3003 (O_3003,N_29690,N_29402);
and UO_3004 (O_3004,N_29762,N_29519);
and UO_3005 (O_3005,N_29597,N_29778);
nand UO_3006 (O_3006,N_29434,N_29736);
nand UO_3007 (O_3007,N_29764,N_29836);
nand UO_3008 (O_3008,N_29629,N_29403);
nand UO_3009 (O_3009,N_29670,N_29953);
nand UO_3010 (O_3010,N_29577,N_29479);
nand UO_3011 (O_3011,N_29463,N_29407);
nor UO_3012 (O_3012,N_29900,N_29815);
or UO_3013 (O_3013,N_29666,N_29631);
xor UO_3014 (O_3014,N_29413,N_29867);
xnor UO_3015 (O_3015,N_29916,N_29861);
nor UO_3016 (O_3016,N_29800,N_29947);
or UO_3017 (O_3017,N_29800,N_29596);
xnor UO_3018 (O_3018,N_29857,N_29866);
and UO_3019 (O_3019,N_29570,N_29880);
nand UO_3020 (O_3020,N_29816,N_29563);
and UO_3021 (O_3021,N_29820,N_29602);
or UO_3022 (O_3022,N_29464,N_29449);
nand UO_3023 (O_3023,N_29965,N_29625);
or UO_3024 (O_3024,N_29417,N_29864);
xnor UO_3025 (O_3025,N_29485,N_29559);
nor UO_3026 (O_3026,N_29804,N_29587);
or UO_3027 (O_3027,N_29490,N_29723);
and UO_3028 (O_3028,N_29722,N_29932);
and UO_3029 (O_3029,N_29630,N_29891);
nor UO_3030 (O_3030,N_29448,N_29803);
and UO_3031 (O_3031,N_29467,N_29415);
and UO_3032 (O_3032,N_29687,N_29564);
or UO_3033 (O_3033,N_29751,N_29560);
and UO_3034 (O_3034,N_29737,N_29614);
nor UO_3035 (O_3035,N_29675,N_29646);
nand UO_3036 (O_3036,N_29651,N_29782);
and UO_3037 (O_3037,N_29998,N_29936);
nand UO_3038 (O_3038,N_29891,N_29900);
or UO_3039 (O_3039,N_29515,N_29912);
nand UO_3040 (O_3040,N_29910,N_29829);
xnor UO_3041 (O_3041,N_29883,N_29545);
or UO_3042 (O_3042,N_29774,N_29561);
nand UO_3043 (O_3043,N_29917,N_29710);
nand UO_3044 (O_3044,N_29791,N_29876);
nand UO_3045 (O_3045,N_29914,N_29923);
nand UO_3046 (O_3046,N_29864,N_29660);
and UO_3047 (O_3047,N_29959,N_29549);
or UO_3048 (O_3048,N_29869,N_29522);
nor UO_3049 (O_3049,N_29915,N_29764);
nor UO_3050 (O_3050,N_29887,N_29474);
nand UO_3051 (O_3051,N_29873,N_29420);
xor UO_3052 (O_3052,N_29748,N_29512);
and UO_3053 (O_3053,N_29695,N_29587);
nor UO_3054 (O_3054,N_29757,N_29433);
xor UO_3055 (O_3055,N_29752,N_29623);
nand UO_3056 (O_3056,N_29489,N_29817);
nand UO_3057 (O_3057,N_29997,N_29636);
xnor UO_3058 (O_3058,N_29652,N_29679);
and UO_3059 (O_3059,N_29581,N_29502);
and UO_3060 (O_3060,N_29826,N_29682);
nand UO_3061 (O_3061,N_29409,N_29826);
nor UO_3062 (O_3062,N_29742,N_29653);
or UO_3063 (O_3063,N_29753,N_29642);
or UO_3064 (O_3064,N_29449,N_29859);
xor UO_3065 (O_3065,N_29650,N_29463);
or UO_3066 (O_3066,N_29742,N_29655);
and UO_3067 (O_3067,N_29806,N_29654);
xor UO_3068 (O_3068,N_29864,N_29599);
nand UO_3069 (O_3069,N_29432,N_29703);
nor UO_3070 (O_3070,N_29527,N_29786);
nand UO_3071 (O_3071,N_29661,N_29586);
and UO_3072 (O_3072,N_29677,N_29807);
and UO_3073 (O_3073,N_29966,N_29409);
nor UO_3074 (O_3074,N_29523,N_29887);
xor UO_3075 (O_3075,N_29529,N_29659);
or UO_3076 (O_3076,N_29472,N_29732);
xor UO_3077 (O_3077,N_29801,N_29555);
and UO_3078 (O_3078,N_29484,N_29737);
nand UO_3079 (O_3079,N_29614,N_29964);
or UO_3080 (O_3080,N_29810,N_29945);
nand UO_3081 (O_3081,N_29551,N_29430);
nor UO_3082 (O_3082,N_29781,N_29881);
and UO_3083 (O_3083,N_29660,N_29987);
or UO_3084 (O_3084,N_29949,N_29509);
nor UO_3085 (O_3085,N_29532,N_29479);
xnor UO_3086 (O_3086,N_29574,N_29799);
nor UO_3087 (O_3087,N_29434,N_29927);
nor UO_3088 (O_3088,N_29715,N_29764);
nand UO_3089 (O_3089,N_29675,N_29961);
xor UO_3090 (O_3090,N_29570,N_29845);
nor UO_3091 (O_3091,N_29675,N_29828);
and UO_3092 (O_3092,N_29480,N_29909);
nor UO_3093 (O_3093,N_29868,N_29980);
or UO_3094 (O_3094,N_29867,N_29888);
and UO_3095 (O_3095,N_29478,N_29933);
and UO_3096 (O_3096,N_29998,N_29463);
or UO_3097 (O_3097,N_29577,N_29915);
xor UO_3098 (O_3098,N_29793,N_29940);
nor UO_3099 (O_3099,N_29480,N_29436);
nor UO_3100 (O_3100,N_29535,N_29561);
xor UO_3101 (O_3101,N_29644,N_29901);
nand UO_3102 (O_3102,N_29567,N_29576);
xor UO_3103 (O_3103,N_29553,N_29878);
nand UO_3104 (O_3104,N_29569,N_29528);
nand UO_3105 (O_3105,N_29557,N_29991);
xnor UO_3106 (O_3106,N_29528,N_29822);
xor UO_3107 (O_3107,N_29428,N_29689);
and UO_3108 (O_3108,N_29786,N_29489);
xnor UO_3109 (O_3109,N_29687,N_29933);
or UO_3110 (O_3110,N_29574,N_29846);
xnor UO_3111 (O_3111,N_29959,N_29933);
nand UO_3112 (O_3112,N_29558,N_29655);
xnor UO_3113 (O_3113,N_29664,N_29945);
or UO_3114 (O_3114,N_29627,N_29659);
nor UO_3115 (O_3115,N_29522,N_29676);
nor UO_3116 (O_3116,N_29591,N_29498);
nor UO_3117 (O_3117,N_29949,N_29578);
and UO_3118 (O_3118,N_29878,N_29902);
nand UO_3119 (O_3119,N_29621,N_29767);
and UO_3120 (O_3120,N_29572,N_29938);
and UO_3121 (O_3121,N_29985,N_29700);
or UO_3122 (O_3122,N_29505,N_29704);
and UO_3123 (O_3123,N_29888,N_29598);
nand UO_3124 (O_3124,N_29425,N_29778);
and UO_3125 (O_3125,N_29551,N_29532);
or UO_3126 (O_3126,N_29517,N_29922);
and UO_3127 (O_3127,N_29402,N_29611);
or UO_3128 (O_3128,N_29607,N_29858);
nand UO_3129 (O_3129,N_29478,N_29572);
nor UO_3130 (O_3130,N_29595,N_29815);
or UO_3131 (O_3131,N_29696,N_29917);
nand UO_3132 (O_3132,N_29946,N_29811);
or UO_3133 (O_3133,N_29952,N_29711);
or UO_3134 (O_3134,N_29597,N_29669);
nor UO_3135 (O_3135,N_29713,N_29684);
nor UO_3136 (O_3136,N_29469,N_29573);
nor UO_3137 (O_3137,N_29489,N_29420);
nor UO_3138 (O_3138,N_29688,N_29974);
nor UO_3139 (O_3139,N_29880,N_29609);
nand UO_3140 (O_3140,N_29649,N_29622);
or UO_3141 (O_3141,N_29620,N_29691);
nor UO_3142 (O_3142,N_29521,N_29561);
nor UO_3143 (O_3143,N_29725,N_29995);
xor UO_3144 (O_3144,N_29874,N_29736);
nand UO_3145 (O_3145,N_29697,N_29968);
or UO_3146 (O_3146,N_29779,N_29501);
or UO_3147 (O_3147,N_29810,N_29692);
xnor UO_3148 (O_3148,N_29567,N_29935);
xnor UO_3149 (O_3149,N_29417,N_29618);
nor UO_3150 (O_3150,N_29880,N_29708);
xor UO_3151 (O_3151,N_29779,N_29658);
nand UO_3152 (O_3152,N_29803,N_29585);
nand UO_3153 (O_3153,N_29946,N_29563);
nand UO_3154 (O_3154,N_29737,N_29559);
nand UO_3155 (O_3155,N_29412,N_29985);
or UO_3156 (O_3156,N_29947,N_29788);
nor UO_3157 (O_3157,N_29837,N_29820);
nor UO_3158 (O_3158,N_29650,N_29589);
or UO_3159 (O_3159,N_29923,N_29480);
nor UO_3160 (O_3160,N_29657,N_29887);
and UO_3161 (O_3161,N_29548,N_29887);
xor UO_3162 (O_3162,N_29777,N_29974);
xor UO_3163 (O_3163,N_29681,N_29492);
xor UO_3164 (O_3164,N_29436,N_29613);
and UO_3165 (O_3165,N_29540,N_29910);
and UO_3166 (O_3166,N_29627,N_29829);
xor UO_3167 (O_3167,N_29847,N_29895);
or UO_3168 (O_3168,N_29541,N_29942);
xnor UO_3169 (O_3169,N_29670,N_29668);
nor UO_3170 (O_3170,N_29851,N_29494);
xor UO_3171 (O_3171,N_29416,N_29978);
nor UO_3172 (O_3172,N_29860,N_29903);
nor UO_3173 (O_3173,N_29660,N_29942);
xor UO_3174 (O_3174,N_29766,N_29809);
xnor UO_3175 (O_3175,N_29757,N_29493);
nor UO_3176 (O_3176,N_29652,N_29584);
or UO_3177 (O_3177,N_29936,N_29740);
nand UO_3178 (O_3178,N_29445,N_29688);
nor UO_3179 (O_3179,N_29429,N_29482);
nor UO_3180 (O_3180,N_29781,N_29410);
xor UO_3181 (O_3181,N_29756,N_29401);
xnor UO_3182 (O_3182,N_29742,N_29570);
or UO_3183 (O_3183,N_29838,N_29523);
nand UO_3184 (O_3184,N_29814,N_29616);
nor UO_3185 (O_3185,N_29492,N_29892);
or UO_3186 (O_3186,N_29632,N_29611);
and UO_3187 (O_3187,N_29718,N_29929);
nand UO_3188 (O_3188,N_29491,N_29615);
nand UO_3189 (O_3189,N_29401,N_29479);
nor UO_3190 (O_3190,N_29832,N_29971);
or UO_3191 (O_3191,N_29430,N_29872);
and UO_3192 (O_3192,N_29771,N_29590);
and UO_3193 (O_3193,N_29510,N_29985);
nor UO_3194 (O_3194,N_29853,N_29939);
nor UO_3195 (O_3195,N_29812,N_29903);
nand UO_3196 (O_3196,N_29408,N_29427);
nand UO_3197 (O_3197,N_29759,N_29568);
or UO_3198 (O_3198,N_29983,N_29776);
and UO_3199 (O_3199,N_29669,N_29435);
nor UO_3200 (O_3200,N_29954,N_29461);
xor UO_3201 (O_3201,N_29763,N_29662);
and UO_3202 (O_3202,N_29890,N_29712);
xor UO_3203 (O_3203,N_29707,N_29427);
nand UO_3204 (O_3204,N_29546,N_29563);
and UO_3205 (O_3205,N_29552,N_29408);
xnor UO_3206 (O_3206,N_29537,N_29634);
and UO_3207 (O_3207,N_29567,N_29518);
and UO_3208 (O_3208,N_29660,N_29912);
nor UO_3209 (O_3209,N_29490,N_29919);
xor UO_3210 (O_3210,N_29607,N_29915);
nand UO_3211 (O_3211,N_29420,N_29803);
nand UO_3212 (O_3212,N_29526,N_29484);
nand UO_3213 (O_3213,N_29734,N_29998);
xor UO_3214 (O_3214,N_29756,N_29721);
and UO_3215 (O_3215,N_29466,N_29586);
and UO_3216 (O_3216,N_29759,N_29777);
and UO_3217 (O_3217,N_29685,N_29653);
or UO_3218 (O_3218,N_29762,N_29787);
or UO_3219 (O_3219,N_29501,N_29791);
or UO_3220 (O_3220,N_29873,N_29600);
nand UO_3221 (O_3221,N_29864,N_29556);
nand UO_3222 (O_3222,N_29545,N_29417);
and UO_3223 (O_3223,N_29942,N_29739);
nand UO_3224 (O_3224,N_29454,N_29980);
or UO_3225 (O_3225,N_29904,N_29493);
nor UO_3226 (O_3226,N_29446,N_29944);
nand UO_3227 (O_3227,N_29432,N_29571);
nor UO_3228 (O_3228,N_29872,N_29843);
nor UO_3229 (O_3229,N_29483,N_29979);
or UO_3230 (O_3230,N_29839,N_29841);
nor UO_3231 (O_3231,N_29803,N_29882);
or UO_3232 (O_3232,N_29508,N_29875);
xor UO_3233 (O_3233,N_29412,N_29876);
or UO_3234 (O_3234,N_29638,N_29559);
or UO_3235 (O_3235,N_29836,N_29628);
xor UO_3236 (O_3236,N_29568,N_29472);
xnor UO_3237 (O_3237,N_29424,N_29401);
and UO_3238 (O_3238,N_29923,N_29633);
nor UO_3239 (O_3239,N_29885,N_29548);
nand UO_3240 (O_3240,N_29742,N_29431);
and UO_3241 (O_3241,N_29475,N_29432);
xnor UO_3242 (O_3242,N_29830,N_29871);
xor UO_3243 (O_3243,N_29796,N_29852);
nand UO_3244 (O_3244,N_29823,N_29532);
nand UO_3245 (O_3245,N_29614,N_29859);
and UO_3246 (O_3246,N_29792,N_29655);
xnor UO_3247 (O_3247,N_29646,N_29462);
nand UO_3248 (O_3248,N_29729,N_29884);
and UO_3249 (O_3249,N_29453,N_29765);
nand UO_3250 (O_3250,N_29486,N_29995);
nor UO_3251 (O_3251,N_29763,N_29454);
nand UO_3252 (O_3252,N_29923,N_29534);
nor UO_3253 (O_3253,N_29544,N_29961);
nand UO_3254 (O_3254,N_29746,N_29791);
or UO_3255 (O_3255,N_29798,N_29845);
nor UO_3256 (O_3256,N_29490,N_29994);
nor UO_3257 (O_3257,N_29530,N_29953);
nand UO_3258 (O_3258,N_29489,N_29597);
nor UO_3259 (O_3259,N_29557,N_29977);
xor UO_3260 (O_3260,N_29489,N_29788);
nor UO_3261 (O_3261,N_29508,N_29973);
nor UO_3262 (O_3262,N_29640,N_29587);
or UO_3263 (O_3263,N_29791,N_29433);
or UO_3264 (O_3264,N_29577,N_29469);
nor UO_3265 (O_3265,N_29858,N_29965);
nand UO_3266 (O_3266,N_29622,N_29861);
nand UO_3267 (O_3267,N_29994,N_29497);
xnor UO_3268 (O_3268,N_29465,N_29562);
nand UO_3269 (O_3269,N_29850,N_29876);
nand UO_3270 (O_3270,N_29644,N_29910);
nand UO_3271 (O_3271,N_29673,N_29999);
and UO_3272 (O_3272,N_29586,N_29955);
or UO_3273 (O_3273,N_29786,N_29637);
nor UO_3274 (O_3274,N_29410,N_29826);
nor UO_3275 (O_3275,N_29715,N_29988);
or UO_3276 (O_3276,N_29762,N_29935);
nor UO_3277 (O_3277,N_29717,N_29767);
xor UO_3278 (O_3278,N_29897,N_29686);
or UO_3279 (O_3279,N_29754,N_29760);
xnor UO_3280 (O_3280,N_29673,N_29582);
xor UO_3281 (O_3281,N_29893,N_29668);
and UO_3282 (O_3282,N_29776,N_29810);
xor UO_3283 (O_3283,N_29744,N_29428);
and UO_3284 (O_3284,N_29809,N_29601);
and UO_3285 (O_3285,N_29811,N_29464);
xor UO_3286 (O_3286,N_29880,N_29720);
and UO_3287 (O_3287,N_29949,N_29558);
and UO_3288 (O_3288,N_29817,N_29560);
or UO_3289 (O_3289,N_29948,N_29772);
nand UO_3290 (O_3290,N_29822,N_29892);
and UO_3291 (O_3291,N_29414,N_29595);
nand UO_3292 (O_3292,N_29848,N_29949);
or UO_3293 (O_3293,N_29720,N_29637);
nor UO_3294 (O_3294,N_29670,N_29891);
xnor UO_3295 (O_3295,N_29825,N_29612);
and UO_3296 (O_3296,N_29478,N_29855);
xor UO_3297 (O_3297,N_29986,N_29687);
nand UO_3298 (O_3298,N_29926,N_29484);
or UO_3299 (O_3299,N_29420,N_29773);
or UO_3300 (O_3300,N_29660,N_29894);
or UO_3301 (O_3301,N_29408,N_29773);
nand UO_3302 (O_3302,N_29776,N_29897);
nor UO_3303 (O_3303,N_29908,N_29717);
nand UO_3304 (O_3304,N_29581,N_29861);
and UO_3305 (O_3305,N_29675,N_29742);
xnor UO_3306 (O_3306,N_29840,N_29869);
nor UO_3307 (O_3307,N_29483,N_29786);
and UO_3308 (O_3308,N_29447,N_29749);
nand UO_3309 (O_3309,N_29739,N_29408);
xnor UO_3310 (O_3310,N_29508,N_29527);
nand UO_3311 (O_3311,N_29812,N_29506);
nand UO_3312 (O_3312,N_29500,N_29947);
or UO_3313 (O_3313,N_29618,N_29543);
xor UO_3314 (O_3314,N_29577,N_29919);
or UO_3315 (O_3315,N_29657,N_29403);
xor UO_3316 (O_3316,N_29574,N_29766);
nor UO_3317 (O_3317,N_29471,N_29901);
nor UO_3318 (O_3318,N_29592,N_29783);
and UO_3319 (O_3319,N_29918,N_29971);
xor UO_3320 (O_3320,N_29624,N_29498);
nand UO_3321 (O_3321,N_29741,N_29902);
nand UO_3322 (O_3322,N_29986,N_29940);
and UO_3323 (O_3323,N_29639,N_29879);
and UO_3324 (O_3324,N_29554,N_29862);
and UO_3325 (O_3325,N_29976,N_29910);
xnor UO_3326 (O_3326,N_29453,N_29771);
nor UO_3327 (O_3327,N_29772,N_29874);
nand UO_3328 (O_3328,N_29658,N_29536);
nand UO_3329 (O_3329,N_29883,N_29403);
xnor UO_3330 (O_3330,N_29798,N_29595);
and UO_3331 (O_3331,N_29738,N_29573);
nor UO_3332 (O_3332,N_29599,N_29961);
or UO_3333 (O_3333,N_29786,N_29474);
and UO_3334 (O_3334,N_29956,N_29881);
or UO_3335 (O_3335,N_29679,N_29931);
and UO_3336 (O_3336,N_29714,N_29489);
or UO_3337 (O_3337,N_29519,N_29552);
nand UO_3338 (O_3338,N_29556,N_29430);
xnor UO_3339 (O_3339,N_29838,N_29810);
and UO_3340 (O_3340,N_29522,N_29781);
nand UO_3341 (O_3341,N_29896,N_29643);
or UO_3342 (O_3342,N_29957,N_29781);
nand UO_3343 (O_3343,N_29805,N_29886);
and UO_3344 (O_3344,N_29707,N_29640);
nand UO_3345 (O_3345,N_29846,N_29828);
nand UO_3346 (O_3346,N_29454,N_29554);
and UO_3347 (O_3347,N_29556,N_29581);
nor UO_3348 (O_3348,N_29596,N_29673);
nand UO_3349 (O_3349,N_29885,N_29798);
xnor UO_3350 (O_3350,N_29838,N_29936);
and UO_3351 (O_3351,N_29994,N_29997);
and UO_3352 (O_3352,N_29835,N_29759);
nand UO_3353 (O_3353,N_29713,N_29674);
and UO_3354 (O_3354,N_29831,N_29941);
and UO_3355 (O_3355,N_29594,N_29445);
nand UO_3356 (O_3356,N_29698,N_29963);
nand UO_3357 (O_3357,N_29492,N_29930);
or UO_3358 (O_3358,N_29989,N_29860);
or UO_3359 (O_3359,N_29968,N_29816);
or UO_3360 (O_3360,N_29871,N_29733);
xnor UO_3361 (O_3361,N_29640,N_29457);
nor UO_3362 (O_3362,N_29587,N_29445);
xnor UO_3363 (O_3363,N_29918,N_29665);
or UO_3364 (O_3364,N_29850,N_29639);
xor UO_3365 (O_3365,N_29915,N_29442);
or UO_3366 (O_3366,N_29834,N_29547);
nor UO_3367 (O_3367,N_29478,N_29442);
nand UO_3368 (O_3368,N_29655,N_29779);
xnor UO_3369 (O_3369,N_29989,N_29430);
nor UO_3370 (O_3370,N_29578,N_29866);
or UO_3371 (O_3371,N_29806,N_29773);
or UO_3372 (O_3372,N_29682,N_29470);
or UO_3373 (O_3373,N_29896,N_29579);
xor UO_3374 (O_3374,N_29650,N_29405);
nor UO_3375 (O_3375,N_29521,N_29416);
and UO_3376 (O_3376,N_29940,N_29683);
xnor UO_3377 (O_3377,N_29918,N_29909);
nor UO_3378 (O_3378,N_29528,N_29508);
or UO_3379 (O_3379,N_29851,N_29472);
xnor UO_3380 (O_3380,N_29883,N_29537);
nand UO_3381 (O_3381,N_29732,N_29470);
and UO_3382 (O_3382,N_29527,N_29526);
and UO_3383 (O_3383,N_29450,N_29967);
nor UO_3384 (O_3384,N_29418,N_29994);
and UO_3385 (O_3385,N_29774,N_29845);
and UO_3386 (O_3386,N_29626,N_29662);
xor UO_3387 (O_3387,N_29459,N_29687);
nor UO_3388 (O_3388,N_29703,N_29527);
or UO_3389 (O_3389,N_29923,N_29662);
or UO_3390 (O_3390,N_29743,N_29510);
nand UO_3391 (O_3391,N_29417,N_29690);
nand UO_3392 (O_3392,N_29936,N_29995);
nand UO_3393 (O_3393,N_29702,N_29945);
xor UO_3394 (O_3394,N_29549,N_29565);
xor UO_3395 (O_3395,N_29831,N_29549);
and UO_3396 (O_3396,N_29518,N_29560);
and UO_3397 (O_3397,N_29974,N_29721);
nand UO_3398 (O_3398,N_29429,N_29929);
and UO_3399 (O_3399,N_29610,N_29704);
and UO_3400 (O_3400,N_29781,N_29757);
xor UO_3401 (O_3401,N_29439,N_29774);
nor UO_3402 (O_3402,N_29734,N_29544);
and UO_3403 (O_3403,N_29880,N_29874);
nand UO_3404 (O_3404,N_29573,N_29827);
nor UO_3405 (O_3405,N_29682,N_29943);
or UO_3406 (O_3406,N_29897,N_29570);
xnor UO_3407 (O_3407,N_29889,N_29623);
xnor UO_3408 (O_3408,N_29824,N_29456);
nor UO_3409 (O_3409,N_29660,N_29522);
nand UO_3410 (O_3410,N_29805,N_29606);
or UO_3411 (O_3411,N_29536,N_29945);
nand UO_3412 (O_3412,N_29620,N_29677);
and UO_3413 (O_3413,N_29610,N_29909);
nor UO_3414 (O_3414,N_29668,N_29635);
xnor UO_3415 (O_3415,N_29541,N_29857);
xnor UO_3416 (O_3416,N_29733,N_29903);
or UO_3417 (O_3417,N_29766,N_29441);
nand UO_3418 (O_3418,N_29695,N_29467);
nor UO_3419 (O_3419,N_29575,N_29922);
xnor UO_3420 (O_3420,N_29926,N_29572);
nor UO_3421 (O_3421,N_29526,N_29452);
xor UO_3422 (O_3422,N_29560,N_29491);
and UO_3423 (O_3423,N_29965,N_29736);
nor UO_3424 (O_3424,N_29469,N_29870);
xnor UO_3425 (O_3425,N_29498,N_29899);
xor UO_3426 (O_3426,N_29834,N_29825);
nand UO_3427 (O_3427,N_29848,N_29766);
xor UO_3428 (O_3428,N_29583,N_29654);
nor UO_3429 (O_3429,N_29796,N_29698);
or UO_3430 (O_3430,N_29446,N_29723);
and UO_3431 (O_3431,N_29523,N_29656);
xnor UO_3432 (O_3432,N_29448,N_29748);
and UO_3433 (O_3433,N_29806,N_29587);
xnor UO_3434 (O_3434,N_29935,N_29640);
nand UO_3435 (O_3435,N_29564,N_29712);
or UO_3436 (O_3436,N_29758,N_29655);
and UO_3437 (O_3437,N_29761,N_29774);
or UO_3438 (O_3438,N_29786,N_29661);
nand UO_3439 (O_3439,N_29878,N_29644);
and UO_3440 (O_3440,N_29770,N_29490);
or UO_3441 (O_3441,N_29686,N_29813);
and UO_3442 (O_3442,N_29840,N_29681);
nor UO_3443 (O_3443,N_29617,N_29620);
and UO_3444 (O_3444,N_29802,N_29662);
xnor UO_3445 (O_3445,N_29838,N_29640);
xor UO_3446 (O_3446,N_29805,N_29689);
nand UO_3447 (O_3447,N_29710,N_29524);
nor UO_3448 (O_3448,N_29478,N_29863);
nor UO_3449 (O_3449,N_29844,N_29625);
xor UO_3450 (O_3450,N_29722,N_29681);
and UO_3451 (O_3451,N_29412,N_29822);
xnor UO_3452 (O_3452,N_29689,N_29510);
or UO_3453 (O_3453,N_29887,N_29930);
nor UO_3454 (O_3454,N_29494,N_29585);
nand UO_3455 (O_3455,N_29687,N_29775);
xor UO_3456 (O_3456,N_29752,N_29413);
or UO_3457 (O_3457,N_29596,N_29408);
nand UO_3458 (O_3458,N_29524,N_29830);
or UO_3459 (O_3459,N_29830,N_29975);
nor UO_3460 (O_3460,N_29466,N_29706);
or UO_3461 (O_3461,N_29544,N_29656);
nand UO_3462 (O_3462,N_29509,N_29855);
xnor UO_3463 (O_3463,N_29744,N_29554);
or UO_3464 (O_3464,N_29616,N_29982);
xor UO_3465 (O_3465,N_29811,N_29565);
xor UO_3466 (O_3466,N_29706,N_29695);
xor UO_3467 (O_3467,N_29537,N_29940);
xor UO_3468 (O_3468,N_29580,N_29834);
and UO_3469 (O_3469,N_29482,N_29768);
xnor UO_3470 (O_3470,N_29440,N_29597);
nand UO_3471 (O_3471,N_29540,N_29931);
and UO_3472 (O_3472,N_29879,N_29693);
and UO_3473 (O_3473,N_29796,N_29629);
nor UO_3474 (O_3474,N_29401,N_29822);
or UO_3475 (O_3475,N_29423,N_29941);
nor UO_3476 (O_3476,N_29669,N_29646);
xnor UO_3477 (O_3477,N_29440,N_29474);
nor UO_3478 (O_3478,N_29990,N_29921);
xnor UO_3479 (O_3479,N_29863,N_29720);
or UO_3480 (O_3480,N_29900,N_29464);
and UO_3481 (O_3481,N_29807,N_29931);
nor UO_3482 (O_3482,N_29552,N_29602);
nand UO_3483 (O_3483,N_29699,N_29927);
xor UO_3484 (O_3484,N_29874,N_29674);
and UO_3485 (O_3485,N_29705,N_29937);
or UO_3486 (O_3486,N_29480,N_29693);
and UO_3487 (O_3487,N_29606,N_29750);
nor UO_3488 (O_3488,N_29772,N_29942);
nor UO_3489 (O_3489,N_29467,N_29487);
xor UO_3490 (O_3490,N_29472,N_29910);
and UO_3491 (O_3491,N_29939,N_29547);
or UO_3492 (O_3492,N_29976,N_29631);
or UO_3493 (O_3493,N_29411,N_29467);
nor UO_3494 (O_3494,N_29682,N_29993);
or UO_3495 (O_3495,N_29508,N_29497);
nor UO_3496 (O_3496,N_29610,N_29854);
or UO_3497 (O_3497,N_29879,N_29910);
xnor UO_3498 (O_3498,N_29903,N_29950);
nand UO_3499 (O_3499,N_29418,N_29835);
endmodule