module basic_2000_20000_2500_25_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1554,In_1814);
xnor U1 (N_1,In_200,In_1037);
or U2 (N_2,In_1039,In_294);
xnor U3 (N_3,In_1375,In_631);
or U4 (N_4,In_1608,In_1316);
xnor U5 (N_5,In_10,In_1582);
xor U6 (N_6,In_1544,In_133);
and U7 (N_7,In_965,In_140);
or U8 (N_8,In_728,In_1597);
nand U9 (N_9,In_1782,In_74);
nor U10 (N_10,In_1270,In_1194);
or U11 (N_11,In_967,In_1163);
and U12 (N_12,In_1502,In_28);
nand U13 (N_13,In_1897,In_1241);
and U14 (N_14,In_1804,In_1747);
xnor U15 (N_15,In_1351,In_1954);
or U16 (N_16,In_1570,In_263);
nor U17 (N_17,In_221,In_1882);
nor U18 (N_18,In_339,In_954);
or U19 (N_19,In_1235,In_218);
nor U20 (N_20,In_86,In_962);
and U21 (N_21,In_1165,In_809);
or U22 (N_22,In_1817,In_1801);
nand U23 (N_23,In_59,In_298);
and U24 (N_24,In_734,In_1064);
nor U25 (N_25,In_454,In_644);
or U26 (N_26,In_771,In_1397);
nand U27 (N_27,In_1896,In_102);
xnor U28 (N_28,In_916,In_742);
and U29 (N_29,In_1991,In_1298);
or U30 (N_30,In_562,In_401);
nor U31 (N_31,In_301,In_7);
and U32 (N_32,In_1996,In_1602);
or U33 (N_33,In_261,In_1259);
xnor U34 (N_34,In_1202,In_1657);
nand U35 (N_35,In_286,In_2);
and U36 (N_36,In_947,In_1403);
nand U37 (N_37,In_1861,In_941);
nor U38 (N_38,In_109,In_1154);
nand U39 (N_39,In_970,In_978);
nor U40 (N_40,In_1084,In_1052);
or U41 (N_41,In_800,In_1355);
and U42 (N_42,In_876,In_313);
or U43 (N_43,In_1646,In_212);
xor U44 (N_44,In_670,In_95);
nor U45 (N_45,In_1419,In_1106);
nand U46 (N_46,In_283,In_1457);
and U47 (N_47,In_1871,In_746);
and U48 (N_48,In_1062,In_1234);
xor U49 (N_49,In_482,In_1123);
and U50 (N_50,In_688,In_1237);
or U51 (N_51,In_429,In_654);
xnor U52 (N_52,In_1886,In_1576);
xnor U53 (N_53,In_126,In_70);
and U54 (N_54,In_91,In_1470);
nand U55 (N_55,In_1126,In_1200);
or U56 (N_56,In_651,In_1127);
xnor U57 (N_57,In_340,In_1409);
and U58 (N_58,In_616,In_696);
and U59 (N_59,In_323,In_289);
nor U60 (N_60,In_972,In_1056);
and U61 (N_61,In_1494,In_1310);
or U62 (N_62,In_1447,In_1515);
and U63 (N_63,In_1045,In_1505);
or U64 (N_64,In_1769,In_1044);
nand U65 (N_65,In_1158,In_216);
or U66 (N_66,In_1577,In_1752);
or U67 (N_67,In_1150,In_1253);
nand U68 (N_68,In_462,In_1879);
nor U69 (N_69,In_1124,In_117);
or U70 (N_70,In_1803,In_1219);
nand U71 (N_71,In_814,In_668);
nor U72 (N_72,In_1247,In_1584);
xnor U73 (N_73,In_1585,In_1443);
nand U74 (N_74,In_657,In_1361);
and U75 (N_75,In_1199,In_1797);
or U76 (N_76,In_1474,In_1408);
xnor U77 (N_77,In_1128,In_355);
xnor U78 (N_78,In_421,In_1710);
xnor U79 (N_79,In_1995,In_418);
nor U80 (N_80,In_1796,In_1183);
or U81 (N_81,In_1012,In_195);
nand U82 (N_82,In_428,In_88);
and U83 (N_83,In_1902,In_1016);
and U84 (N_84,In_1174,In_1853);
xor U85 (N_85,In_763,In_1700);
nand U86 (N_86,In_956,In_1628);
nand U87 (N_87,In_1347,In_567);
nand U88 (N_88,In_740,In_1907);
and U89 (N_89,In_1178,In_624);
xor U90 (N_90,In_394,In_1468);
and U91 (N_91,In_1566,In_1020);
xnor U92 (N_92,In_460,In_1812);
xnor U93 (N_93,In_1824,In_598);
nor U94 (N_94,In_1878,In_344);
nand U95 (N_95,In_1483,In_159);
nor U96 (N_96,In_958,In_123);
nor U97 (N_97,In_539,In_191);
nor U98 (N_98,In_158,In_1831);
and U99 (N_99,In_867,In_1737);
nor U100 (N_100,In_68,In_1077);
nand U101 (N_101,In_1673,In_773);
or U102 (N_102,In_1181,In_781);
xnor U103 (N_103,In_755,In_500);
and U104 (N_104,In_757,In_1192);
nand U105 (N_105,In_1205,In_107);
nor U106 (N_106,In_730,In_1724);
nand U107 (N_107,In_1810,In_1644);
and U108 (N_108,In_1023,In_292);
nand U109 (N_109,In_1645,In_1445);
nor U110 (N_110,In_1435,In_1735);
or U111 (N_111,In_1667,In_1004);
or U112 (N_112,In_503,In_424);
nand U113 (N_113,In_1155,In_78);
nand U114 (N_114,In_177,In_820);
nand U115 (N_115,In_264,In_186);
and U116 (N_116,In_1232,In_1627);
or U117 (N_117,In_1263,In_1706);
nor U118 (N_118,In_367,In_1481);
nor U119 (N_119,In_1327,In_165);
nand U120 (N_120,In_945,In_278);
xor U121 (N_121,In_1042,In_1742);
or U122 (N_122,In_853,In_439);
or U123 (N_123,In_173,In_402);
xnor U124 (N_124,In_134,In_1449);
nand U125 (N_125,In_903,In_1066);
and U126 (N_126,In_957,In_618);
or U127 (N_127,In_214,In_625);
xnor U128 (N_128,In_994,In_217);
or U129 (N_129,In_1252,In_1957);
and U130 (N_130,In_284,In_1081);
and U131 (N_131,In_331,In_1371);
or U132 (N_132,In_1575,In_735);
and U133 (N_133,In_101,In_921);
xnor U134 (N_134,In_891,In_341);
xor U135 (N_135,In_547,In_675);
or U136 (N_136,In_733,In_1619);
and U137 (N_137,In_67,In_1731);
nor U138 (N_138,In_12,In_1143);
xnor U139 (N_139,In_1523,In_1137);
nand U140 (N_140,In_1607,In_1911);
nand U141 (N_141,In_219,In_1388);
and U142 (N_142,In_443,In_1217);
nand U143 (N_143,In_1763,In_416);
nand U144 (N_144,In_775,In_1373);
nor U145 (N_145,In_606,In_1758);
and U146 (N_146,In_432,In_1663);
nor U147 (N_147,In_1550,In_1190);
nor U148 (N_148,In_1671,In_655);
and U149 (N_149,In_1580,In_119);
nand U150 (N_150,In_351,In_472);
or U151 (N_151,In_113,In_659);
nand U152 (N_152,In_1416,In_139);
or U153 (N_153,In_122,In_1276);
nand U154 (N_154,In_577,In_556);
xnor U155 (N_155,In_1959,In_155);
nand U156 (N_156,In_1581,In_1227);
nand U157 (N_157,In_1287,In_1753);
or U158 (N_158,In_437,In_1631);
nand U159 (N_159,In_727,In_1255);
nor U160 (N_160,In_1406,In_8);
nor U161 (N_161,In_1212,In_1517);
nand U162 (N_162,In_744,In_745);
nor U163 (N_163,In_1977,In_1510);
or U164 (N_164,In_810,In_1041);
or U165 (N_165,In_364,In_1475);
and U166 (N_166,In_234,In_441);
nor U167 (N_167,In_1551,In_300);
and U168 (N_168,In_888,In_1305);
and U169 (N_169,In_1153,In_1808);
nor U170 (N_170,In_1069,In_878);
and U171 (N_171,In_1083,In_1152);
nor U172 (N_172,In_20,In_1637);
nor U173 (N_173,In_1345,In_1442);
nor U174 (N_174,In_132,In_148);
or U175 (N_175,In_1650,In_619);
nand U176 (N_176,In_1132,In_789);
and U177 (N_177,In_1617,In_1144);
and U178 (N_178,In_373,In_1257);
nand U179 (N_179,In_188,In_581);
or U180 (N_180,In_1620,In_984);
nand U181 (N_181,In_1961,In_150);
xor U182 (N_182,In_321,In_807);
or U183 (N_183,In_386,In_266);
nor U184 (N_184,In_1433,In_1821);
and U185 (N_185,In_1177,In_1883);
or U186 (N_186,In_152,In_345);
nand U187 (N_187,In_1254,In_516);
or U188 (N_188,In_1337,In_365);
or U189 (N_189,In_1010,In_1989);
nand U190 (N_190,In_1778,In_719);
nor U191 (N_191,In_1353,In_739);
nand U192 (N_192,In_143,In_1071);
or U193 (N_193,In_580,In_988);
nor U194 (N_194,In_538,In_812);
xor U195 (N_195,In_1203,In_1274);
and U196 (N_196,In_517,In_633);
nand U197 (N_197,In_447,In_1262);
and U198 (N_198,In_1036,In_1526);
nand U199 (N_199,In_377,In_950);
xor U200 (N_200,In_1591,In_1895);
xor U201 (N_201,In_642,In_1198);
nand U202 (N_202,In_1926,In_783);
xor U203 (N_203,In_1113,In_667);
xnor U204 (N_204,In_1809,In_1221);
nor U205 (N_205,In_1962,In_1107);
or U206 (N_206,In_981,In_1011);
nand U207 (N_207,In_130,In_845);
nand U208 (N_208,In_6,In_1890);
nand U209 (N_209,In_1556,In_259);
nor U210 (N_210,In_378,In_720);
and U211 (N_211,In_1691,In_1649);
nor U212 (N_212,In_494,In_1430);
nor U213 (N_213,In_1857,In_1389);
and U214 (N_214,In_393,In_290);
nand U215 (N_215,In_647,In_1102);
nor U216 (N_216,In_1451,In_1988);
nand U217 (N_217,In_1944,In_1592);
nor U218 (N_218,In_382,In_430);
or U219 (N_219,In_1208,In_699);
xnor U220 (N_220,In_174,In_162);
or U221 (N_221,In_963,In_678);
or U222 (N_222,In_198,In_1324);
or U223 (N_223,In_1354,In_1394);
or U224 (N_224,In_453,In_1296);
nor U225 (N_225,In_1937,In_1231);
xnor U226 (N_226,In_834,In_164);
nor U227 (N_227,In_49,In_293);
or U228 (N_228,In_765,In_1586);
nand U229 (N_229,In_1372,In_395);
and U230 (N_230,In_1643,In_1967);
or U231 (N_231,In_1846,In_163);
xor U232 (N_232,In_566,In_1173);
nand U233 (N_233,In_1067,In_672);
nor U234 (N_234,In_1424,In_1176);
nor U235 (N_235,In_1286,In_523);
or U236 (N_236,In_711,In_752);
or U237 (N_237,In_767,In_1518);
xnor U238 (N_238,In_1930,In_1179);
nor U239 (N_239,In_1462,In_388);
or U240 (N_240,In_1079,In_229);
or U241 (N_241,In_451,In_248);
and U242 (N_242,In_872,In_885);
xor U243 (N_243,In_1877,In_1514);
and U244 (N_244,In_1716,In_1788);
nor U245 (N_245,In_26,In_1000);
xnor U246 (N_246,In_125,In_1754);
xor U247 (N_247,In_1683,In_305);
nand U248 (N_248,In_759,In_1486);
nand U249 (N_249,In_1032,In_37);
and U250 (N_250,In_1065,In_960);
nand U251 (N_251,In_934,In_729);
or U252 (N_252,In_156,In_1794);
xor U253 (N_253,In_1479,In_721);
or U254 (N_254,In_1463,In_1686);
nand U255 (N_255,In_1238,In_1315);
xor U256 (N_256,In_223,In_1530);
nor U257 (N_257,In_1903,In_483);
nand U258 (N_258,In_1215,In_1674);
xnor U259 (N_259,In_435,In_705);
xnor U260 (N_260,In_1312,In_491);
nand U261 (N_261,In_80,In_652);
nor U262 (N_262,In_732,In_1555);
nor U263 (N_263,In_777,In_222);
nor U264 (N_264,In_1987,In_1539);
nand U265 (N_265,In_1092,In_1822);
and U266 (N_266,In_875,In_1135);
or U267 (N_267,In_330,In_154);
nand U268 (N_268,In_1418,In_239);
nand U269 (N_269,In_179,In_1832);
nor U270 (N_270,In_477,In_1516);
xnor U271 (N_271,In_142,In_1851);
or U272 (N_272,In_1080,In_1059);
nor U273 (N_273,In_1367,In_816);
or U274 (N_274,In_1326,In_1058);
and U275 (N_275,In_683,In_992);
nand U276 (N_276,In_1201,In_748);
nand U277 (N_277,In_509,In_691);
xnor U278 (N_278,In_622,In_660);
nor U279 (N_279,In_1171,In_533);
or U280 (N_280,In_400,In_227);
xor U281 (N_281,In_1746,In_1913);
nor U282 (N_282,In_1090,In_641);
nand U283 (N_283,In_1019,In_852);
xor U284 (N_284,In_1999,In_948);
nand U285 (N_285,In_325,In_209);
nand U286 (N_286,In_192,In_907);
xnor U287 (N_287,In_35,In_27);
or U288 (N_288,In_955,In_1715);
or U289 (N_289,In_1444,In_207);
and U290 (N_290,In_1701,In_1151);
and U291 (N_291,In_1185,In_1960);
nor U292 (N_292,In_1112,In_111);
and U293 (N_293,In_927,In_635);
or U294 (N_294,In_1393,In_228);
or U295 (N_295,In_1348,In_610);
and U296 (N_296,In_1108,In_342);
and U297 (N_297,In_1751,In_793);
nor U298 (N_298,In_1148,In_1615);
xnor U299 (N_299,In_66,In_495);
xnor U300 (N_300,In_784,In_846);
nor U301 (N_301,In_1705,In_361);
or U302 (N_302,In_11,In_564);
xor U303 (N_303,In_436,In_178);
and U304 (N_304,In_1626,In_1209);
or U305 (N_305,In_913,In_1888);
nor U306 (N_306,In_1230,In_674);
nand U307 (N_307,In_986,In_138);
or U308 (N_308,In_206,In_1014);
and U309 (N_309,In_1325,In_1986);
and U310 (N_310,In_480,In_1480);
and U311 (N_311,In_684,In_1780);
nand U312 (N_312,In_1269,In_1495);
nand U313 (N_313,In_605,In_1792);
and U314 (N_314,In_1411,In_1594);
nand U315 (N_315,In_1546,In_1425);
or U316 (N_316,In_1980,In_90);
nor U317 (N_317,In_1867,In_584);
nand U318 (N_318,In_1893,In_1501);
or U319 (N_319,In_458,In_1121);
xor U320 (N_320,In_609,In_1122);
nor U321 (N_321,In_1417,In_1027);
or U322 (N_322,In_1811,In_521);
xor U323 (N_323,In_1918,In_1382);
xor U324 (N_324,In_1119,In_1309);
and U325 (N_325,In_57,In_1826);
or U326 (N_326,In_1161,In_1740);
and U327 (N_327,In_303,In_842);
and U328 (N_328,In_1346,In_1783);
or U329 (N_329,In_1929,In_1224);
xor U330 (N_330,In_116,In_1454);
and U331 (N_331,In_1243,In_700);
nand U332 (N_332,In_724,In_354);
or U333 (N_333,In_362,In_285);
nor U334 (N_334,In_679,In_526);
or U335 (N_335,In_717,In_985);
and U336 (N_336,In_79,In_1665);
or U337 (N_337,In_316,In_24);
xnor U338 (N_338,In_136,In_637);
xor U339 (N_339,In_1789,In_1549);
or U340 (N_340,In_1927,In_1864);
nand U341 (N_341,In_829,In_1750);
nand U342 (N_342,In_1025,In_270);
nand U343 (N_343,In_1170,In_894);
or U344 (N_344,In_1698,In_1146);
and U345 (N_345,In_302,In_998);
nor U346 (N_346,In_244,In_589);
or U347 (N_347,In_1304,In_1050);
nand U348 (N_348,In_1914,In_1847);
nand U349 (N_349,In_1567,In_1129);
and U350 (N_350,In_1116,In_245);
and U351 (N_351,In_258,In_1815);
nand U352 (N_352,In_1855,In_1924);
and U353 (N_353,In_1689,In_1806);
nand U354 (N_354,In_336,In_695);
nor U355 (N_355,In_525,In_385);
xor U356 (N_356,In_201,In_1975);
nor U357 (N_357,In_280,In_249);
nor U358 (N_358,In_1362,In_230);
nand U359 (N_359,In_318,In_979);
or U360 (N_360,In_836,In_358);
nand U361 (N_361,In_1863,In_1755);
xnor U362 (N_362,In_128,In_1876);
xnor U363 (N_363,In_764,In_1708);
or U364 (N_364,In_455,In_706);
or U365 (N_365,In_1917,In_236);
or U366 (N_366,In_596,In_1568);
or U367 (N_367,In_1819,In_976);
or U368 (N_368,In_1484,In_1082);
nor U369 (N_369,In_1078,In_808);
xor U370 (N_370,In_912,In_1563);
nor U371 (N_371,In_1035,In_1175);
nand U372 (N_372,In_1574,In_260);
nand U373 (N_373,In_750,In_1509);
nor U374 (N_374,In_99,In_61);
nor U375 (N_375,In_1384,In_1095);
and U376 (N_376,In_1068,In_64);
or U377 (N_377,In_127,In_1328);
nor U378 (N_378,In_928,In_528);
or U379 (N_379,In_1557,In_1965);
xnor U380 (N_380,In_213,In_1005);
and U381 (N_381,In_1843,In_648);
or U382 (N_382,In_1653,In_54);
or U383 (N_383,In_1820,In_508);
xor U384 (N_384,In_1464,In_131);
nor U385 (N_385,In_1997,In_1642);
nor U386 (N_386,In_1497,In_55);
and U387 (N_387,In_1094,In_1168);
and U388 (N_388,In_1900,In_553);
or U389 (N_389,In_881,In_1765);
nor U390 (N_390,In_89,In_1038);
and U391 (N_391,In_287,In_936);
nor U392 (N_392,In_1640,In_1603);
xnor U393 (N_393,In_1402,In_1441);
nand U394 (N_394,In_1491,In_43);
nor U395 (N_395,In_268,In_319);
nor U396 (N_396,In_621,In_1839);
and U397 (N_397,In_628,In_1489);
and U398 (N_398,In_357,In_1834);
xor U399 (N_399,In_604,In_1983);
nor U400 (N_400,In_53,In_271);
and U401 (N_401,In_1682,In_576);
xor U402 (N_402,In_1429,In_1955);
and U403 (N_403,In_1320,In_81);
nand U404 (N_404,In_1541,In_1376);
and U405 (N_405,In_1508,In_1452);
xnor U406 (N_406,In_833,In_1573);
nor U407 (N_407,In_1048,In_1450);
xnor U408 (N_408,In_1422,In_623);
xnor U409 (N_409,In_1164,In_1085);
xor U410 (N_410,In_1725,In_1629);
nand U411 (N_411,In_1786,In_1841);
or U412 (N_412,In_1115,In_368);
nor U413 (N_413,In_895,In_1958);
or U414 (N_414,In_1726,In_1942);
xnor U415 (N_415,In_1934,In_1404);
nor U416 (N_416,In_1003,In_524);
nor U417 (N_417,In_1558,In_277);
and U418 (N_418,In_692,In_519);
and U419 (N_419,In_419,In_1856);
xor U420 (N_420,In_1736,In_308);
and U421 (N_421,In_502,In_663);
or U422 (N_422,In_1340,In_44);
xnor U423 (N_423,In_1941,In_82);
nor U424 (N_424,In_1933,In_431);
or U425 (N_425,In_937,In_993);
nor U426 (N_426,In_1828,In_532);
xnor U427 (N_427,In_1350,In_426);
xor U428 (N_428,In_1264,In_1378);
and U429 (N_429,In_1676,In_681);
and U430 (N_430,In_1721,In_499);
or U431 (N_431,In_1915,In_702);
nand U432 (N_432,In_1172,In_1912);
nand U433 (N_433,In_788,In_756);
nand U434 (N_434,In_738,In_1583);
or U435 (N_435,In_369,In_473);
or U436 (N_436,In_1157,In_1842);
nand U437 (N_437,In_1459,In_1145);
or U438 (N_438,In_1836,In_17);
nor U439 (N_439,In_1992,In_886);
nand U440 (N_440,In_22,In_5);
or U441 (N_441,In_1482,In_574);
nand U442 (N_442,In_1687,In_487);
nor U443 (N_443,In_791,In_1948);
nand U444 (N_444,In_1825,In_1935);
nand U445 (N_445,In_1385,In_327);
and U446 (N_446,In_243,In_396);
and U447 (N_447,In_1428,In_1225);
xor U448 (N_448,In_1823,In_841);
or U449 (N_449,In_507,In_685);
xnor U450 (N_450,In_815,In_1311);
and U451 (N_451,In_1777,In_1141);
nor U452 (N_452,In_422,In_1471);
nand U453 (N_453,In_1297,In_1946);
and U454 (N_454,In_819,In_1655);
and U455 (N_455,In_896,In_1600);
or U456 (N_456,In_922,In_40);
and U457 (N_457,In_1533,In_247);
and U458 (N_458,In_558,In_1981);
and U459 (N_459,In_1446,In_1290);
nor U460 (N_460,In_1887,In_1030);
nand U461 (N_461,In_1921,In_626);
nor U462 (N_462,In_1859,In_1307);
and U463 (N_463,In_38,In_1791);
nor U464 (N_464,In_1002,In_105);
nand U465 (N_465,In_62,In_1195);
or U466 (N_466,In_890,In_786);
nor U467 (N_467,In_1420,In_1054);
nand U468 (N_468,In_1938,In_1432);
xnor U469 (N_469,In_726,In_1985);
and U470 (N_470,In_1816,In_559);
or U471 (N_471,In_1493,In_1246);
nor U472 (N_472,In_952,In_1381);
and U473 (N_473,In_1873,In_1538);
nand U474 (N_474,In_1668,In_1009);
xor U475 (N_475,In_1739,In_1738);
xor U476 (N_476,In_1291,In_982);
xnor U477 (N_477,In_1399,In_599);
or U478 (N_478,In_463,In_32);
nand U479 (N_479,In_639,In_794);
or U480 (N_480,In_18,In_411);
or U481 (N_481,In_238,In_172);
and U482 (N_482,In_1216,In_792);
nor U483 (N_483,In_255,In_1461);
xnor U484 (N_484,In_632,In_1063);
nand U485 (N_485,In_13,In_1971);
or U486 (N_486,In_701,In_1073);
nand U487 (N_487,In_3,In_202);
or U488 (N_488,In_629,In_1017);
nor U489 (N_489,In_1018,In_935);
nand U490 (N_490,In_811,In_909);
and U491 (N_491,In_827,In_1322);
and U492 (N_492,In_310,In_1271);
or U493 (N_493,In_1537,In_215);
nand U494 (N_494,In_157,In_1970);
and U495 (N_495,In_680,In_1395);
nand U496 (N_496,In_546,In_1414);
xnor U497 (N_497,In_1329,In_1249);
nor U498 (N_498,In_1953,In_446);
nand U499 (N_499,In_656,In_1616);
or U500 (N_500,In_1460,In_1245);
nor U501 (N_501,In_1097,In_1734);
or U502 (N_502,In_92,In_571);
nor U503 (N_503,In_504,In_1720);
nand U504 (N_504,In_554,In_366);
or U505 (N_505,In_1256,In_669);
and U506 (N_506,In_870,In_1308);
xnor U507 (N_507,In_687,In_415);
xnor U508 (N_508,In_1605,In_762);
and U509 (N_509,In_135,In_391);
xor U510 (N_510,In_1588,In_1284);
nand U511 (N_511,In_1401,In_1110);
or U512 (N_512,In_1519,In_288);
nor U513 (N_513,In_718,In_475);
nand U514 (N_514,In_1940,In_552);
xor U515 (N_515,In_592,In_594);
nand U516 (N_516,In_1952,In_898);
xnor U517 (N_517,In_796,In_501);
and U518 (N_518,In_995,In_1661);
and U519 (N_519,In_1265,In_1439);
or U520 (N_520,In_689,In_860);
xnor U521 (N_521,In_1169,In_295);
xor U522 (N_522,In_39,In_1579);
and U523 (N_523,In_1436,In_1167);
nor U524 (N_524,In_1507,In_1524);
or U525 (N_525,In_1838,In_1850);
nand U526 (N_526,In_1542,In_1596);
and U527 (N_527,In_543,In_118);
nand U528 (N_528,In_779,In_1438);
or U529 (N_529,In_866,In_1885);
and U530 (N_530,In_1207,In_944);
nand U531 (N_531,In_1105,In_953);
xor U532 (N_532,In_601,In_1595);
nand U533 (N_533,In_863,In_591);
or U534 (N_534,In_1976,In_1894);
xnor U535 (N_535,In_1680,In_1651);
xnor U536 (N_536,In_1511,In_1088);
nor U537 (N_537,In_274,In_1852);
nor U538 (N_538,In_1624,In_1660);
and U539 (N_539,In_1390,In_448);
and U540 (N_540,In_946,In_203);
nor U541 (N_541,In_906,In_1761);
nand U542 (N_542,In_1488,In_1670);
xor U543 (N_543,In_476,In_661);
and U544 (N_544,In_208,In_1904);
xor U545 (N_545,In_990,In_1781);
nor U546 (N_546,In_50,In_555);
or U547 (N_547,In_858,In_918);
nand U548 (N_548,In_297,In_464);
and U549 (N_549,In_1380,In_199);
and U550 (N_550,In_1260,In_557);
or U551 (N_551,In_693,In_1866);
nand U552 (N_552,In_1741,In_1131);
or U553 (N_553,In_124,In_1248);
nand U554 (N_554,In_404,In_1210);
or U555 (N_555,In_1982,In_645);
nand U556 (N_556,In_406,In_1331);
or U557 (N_557,In_511,In_1969);
nand U558 (N_558,In_108,In_231);
nand U559 (N_559,In_370,In_376);
or U560 (N_560,In_823,In_1335);
nor U561 (N_561,In_1278,In_1344);
nand U562 (N_562,In_1748,In_232);
nor U563 (N_563,In_1678,In_780);
xnor U564 (N_564,In_1925,In_880);
and U565 (N_565,In_991,In_1572);
and U566 (N_566,In_714,In_256);
and U567 (N_567,In_877,In_1717);
and U568 (N_568,In_795,In_241);
or U569 (N_569,In_1766,In_42);
nand U570 (N_570,In_837,In_1244);
nand U571 (N_571,In_1364,In_749);
and U572 (N_572,In_1696,In_686);
nand U573 (N_573,In_1881,In_1898);
nor U574 (N_574,In_931,In_56);
and U575 (N_575,In_1949,In_551);
and U576 (N_576,In_1529,In_452);
or U577 (N_577,In_578,In_1267);
or U578 (N_578,In_237,In_817);
nor U579 (N_579,In_1652,In_787);
nand U580 (N_580,In_1076,In_112);
or U581 (N_581,In_1314,In_1188);
nand U582 (N_582,In_856,In_1854);
nand U583 (N_583,In_1339,In_493);
xor U584 (N_584,In_183,In_1302);
nor U585 (N_585,In_346,In_1695);
or U586 (N_586,In_704,In_1049);
and U587 (N_587,In_465,In_634);
and U588 (N_588,In_1589,In_772);
xor U589 (N_589,In_193,In_1487);
xnor U590 (N_590,In_1101,In_568);
or U591 (N_591,In_225,In_1046);
nor U592 (N_592,In_315,In_347);
or U593 (N_593,In_813,In_144);
and U594 (N_594,In_246,In_1901);
or U595 (N_595,In_843,In_973);
and U596 (N_596,In_1702,In_168);
or U597 (N_597,In_1300,In_85);
or U598 (N_598,In_1552,In_760);
nand U599 (N_599,In_925,In_676);
xnor U600 (N_600,In_488,In_868);
or U601 (N_601,In_531,In_869);
xor U602 (N_602,In_1391,In_910);
nand U603 (N_603,In_170,In_1086);
nand U604 (N_604,In_1675,In_1333);
and U605 (N_605,In_337,In_999);
and U606 (N_606,In_299,In_1366);
nand U607 (N_607,In_600,In_897);
nor U608 (N_608,In_71,In_1679);
nand U609 (N_609,In_636,In_1956);
and U610 (N_610,In_971,In_514);
xor U611 (N_611,In_1684,In_1047);
xor U612 (N_612,In_384,In_196);
nor U613 (N_613,In_110,In_939);
and U614 (N_614,In_1978,In_1499);
and U615 (N_615,In_1437,In_1635);
nor U616 (N_616,In_1279,In_176);
nand U617 (N_617,In_798,In_1609);
xor U618 (N_618,In_72,In_864);
or U619 (N_619,In_854,In_36);
and U620 (N_620,In_908,In_1273);
and U621 (N_621,In_349,In_282);
nand U622 (N_622,In_797,In_1392);
nor U623 (N_623,In_920,In_121);
or U624 (N_624,In_343,In_1109);
or U625 (N_625,In_169,In_803);
and U626 (N_626,In_904,In_515);
xnor U627 (N_627,In_1166,In_360);
nand U628 (N_628,In_1213,In_326);
nand U629 (N_629,In_530,In_332);
or U630 (N_630,In_1415,In_1964);
and U631 (N_631,In_1332,In_996);
or U632 (N_632,In_1013,In_1440);
xor U633 (N_633,In_1317,In_1939);
nor U634 (N_634,In_997,In_1184);
nor U635 (N_635,In_272,In_1703);
or U636 (N_636,In_363,In_390);
and U637 (N_637,In_1984,In_1469);
nand U638 (N_638,In_1026,In_235);
xor U639 (N_639,In_1553,In_1564);
or U640 (N_640,In_1147,In_1621);
nand U641 (N_641,In_1531,In_87);
xnor U642 (N_642,In_16,In_1156);
nand U643 (N_643,In_490,In_1467);
xnor U644 (N_644,In_1560,In_1759);
xor U645 (N_645,In_905,In_1294);
or U646 (N_646,In_1053,In_611);
or U647 (N_647,In_23,In_470);
and U648 (N_648,In_1099,In_505);
xnor U649 (N_649,In_650,In_1140);
and U650 (N_650,In_474,In_1096);
and U651 (N_651,In_1528,In_1139);
nor U652 (N_652,In_1220,In_324);
or U653 (N_653,In_1535,In_1001);
nor U654 (N_654,In_915,In_573);
nand U655 (N_655,In_1562,In_1945);
or U656 (N_656,In_537,In_1707);
or U657 (N_657,In_296,In_1659);
and U658 (N_658,In_445,In_534);
xor U659 (N_659,In_413,In_1920);
nand U660 (N_660,In_716,In_917);
nor U661 (N_661,In_1386,In_1500);
and U662 (N_662,In_713,In_1875);
xnor U663 (N_663,In_420,In_252);
nand U664 (N_664,In_804,In_83);
nor U665 (N_665,In_58,In_1543);
or U666 (N_666,In_1973,In_1862);
or U667 (N_667,In_983,In_114);
xor U668 (N_668,In_506,In_1222);
nor U669 (N_669,In_1634,In_838);
and U670 (N_670,In_334,In_929);
nor U671 (N_671,In_312,In_968);
nor U672 (N_672,In_1547,In_73);
nor U673 (N_673,In_459,In_1943);
nor U674 (N_674,In_96,In_1377);
xor U675 (N_675,In_1599,In_840);
xnor U676 (N_676,In_389,In_1732);
nand U677 (N_677,In_262,In_1601);
and U678 (N_678,In_1319,In_359);
nand U679 (N_679,In_640,In_1923);
nor U680 (N_680,In_1341,In_671);
xor U681 (N_681,In_1756,In_1614);
nor U682 (N_682,In_627,In_1623);
nor U683 (N_683,In_1767,In_31);
or U684 (N_684,In_653,In_311);
nor U685 (N_685,In_1704,In_1204);
or U686 (N_686,In_1357,In_1880);
nor U687 (N_687,In_1149,In_587);
or U688 (N_688,In_1028,In_1906);
nor U689 (N_689,In_1534,In_824);
or U690 (N_690,In_1527,In_1764);
and U691 (N_691,In_1688,In_1611);
nand U692 (N_692,In_1908,In_1138);
nand U693 (N_693,In_279,In_964);
xor U694 (N_694,In_1196,In_1830);
or U695 (N_695,In_1288,In_1021);
nand U696 (N_696,In_930,In_25);
or U697 (N_697,In_751,In_1087);
and U698 (N_698,In_408,In_291);
nor U699 (N_699,In_211,In_643);
nor U700 (N_700,In_1496,In_563);
nand U701 (N_701,In_251,In_575);
and U702 (N_702,In_1261,In_1837);
nor U703 (N_703,In_1770,In_1303);
nor U704 (N_704,In_826,In_1360);
nand U705 (N_705,In_469,In_1292);
nor U706 (N_706,In_549,In_141);
xor U707 (N_707,In_1598,In_322);
nand U708 (N_708,In_253,In_1033);
nand U709 (N_709,In_1947,In_1711);
nor U710 (N_710,In_1472,In_873);
nor U711 (N_711,In_1162,In_166);
nor U712 (N_712,In_21,In_19);
nor U713 (N_713,In_673,In_1762);
and U714 (N_714,In_1677,In_708);
or U715 (N_715,In_617,In_1072);
xnor U716 (N_716,In_1972,In_1666);
or U717 (N_717,In_309,In_1299);
nor U718 (N_718,In_1936,In_1833);
nor U719 (N_719,In_1318,In_1681);
and U720 (N_720,In_46,In_348);
and U721 (N_721,In_387,In_542);
nand U722 (N_722,In_602,In_1692);
or U723 (N_723,In_47,In_690);
or U724 (N_724,In_1633,In_374);
xor U725 (N_725,In_522,In_276);
nor U726 (N_726,In_479,In_940);
or U727 (N_727,In_467,In_1396);
xnor U728 (N_728,In_747,In_1757);
nand U729 (N_729,In_1295,In_1790);
xor U730 (N_730,In_1690,In_932);
and U731 (N_731,In_879,In_1928);
or U732 (N_732,In_1473,In_649);
xnor U733 (N_733,In_1277,In_1272);
xnor U734 (N_734,In_1187,In_1979);
nor U735 (N_735,In_267,In_709);
nand U736 (N_736,In_847,In_182);
nor U737 (N_737,In_1186,In_1359);
and U738 (N_738,In_1503,In_862);
or U739 (N_739,In_161,In_1569);
nor U740 (N_740,In_1434,In_254);
nand U741 (N_741,In_1343,In_1398);
or U742 (N_742,In_1379,In_1648);
xor U743 (N_743,In_1829,In_1521);
and U744 (N_744,In_901,In_189);
and U745 (N_745,In_828,In_588);
xnor U746 (N_746,In_806,In_565);
nor U747 (N_747,In_275,In_1849);
nor U748 (N_748,In_33,In_1730);
nand U749 (N_749,In_220,In_1476);
nor U750 (N_750,In_664,In_975);
or U751 (N_751,In_933,In_204);
nand U752 (N_752,In_153,In_1358);
and U753 (N_753,In_899,In_1120);
and U754 (N_754,In_449,In_1197);
nand U755 (N_755,In_919,In_1431);
and U756 (N_756,In_741,In_969);
nor U757 (N_757,In_69,In_471);
nor U758 (N_758,In_582,In_1352);
nand U759 (N_759,In_1282,In_1593);
and U760 (N_760,In_902,In_871);
nor U761 (N_761,In_1251,In_1745);
nand U762 (N_762,In_1407,In_84);
and U763 (N_763,In_989,In_1775);
or U764 (N_764,In_94,In_65);
or U765 (N_765,In_492,In_825);
xor U766 (N_766,In_512,In_725);
and U767 (N_767,In_4,In_1891);
nand U768 (N_768,In_1250,In_1306);
nand U769 (N_769,In_306,In_433);
and U770 (N_770,In_1874,In_801);
or U771 (N_771,In_184,In_1793);
and U772 (N_772,In_923,In_924);
xnor U773 (N_773,In_1142,In_620);
and U774 (N_774,In_405,In_535);
nand U775 (N_775,In_1536,In_461);
xor U776 (N_776,In_1641,In_1498);
and U777 (N_777,In_615,In_1919);
xor U778 (N_778,In_1540,In_147);
nand U779 (N_779,In_1884,In_160);
or U780 (N_780,In_1034,In_614);
nor U781 (N_781,In_29,In_743);
nand U782 (N_782,In_1427,In_938);
nand U783 (N_783,In_1374,In_1743);
xnor U784 (N_784,In_540,In_1075);
xnor U785 (N_785,In_379,In_1571);
xnor U786 (N_786,In_1125,In_722);
or U787 (N_787,In_129,In_1694);
or U788 (N_788,In_603,In_770);
or U789 (N_789,In_1712,In_1280);
nor U790 (N_790,In_1870,In_857);
and U791 (N_791,In_1916,In_1301);
xnor U792 (N_792,In_317,In_423);
nor U793 (N_793,In_1387,In_520);
xor U794 (N_794,In_1114,In_1134);
xnor U795 (N_795,In_1779,In_851);
xor U796 (N_796,In_892,In_77);
nor U797 (N_797,In_1827,In_1513);
or U798 (N_798,In_712,In_1313);
xor U799 (N_799,In_1465,In_1336);
and U800 (N_800,In_381,In_1578);
nor U801 (N_801,N_552,N_615);
nor U802 (N_802,N_273,N_621);
nand U803 (N_803,N_74,N_284);
nor U804 (N_804,In_1805,N_163);
nor U805 (N_805,N_763,N_712);
xnor U806 (N_806,N_317,N_183);
nand U807 (N_807,N_59,N_41);
or U808 (N_808,N_351,In_180);
or U809 (N_809,N_504,N_334);
nand U810 (N_810,N_745,N_409);
nand U811 (N_811,N_216,N_397);
nor U812 (N_812,N_398,N_758);
xnor U813 (N_813,N_111,In_410);
and U814 (N_814,In_1993,N_90);
nor U815 (N_815,N_446,N_270);
and U816 (N_816,N_73,N_707);
xnor U817 (N_817,N_139,N_45);
nor U818 (N_818,N_102,N_61);
nand U819 (N_819,N_31,N_765);
nor U820 (N_820,In_593,N_126);
nor U821 (N_821,N_248,N_116);
or U822 (N_822,N_452,N_283);
and U823 (N_823,N_559,N_637);
xnor U824 (N_824,N_201,N_750);
nor U825 (N_825,N_547,N_88);
nand U826 (N_826,N_115,In_338);
nand U827 (N_827,N_239,In_987);
xor U828 (N_828,N_144,N_186);
or U829 (N_829,N_301,In_240);
nand U830 (N_830,N_87,N_214);
nor U831 (N_831,In_1845,In_658);
or U832 (N_832,In_1905,N_612);
xnor U833 (N_833,In_758,N_225);
nor U834 (N_834,In_438,In_1093);
and U835 (N_835,In_1051,N_483);
xnor U836 (N_836,In_1722,N_625);
or U837 (N_837,In_1587,N_303);
xor U838 (N_838,N_647,In_1848);
and U839 (N_839,In_1061,In_774);
xor U840 (N_840,In_1749,N_674);
or U841 (N_841,N_319,N_282);
and U842 (N_842,In_1714,N_480);
xnor U843 (N_843,N_627,N_222);
nand U844 (N_844,N_584,N_749);
or U845 (N_845,N_434,N_680);
xnor U846 (N_846,In_145,N_691);
nand U847 (N_847,In_1525,In_403);
nor U848 (N_848,N_292,N_243);
xor U849 (N_849,In_597,In_832);
and U850 (N_850,N_320,N_436);
nand U851 (N_851,In_723,In_466);
or U852 (N_852,N_729,N_510);
nand U853 (N_853,N_575,N_205);
nor U854 (N_854,In_1813,N_390);
and U855 (N_855,N_422,N_375);
xor U856 (N_856,In_328,N_230);
nor U857 (N_857,In_171,N_541);
xnor U858 (N_858,N_98,N_596);
nand U859 (N_859,N_196,N_240);
and U860 (N_860,N_394,N_178);
and U861 (N_861,In_1768,N_356);
and U862 (N_862,N_302,In_1685);
and U863 (N_863,N_556,N_430);
or U864 (N_864,In_1006,N_4);
or U865 (N_865,N_700,In_1559);
and U866 (N_866,N_259,N_321);
xor U867 (N_867,In_1206,N_340);
or U868 (N_868,N_215,N_221);
or U869 (N_869,N_384,In_1365);
nor U870 (N_870,N_734,In_638);
xor U871 (N_871,N_56,In_265);
nand U872 (N_872,N_413,In_1323);
nor U873 (N_873,N_453,In_1159);
or U874 (N_874,In_75,N_162);
nand U875 (N_875,N_253,N_173);
xnor U876 (N_876,In_761,N_553);
or U877 (N_877,N_412,N_92);
and U878 (N_878,N_79,In_1117);
nand U879 (N_879,In_478,In_106);
nor U880 (N_880,N_120,N_437);
and U881 (N_881,N_523,N_258);
or U882 (N_882,N_330,In_961);
or U883 (N_883,N_264,N_508);
or U884 (N_884,N_166,N_439);
and U885 (N_885,In_224,In_1776);
nor U886 (N_886,N_269,N_193);
and U887 (N_887,N_445,In_1456);
xor U888 (N_888,In_1658,In_665);
or U889 (N_889,N_316,In_822);
or U890 (N_890,N_308,N_160);
or U891 (N_891,N_313,In_45);
nand U892 (N_892,In_371,N_684);
nor U893 (N_893,In_98,N_624);
nor U894 (N_894,N_641,N_677);
and U895 (N_895,N_488,N_311);
nor U896 (N_896,N_156,In_1029);
nand U897 (N_897,N_668,N_479);
xor U898 (N_898,N_753,In_1040);
and U899 (N_899,N_325,N_182);
and U900 (N_900,N_14,In_510);
nand U901 (N_901,N_223,N_507);
or U902 (N_902,In_646,In_737);
or U903 (N_903,N_326,N_564);
nand U904 (N_904,In_1242,In_1492);
and U905 (N_905,N_318,In_1618);
and U906 (N_906,In_1872,N_286);
nor U907 (N_907,In_425,In_1211);
nand U908 (N_908,In_210,N_477);
or U909 (N_909,N_227,N_371);
nor U910 (N_910,N_337,N_678);
nor U911 (N_911,N_352,N_295);
and U912 (N_912,N_212,N_535);
xor U913 (N_913,In_60,N_457);
nand U914 (N_914,In_560,N_487);
nor U915 (N_915,In_51,In_850);
or U916 (N_916,N_148,N_154);
nand U917 (N_917,N_406,N_796);
xor U918 (N_918,In_1860,N_360);
or U919 (N_919,N_611,In_682);
xor U920 (N_920,In_450,N_26);
or U921 (N_921,In_1289,N_66);
or U922 (N_922,In_175,N_517);
or U923 (N_923,In_398,N_592);
or U924 (N_924,N_132,In_383);
and U925 (N_925,In_52,N_601);
and U926 (N_926,In_1889,N_312);
and U927 (N_927,N_27,In_1283);
and U928 (N_928,N_172,N_123);
or U929 (N_929,In_544,N_521);
or U930 (N_930,N_107,In_1410);
or U931 (N_931,N_792,N_599);
xnor U932 (N_932,N_623,N_181);
xor U933 (N_933,In_1664,N_95);
nand U934 (N_934,In_185,N_786);
or U935 (N_935,In_1545,N_714);
and U936 (N_936,In_434,N_702);
and U937 (N_937,N_235,N_708);
or U938 (N_938,N_81,N_490);
xnor U939 (N_939,In_233,In_889);
nor U940 (N_940,N_538,N_137);
and U941 (N_941,N_261,N_471);
or U942 (N_942,N_740,N_22);
or U943 (N_943,N_660,N_654);
nand U944 (N_944,N_83,In_427);
xor U945 (N_945,N_768,N_444);
nand U946 (N_946,In_486,N_285);
or U947 (N_947,N_739,N_664);
or U948 (N_948,N_676,In_1522);
and U949 (N_949,N_722,N_287);
and U950 (N_950,In_859,N_655);
nand U951 (N_951,N_733,In_1622);
nand U952 (N_952,N_373,N_233);
nand U953 (N_953,N_28,In_352);
nor U954 (N_954,N_419,N_544);
and U955 (N_955,In_914,In_1293);
nor U956 (N_956,N_590,N_131);
xor U957 (N_957,In_790,In_782);
xor U958 (N_958,N_701,In_34);
or U959 (N_959,N_299,In_1639);
or U960 (N_960,In_579,In_1031);
or U961 (N_961,N_401,In_414);
nor U962 (N_962,N_392,N_728);
nor U963 (N_963,N_628,In_778);
xnor U964 (N_964,In_677,N_494);
nor U965 (N_965,In_818,In_187);
xnor U966 (N_966,N_595,In_776);
xnor U967 (N_967,In_14,N_11);
xnor U968 (N_968,N_774,In_226);
or U969 (N_969,In_1426,N_602);
nand U970 (N_970,N_463,In_613);
xnor U971 (N_971,N_78,N_106);
nand U972 (N_972,N_638,N_32);
xor U973 (N_973,N_242,In_548);
or U974 (N_974,N_249,N_208);
xor U975 (N_975,N_607,N_174);
nand U976 (N_976,N_353,N_626);
xnor U977 (N_977,N_686,N_291);
and U978 (N_978,N_403,N_161);
xor U979 (N_979,N_688,N_766);
nor U980 (N_980,N_109,N_498);
nor U981 (N_981,N_656,N_263);
and U982 (N_982,N_369,N_555);
xnor U983 (N_983,N_527,N_579);
and U984 (N_984,N_128,N_531);
or U985 (N_985,In_489,N_55);
nor U986 (N_986,In_409,In_1485);
and U987 (N_987,N_606,N_277);
nand U988 (N_988,N_683,N_168);
nor U989 (N_989,N_153,In_883);
or U990 (N_990,N_194,In_1338);
and U991 (N_991,In_1008,N_10);
and U992 (N_992,In_513,N_561);
and U993 (N_993,N_730,In_1565);
and U994 (N_994,N_526,In_1413);
xor U995 (N_995,In_190,In_1334);
nor U996 (N_996,N_666,N_228);
xnor U997 (N_997,In_550,N_587);
and U998 (N_998,N_448,N_591);
xnor U999 (N_999,N_617,In_1478);
nor U1000 (N_1000,In_849,In_1370);
nor U1001 (N_1001,In_736,N_57);
and U1002 (N_1002,N_557,N_505);
nor U1003 (N_1003,N_634,In_1285);
nand U1004 (N_1004,In_104,N_140);
xnor U1005 (N_1005,In_1771,In_893);
nand U1006 (N_1006,N_349,In_831);
nor U1007 (N_1007,N_35,N_776);
xor U1008 (N_1008,In_1421,N_49);
or U1009 (N_1009,In_48,N_715);
and U1010 (N_1010,In_468,N_735);
nand U1011 (N_1011,In_1342,In_15);
and U1012 (N_1012,In_329,N_489);
nand U1013 (N_1013,N_455,In_1532);
nand U1014 (N_1014,In_799,In_666);
nor U1015 (N_1015,In_884,N_779);
nand U1016 (N_1016,In_1055,In_607);
nor U1017 (N_1017,In_1015,N_211);
nand U1018 (N_1018,In_392,N_53);
xor U1019 (N_1019,In_314,N_593);
and U1020 (N_1020,In_1733,N_657);
xnor U1021 (N_1021,N_71,In_1963);
or U1022 (N_1022,In_1504,In_1103);
nand U1023 (N_1023,In_1100,N_577);
nand U1024 (N_1024,N_458,N_450);
or U1025 (N_1025,N_549,N_343);
xor U1026 (N_1026,In_1240,N_548);
xnor U1027 (N_1027,N_703,N_234);
and U1028 (N_1028,N_147,N_781);
nor U1029 (N_1029,N_103,N_206);
nor U1030 (N_1030,N_777,In_399);
or U1031 (N_1031,N_512,N_246);
nor U1032 (N_1032,N_378,N_440);
nand U1033 (N_1033,In_250,N_50);
nand U1034 (N_1034,N_276,N_151);
nand U1035 (N_1035,N_632,In_1275);
xor U1036 (N_1036,N_472,N_408);
nor U1037 (N_1037,N_145,N_323);
nand U1038 (N_1038,In_769,N_399);
xnor U1039 (N_1039,N_359,In_1466);
nand U1040 (N_1040,In_1520,N_608);
nand U1041 (N_1041,In_1910,N_25);
nor U1042 (N_1042,In_1214,N_255);
nor U1043 (N_1043,N_610,In_900);
nor U1044 (N_1044,N_639,N_187);
or U1045 (N_1045,N_335,N_619);
xnor U1046 (N_1046,N_699,In_1994);
nor U1047 (N_1047,In_1899,N_697);
or U1048 (N_1048,N_665,In_412);
or U1049 (N_1049,N_659,N_645);
nor U1050 (N_1050,N_603,N_640);
and U1051 (N_1051,N_60,In_1258);
and U1052 (N_1052,N_769,In_1729);
nand U1053 (N_1053,N_195,In_1133);
nand U1054 (N_1054,N_257,N_755);
nand U1055 (N_1055,N_574,N_185);
xnor U1056 (N_1056,N_164,N_30);
and U1057 (N_1057,N_372,N_345);
xnor U1058 (N_1058,N_719,In_865);
xnor U1059 (N_1059,In_608,In_766);
nor U1060 (N_1060,N_149,N_662);
or U1061 (N_1061,N_377,N_105);
and U1062 (N_1062,N_798,N_388);
and U1063 (N_1063,In_375,N_533);
or U1064 (N_1064,N_100,N_696);
nor U1065 (N_1065,N_773,In_527);
nand U1066 (N_1066,N_476,N_672);
nand U1067 (N_1067,N_784,In_1218);
nand U1068 (N_1068,N_721,In_570);
xor U1069 (N_1069,In_1118,N_536);
nor U1070 (N_1070,N_720,In_1844);
xnor U1071 (N_1071,In_1654,N_244);
xnor U1072 (N_1072,In_1383,In_887);
nand U1073 (N_1073,N_329,In_1223);
and U1074 (N_1074,In_1239,N_761);
nor U1075 (N_1075,N_475,N_442);
xnor U1076 (N_1076,N_89,N_690);
and U1077 (N_1077,N_514,In_926);
nand U1078 (N_1078,N_40,N_67);
xnor U1079 (N_1079,N_509,N_613);
or U1080 (N_1080,N_661,N_795);
nor U1081 (N_1081,In_320,N_93);
nor U1082 (N_1082,N_129,N_367);
nand U1083 (N_1083,N_2,In_1922);
nor U1084 (N_1084,In_966,In_1180);
or U1085 (N_1085,N_609,In_440);
xor U1086 (N_1086,N_418,In_1723);
nor U1087 (N_1087,In_861,N_247);
xnor U1088 (N_1088,N_379,In_1656);
nor U1089 (N_1089,In_1321,N_364);
or U1090 (N_1090,N_338,N_717);
xor U1091 (N_1091,In_1057,In_844);
xor U1092 (N_1092,In_1104,N_29);
nand U1093 (N_1093,In_1136,In_518);
nand U1094 (N_1094,N_542,N_404);
or U1095 (N_1095,N_767,In_1773);
nor U1096 (N_1096,N_13,In_1610);
nand U1097 (N_1097,N_347,N_464);
or U1098 (N_1098,N_529,In_63);
or U1099 (N_1099,In_1787,In_586);
and U1100 (N_1100,N_692,N_365);
or U1101 (N_1101,In_1236,In_753);
nand U1102 (N_1102,In_1974,In_1774);
and U1103 (N_1103,N_218,N_113);
and U1104 (N_1104,N_289,In_1818);
or U1105 (N_1105,N_315,N_582);
or U1106 (N_1106,In_1477,N_110);
or U1107 (N_1107,In_1455,In_662);
or U1108 (N_1108,N_54,N_237);
or U1109 (N_1109,In_1606,In_1281);
nand U1110 (N_1110,N_426,N_503);
and U1111 (N_1111,N_17,N_482);
nor U1112 (N_1112,N_328,N_42);
or U1113 (N_1113,N_354,In_715);
nor U1114 (N_1114,N_622,In_442);
or U1115 (N_1115,N_554,In_1632);
nand U1116 (N_1116,N_679,N_381);
or U1117 (N_1117,In_980,N_152);
nor U1118 (N_1118,N_69,In_802);
nor U1119 (N_1119,N_578,In_848);
or U1120 (N_1120,N_34,N_576);
or U1121 (N_1121,N_191,In_1807);
nor U1122 (N_1122,N_85,N_72);
nand U1123 (N_1123,N_569,In_457);
and U1124 (N_1124,N_771,N_420);
xnor U1125 (N_1125,N_204,N_646);
nand U1126 (N_1126,In_444,In_1356);
nor U1127 (N_1127,N_304,N_82);
and U1128 (N_1128,N_764,N_217);
xor U1129 (N_1129,N_122,N_250);
nand U1130 (N_1130,N_175,N_713);
and U1131 (N_1131,N_272,N_275);
nor U1132 (N_1132,In_572,N_522);
or U1133 (N_1133,In_257,N_91);
nor U1134 (N_1134,N_20,N_76);
or U1135 (N_1135,N_314,N_376);
nor U1136 (N_1136,N_271,In_1060);
or U1137 (N_1137,N_754,N_118);
nand U1138 (N_1138,N_562,In_146);
or U1139 (N_1139,In_1662,In_1966);
and U1140 (N_1140,N_358,N_485);
nand U1141 (N_1141,N_238,N_184);
and U1142 (N_1142,N_158,N_68);
or U1143 (N_1143,In_1400,In_1784);
xnor U1144 (N_1144,N_135,In_1229);
nor U1145 (N_1145,N_229,In_1909);
nand U1146 (N_1146,N_21,N_189);
and U1147 (N_1147,N_37,N_685);
xor U1148 (N_1148,N_629,N_133);
xor U1149 (N_1149,N_220,N_251);
nand U1150 (N_1150,In_1613,N_644);
or U1151 (N_1151,N_528,In_754);
and U1152 (N_1152,In_1799,In_1458);
nand U1153 (N_1153,N_298,N_18);
nand U1154 (N_1154,N_663,N_492);
xor U1155 (N_1155,N_262,N_62);
xor U1156 (N_1156,N_760,In_485);
and U1157 (N_1157,In_1548,In_1226);
nor U1158 (N_1158,N_558,N_23);
nand U1159 (N_1159,N_497,In_1506);
nor U1160 (N_1160,N_63,In_1349);
and U1161 (N_1161,N_6,N_451);
nor U1162 (N_1162,In_805,In_1795);
nor U1163 (N_1163,In_949,N_213);
nand U1164 (N_1164,N_747,N_704);
or U1165 (N_1165,N_675,N_757);
or U1166 (N_1166,N_746,In_1368);
nor U1167 (N_1167,In_1630,In_835);
nor U1168 (N_1168,N_202,N_405);
nand U1169 (N_1169,N_77,N_306);
nor U1170 (N_1170,N_631,N_327);
and U1171 (N_1171,N_642,In_545);
xnor U1172 (N_1172,N_429,N_456);
and U1173 (N_1173,N_254,N_355);
nand U1174 (N_1174,N_513,N_197);
nor U1175 (N_1175,N_778,In_1266);
and U1176 (N_1176,N_188,N_571);
xor U1177 (N_1177,N_589,In_30);
nor U1178 (N_1178,N_210,N_423);
and U1179 (N_1179,N_124,N_432);
nand U1180 (N_1180,N_687,In_407);
nor U1181 (N_1181,N_794,N_305);
nand U1182 (N_1182,In_481,N_142);
nand U1183 (N_1183,N_278,N_64);
and U1184 (N_1184,N_382,N_363);
or U1185 (N_1185,In_1672,N_793);
nor U1186 (N_1186,In_1968,N_39);
and U1187 (N_1187,In_1330,N_543);
nor U1188 (N_1188,N_48,N_16);
nand U1189 (N_1189,N_130,N_709);
nand U1190 (N_1190,In_137,N_518);
and U1191 (N_1191,N_441,In_1612);
and U1192 (N_1192,N_573,N_724);
nor U1193 (N_1193,N_519,N_525);
nor U1194 (N_1194,N_350,N_736);
and U1195 (N_1195,In_1858,N_534);
nand U1196 (N_1196,N_484,In_115);
nand U1197 (N_1197,N_473,N_461);
xor U1198 (N_1198,N_209,In_97);
xor U1199 (N_1199,In_1990,N_198);
nand U1200 (N_1200,N_24,In_1869);
nor U1201 (N_1201,N_770,N_718);
and U1202 (N_1202,In_181,N_443);
and U1203 (N_1203,In_1448,N_651);
nor U1204 (N_1204,N_435,In_974);
and U1205 (N_1205,N_500,In_167);
and U1206 (N_1206,In_335,In_1111);
or U1207 (N_1207,N_266,N_362);
xor U1208 (N_1208,N_9,N_138);
and U1209 (N_1209,N_785,N_428);
nor U1210 (N_1210,In_1713,N_648);
xor U1211 (N_1211,N_653,N_177);
xor U1212 (N_1212,N_179,In_1590);
nand U1213 (N_1213,N_176,In_333);
nand U1214 (N_1214,N_705,In_1043);
nand U1215 (N_1215,N_307,N_775);
or U1216 (N_1216,N_51,N_431);
nor U1217 (N_1217,In_703,N_159);
or U1218 (N_1218,N_600,N_737);
or U1219 (N_1219,N_279,N_491);
and U1220 (N_1220,In_1669,In_785);
xnor U1221 (N_1221,N_597,In_456);
nor U1222 (N_1222,N_58,In_1625);
nand U1223 (N_1223,In_273,N_331);
nor U1224 (N_1224,N_300,In_1693);
or U1225 (N_1225,N_324,N_465);
nor U1226 (N_1226,N_125,In_1998);
and U1227 (N_1227,N_296,In_874);
and U1228 (N_1228,N_336,In_839);
nor U1229 (N_1229,N_466,N_411);
and U1230 (N_1230,N_586,In_1931);
nor U1231 (N_1231,In_1228,N_385);
and U1232 (N_1232,N_563,N_361);
and U1233 (N_1233,N_236,N_96);
or U1234 (N_1234,N_459,N_604);
xnor U1235 (N_1235,N_245,N_200);
xor U1236 (N_1236,N_671,N_167);
and U1237 (N_1237,N_667,In_1785);
or U1238 (N_1238,N_673,In_1719);
and U1239 (N_1239,N_669,N_652);
xor U1240 (N_1240,In_242,In_1604);
xnor U1241 (N_1241,N_616,N_281);
nand U1242 (N_1242,In_1727,N_635);
and U1243 (N_1243,N_447,N_620);
nand U1244 (N_1244,In_1233,N_572);
or U1245 (N_1245,In_1951,N_546);
nand U1246 (N_1246,N_501,N_80);
xor U1247 (N_1247,N_711,In_1800);
or U1248 (N_1248,N_36,N_649);
or U1249 (N_1249,N_169,In_372);
or U1250 (N_1250,N_567,N_742);
nor U1251 (N_1251,N_605,In_707);
xor U1252 (N_1252,N_658,In_1744);
nor U1253 (N_1253,N_274,N_493);
nand U1254 (N_1254,N_693,N_417);
nor U1255 (N_1255,N_520,N_468);
nand U1256 (N_1256,N_309,In_855);
and U1257 (N_1257,In_1709,N_101);
or U1258 (N_1258,N_726,N_583);
nand U1259 (N_1259,In_1191,In_1070);
nand U1260 (N_1260,In_151,In_1007);
or U1261 (N_1261,N_524,N_165);
and U1262 (N_1262,In_1130,N_759);
nor U1263 (N_1263,N_134,In_630);
nor U1264 (N_1264,N_789,In_269);
and U1265 (N_1265,In_1636,N_732);
xnor U1266 (N_1266,N_425,N_788);
or U1267 (N_1267,N_391,N_537);
and U1268 (N_1268,N_424,N_241);
and U1269 (N_1269,N_127,N_415);
or U1270 (N_1270,N_157,In_710);
or U1271 (N_1271,N_762,N_192);
and U1272 (N_1272,N_414,In_0);
nand U1273 (N_1273,In_821,N_438);
nand U1274 (N_1274,In_1932,N_474);
nand U1275 (N_1275,N_598,In_281);
or U1276 (N_1276,In_496,In_1363);
or U1277 (N_1277,In_536,In_1024);
or U1278 (N_1278,In_951,N_333);
nor U1279 (N_1279,N_386,N_265);
nand U1280 (N_1280,N_670,N_566);
or U1281 (N_1281,In_1802,N_219);
and U1282 (N_1282,N_682,N_43);
nand U1283 (N_1283,N_366,In_694);
and U1284 (N_1284,In_541,In_1193);
or U1285 (N_1285,In_120,In_1022);
and U1286 (N_1286,N_539,N_94);
or U1287 (N_1287,N_146,N_171);
and U1288 (N_1288,N_751,N_515);
nor U1289 (N_1289,N_738,N_339);
nor U1290 (N_1290,In_498,In_1868);
and U1291 (N_1291,N_252,In_1074);
and U1292 (N_1292,In_103,In_149);
xnor U1293 (N_1293,In_497,N_288);
nand U1294 (N_1294,N_112,In_1453);
xnor U1295 (N_1295,N_290,N_470);
or U1296 (N_1296,N_741,N_256);
or U1297 (N_1297,In_882,N_199);
xnor U1298 (N_1298,In_959,In_977);
nand U1299 (N_1299,In_1728,In_397);
nand U1300 (N_1300,N_570,In_1268);
and U1301 (N_1301,N_396,In_830);
nor U1302 (N_1302,N_117,N_47);
and U1303 (N_1303,N_633,In_529);
nand U1304 (N_1304,N_782,N_756);
or U1305 (N_1305,In_353,N_748);
nor U1306 (N_1306,In_1699,In_380);
or U1307 (N_1307,In_356,N_310);
xor U1308 (N_1308,N_502,N_731);
xnor U1309 (N_1309,N_630,In_1412);
nand U1310 (N_1310,In_1772,N_706);
or U1311 (N_1311,In_417,N_97);
nand U1312 (N_1312,In_590,N_260);
or U1313 (N_1313,N_694,N_545);
and U1314 (N_1314,In_1160,N_496);
and U1315 (N_1315,N_743,In_1638);
xor U1316 (N_1316,In_1697,N_551);
nor U1317 (N_1317,N_294,In_1798);
nand U1318 (N_1318,N_400,In_1835);
and U1319 (N_1319,N_15,N_180);
or U1320 (N_1320,N_224,N_370);
or U1321 (N_1321,N_772,N_33);
xor U1322 (N_1322,N_725,N_342);
or U1323 (N_1323,N_506,N_70);
and U1324 (N_1324,In_304,In_1490);
nand U1325 (N_1325,In_1647,In_1718);
nand U1326 (N_1326,N_421,N_280);
nand U1327 (N_1327,N_454,N_322);
nand U1328 (N_1328,N_268,N_65);
and U1329 (N_1329,In_1840,N_681);
or U1330 (N_1330,In_1950,N_540);
nand U1331 (N_1331,In_595,N_380);
xnor U1332 (N_1332,In_1405,N_530);
or U1333 (N_1333,N_19,N_150);
or U1334 (N_1334,In_731,N_232);
nor U1335 (N_1335,In_100,N_402);
or U1336 (N_1336,N_689,N_1);
xnor U1337 (N_1337,N_585,N_190);
nor U1338 (N_1338,N_791,In_561);
xor U1339 (N_1339,N_104,N_636);
and U1340 (N_1340,N_511,N_346);
nor U1341 (N_1341,In_1512,In_9);
nor U1342 (N_1342,In_583,N_348);
nand U1343 (N_1343,N_3,In_1091);
and U1344 (N_1344,In_197,N_344);
and U1345 (N_1345,N_594,N_744);
nor U1346 (N_1346,N_790,N_469);
nor U1347 (N_1347,N_643,N_86);
xor U1348 (N_1348,N_486,N_499);
xnor U1349 (N_1349,N_449,N_495);
or U1350 (N_1350,N_155,N_374);
or U1351 (N_1351,N_797,In_1561);
and U1352 (N_1352,In_569,N_752);
or U1353 (N_1353,N_267,N_481);
nor U1354 (N_1354,In_1182,N_44);
or U1355 (N_1355,N_407,In_697);
nor U1356 (N_1356,N_416,N_5);
and U1357 (N_1357,In_1369,N_695);
nor U1358 (N_1358,N_516,N_467);
nor U1359 (N_1359,N_38,N_297);
nand U1360 (N_1360,N_7,In_1892);
nor U1361 (N_1361,N_141,N_710);
nand U1362 (N_1362,In_307,In_194);
xor U1363 (N_1363,N_565,N_478);
nand U1364 (N_1364,N_716,N_341);
nand U1365 (N_1365,In_585,N_119);
nand U1366 (N_1366,In_943,N_293);
or U1367 (N_1367,N_332,In_942);
xnor U1368 (N_1368,In_768,N_650);
or U1369 (N_1369,N_799,N_580);
nand U1370 (N_1370,In_1865,In_1);
and U1371 (N_1371,N_698,N_581);
nor U1372 (N_1372,In_1189,N_395);
and U1373 (N_1373,N_433,In_698);
nor U1374 (N_1374,N_389,N_8);
and U1375 (N_1375,N_52,N_568);
xnor U1376 (N_1376,N_0,N_84);
or U1377 (N_1377,N_780,N_618);
or U1378 (N_1378,N_614,N_532);
nand U1379 (N_1379,In_350,N_226);
and U1380 (N_1380,N_462,N_108);
and U1381 (N_1381,In_205,N_143);
xnor U1382 (N_1382,In_93,In_612);
nor U1383 (N_1383,N_427,N_393);
and U1384 (N_1384,N_368,In_484);
xor U1385 (N_1385,In_76,N_550);
xnor U1386 (N_1386,N_357,N_99);
nor U1387 (N_1387,In_41,N_136);
or U1388 (N_1388,N_383,In_1423);
or U1389 (N_1389,N_588,N_121);
nand U1390 (N_1390,N_12,N_387);
nand U1391 (N_1391,N_203,N_231);
xnor U1392 (N_1392,N_783,In_911);
and U1393 (N_1393,N_46,N_114);
nand U1394 (N_1394,N_560,In_1760);
and U1395 (N_1395,In_1089,N_727);
or U1396 (N_1396,N_170,N_410);
nand U1397 (N_1397,N_207,In_1098);
nor U1398 (N_1398,N_460,N_723);
or U1399 (N_1399,N_75,N_787);
xnor U1400 (N_1400,N_729,N_220);
nor U1401 (N_1401,N_9,In_1858);
nor U1402 (N_1402,In_427,In_1421);
and U1403 (N_1403,In_1015,In_444);
nor U1404 (N_1404,In_1813,N_253);
nor U1405 (N_1405,N_162,N_436);
nor U1406 (N_1406,N_692,In_830);
nand U1407 (N_1407,N_354,N_147);
nand U1408 (N_1408,N_568,In_52);
and U1409 (N_1409,N_314,N_76);
nor U1410 (N_1410,N_309,In_884);
nand U1411 (N_1411,N_717,N_642);
or U1412 (N_1412,N_222,N_271);
xor U1413 (N_1413,N_323,N_325);
nor U1414 (N_1414,N_74,N_128);
nand U1415 (N_1415,In_486,N_223);
and U1416 (N_1416,N_304,N_743);
nand U1417 (N_1417,N_464,N_411);
xnor U1418 (N_1418,N_399,In_569);
nor U1419 (N_1419,N_665,N_300);
and U1420 (N_1420,N_124,In_774);
or U1421 (N_1421,In_527,In_1868);
or U1422 (N_1422,N_585,N_20);
nand U1423 (N_1423,In_226,N_769);
xor U1424 (N_1424,N_362,In_1966);
and U1425 (N_1425,In_855,In_758);
nor U1426 (N_1426,N_500,In_914);
xnor U1427 (N_1427,N_655,N_167);
and U1428 (N_1428,N_126,In_1182);
and U1429 (N_1429,N_413,N_419);
xnor U1430 (N_1430,N_207,N_153);
or U1431 (N_1431,In_966,N_535);
xnor U1432 (N_1432,N_126,N_584);
xor U1433 (N_1433,N_47,In_1103);
or U1434 (N_1434,N_404,N_560);
or U1435 (N_1435,N_578,In_1400);
nor U1436 (N_1436,In_1719,N_219);
xnor U1437 (N_1437,N_114,In_1618);
or U1438 (N_1438,N_760,In_541);
xnor U1439 (N_1439,N_89,N_203);
or U1440 (N_1440,N_335,N_610);
or U1441 (N_1441,N_366,In_171);
or U1442 (N_1442,N_754,N_212);
xnor U1443 (N_1443,In_1022,N_622);
nor U1444 (N_1444,N_618,N_390);
or U1445 (N_1445,N_457,In_1922);
nand U1446 (N_1446,N_449,N_401);
xor U1447 (N_1447,N_725,N_520);
nand U1448 (N_1448,In_1910,N_389);
and U1449 (N_1449,N_494,In_1968);
nand U1450 (N_1450,N_374,In_1369);
nor U1451 (N_1451,N_88,N_377);
or U1452 (N_1452,N_546,In_1008);
xor U1453 (N_1453,In_1117,N_609);
xnor U1454 (N_1454,N_153,In_481);
nand U1455 (N_1455,N_208,N_702);
nor U1456 (N_1456,N_7,In_1813);
xor U1457 (N_1457,In_1728,In_1848);
xor U1458 (N_1458,N_621,In_1007);
xnor U1459 (N_1459,In_307,N_593);
xnor U1460 (N_1460,In_1405,N_500);
xnor U1461 (N_1461,In_1365,N_93);
xor U1462 (N_1462,N_362,In_1410);
and U1463 (N_1463,N_499,N_403);
and U1464 (N_1464,N_151,N_377);
and U1465 (N_1465,N_626,N_703);
or U1466 (N_1466,In_1104,N_706);
and U1467 (N_1467,N_605,N_445);
nor U1468 (N_1468,In_980,N_385);
xnor U1469 (N_1469,N_723,N_228);
xnor U1470 (N_1470,N_345,N_183);
xor U1471 (N_1471,N_107,N_504);
nand U1472 (N_1472,N_88,In_769);
nor U1473 (N_1473,N_703,N_430);
or U1474 (N_1474,N_391,N_532);
or U1475 (N_1475,N_723,N_261);
nand U1476 (N_1476,N_561,N_474);
xnor U1477 (N_1477,N_679,In_541);
or U1478 (N_1478,N_33,N_756);
and U1479 (N_1479,N_328,N_222);
and U1480 (N_1480,In_1578,N_217);
and U1481 (N_1481,N_729,N_400);
and U1482 (N_1482,N_667,N_665);
or U1483 (N_1483,N_557,N_377);
nor U1484 (N_1484,In_821,In_1093);
xor U1485 (N_1485,N_627,N_268);
nor U1486 (N_1486,N_729,N_641);
nor U1487 (N_1487,N_384,In_414);
nor U1488 (N_1488,In_1522,In_703);
xnor U1489 (N_1489,N_462,N_278);
or U1490 (N_1490,In_34,N_662);
xnor U1491 (N_1491,N_60,In_737);
and U1492 (N_1492,N_105,In_1070);
nor U1493 (N_1493,N_712,N_440);
or U1494 (N_1494,In_304,N_465);
and U1495 (N_1495,N_743,N_215);
and U1496 (N_1496,N_552,In_1289);
nand U1497 (N_1497,N_610,N_346);
or U1498 (N_1498,N_192,N_403);
xor U1499 (N_1499,N_417,N_763);
nor U1500 (N_1500,N_581,N_349);
or U1501 (N_1501,N_537,N_46);
and U1502 (N_1502,In_949,N_796);
nand U1503 (N_1503,N_777,In_9);
nor U1504 (N_1504,In_409,N_324);
and U1505 (N_1505,N_165,N_268);
or U1506 (N_1506,N_684,N_57);
and U1507 (N_1507,In_1858,N_628);
nand U1508 (N_1508,In_1905,N_225);
or U1509 (N_1509,N_308,N_283);
or U1510 (N_1510,N_409,In_417);
or U1511 (N_1511,N_233,N_769);
xnor U1512 (N_1512,N_358,In_1455);
nor U1513 (N_1513,N_334,N_64);
and U1514 (N_1514,N_181,N_703);
nand U1515 (N_1515,N_396,In_569);
nor U1516 (N_1516,N_90,In_839);
or U1517 (N_1517,In_1909,N_749);
nand U1518 (N_1518,N_75,N_729);
and U1519 (N_1519,In_666,N_50);
nor U1520 (N_1520,In_1160,In_149);
or U1521 (N_1521,In_1368,In_1024);
nand U1522 (N_1522,N_157,N_690);
nand U1523 (N_1523,N_224,N_554);
xnor U1524 (N_1524,N_792,In_498);
nor U1525 (N_1525,N_339,In_1950);
and U1526 (N_1526,N_776,N_564);
nor U1527 (N_1527,N_610,N_399);
nor U1528 (N_1528,N_412,In_304);
and U1529 (N_1529,N_8,N_476);
or U1530 (N_1530,N_445,In_1423);
nor U1531 (N_1531,N_657,N_32);
nand U1532 (N_1532,N_332,N_360);
nand U1533 (N_1533,N_668,In_1578);
nor U1534 (N_1534,N_713,N_567);
and U1535 (N_1535,N_575,N_42);
nor U1536 (N_1536,N_401,N_47);
xnor U1537 (N_1537,N_485,N_70);
nand U1538 (N_1538,N_623,N_339);
nor U1539 (N_1539,N_583,N_503);
nor U1540 (N_1540,N_735,N_475);
and U1541 (N_1541,N_561,N_420);
xnor U1542 (N_1542,N_241,N_432);
and U1543 (N_1543,N_326,In_959);
and U1544 (N_1544,N_349,N_601);
nand U1545 (N_1545,N_553,N_55);
or U1546 (N_1546,N_94,N_575);
or U1547 (N_1547,In_250,N_335);
nand U1548 (N_1548,In_1040,N_351);
and U1549 (N_1549,N_615,In_100);
or U1550 (N_1550,N_659,N_281);
or U1551 (N_1551,In_1784,N_620);
or U1552 (N_1552,N_309,N_244);
or U1553 (N_1553,N_156,N_57);
nor U1554 (N_1554,N_522,N_31);
and U1555 (N_1555,In_265,N_452);
or U1556 (N_1556,N_739,N_512);
nand U1557 (N_1557,N_553,In_1061);
or U1558 (N_1558,In_1772,N_437);
nor U1559 (N_1559,N_679,N_160);
and U1560 (N_1560,In_304,N_143);
xor U1561 (N_1561,In_1236,In_883);
and U1562 (N_1562,N_350,In_698);
or U1563 (N_1563,N_673,N_291);
xnor U1564 (N_1564,N_630,In_774);
or U1565 (N_1565,N_681,In_1100);
xor U1566 (N_1566,N_613,N_293);
or U1567 (N_1567,N_785,In_1423);
or U1568 (N_1568,N_214,N_1);
or U1569 (N_1569,N_151,N_336);
nor U1570 (N_1570,N_390,In_320);
and U1571 (N_1571,N_763,N_306);
nand U1572 (N_1572,In_167,N_98);
or U1573 (N_1573,In_329,In_1844);
and U1574 (N_1574,In_883,In_265);
and U1575 (N_1575,In_1060,N_282);
nor U1576 (N_1576,N_445,N_284);
nand U1577 (N_1577,N_132,In_444);
or U1578 (N_1578,In_822,N_313);
xor U1579 (N_1579,N_250,N_420);
or U1580 (N_1580,N_92,N_567);
nor U1581 (N_1581,N_394,N_627);
nor U1582 (N_1582,N_312,N_265);
nand U1583 (N_1583,N_680,In_1055);
nand U1584 (N_1584,N_698,In_1664);
nor U1585 (N_1585,In_410,N_396);
or U1586 (N_1586,N_573,N_134);
and U1587 (N_1587,In_1931,In_1799);
and U1588 (N_1588,N_150,In_1229);
or U1589 (N_1589,N_494,N_172);
nor U1590 (N_1590,N_796,In_1733);
nor U1591 (N_1591,N_172,N_124);
nor U1592 (N_1592,N_489,In_1799);
nor U1593 (N_1593,N_626,In_1774);
nand U1594 (N_1594,In_51,N_99);
xor U1595 (N_1595,In_595,N_166);
nand U1596 (N_1596,N_121,In_412);
or U1597 (N_1597,N_525,In_1899);
xor U1598 (N_1598,N_68,N_767);
and U1599 (N_1599,N_344,In_1800);
and U1600 (N_1600,N_949,N_902);
and U1601 (N_1601,N_1084,N_824);
xor U1602 (N_1602,N_1559,N_957);
xnor U1603 (N_1603,N_1260,N_948);
or U1604 (N_1604,N_1379,N_1355);
xor U1605 (N_1605,N_1539,N_998);
nor U1606 (N_1606,N_1057,N_995);
or U1607 (N_1607,N_1536,N_1107);
xor U1608 (N_1608,N_1284,N_1129);
nand U1609 (N_1609,N_1207,N_1576);
xor U1610 (N_1610,N_1186,N_1088);
and U1611 (N_1611,N_927,N_1486);
xor U1612 (N_1612,N_1155,N_1202);
nand U1613 (N_1613,N_1450,N_1393);
nor U1614 (N_1614,N_1430,N_940);
and U1615 (N_1615,N_973,N_1052);
nand U1616 (N_1616,N_1425,N_880);
and U1617 (N_1617,N_1037,N_1327);
or U1618 (N_1618,N_1347,N_946);
and U1619 (N_1619,N_1521,N_1172);
and U1620 (N_1620,N_853,N_1546);
xnor U1621 (N_1621,N_1015,N_1116);
and U1622 (N_1622,N_1376,N_1526);
nor U1623 (N_1623,N_823,N_1404);
xnor U1624 (N_1624,N_1312,N_1293);
and U1625 (N_1625,N_1375,N_1268);
or U1626 (N_1626,N_1512,N_1493);
xor U1627 (N_1627,N_1326,N_1089);
xnor U1628 (N_1628,N_1003,N_867);
nand U1629 (N_1629,N_1227,N_1416);
nand U1630 (N_1630,N_1205,N_1018);
nor U1631 (N_1631,N_1201,N_992);
xor U1632 (N_1632,N_1577,N_1456);
nand U1633 (N_1633,N_829,N_1535);
and U1634 (N_1634,N_1215,N_1511);
or U1635 (N_1635,N_1256,N_999);
xnor U1636 (N_1636,N_846,N_972);
and U1637 (N_1637,N_1438,N_873);
nand U1638 (N_1638,N_920,N_1157);
nor U1639 (N_1639,N_1406,N_1074);
or U1640 (N_1640,N_1304,N_1253);
or U1641 (N_1641,N_1023,N_1542);
nor U1642 (N_1642,N_907,N_1458);
or U1643 (N_1643,N_901,N_919);
nor U1644 (N_1644,N_1342,N_1285);
nand U1645 (N_1645,N_898,N_1498);
or U1646 (N_1646,N_1453,N_1179);
nor U1647 (N_1647,N_1586,N_1318);
and U1648 (N_1648,N_1032,N_974);
nor U1649 (N_1649,N_1206,N_1166);
nand U1650 (N_1650,N_1209,N_1006);
xor U1651 (N_1651,N_872,N_1001);
or U1652 (N_1652,N_1282,N_1027);
nor U1653 (N_1653,N_1581,N_1353);
xnor U1654 (N_1654,N_1358,N_1529);
nor U1655 (N_1655,N_1403,N_1047);
and U1656 (N_1656,N_1275,N_1570);
nor U1657 (N_1657,N_816,N_819);
xor U1658 (N_1658,N_1385,N_1017);
nor U1659 (N_1659,N_1504,N_1171);
and U1660 (N_1660,N_960,N_848);
nor U1661 (N_1661,N_1051,N_1295);
nor U1662 (N_1662,N_1587,N_1560);
nor U1663 (N_1663,N_850,N_1468);
and U1664 (N_1664,N_1123,N_887);
xor U1665 (N_1665,N_1121,N_1176);
nand U1666 (N_1666,N_1109,N_1432);
nand U1667 (N_1667,N_1154,N_1200);
xnor U1668 (N_1668,N_1263,N_1354);
nor U1669 (N_1669,N_1483,N_1218);
or U1670 (N_1670,N_1269,N_956);
xor U1671 (N_1671,N_1046,N_1502);
nand U1672 (N_1672,N_1296,N_1214);
nand U1673 (N_1673,N_1050,N_947);
and U1674 (N_1674,N_879,N_1035);
nor U1675 (N_1675,N_1055,N_1356);
nand U1676 (N_1676,N_881,N_1044);
xor U1677 (N_1677,N_945,N_1558);
xnor U1678 (N_1678,N_1122,N_942);
and U1679 (N_1679,N_978,N_833);
nand U1680 (N_1680,N_843,N_1224);
nor U1681 (N_1681,N_1593,N_1369);
nor U1682 (N_1682,N_1597,N_1141);
nor U1683 (N_1683,N_968,N_1307);
or U1684 (N_1684,N_1437,N_1064);
or U1685 (N_1685,N_1026,N_1213);
and U1686 (N_1686,N_821,N_923);
or U1687 (N_1687,N_842,N_921);
xnor U1688 (N_1688,N_1241,N_1520);
or U1689 (N_1689,N_812,N_1034);
or U1690 (N_1690,N_1422,N_1408);
nand U1691 (N_1691,N_1411,N_985);
xor U1692 (N_1692,N_1451,N_807);
or U1693 (N_1693,N_1565,N_1135);
xnor U1694 (N_1694,N_884,N_1501);
nor U1695 (N_1695,N_1232,N_1271);
nand U1696 (N_1696,N_882,N_925);
nand U1697 (N_1697,N_1567,N_1329);
nand U1698 (N_1698,N_1447,N_1277);
or U1699 (N_1699,N_871,N_1158);
and U1700 (N_1700,N_917,N_1211);
nor U1701 (N_1701,N_938,N_1522);
or U1702 (N_1702,N_1324,N_1040);
or U1703 (N_1703,N_966,N_1181);
nor U1704 (N_1704,N_1175,N_1196);
and U1705 (N_1705,N_1281,N_1194);
or U1706 (N_1706,N_987,N_1002);
or U1707 (N_1707,N_1485,N_864);
or U1708 (N_1708,N_1407,N_1273);
nand U1709 (N_1709,N_1428,N_1087);
nor U1710 (N_1710,N_1462,N_1114);
nand U1711 (N_1711,N_986,N_1221);
xnor U1712 (N_1712,N_1070,N_1575);
or U1713 (N_1713,N_1279,N_1195);
nor U1714 (N_1714,N_1431,N_1484);
and U1715 (N_1715,N_1106,N_813);
or U1716 (N_1716,N_1383,N_851);
and U1717 (N_1717,N_804,N_1477);
nand U1718 (N_1718,N_828,N_1076);
or U1719 (N_1719,N_1149,N_1569);
nor U1720 (N_1720,N_1170,N_1243);
nand U1721 (N_1721,N_994,N_814);
nor U1722 (N_1722,N_1152,N_1153);
nand U1723 (N_1723,N_1454,N_859);
and U1724 (N_1724,N_891,N_1573);
xnor U1725 (N_1725,N_1165,N_1523);
nand U1726 (N_1726,N_903,N_991);
xnor U1727 (N_1727,N_932,N_1506);
and U1728 (N_1728,N_890,N_941);
nor U1729 (N_1729,N_861,N_1473);
nand U1730 (N_1730,N_1497,N_1212);
xor U1731 (N_1731,N_854,N_841);
nand U1732 (N_1732,N_1125,N_1457);
and U1733 (N_1733,N_1097,N_1306);
nor U1734 (N_1734,N_976,N_1334);
or U1735 (N_1735,N_1313,N_1083);
and U1736 (N_1736,N_1478,N_1138);
nor U1737 (N_1737,N_1496,N_1156);
or U1738 (N_1738,N_1427,N_1148);
nand U1739 (N_1739,N_1240,N_837);
xnor U1740 (N_1740,N_822,N_1352);
and U1741 (N_1741,N_1530,N_983);
xor U1742 (N_1742,N_1549,N_1548);
nor U1743 (N_1743,N_1231,N_1596);
nand U1744 (N_1744,N_1139,N_1096);
nand U1745 (N_1745,N_1386,N_1305);
or U1746 (N_1746,N_1262,N_805);
and U1747 (N_1747,N_868,N_1012);
nand U1748 (N_1748,N_835,N_1441);
nand U1749 (N_1749,N_965,N_1345);
nor U1750 (N_1750,N_1599,N_1225);
and U1751 (N_1751,N_1359,N_1585);
nand U1752 (N_1752,N_1259,N_1161);
xor U1753 (N_1753,N_888,N_1553);
nor U1754 (N_1754,N_1086,N_809);
nand U1755 (N_1755,N_831,N_1019);
nor U1756 (N_1756,N_1563,N_870);
nor U1757 (N_1757,N_1366,N_915);
nand U1758 (N_1758,N_1024,N_1402);
nand U1759 (N_1759,N_869,N_1412);
or U1760 (N_1760,N_1311,N_1409);
nand U1761 (N_1761,N_1405,N_1444);
xnor U1762 (N_1762,N_1338,N_1474);
nand U1763 (N_1763,N_1067,N_1490);
nand U1764 (N_1764,N_806,N_1397);
nor U1765 (N_1765,N_862,N_844);
and U1766 (N_1766,N_1102,N_1487);
nand U1767 (N_1767,N_1020,N_953);
or U1768 (N_1768,N_1361,N_1391);
and U1769 (N_1769,N_1180,N_904);
nand U1770 (N_1770,N_1128,N_1399);
or U1771 (N_1771,N_1488,N_893);
or U1772 (N_1772,N_1025,N_906);
or U1773 (N_1773,N_1120,N_1396);
or U1774 (N_1774,N_984,N_857);
xnor U1775 (N_1775,N_989,N_1499);
and U1776 (N_1776,N_1317,N_1081);
or U1777 (N_1777,N_1278,N_1467);
or U1778 (N_1778,N_1042,N_1339);
nor U1779 (N_1779,N_1532,N_895);
nand U1780 (N_1780,N_1518,N_849);
and U1781 (N_1781,N_918,N_1235);
nand U1782 (N_1782,N_1413,N_1142);
nor U1783 (N_1783,N_1092,N_914);
nand U1784 (N_1784,N_1442,N_1028);
or U1785 (N_1785,N_1579,N_1566);
nand U1786 (N_1786,N_931,N_1079);
and U1787 (N_1787,N_1325,N_990);
nand U1788 (N_1788,N_1346,N_1300);
nand U1789 (N_1789,N_1330,N_979);
and U1790 (N_1790,N_1013,N_1443);
xor U1791 (N_1791,N_997,N_1054);
or U1792 (N_1792,N_961,N_1541);
xnor U1793 (N_1793,N_1140,N_889);
xnor U1794 (N_1794,N_900,N_1133);
and U1795 (N_1795,N_1545,N_969);
and U1796 (N_1796,N_1384,N_1117);
nor U1797 (N_1797,N_1189,N_1350);
nor U1798 (N_1798,N_1555,N_1315);
and U1799 (N_1799,N_1100,N_1528);
xnor U1800 (N_1800,N_1434,N_1564);
nor U1801 (N_1801,N_943,N_855);
nor U1802 (N_1802,N_1340,N_1582);
or U1803 (N_1803,N_1400,N_1460);
xor U1804 (N_1804,N_1137,N_1078);
nand U1805 (N_1805,N_1544,N_1261);
xor U1806 (N_1806,N_1198,N_1222);
and U1807 (N_1807,N_1316,N_937);
or U1808 (N_1808,N_1029,N_912);
and U1809 (N_1809,N_820,N_1455);
xnor U1810 (N_1810,N_1418,N_1127);
and U1811 (N_1811,N_1491,N_1435);
or U1812 (N_1812,N_1093,N_1159);
and U1813 (N_1813,N_886,N_1174);
nand U1814 (N_1814,N_1531,N_1517);
nand U1815 (N_1815,N_1303,N_993);
nor U1816 (N_1816,N_1415,N_1410);
xnor U1817 (N_1817,N_1217,N_1192);
and U1818 (N_1818,N_1124,N_1562);
nand U1819 (N_1819,N_1101,N_1115);
and U1820 (N_1820,N_1348,N_967);
or U1821 (N_1821,N_1131,N_1515);
xor U1822 (N_1822,N_1594,N_874);
and U1823 (N_1823,N_1004,N_1381);
nand U1824 (N_1824,N_939,N_1446);
xor U1825 (N_1825,N_1465,N_1203);
nor U1826 (N_1826,N_1264,N_858);
and U1827 (N_1827,N_908,N_811);
nor U1828 (N_1828,N_1367,N_1463);
nor U1829 (N_1829,N_1533,N_1561);
nor U1830 (N_1830,N_962,N_910);
or U1831 (N_1831,N_1314,N_1077);
xnor U1832 (N_1832,N_988,N_896);
xor U1833 (N_1833,N_832,N_1049);
nand U1834 (N_1834,N_909,N_1229);
xnor U1835 (N_1835,N_1426,N_803);
and U1836 (N_1836,N_1395,N_1053);
nand U1837 (N_1837,N_834,N_1072);
or U1838 (N_1838,N_1045,N_1111);
nand U1839 (N_1839,N_1238,N_1507);
nand U1840 (N_1840,N_950,N_1583);
nor U1841 (N_1841,N_1362,N_1119);
nand U1842 (N_1842,N_1349,N_1481);
nor U1843 (N_1843,N_1372,N_1233);
or U1844 (N_1844,N_1322,N_1147);
or U1845 (N_1845,N_1254,N_970);
or U1846 (N_1846,N_1219,N_863);
nor U1847 (N_1847,N_1065,N_1302);
or U1848 (N_1848,N_1389,N_1080);
xnor U1849 (N_1849,N_1288,N_1373);
or U1850 (N_1850,N_933,N_1056);
nand U1851 (N_1851,N_818,N_1557);
xnor U1852 (N_1852,N_1370,N_1363);
and U1853 (N_1853,N_801,N_1323);
and U1854 (N_1854,N_1445,N_1062);
and U1855 (N_1855,N_911,N_1503);
nand U1856 (N_1856,N_817,N_1103);
or U1857 (N_1857,N_1104,N_958);
nand U1858 (N_1858,N_1274,N_1160);
xnor U1859 (N_1859,N_955,N_1572);
and U1860 (N_1860,N_1151,N_1505);
nor U1861 (N_1861,N_1598,N_981);
and U1862 (N_1862,N_1509,N_930);
or U1863 (N_1863,N_1333,N_825);
nor U1864 (N_1864,N_1237,N_1150);
xor U1865 (N_1865,N_1041,N_1534);
nand U1866 (N_1866,N_1368,N_1132);
nor U1867 (N_1867,N_1439,N_1344);
or U1868 (N_1868,N_1245,N_1134);
nor U1869 (N_1869,N_1190,N_1479);
nand U1870 (N_1870,N_1164,N_905);
and U1871 (N_1871,N_936,N_1095);
or U1872 (N_1872,N_1270,N_1464);
nand U1873 (N_1873,N_1500,N_1038);
nor U1874 (N_1874,N_996,N_826);
xnor U1875 (N_1875,N_875,N_1014);
nor U1876 (N_1876,N_1357,N_977);
nand U1877 (N_1877,N_876,N_1091);
xor U1878 (N_1878,N_1291,N_1005);
or U1879 (N_1879,N_1230,N_1440);
and U1880 (N_1880,N_1414,N_1592);
nor U1881 (N_1881,N_845,N_1398);
nor U1882 (N_1882,N_1255,N_1173);
nand U1883 (N_1883,N_1328,N_808);
or U1884 (N_1884,N_1031,N_1554);
nor U1885 (N_1885,N_1226,N_971);
nand U1886 (N_1886,N_1290,N_1112);
and U1887 (N_1887,N_982,N_1387);
nand U1888 (N_1888,N_885,N_1061);
or U1889 (N_1889,N_1420,N_1547);
and U1890 (N_1890,N_1033,N_1223);
nand U1891 (N_1891,N_1336,N_1287);
nand U1892 (N_1892,N_1371,N_1489);
or U1893 (N_1893,N_1280,N_1514);
xor U1894 (N_1894,N_1251,N_1543);
nor U1895 (N_1895,N_1394,N_1130);
nand U1896 (N_1896,N_1178,N_1169);
nand U1897 (N_1897,N_1183,N_1424);
nor U1898 (N_1898,N_1286,N_847);
or U1899 (N_1899,N_1508,N_1429);
and U1900 (N_1900,N_954,N_840);
xnor U1901 (N_1901,N_935,N_1331);
xnor U1902 (N_1902,N_1250,N_865);
or U1903 (N_1903,N_1309,N_1292);
xor U1904 (N_1904,N_1162,N_1510);
nand U1905 (N_1905,N_1187,N_1294);
nor U1906 (N_1906,N_1094,N_1085);
nor U1907 (N_1907,N_1556,N_836);
xor U1908 (N_1908,N_1252,N_1419);
nor U1909 (N_1909,N_802,N_1191);
and U1910 (N_1910,N_1216,N_916);
and U1911 (N_1911,N_1043,N_1421);
nand U1912 (N_1912,N_1071,N_1364);
or U1913 (N_1913,N_894,N_1589);
or U1914 (N_1914,N_1184,N_1082);
nand U1915 (N_1915,N_1433,N_952);
nor U1916 (N_1916,N_1471,N_1126);
and U1917 (N_1917,N_1022,N_1476);
nor U1918 (N_1918,N_1118,N_852);
nor U1919 (N_1919,N_1208,N_1475);
xnor U1920 (N_1920,N_897,N_1000);
xnor U1921 (N_1921,N_1283,N_1069);
xor U1922 (N_1922,N_899,N_1301);
and U1923 (N_1923,N_1571,N_1234);
nand U1924 (N_1924,N_1568,N_1058);
xor U1925 (N_1925,N_1516,N_1423);
nand U1926 (N_1926,N_1167,N_963);
nor U1927 (N_1927,N_1320,N_1584);
nand U1928 (N_1928,N_1524,N_878);
or U1929 (N_1929,N_1066,N_1257);
xnor U1930 (N_1930,N_856,N_1099);
and U1931 (N_1931,N_1537,N_1452);
or U1932 (N_1932,N_1060,N_860);
xnor U1933 (N_1933,N_980,N_1382);
xnor U1934 (N_1934,N_924,N_1377);
xor U1935 (N_1935,N_883,N_1039);
nor U1936 (N_1936,N_1193,N_1449);
xnor U1937 (N_1937,N_1016,N_1244);
or U1938 (N_1938,N_1008,N_1063);
xor U1939 (N_1939,N_1247,N_1550);
or U1940 (N_1940,N_1459,N_1365);
nor U1941 (N_1941,N_1146,N_1110);
or U1942 (N_1942,N_1297,N_1401);
xnor U1943 (N_1943,N_951,N_929);
nand U1944 (N_1944,N_1258,N_1210);
or U1945 (N_1945,N_1144,N_1177);
or U1946 (N_1946,N_1436,N_1249);
and U1947 (N_1947,N_1030,N_1036);
xnor U1948 (N_1948,N_1242,N_1472);
and U1949 (N_1949,N_810,N_1591);
and U1950 (N_1950,N_1136,N_1266);
nand U1951 (N_1951,N_1590,N_1105);
nor U1952 (N_1952,N_1332,N_1228);
and U1953 (N_1953,N_1574,N_1540);
nor U1954 (N_1954,N_1098,N_1276);
xor U1955 (N_1955,N_1513,N_1319);
nand U1956 (N_1956,N_1145,N_1021);
nand U1957 (N_1957,N_1482,N_800);
nand U1958 (N_1958,N_1417,N_1289);
and U1959 (N_1959,N_1392,N_1048);
nor U1960 (N_1960,N_1199,N_1492);
or U1961 (N_1961,N_1321,N_928);
nor U1962 (N_1962,N_1298,N_892);
or U1963 (N_1963,N_975,N_1108);
and U1964 (N_1964,N_1494,N_830);
and U1965 (N_1965,N_839,N_1337);
nand U1966 (N_1966,N_1059,N_1090);
nor U1967 (N_1967,N_1525,N_1272);
xnor U1968 (N_1968,N_1299,N_934);
and U1969 (N_1969,N_1236,N_1220);
nand U1970 (N_1970,N_1374,N_922);
nand U1971 (N_1971,N_1075,N_1010);
or U1972 (N_1972,N_1009,N_1578);
nor U1973 (N_1973,N_1466,N_1239);
and U1974 (N_1974,N_1068,N_1448);
or U1975 (N_1975,N_1538,N_1341);
and U1976 (N_1976,N_926,N_913);
xnor U1977 (N_1977,N_1007,N_1552);
or U1978 (N_1978,N_1461,N_1480);
nor U1979 (N_1979,N_1113,N_1360);
nor U1980 (N_1980,N_1495,N_866);
nand U1981 (N_1981,N_1390,N_838);
and U1982 (N_1982,N_1378,N_1185);
nor U1983 (N_1983,N_964,N_1343);
xor U1984 (N_1984,N_1246,N_1073);
and U1985 (N_1985,N_1163,N_1143);
or U1986 (N_1986,N_959,N_1380);
or U1987 (N_1987,N_1470,N_1188);
or U1988 (N_1988,N_944,N_827);
and U1989 (N_1989,N_1580,N_1588);
nand U1990 (N_1990,N_1248,N_1265);
nor U1991 (N_1991,N_1267,N_1204);
or U1992 (N_1992,N_815,N_1595);
or U1993 (N_1993,N_1469,N_1351);
nand U1994 (N_1994,N_1388,N_1197);
xor U1995 (N_1995,N_877,N_1335);
or U1996 (N_1996,N_1308,N_1310);
or U1997 (N_1997,N_1011,N_1519);
xnor U1998 (N_1998,N_1182,N_1168);
and U1999 (N_1999,N_1551,N_1527);
or U2000 (N_2000,N_1541,N_936);
or U2001 (N_2001,N_878,N_1327);
xnor U2002 (N_2002,N_840,N_1513);
or U2003 (N_2003,N_947,N_951);
nor U2004 (N_2004,N_974,N_1173);
nand U2005 (N_2005,N_1019,N_847);
or U2006 (N_2006,N_1319,N_1152);
nand U2007 (N_2007,N_1507,N_1376);
nor U2008 (N_2008,N_1470,N_1099);
xnor U2009 (N_2009,N_1040,N_961);
or U2010 (N_2010,N_890,N_1031);
or U2011 (N_2011,N_1027,N_816);
nor U2012 (N_2012,N_1457,N_1242);
or U2013 (N_2013,N_1519,N_1395);
or U2014 (N_2014,N_1522,N_1506);
or U2015 (N_2015,N_1429,N_946);
nor U2016 (N_2016,N_1270,N_1407);
or U2017 (N_2017,N_1066,N_1268);
or U2018 (N_2018,N_1042,N_1537);
nor U2019 (N_2019,N_1397,N_982);
xnor U2020 (N_2020,N_1453,N_1421);
and U2021 (N_2021,N_1379,N_1201);
or U2022 (N_2022,N_1442,N_1119);
nand U2023 (N_2023,N_927,N_958);
nor U2024 (N_2024,N_1263,N_1377);
xor U2025 (N_2025,N_954,N_1238);
and U2026 (N_2026,N_866,N_1529);
and U2027 (N_2027,N_892,N_1315);
xnor U2028 (N_2028,N_1076,N_1261);
xnor U2029 (N_2029,N_1470,N_1324);
nand U2030 (N_2030,N_971,N_823);
and U2031 (N_2031,N_1322,N_1251);
or U2032 (N_2032,N_1123,N_829);
or U2033 (N_2033,N_856,N_927);
or U2034 (N_2034,N_1570,N_1125);
xor U2035 (N_2035,N_1219,N_1291);
nand U2036 (N_2036,N_1227,N_1071);
nor U2037 (N_2037,N_1030,N_802);
nor U2038 (N_2038,N_1137,N_1169);
nand U2039 (N_2039,N_1335,N_1215);
nor U2040 (N_2040,N_1584,N_1059);
nor U2041 (N_2041,N_1470,N_1466);
xor U2042 (N_2042,N_1179,N_912);
nor U2043 (N_2043,N_1284,N_1061);
or U2044 (N_2044,N_1209,N_1023);
nor U2045 (N_2045,N_959,N_935);
nor U2046 (N_2046,N_1472,N_1351);
nand U2047 (N_2047,N_1076,N_1457);
nor U2048 (N_2048,N_1280,N_1259);
nor U2049 (N_2049,N_1223,N_932);
xor U2050 (N_2050,N_1583,N_1313);
xor U2051 (N_2051,N_963,N_1324);
nor U2052 (N_2052,N_1369,N_966);
nand U2053 (N_2053,N_986,N_1207);
xnor U2054 (N_2054,N_851,N_1403);
nand U2055 (N_2055,N_1093,N_953);
xnor U2056 (N_2056,N_1300,N_1070);
and U2057 (N_2057,N_1374,N_993);
and U2058 (N_2058,N_1499,N_1497);
and U2059 (N_2059,N_1121,N_1579);
nor U2060 (N_2060,N_1127,N_833);
xor U2061 (N_2061,N_1114,N_1579);
nand U2062 (N_2062,N_1323,N_1569);
xor U2063 (N_2063,N_1216,N_804);
nand U2064 (N_2064,N_1557,N_970);
nand U2065 (N_2065,N_1171,N_1501);
and U2066 (N_2066,N_1171,N_837);
nand U2067 (N_2067,N_1564,N_1337);
nor U2068 (N_2068,N_1493,N_1243);
and U2069 (N_2069,N_971,N_1183);
xor U2070 (N_2070,N_1249,N_1561);
nor U2071 (N_2071,N_1553,N_1599);
or U2072 (N_2072,N_816,N_1490);
nor U2073 (N_2073,N_1502,N_1497);
and U2074 (N_2074,N_1453,N_1042);
or U2075 (N_2075,N_879,N_1229);
and U2076 (N_2076,N_1592,N_1541);
or U2077 (N_2077,N_1368,N_1355);
nand U2078 (N_2078,N_1350,N_1126);
and U2079 (N_2079,N_1227,N_1175);
or U2080 (N_2080,N_1324,N_1321);
nor U2081 (N_2081,N_1239,N_1556);
and U2082 (N_2082,N_979,N_1280);
nor U2083 (N_2083,N_1045,N_1464);
nor U2084 (N_2084,N_1235,N_820);
or U2085 (N_2085,N_1384,N_1330);
xnor U2086 (N_2086,N_909,N_1490);
and U2087 (N_2087,N_1450,N_1272);
nor U2088 (N_2088,N_1118,N_992);
nor U2089 (N_2089,N_1318,N_1131);
nor U2090 (N_2090,N_1313,N_1130);
xor U2091 (N_2091,N_800,N_1203);
or U2092 (N_2092,N_1018,N_1480);
nand U2093 (N_2093,N_1362,N_1402);
or U2094 (N_2094,N_817,N_1360);
and U2095 (N_2095,N_1424,N_1279);
or U2096 (N_2096,N_922,N_954);
xnor U2097 (N_2097,N_1309,N_947);
and U2098 (N_2098,N_1531,N_1125);
or U2099 (N_2099,N_1303,N_906);
and U2100 (N_2100,N_1404,N_942);
xnor U2101 (N_2101,N_1541,N_1058);
or U2102 (N_2102,N_1505,N_1570);
xnor U2103 (N_2103,N_1451,N_1178);
nand U2104 (N_2104,N_1322,N_828);
nor U2105 (N_2105,N_803,N_1402);
nor U2106 (N_2106,N_1131,N_1277);
nor U2107 (N_2107,N_1283,N_1128);
nand U2108 (N_2108,N_1062,N_1542);
or U2109 (N_2109,N_1181,N_1301);
nor U2110 (N_2110,N_927,N_1027);
or U2111 (N_2111,N_994,N_1112);
xnor U2112 (N_2112,N_971,N_1418);
or U2113 (N_2113,N_1515,N_1083);
and U2114 (N_2114,N_1178,N_1429);
nor U2115 (N_2115,N_912,N_1041);
nand U2116 (N_2116,N_1592,N_1478);
or U2117 (N_2117,N_1539,N_1391);
and U2118 (N_2118,N_1325,N_1184);
nor U2119 (N_2119,N_1482,N_1518);
xnor U2120 (N_2120,N_1426,N_1087);
xor U2121 (N_2121,N_869,N_800);
xor U2122 (N_2122,N_1003,N_1453);
or U2123 (N_2123,N_1161,N_1499);
nand U2124 (N_2124,N_1132,N_1169);
nand U2125 (N_2125,N_1056,N_1390);
nand U2126 (N_2126,N_960,N_1272);
or U2127 (N_2127,N_990,N_1183);
nor U2128 (N_2128,N_1522,N_1370);
nand U2129 (N_2129,N_1237,N_1236);
or U2130 (N_2130,N_841,N_1588);
nor U2131 (N_2131,N_1218,N_1461);
nand U2132 (N_2132,N_1060,N_1423);
nor U2133 (N_2133,N_987,N_1384);
or U2134 (N_2134,N_1038,N_1000);
or U2135 (N_2135,N_810,N_1142);
xor U2136 (N_2136,N_969,N_1005);
and U2137 (N_2137,N_826,N_1564);
nand U2138 (N_2138,N_1428,N_1538);
nor U2139 (N_2139,N_972,N_891);
nand U2140 (N_2140,N_1141,N_1058);
nor U2141 (N_2141,N_945,N_1494);
or U2142 (N_2142,N_1132,N_830);
nand U2143 (N_2143,N_1107,N_1492);
nand U2144 (N_2144,N_1067,N_1494);
nand U2145 (N_2145,N_974,N_1244);
nor U2146 (N_2146,N_1148,N_1268);
xnor U2147 (N_2147,N_882,N_875);
nor U2148 (N_2148,N_835,N_1262);
nor U2149 (N_2149,N_1326,N_1108);
or U2150 (N_2150,N_897,N_1099);
nor U2151 (N_2151,N_1044,N_1576);
nor U2152 (N_2152,N_1416,N_1509);
or U2153 (N_2153,N_901,N_1485);
xnor U2154 (N_2154,N_844,N_1167);
xor U2155 (N_2155,N_970,N_1386);
and U2156 (N_2156,N_1274,N_937);
nor U2157 (N_2157,N_1238,N_1491);
nor U2158 (N_2158,N_939,N_1514);
nand U2159 (N_2159,N_897,N_918);
or U2160 (N_2160,N_1191,N_1044);
or U2161 (N_2161,N_1319,N_966);
and U2162 (N_2162,N_1433,N_1090);
and U2163 (N_2163,N_1026,N_1135);
or U2164 (N_2164,N_1095,N_1436);
nor U2165 (N_2165,N_1070,N_824);
or U2166 (N_2166,N_1537,N_1523);
and U2167 (N_2167,N_1460,N_994);
or U2168 (N_2168,N_1100,N_1127);
or U2169 (N_2169,N_809,N_1437);
or U2170 (N_2170,N_882,N_1037);
or U2171 (N_2171,N_1003,N_1169);
nor U2172 (N_2172,N_1051,N_1222);
xnor U2173 (N_2173,N_847,N_1402);
nand U2174 (N_2174,N_990,N_1368);
nor U2175 (N_2175,N_888,N_823);
or U2176 (N_2176,N_883,N_1078);
xnor U2177 (N_2177,N_1304,N_971);
and U2178 (N_2178,N_1135,N_1149);
nor U2179 (N_2179,N_932,N_862);
nor U2180 (N_2180,N_948,N_1178);
or U2181 (N_2181,N_1277,N_958);
nand U2182 (N_2182,N_1194,N_1594);
and U2183 (N_2183,N_1533,N_1150);
nand U2184 (N_2184,N_1548,N_1541);
xnor U2185 (N_2185,N_1458,N_1137);
nand U2186 (N_2186,N_1334,N_1594);
xnor U2187 (N_2187,N_826,N_987);
or U2188 (N_2188,N_1164,N_1305);
xnor U2189 (N_2189,N_1364,N_1543);
or U2190 (N_2190,N_1446,N_1242);
and U2191 (N_2191,N_1553,N_1062);
nor U2192 (N_2192,N_962,N_1458);
and U2193 (N_2193,N_1190,N_813);
nand U2194 (N_2194,N_918,N_1214);
xor U2195 (N_2195,N_1577,N_1042);
nand U2196 (N_2196,N_1386,N_1546);
and U2197 (N_2197,N_1367,N_1450);
nor U2198 (N_2198,N_1267,N_1298);
or U2199 (N_2199,N_1347,N_1398);
xnor U2200 (N_2200,N_1448,N_1454);
nor U2201 (N_2201,N_1463,N_1339);
or U2202 (N_2202,N_1542,N_1577);
xnor U2203 (N_2203,N_954,N_1032);
and U2204 (N_2204,N_1253,N_810);
or U2205 (N_2205,N_1537,N_1274);
and U2206 (N_2206,N_1401,N_816);
nor U2207 (N_2207,N_1056,N_1463);
nand U2208 (N_2208,N_1150,N_1014);
nand U2209 (N_2209,N_1059,N_1002);
nand U2210 (N_2210,N_1115,N_1124);
or U2211 (N_2211,N_1508,N_1287);
and U2212 (N_2212,N_1200,N_1475);
xor U2213 (N_2213,N_1163,N_1289);
xor U2214 (N_2214,N_1097,N_1167);
xnor U2215 (N_2215,N_1413,N_920);
xnor U2216 (N_2216,N_1413,N_1073);
nor U2217 (N_2217,N_1303,N_1359);
xnor U2218 (N_2218,N_1224,N_1463);
nor U2219 (N_2219,N_1002,N_870);
xnor U2220 (N_2220,N_905,N_857);
or U2221 (N_2221,N_1055,N_1022);
nor U2222 (N_2222,N_935,N_873);
xor U2223 (N_2223,N_1311,N_1186);
nand U2224 (N_2224,N_1446,N_947);
nor U2225 (N_2225,N_1335,N_1350);
nor U2226 (N_2226,N_1267,N_847);
nand U2227 (N_2227,N_972,N_1589);
xnor U2228 (N_2228,N_808,N_1509);
xnor U2229 (N_2229,N_1075,N_1132);
and U2230 (N_2230,N_1246,N_1342);
and U2231 (N_2231,N_1349,N_1163);
or U2232 (N_2232,N_930,N_1036);
xnor U2233 (N_2233,N_1065,N_969);
nand U2234 (N_2234,N_1423,N_1041);
nor U2235 (N_2235,N_1134,N_1044);
nor U2236 (N_2236,N_1316,N_1282);
nand U2237 (N_2237,N_1358,N_857);
or U2238 (N_2238,N_894,N_1308);
nor U2239 (N_2239,N_1588,N_1160);
nand U2240 (N_2240,N_1434,N_1513);
xor U2241 (N_2241,N_1163,N_1133);
or U2242 (N_2242,N_1574,N_1143);
and U2243 (N_2243,N_1414,N_1127);
and U2244 (N_2244,N_828,N_1342);
nand U2245 (N_2245,N_1066,N_1267);
nor U2246 (N_2246,N_1056,N_956);
or U2247 (N_2247,N_1046,N_850);
xnor U2248 (N_2248,N_1194,N_1329);
or U2249 (N_2249,N_1299,N_1365);
nand U2250 (N_2250,N_1346,N_940);
xnor U2251 (N_2251,N_1111,N_1170);
nor U2252 (N_2252,N_1586,N_1478);
nand U2253 (N_2253,N_1117,N_1452);
xnor U2254 (N_2254,N_956,N_1396);
nor U2255 (N_2255,N_995,N_1544);
and U2256 (N_2256,N_1350,N_1256);
xor U2257 (N_2257,N_1174,N_1393);
and U2258 (N_2258,N_907,N_1010);
or U2259 (N_2259,N_1387,N_1493);
xnor U2260 (N_2260,N_1241,N_1481);
xnor U2261 (N_2261,N_1174,N_1024);
nor U2262 (N_2262,N_1487,N_1503);
nand U2263 (N_2263,N_1457,N_1351);
and U2264 (N_2264,N_1286,N_1440);
nand U2265 (N_2265,N_1118,N_1474);
nor U2266 (N_2266,N_937,N_1586);
xor U2267 (N_2267,N_1468,N_1075);
nor U2268 (N_2268,N_811,N_1220);
nand U2269 (N_2269,N_1094,N_1584);
or U2270 (N_2270,N_1529,N_1159);
nand U2271 (N_2271,N_843,N_1277);
and U2272 (N_2272,N_1372,N_1135);
xor U2273 (N_2273,N_854,N_869);
nor U2274 (N_2274,N_1569,N_1004);
or U2275 (N_2275,N_855,N_828);
xor U2276 (N_2276,N_1341,N_1417);
or U2277 (N_2277,N_903,N_942);
and U2278 (N_2278,N_1349,N_1170);
or U2279 (N_2279,N_1584,N_996);
nor U2280 (N_2280,N_857,N_1178);
and U2281 (N_2281,N_1280,N_1534);
and U2282 (N_2282,N_1165,N_1277);
nand U2283 (N_2283,N_1187,N_1052);
and U2284 (N_2284,N_918,N_1520);
nand U2285 (N_2285,N_1566,N_978);
nor U2286 (N_2286,N_1249,N_1262);
nand U2287 (N_2287,N_1403,N_1226);
nor U2288 (N_2288,N_1229,N_817);
xor U2289 (N_2289,N_801,N_925);
xnor U2290 (N_2290,N_1353,N_1543);
or U2291 (N_2291,N_1110,N_1016);
xor U2292 (N_2292,N_919,N_1147);
nand U2293 (N_2293,N_1582,N_1163);
nand U2294 (N_2294,N_1425,N_1068);
nand U2295 (N_2295,N_1594,N_1460);
nand U2296 (N_2296,N_1559,N_1339);
xor U2297 (N_2297,N_1097,N_1195);
nor U2298 (N_2298,N_1229,N_1498);
nand U2299 (N_2299,N_1320,N_1053);
xnor U2300 (N_2300,N_909,N_1205);
or U2301 (N_2301,N_912,N_1150);
and U2302 (N_2302,N_1568,N_879);
nor U2303 (N_2303,N_1334,N_1069);
or U2304 (N_2304,N_1003,N_1112);
nor U2305 (N_2305,N_1210,N_1063);
nor U2306 (N_2306,N_999,N_1425);
and U2307 (N_2307,N_849,N_1186);
xor U2308 (N_2308,N_1115,N_1129);
and U2309 (N_2309,N_834,N_1436);
nor U2310 (N_2310,N_1468,N_875);
xnor U2311 (N_2311,N_1098,N_1278);
nand U2312 (N_2312,N_837,N_1202);
or U2313 (N_2313,N_1323,N_1470);
and U2314 (N_2314,N_1340,N_1305);
and U2315 (N_2315,N_1267,N_896);
or U2316 (N_2316,N_864,N_848);
xor U2317 (N_2317,N_895,N_1574);
nand U2318 (N_2318,N_1417,N_1174);
nor U2319 (N_2319,N_1040,N_1155);
nand U2320 (N_2320,N_1490,N_1357);
nor U2321 (N_2321,N_1186,N_1508);
or U2322 (N_2322,N_1360,N_1392);
xnor U2323 (N_2323,N_1433,N_1190);
or U2324 (N_2324,N_1506,N_1435);
and U2325 (N_2325,N_1163,N_1589);
xor U2326 (N_2326,N_1396,N_1013);
and U2327 (N_2327,N_1197,N_1306);
nor U2328 (N_2328,N_1452,N_965);
nor U2329 (N_2329,N_889,N_1022);
nor U2330 (N_2330,N_1424,N_1443);
xnor U2331 (N_2331,N_915,N_1190);
or U2332 (N_2332,N_1175,N_1176);
and U2333 (N_2333,N_958,N_1159);
xor U2334 (N_2334,N_985,N_851);
xnor U2335 (N_2335,N_1160,N_1319);
or U2336 (N_2336,N_1473,N_1027);
and U2337 (N_2337,N_1171,N_1099);
or U2338 (N_2338,N_1195,N_1189);
and U2339 (N_2339,N_1080,N_930);
xor U2340 (N_2340,N_1064,N_1543);
nor U2341 (N_2341,N_1171,N_1372);
xor U2342 (N_2342,N_1455,N_1165);
and U2343 (N_2343,N_1205,N_932);
and U2344 (N_2344,N_862,N_1528);
xor U2345 (N_2345,N_1398,N_1028);
or U2346 (N_2346,N_964,N_1571);
nor U2347 (N_2347,N_1038,N_852);
nand U2348 (N_2348,N_1095,N_1519);
xnor U2349 (N_2349,N_1537,N_1058);
xor U2350 (N_2350,N_1119,N_1256);
or U2351 (N_2351,N_1211,N_1260);
and U2352 (N_2352,N_1388,N_913);
nand U2353 (N_2353,N_1475,N_865);
nor U2354 (N_2354,N_1395,N_898);
or U2355 (N_2355,N_836,N_895);
nand U2356 (N_2356,N_1053,N_920);
and U2357 (N_2357,N_1181,N_1149);
nand U2358 (N_2358,N_1477,N_1261);
xnor U2359 (N_2359,N_1243,N_1226);
nor U2360 (N_2360,N_998,N_1520);
nand U2361 (N_2361,N_973,N_1421);
xnor U2362 (N_2362,N_872,N_1158);
or U2363 (N_2363,N_1495,N_1060);
and U2364 (N_2364,N_1277,N_1377);
and U2365 (N_2365,N_1071,N_983);
nor U2366 (N_2366,N_1406,N_1068);
and U2367 (N_2367,N_1587,N_1552);
xnor U2368 (N_2368,N_1510,N_987);
nor U2369 (N_2369,N_1431,N_1103);
or U2370 (N_2370,N_1238,N_962);
xor U2371 (N_2371,N_1271,N_1473);
nand U2372 (N_2372,N_1529,N_1103);
nand U2373 (N_2373,N_1567,N_1134);
nor U2374 (N_2374,N_1423,N_1369);
and U2375 (N_2375,N_1583,N_1184);
nand U2376 (N_2376,N_1122,N_1581);
and U2377 (N_2377,N_1512,N_1032);
nor U2378 (N_2378,N_876,N_1223);
or U2379 (N_2379,N_1278,N_1436);
or U2380 (N_2380,N_1018,N_1526);
nand U2381 (N_2381,N_1253,N_1543);
xor U2382 (N_2382,N_1006,N_1000);
or U2383 (N_2383,N_1254,N_1498);
or U2384 (N_2384,N_1198,N_961);
nor U2385 (N_2385,N_1403,N_953);
or U2386 (N_2386,N_857,N_1141);
xor U2387 (N_2387,N_1162,N_1483);
xnor U2388 (N_2388,N_1254,N_1591);
nand U2389 (N_2389,N_1399,N_910);
nand U2390 (N_2390,N_1451,N_1557);
nor U2391 (N_2391,N_1052,N_834);
nand U2392 (N_2392,N_951,N_1212);
or U2393 (N_2393,N_834,N_1196);
or U2394 (N_2394,N_1030,N_1119);
xor U2395 (N_2395,N_1164,N_972);
xor U2396 (N_2396,N_1548,N_1432);
nor U2397 (N_2397,N_1347,N_1192);
or U2398 (N_2398,N_950,N_1520);
or U2399 (N_2399,N_1158,N_1349);
and U2400 (N_2400,N_2003,N_2163);
nand U2401 (N_2401,N_2209,N_1946);
xnor U2402 (N_2402,N_1935,N_2284);
nor U2403 (N_2403,N_2008,N_2353);
nand U2404 (N_2404,N_2026,N_2208);
nor U2405 (N_2405,N_1980,N_2350);
nor U2406 (N_2406,N_2255,N_2357);
or U2407 (N_2407,N_2153,N_2313);
nand U2408 (N_2408,N_1763,N_1627);
or U2409 (N_2409,N_2343,N_2286);
xnor U2410 (N_2410,N_1971,N_1717);
nor U2411 (N_2411,N_1728,N_1642);
or U2412 (N_2412,N_1911,N_2365);
or U2413 (N_2413,N_2278,N_2063);
or U2414 (N_2414,N_1932,N_2193);
xnor U2415 (N_2415,N_2356,N_1606);
or U2416 (N_2416,N_2273,N_2188);
nor U2417 (N_2417,N_2174,N_1989);
xor U2418 (N_2418,N_2261,N_2075);
and U2419 (N_2419,N_2245,N_1873);
nand U2420 (N_2420,N_1698,N_1725);
nand U2421 (N_2421,N_1770,N_2029);
nor U2422 (N_2422,N_2253,N_2056);
and U2423 (N_2423,N_1856,N_1679);
and U2424 (N_2424,N_1715,N_2220);
and U2425 (N_2425,N_1791,N_2123);
and U2426 (N_2426,N_1726,N_2215);
and U2427 (N_2427,N_2359,N_1978);
or U2428 (N_2428,N_1951,N_1991);
nor U2429 (N_2429,N_1927,N_1787);
nor U2430 (N_2430,N_1822,N_1943);
and U2431 (N_2431,N_1781,N_2006);
nand U2432 (N_2432,N_1904,N_1879);
nor U2433 (N_2433,N_2371,N_1967);
xor U2434 (N_2434,N_2324,N_2305);
xor U2435 (N_2435,N_1891,N_1814);
nand U2436 (N_2436,N_2079,N_1795);
nor U2437 (N_2437,N_2165,N_1802);
nor U2438 (N_2438,N_2272,N_2391);
and U2439 (N_2439,N_1643,N_1645);
or U2440 (N_2440,N_2111,N_2173);
xor U2441 (N_2441,N_1656,N_2190);
nor U2442 (N_2442,N_1972,N_1664);
nand U2443 (N_2443,N_2268,N_1719);
nand U2444 (N_2444,N_1687,N_1695);
nor U2445 (N_2445,N_1753,N_1670);
and U2446 (N_2446,N_1716,N_1961);
nor U2447 (N_2447,N_1844,N_1624);
nor U2448 (N_2448,N_2149,N_1860);
nor U2449 (N_2449,N_2086,N_2069);
nand U2450 (N_2450,N_2399,N_2218);
and U2451 (N_2451,N_2226,N_2099);
nor U2452 (N_2452,N_1906,N_2078);
nor U2453 (N_2453,N_1668,N_2258);
or U2454 (N_2454,N_1865,N_1612);
xnor U2455 (N_2455,N_1644,N_2129);
nor U2456 (N_2456,N_1834,N_1926);
or U2457 (N_2457,N_2125,N_1776);
and U2458 (N_2458,N_2093,N_1647);
and U2459 (N_2459,N_1654,N_1760);
nor U2460 (N_2460,N_1823,N_2348);
or U2461 (N_2461,N_1956,N_1613);
or U2462 (N_2462,N_2339,N_2177);
or U2463 (N_2463,N_1966,N_2335);
nand U2464 (N_2464,N_2297,N_2044);
or U2465 (N_2465,N_2317,N_1863);
xor U2466 (N_2466,N_1677,N_2352);
nand U2467 (N_2467,N_2217,N_2010);
or U2468 (N_2468,N_2050,N_1918);
xor U2469 (N_2469,N_2132,N_1713);
nand U2470 (N_2470,N_1744,N_2027);
nand U2471 (N_2471,N_1621,N_1730);
nand U2472 (N_2472,N_2289,N_1732);
or U2473 (N_2473,N_1736,N_2288);
or U2474 (N_2474,N_2195,N_2394);
nand U2475 (N_2475,N_1700,N_2088);
nand U2476 (N_2476,N_1762,N_2071);
nand U2477 (N_2477,N_1742,N_1707);
nand U2478 (N_2478,N_2119,N_2200);
or U2479 (N_2479,N_1907,N_1632);
or U2480 (N_2480,N_1960,N_2247);
xor U2481 (N_2481,N_2130,N_2304);
nand U2482 (N_2482,N_1761,N_1747);
xnor U2483 (N_2483,N_2176,N_2332);
and U2484 (N_2484,N_2227,N_1875);
and U2485 (N_2485,N_2228,N_2147);
or U2486 (N_2486,N_2368,N_1618);
and U2487 (N_2487,N_2128,N_2347);
xor U2488 (N_2488,N_1908,N_2376);
or U2489 (N_2489,N_1866,N_2393);
and U2490 (N_2490,N_1712,N_2275);
and U2491 (N_2491,N_2291,N_1758);
nand U2492 (N_2492,N_2315,N_2386);
nand U2493 (N_2493,N_1626,N_2095);
and U2494 (N_2494,N_1601,N_1925);
xor U2495 (N_2495,N_1714,N_2282);
and U2496 (N_2496,N_1815,N_1958);
nand U2497 (N_2497,N_1604,N_1779);
nor U2498 (N_2498,N_2201,N_2028);
nor U2499 (N_2499,N_2229,N_2156);
and U2500 (N_2500,N_2197,N_1636);
xnor U2501 (N_2501,N_2096,N_2169);
xor U2502 (N_2502,N_1916,N_2043);
nand U2503 (N_2503,N_1688,N_2280);
and U2504 (N_2504,N_2392,N_1709);
nand U2505 (N_2505,N_1705,N_1962);
nor U2506 (N_2506,N_1658,N_2054);
and U2507 (N_2507,N_1765,N_1724);
nand U2508 (N_2508,N_2113,N_1862);
xnor U2509 (N_2509,N_2293,N_2144);
and U2510 (N_2510,N_1885,N_2005);
nor U2511 (N_2511,N_1818,N_2294);
or U2512 (N_2512,N_1970,N_1859);
and U2513 (N_2513,N_2047,N_1871);
and U2514 (N_2514,N_2387,N_1775);
nand U2515 (N_2515,N_1843,N_2023);
nor U2516 (N_2516,N_1693,N_2384);
nand U2517 (N_2517,N_1741,N_2222);
nor U2518 (N_2518,N_2342,N_1832);
xor U2519 (N_2519,N_2326,N_1796);
or U2520 (N_2520,N_1740,N_1888);
xnor U2521 (N_2521,N_1901,N_1799);
and U2522 (N_2522,N_2072,N_1727);
xnor U2523 (N_2523,N_2180,N_1996);
nand U2524 (N_2524,N_1640,N_2328);
and U2525 (N_2525,N_1905,N_2112);
nand U2526 (N_2526,N_2249,N_1772);
and U2527 (N_2527,N_1826,N_1833);
nand U2528 (N_2528,N_1667,N_1820);
and U2529 (N_2529,N_1910,N_1939);
or U2530 (N_2530,N_2181,N_1630);
and U2531 (N_2531,N_1735,N_2066);
and U2532 (N_2532,N_1917,N_1778);
xnor U2533 (N_2533,N_2207,N_2016);
and U2534 (N_2534,N_2135,N_2115);
nand U2535 (N_2535,N_2299,N_1985);
nor U2536 (N_2536,N_2118,N_1987);
xnor U2537 (N_2537,N_2062,N_1824);
nor U2538 (N_2538,N_2308,N_2320);
or U2539 (N_2539,N_1811,N_1648);
or U2540 (N_2540,N_1652,N_2267);
nor U2541 (N_2541,N_2231,N_2212);
nand U2542 (N_2542,N_2061,N_2141);
or U2543 (N_2543,N_1783,N_2341);
xnor U2544 (N_2544,N_2240,N_1831);
nor U2545 (N_2545,N_1738,N_1973);
xnor U2546 (N_2546,N_2007,N_2051);
or U2547 (N_2547,N_1982,N_2285);
nand U2548 (N_2548,N_1890,N_2198);
nor U2549 (N_2549,N_2360,N_1649);
nand U2550 (N_2550,N_2307,N_1773);
nand U2551 (N_2551,N_2367,N_2355);
and U2552 (N_2552,N_1701,N_1858);
nand U2553 (N_2553,N_1754,N_2224);
nand U2554 (N_2554,N_1768,N_2065);
nand U2555 (N_2555,N_1611,N_1681);
xor U2556 (N_2556,N_1968,N_2358);
and U2557 (N_2557,N_2040,N_1674);
nand U2558 (N_2558,N_1813,N_2379);
nor U2559 (N_2559,N_2298,N_1751);
xnor U2560 (N_2560,N_2155,N_1603);
xor U2561 (N_2561,N_2120,N_2236);
nor U2562 (N_2562,N_2219,N_2131);
and U2563 (N_2563,N_2263,N_2262);
xnor U2564 (N_2564,N_2041,N_1782);
xor U2565 (N_2565,N_2046,N_2036);
nand U2566 (N_2566,N_1828,N_1789);
and U2567 (N_2567,N_2260,N_1948);
nand U2568 (N_2568,N_1756,N_2183);
nor U2569 (N_2569,N_1635,N_2114);
nand U2570 (N_2570,N_2127,N_2389);
nor U2571 (N_2571,N_2187,N_2238);
nand U2572 (N_2572,N_2045,N_1899);
and U2573 (N_2573,N_1706,N_2302);
or U2574 (N_2574,N_2152,N_2378);
nor U2575 (N_2575,N_2203,N_1845);
nand U2576 (N_2576,N_1673,N_2287);
nand U2577 (N_2577,N_2015,N_2170);
nand U2578 (N_2578,N_2312,N_2139);
or U2579 (N_2579,N_1839,N_1825);
and U2580 (N_2580,N_2216,N_1794);
nand U2581 (N_2581,N_2014,N_2038);
and U2582 (N_2582,N_2295,N_2080);
xor U2583 (N_2583,N_2101,N_1861);
or U2584 (N_2584,N_2202,N_1608);
or U2585 (N_2585,N_2084,N_2100);
nand U2586 (N_2586,N_1920,N_2148);
xor U2587 (N_2587,N_1663,N_2091);
xnor U2588 (N_2588,N_1734,N_2162);
or U2589 (N_2589,N_2396,N_1912);
nand U2590 (N_2590,N_2322,N_2001);
and U2591 (N_2591,N_1692,N_2372);
or U2592 (N_2592,N_2191,N_2234);
nand U2593 (N_2593,N_1934,N_2252);
or U2594 (N_2594,N_2158,N_2124);
xor U2595 (N_2595,N_1662,N_2002);
nor U2596 (N_2596,N_2166,N_2048);
and U2597 (N_2597,N_1750,N_1723);
xor U2598 (N_2598,N_1941,N_2107);
nor U2599 (N_2599,N_1855,N_2142);
or U2600 (N_2600,N_1729,N_2381);
and U2601 (N_2601,N_2380,N_2385);
nor U2602 (N_2602,N_2214,N_2035);
and U2603 (N_2603,N_2089,N_1650);
and U2604 (N_2604,N_2087,N_2331);
nand U2605 (N_2605,N_1766,N_1919);
or U2606 (N_2606,N_1610,N_2070);
and U2607 (N_2607,N_1696,N_1748);
and U2608 (N_2608,N_1702,N_1949);
nand U2609 (N_2609,N_1848,N_2186);
and U2610 (N_2610,N_2344,N_1938);
nand U2611 (N_2611,N_2388,N_1684);
nor U2612 (N_2612,N_1864,N_2032);
or U2613 (N_2613,N_1671,N_2037);
nor U2614 (N_2614,N_1805,N_2327);
and U2615 (N_2615,N_1990,N_1721);
nand U2616 (N_2616,N_2345,N_1894);
nor U2617 (N_2617,N_2319,N_2013);
and U2618 (N_2618,N_1857,N_1959);
nand U2619 (N_2619,N_2161,N_1965);
xnor U2620 (N_2620,N_2349,N_1669);
nor U2621 (N_2621,N_2104,N_1836);
nand U2622 (N_2622,N_1981,N_1703);
or U2623 (N_2623,N_2109,N_2138);
or U2624 (N_2624,N_1680,N_2019);
and U2625 (N_2625,N_2271,N_1620);
or U2626 (N_2626,N_1914,N_1922);
nand U2627 (N_2627,N_2254,N_2090);
xor U2628 (N_2628,N_2182,N_2024);
nand U2629 (N_2629,N_1708,N_1937);
and U2630 (N_2630,N_2076,N_2058);
nand U2631 (N_2631,N_2309,N_2117);
or U2632 (N_2632,N_2122,N_2020);
nor U2633 (N_2633,N_1808,N_1997);
and U2634 (N_2634,N_1623,N_2167);
nand U2635 (N_2635,N_1840,N_2338);
xor U2636 (N_2636,N_2073,N_2346);
nand U2637 (N_2637,N_2230,N_2157);
nor U2638 (N_2638,N_1803,N_1685);
xor U2639 (N_2639,N_1876,N_1634);
nor U2640 (N_2640,N_2264,N_1842);
and U2641 (N_2641,N_2323,N_2194);
nand U2642 (N_2642,N_2241,N_2081);
xor U2643 (N_2643,N_2250,N_1957);
nor U2644 (N_2644,N_1812,N_1896);
nor U2645 (N_2645,N_1682,N_2395);
and U2646 (N_2646,N_1979,N_1928);
nand U2647 (N_2647,N_1963,N_1954);
nand U2648 (N_2648,N_1880,N_2143);
and U2649 (N_2649,N_2375,N_2185);
xnor U2650 (N_2650,N_1942,N_1699);
and U2651 (N_2651,N_1913,N_1886);
xor U2652 (N_2652,N_2281,N_1659);
nor U2653 (N_2653,N_1757,N_1950);
or U2654 (N_2654,N_1755,N_1953);
xor U2655 (N_2655,N_1992,N_1945);
xnor U2656 (N_2656,N_2223,N_2042);
xor U2657 (N_2657,N_2325,N_2108);
nor U2658 (N_2658,N_2031,N_1749);
nor U2659 (N_2659,N_1666,N_2351);
and U2660 (N_2660,N_1691,N_1853);
nor U2661 (N_2661,N_1655,N_2397);
nor U2662 (N_2662,N_2004,N_1877);
xnor U2663 (N_2663,N_1752,N_1777);
xnor U2664 (N_2664,N_2232,N_2276);
xor U2665 (N_2665,N_1881,N_1924);
nand U2666 (N_2666,N_1984,N_1902);
nor U2667 (N_2667,N_2094,N_1854);
and U2668 (N_2668,N_2364,N_2009);
and U2669 (N_2669,N_1819,N_2146);
xnor U2670 (N_2670,N_1838,N_2246);
and U2671 (N_2671,N_1852,N_1993);
xnor U2672 (N_2672,N_1974,N_1619);
nand U2673 (N_2673,N_2021,N_1882);
nor U2674 (N_2674,N_2300,N_2172);
xnor U2675 (N_2675,N_1827,N_2192);
or U2676 (N_2676,N_2171,N_2067);
or U2677 (N_2677,N_2103,N_2277);
nand U2678 (N_2678,N_1872,N_1798);
nand U2679 (N_2679,N_2049,N_2092);
nor U2680 (N_2680,N_2098,N_2074);
nor U2681 (N_2681,N_1722,N_1883);
nand U2682 (N_2682,N_2033,N_2204);
nor U2683 (N_2683,N_2097,N_1657);
and U2684 (N_2684,N_2259,N_1887);
or U2685 (N_2685,N_2110,N_2160);
xor U2686 (N_2686,N_1952,N_1923);
and U2687 (N_2687,N_2321,N_1800);
xor U2688 (N_2688,N_1690,N_1785);
nor U2689 (N_2689,N_1651,N_1900);
nand U2690 (N_2690,N_2134,N_1977);
or U2691 (N_2691,N_1683,N_2390);
nor U2692 (N_2692,N_2373,N_2377);
or U2693 (N_2693,N_1994,N_2205);
or U2694 (N_2694,N_1641,N_2316);
and U2695 (N_2695,N_2383,N_2068);
xor U2696 (N_2696,N_1617,N_2085);
xnor U2697 (N_2697,N_2017,N_1637);
and U2698 (N_2698,N_1988,N_1769);
xnor U2699 (N_2699,N_1629,N_2140);
or U2700 (N_2700,N_1884,N_1639);
xor U2701 (N_2701,N_1711,N_2105);
or U2702 (N_2702,N_2059,N_2369);
nand U2703 (N_2703,N_1835,N_2189);
nand U2704 (N_2704,N_2337,N_2057);
nor U2705 (N_2705,N_1807,N_2083);
xor U2706 (N_2706,N_2270,N_1602);
nand U2707 (N_2707,N_1870,N_1737);
and U2708 (N_2708,N_1733,N_2211);
and U2709 (N_2709,N_1929,N_2366);
nor U2710 (N_2710,N_1869,N_2179);
nand U2711 (N_2711,N_2362,N_1646);
nor U2712 (N_2712,N_2082,N_1851);
xor U2713 (N_2713,N_2034,N_2225);
and U2714 (N_2714,N_2196,N_2382);
and U2715 (N_2715,N_1633,N_1676);
xor U2716 (N_2716,N_2336,N_2269);
nor U2717 (N_2717,N_2363,N_2251);
and U2718 (N_2718,N_2334,N_2064);
nor U2719 (N_2719,N_1767,N_1878);
nor U2720 (N_2720,N_1850,N_2303);
nor U2721 (N_2721,N_1731,N_1810);
xnor U2722 (N_2722,N_1816,N_1983);
and U2723 (N_2723,N_2265,N_2022);
nor U2724 (N_2724,N_1874,N_1898);
and U2725 (N_2725,N_1847,N_1976);
nand U2726 (N_2726,N_2012,N_2154);
xor U2727 (N_2727,N_2164,N_2398);
xor U2728 (N_2728,N_1694,N_2077);
xor U2729 (N_2729,N_2374,N_2243);
nor U2730 (N_2730,N_2301,N_2000);
nor U2731 (N_2731,N_2102,N_2184);
or U2732 (N_2732,N_1614,N_1969);
and U2733 (N_2733,N_2340,N_1931);
xor U2734 (N_2734,N_1936,N_2011);
nor U2735 (N_2735,N_1933,N_1660);
nand U2736 (N_2736,N_2311,N_2361);
nand U2737 (N_2737,N_2333,N_1986);
xor U2738 (N_2738,N_1745,N_2178);
nor U2739 (N_2739,N_2290,N_1868);
or U2740 (N_2740,N_1622,N_1909);
xor U2741 (N_2741,N_2283,N_2370);
or U2742 (N_2742,N_2296,N_1955);
nand U2743 (N_2743,N_2060,N_2213);
or U2744 (N_2744,N_2310,N_1944);
xor U2745 (N_2745,N_1915,N_1786);
and U2746 (N_2746,N_2150,N_1631);
xnor U2747 (N_2747,N_2266,N_1788);
xor U2748 (N_2748,N_1998,N_2055);
or U2749 (N_2749,N_2330,N_2030);
and U2750 (N_2750,N_1780,N_2210);
nand U2751 (N_2751,N_1809,N_2239);
nor U2752 (N_2752,N_1759,N_1930);
xnor U2753 (N_2753,N_2133,N_1947);
xor U2754 (N_2754,N_1697,N_1704);
and U2755 (N_2755,N_1903,N_1897);
nor U2756 (N_2756,N_1689,N_1615);
xor U2757 (N_2757,N_1889,N_2116);
nand U2758 (N_2758,N_2145,N_2039);
nor U2759 (N_2759,N_2206,N_1784);
nor U2760 (N_2760,N_1605,N_2151);
xnor U2761 (N_2761,N_1849,N_1841);
nor U2762 (N_2762,N_2256,N_1797);
and U2763 (N_2763,N_2242,N_1771);
nand U2764 (N_2764,N_2354,N_1665);
nor U2765 (N_2765,N_1830,N_1921);
or U2766 (N_2766,N_1964,N_1867);
nor U2767 (N_2767,N_2052,N_1718);
nor U2768 (N_2768,N_1746,N_2175);
and U2769 (N_2769,N_2274,N_1675);
nor U2770 (N_2770,N_1806,N_1710);
and U2771 (N_2771,N_2121,N_2126);
nor U2772 (N_2772,N_2221,N_1846);
nor U2773 (N_2773,N_1999,N_2292);
xnor U2774 (N_2774,N_1720,N_1743);
nand U2775 (N_2775,N_2137,N_1895);
nand U2776 (N_2776,N_1793,N_1817);
nand U2777 (N_2777,N_1821,N_2233);
nand U2778 (N_2778,N_1975,N_1837);
xnor U2779 (N_2779,N_2136,N_1661);
nand U2780 (N_2780,N_1600,N_1829);
nand U2781 (N_2781,N_2199,N_1792);
nor U2782 (N_2782,N_2279,N_2018);
xor U2783 (N_2783,N_1628,N_2159);
nor U2784 (N_2784,N_2237,N_1790);
nand U2785 (N_2785,N_1764,N_2257);
xor U2786 (N_2786,N_1607,N_1616);
nand U2787 (N_2787,N_1625,N_1678);
nor U2788 (N_2788,N_2025,N_2314);
nand U2789 (N_2789,N_2306,N_1940);
xor U2790 (N_2790,N_2106,N_2244);
and U2791 (N_2791,N_1801,N_2318);
and U2792 (N_2792,N_2329,N_1995);
and U2793 (N_2793,N_1638,N_1804);
xnor U2794 (N_2794,N_2168,N_1686);
or U2795 (N_2795,N_1774,N_1672);
and U2796 (N_2796,N_1609,N_2235);
nand U2797 (N_2797,N_1739,N_1653);
nor U2798 (N_2798,N_2248,N_1893);
or U2799 (N_2799,N_1892,N_2053);
or U2800 (N_2800,N_2128,N_2229);
nand U2801 (N_2801,N_1767,N_1936);
nor U2802 (N_2802,N_1745,N_2208);
nand U2803 (N_2803,N_1727,N_1794);
nor U2804 (N_2804,N_2361,N_1922);
or U2805 (N_2805,N_1742,N_2003);
or U2806 (N_2806,N_2066,N_2248);
or U2807 (N_2807,N_1606,N_2102);
or U2808 (N_2808,N_2332,N_1780);
xor U2809 (N_2809,N_2251,N_1618);
or U2810 (N_2810,N_2011,N_1743);
nor U2811 (N_2811,N_2038,N_1724);
and U2812 (N_2812,N_2395,N_1804);
nand U2813 (N_2813,N_2318,N_1808);
or U2814 (N_2814,N_1879,N_2382);
or U2815 (N_2815,N_2133,N_1608);
nand U2816 (N_2816,N_2227,N_1935);
and U2817 (N_2817,N_2183,N_1868);
xnor U2818 (N_2818,N_2215,N_2328);
xnor U2819 (N_2819,N_1804,N_2054);
nand U2820 (N_2820,N_2207,N_1851);
xor U2821 (N_2821,N_1888,N_1904);
and U2822 (N_2822,N_2148,N_1897);
and U2823 (N_2823,N_1871,N_2295);
and U2824 (N_2824,N_1756,N_1921);
xor U2825 (N_2825,N_1832,N_1871);
xnor U2826 (N_2826,N_1960,N_2041);
nor U2827 (N_2827,N_1728,N_1945);
xnor U2828 (N_2828,N_2110,N_1735);
nand U2829 (N_2829,N_2385,N_1661);
or U2830 (N_2830,N_1709,N_2233);
nand U2831 (N_2831,N_1834,N_2303);
and U2832 (N_2832,N_2320,N_2208);
or U2833 (N_2833,N_1707,N_1922);
or U2834 (N_2834,N_1608,N_1617);
or U2835 (N_2835,N_1696,N_2065);
nor U2836 (N_2836,N_2278,N_1866);
xor U2837 (N_2837,N_2270,N_2245);
and U2838 (N_2838,N_2339,N_1844);
nand U2839 (N_2839,N_1711,N_1730);
xnor U2840 (N_2840,N_1650,N_1943);
nor U2841 (N_2841,N_2384,N_1936);
nand U2842 (N_2842,N_1928,N_2188);
xnor U2843 (N_2843,N_2188,N_2120);
nor U2844 (N_2844,N_2251,N_1796);
and U2845 (N_2845,N_2314,N_2122);
nand U2846 (N_2846,N_2211,N_2126);
nand U2847 (N_2847,N_1655,N_1910);
nand U2848 (N_2848,N_1717,N_1889);
nand U2849 (N_2849,N_1910,N_1854);
and U2850 (N_2850,N_2373,N_2037);
or U2851 (N_2851,N_2241,N_1855);
and U2852 (N_2852,N_2024,N_1939);
and U2853 (N_2853,N_2360,N_2268);
xor U2854 (N_2854,N_2295,N_1631);
nor U2855 (N_2855,N_1777,N_1691);
nor U2856 (N_2856,N_2125,N_1663);
nand U2857 (N_2857,N_2075,N_1798);
xnor U2858 (N_2858,N_1601,N_2132);
nor U2859 (N_2859,N_2314,N_2017);
nor U2860 (N_2860,N_1844,N_2384);
and U2861 (N_2861,N_2362,N_1612);
xnor U2862 (N_2862,N_1752,N_1935);
or U2863 (N_2863,N_1864,N_2091);
or U2864 (N_2864,N_1654,N_1862);
and U2865 (N_2865,N_1726,N_2073);
nor U2866 (N_2866,N_2024,N_2207);
nor U2867 (N_2867,N_2034,N_2191);
nor U2868 (N_2868,N_2125,N_2040);
nor U2869 (N_2869,N_2090,N_2374);
or U2870 (N_2870,N_2024,N_1849);
nor U2871 (N_2871,N_1869,N_2105);
or U2872 (N_2872,N_2084,N_1661);
nand U2873 (N_2873,N_1810,N_2051);
xor U2874 (N_2874,N_1959,N_1740);
nor U2875 (N_2875,N_1929,N_2118);
xor U2876 (N_2876,N_2245,N_1839);
and U2877 (N_2877,N_1849,N_2115);
xor U2878 (N_2878,N_1814,N_1802);
or U2879 (N_2879,N_1805,N_1725);
and U2880 (N_2880,N_2363,N_1608);
nor U2881 (N_2881,N_2102,N_1830);
xnor U2882 (N_2882,N_2113,N_2159);
nor U2883 (N_2883,N_1885,N_2272);
or U2884 (N_2884,N_1622,N_1809);
or U2885 (N_2885,N_2053,N_2394);
and U2886 (N_2886,N_2207,N_1819);
nand U2887 (N_2887,N_1732,N_1863);
or U2888 (N_2888,N_2375,N_2292);
xor U2889 (N_2889,N_2180,N_1789);
or U2890 (N_2890,N_1740,N_1631);
xnor U2891 (N_2891,N_2170,N_2237);
nor U2892 (N_2892,N_1747,N_1700);
and U2893 (N_2893,N_1809,N_1653);
or U2894 (N_2894,N_1632,N_2377);
xor U2895 (N_2895,N_2350,N_2191);
nor U2896 (N_2896,N_2145,N_1626);
and U2897 (N_2897,N_2076,N_2143);
and U2898 (N_2898,N_1941,N_1776);
xnor U2899 (N_2899,N_2324,N_1917);
and U2900 (N_2900,N_1678,N_2050);
nor U2901 (N_2901,N_2354,N_1963);
nor U2902 (N_2902,N_2192,N_2036);
and U2903 (N_2903,N_2174,N_2175);
xnor U2904 (N_2904,N_2346,N_2349);
and U2905 (N_2905,N_2392,N_2208);
or U2906 (N_2906,N_2245,N_1788);
nand U2907 (N_2907,N_2180,N_2024);
nor U2908 (N_2908,N_1953,N_2192);
or U2909 (N_2909,N_2355,N_2377);
or U2910 (N_2910,N_1999,N_1672);
nor U2911 (N_2911,N_1674,N_1812);
or U2912 (N_2912,N_2064,N_2169);
and U2913 (N_2913,N_2338,N_1959);
nand U2914 (N_2914,N_1724,N_2172);
xnor U2915 (N_2915,N_2347,N_1675);
and U2916 (N_2916,N_2139,N_1798);
and U2917 (N_2917,N_2164,N_1838);
or U2918 (N_2918,N_1708,N_1700);
or U2919 (N_2919,N_2152,N_2287);
or U2920 (N_2920,N_2104,N_1799);
xnor U2921 (N_2921,N_2237,N_1691);
nand U2922 (N_2922,N_2244,N_2000);
and U2923 (N_2923,N_1658,N_1759);
xor U2924 (N_2924,N_1934,N_1796);
and U2925 (N_2925,N_1654,N_1861);
or U2926 (N_2926,N_2165,N_1918);
or U2927 (N_2927,N_2340,N_1727);
xnor U2928 (N_2928,N_1933,N_1819);
nand U2929 (N_2929,N_1660,N_2060);
and U2930 (N_2930,N_2331,N_2178);
xnor U2931 (N_2931,N_1846,N_2169);
or U2932 (N_2932,N_2267,N_1693);
or U2933 (N_2933,N_1636,N_2370);
xnor U2934 (N_2934,N_1785,N_2224);
or U2935 (N_2935,N_1949,N_1835);
nor U2936 (N_2936,N_1733,N_1825);
xor U2937 (N_2937,N_1758,N_2122);
xor U2938 (N_2938,N_1653,N_1938);
xnor U2939 (N_2939,N_2350,N_1691);
xnor U2940 (N_2940,N_2245,N_2040);
nor U2941 (N_2941,N_1824,N_1711);
xor U2942 (N_2942,N_2108,N_1858);
nor U2943 (N_2943,N_2374,N_1658);
and U2944 (N_2944,N_2147,N_1609);
or U2945 (N_2945,N_1664,N_2211);
and U2946 (N_2946,N_2044,N_2278);
xor U2947 (N_2947,N_2324,N_2277);
nand U2948 (N_2948,N_2011,N_1769);
and U2949 (N_2949,N_1986,N_2270);
nor U2950 (N_2950,N_2128,N_1795);
nand U2951 (N_2951,N_1637,N_1754);
nor U2952 (N_2952,N_1874,N_2096);
and U2953 (N_2953,N_2350,N_1654);
nand U2954 (N_2954,N_1958,N_2331);
nor U2955 (N_2955,N_2233,N_2122);
nor U2956 (N_2956,N_2015,N_2031);
nand U2957 (N_2957,N_1800,N_2335);
nor U2958 (N_2958,N_1911,N_2124);
nand U2959 (N_2959,N_2072,N_1640);
xnor U2960 (N_2960,N_2065,N_1870);
nand U2961 (N_2961,N_1739,N_2138);
nand U2962 (N_2962,N_1982,N_1706);
nand U2963 (N_2963,N_2000,N_2320);
and U2964 (N_2964,N_1852,N_1738);
xnor U2965 (N_2965,N_1916,N_2220);
xor U2966 (N_2966,N_2246,N_2264);
nor U2967 (N_2967,N_2299,N_2381);
nand U2968 (N_2968,N_2022,N_2273);
nor U2969 (N_2969,N_1810,N_1814);
or U2970 (N_2970,N_1987,N_1807);
nor U2971 (N_2971,N_2044,N_1670);
xor U2972 (N_2972,N_2035,N_1798);
or U2973 (N_2973,N_2224,N_1827);
or U2974 (N_2974,N_1832,N_2022);
and U2975 (N_2975,N_2232,N_1847);
nand U2976 (N_2976,N_2261,N_2138);
xnor U2977 (N_2977,N_2271,N_1837);
or U2978 (N_2978,N_1921,N_2158);
or U2979 (N_2979,N_1839,N_1889);
or U2980 (N_2980,N_1740,N_1621);
and U2981 (N_2981,N_1842,N_2364);
and U2982 (N_2982,N_1730,N_2367);
nor U2983 (N_2983,N_2190,N_2212);
xor U2984 (N_2984,N_2045,N_1875);
or U2985 (N_2985,N_1612,N_2167);
xnor U2986 (N_2986,N_2072,N_2303);
nand U2987 (N_2987,N_1659,N_2066);
and U2988 (N_2988,N_2238,N_1869);
nand U2989 (N_2989,N_2313,N_2053);
nor U2990 (N_2990,N_1802,N_1707);
xnor U2991 (N_2991,N_2346,N_2121);
nand U2992 (N_2992,N_1800,N_2251);
nand U2993 (N_2993,N_2218,N_2104);
xor U2994 (N_2994,N_1961,N_2018);
nand U2995 (N_2995,N_2220,N_2204);
nor U2996 (N_2996,N_1651,N_2171);
xnor U2997 (N_2997,N_2133,N_2165);
and U2998 (N_2998,N_1873,N_1817);
nand U2999 (N_2999,N_1692,N_2056);
and U3000 (N_3000,N_1629,N_1910);
nand U3001 (N_3001,N_2237,N_2193);
or U3002 (N_3002,N_2150,N_1714);
and U3003 (N_3003,N_2084,N_2300);
and U3004 (N_3004,N_2375,N_1737);
and U3005 (N_3005,N_2120,N_1914);
or U3006 (N_3006,N_1629,N_1735);
or U3007 (N_3007,N_1665,N_2258);
and U3008 (N_3008,N_1927,N_1827);
and U3009 (N_3009,N_1784,N_1968);
and U3010 (N_3010,N_2268,N_2279);
nand U3011 (N_3011,N_2062,N_2181);
nor U3012 (N_3012,N_2205,N_2275);
xor U3013 (N_3013,N_2381,N_1876);
nand U3014 (N_3014,N_2344,N_2069);
nand U3015 (N_3015,N_1918,N_1890);
nand U3016 (N_3016,N_2225,N_2215);
or U3017 (N_3017,N_2195,N_2324);
and U3018 (N_3018,N_1728,N_2293);
nor U3019 (N_3019,N_2053,N_1773);
and U3020 (N_3020,N_2185,N_1765);
and U3021 (N_3021,N_1809,N_1871);
xor U3022 (N_3022,N_1735,N_1875);
xnor U3023 (N_3023,N_1733,N_1901);
and U3024 (N_3024,N_1842,N_2031);
nand U3025 (N_3025,N_1780,N_1744);
xor U3026 (N_3026,N_1952,N_1960);
xor U3027 (N_3027,N_1616,N_1646);
nor U3028 (N_3028,N_1944,N_1687);
or U3029 (N_3029,N_1957,N_2249);
and U3030 (N_3030,N_2163,N_2185);
or U3031 (N_3031,N_2044,N_1667);
nand U3032 (N_3032,N_2213,N_2135);
and U3033 (N_3033,N_1856,N_2175);
and U3034 (N_3034,N_1985,N_1608);
nand U3035 (N_3035,N_1814,N_2227);
or U3036 (N_3036,N_1921,N_1936);
nor U3037 (N_3037,N_1730,N_1673);
or U3038 (N_3038,N_1857,N_1889);
nor U3039 (N_3039,N_1636,N_1909);
nor U3040 (N_3040,N_2090,N_1789);
nand U3041 (N_3041,N_2195,N_1984);
nand U3042 (N_3042,N_2038,N_1924);
and U3043 (N_3043,N_2226,N_2140);
xor U3044 (N_3044,N_1921,N_2004);
nor U3045 (N_3045,N_2264,N_1916);
and U3046 (N_3046,N_1984,N_2370);
and U3047 (N_3047,N_1847,N_1896);
xnor U3048 (N_3048,N_1639,N_2052);
nor U3049 (N_3049,N_1988,N_1801);
xor U3050 (N_3050,N_1908,N_1990);
nand U3051 (N_3051,N_1911,N_1708);
or U3052 (N_3052,N_1733,N_1613);
xor U3053 (N_3053,N_1772,N_1965);
or U3054 (N_3054,N_1653,N_1661);
nand U3055 (N_3055,N_1886,N_1616);
xor U3056 (N_3056,N_2144,N_2143);
nand U3057 (N_3057,N_2228,N_2195);
xnor U3058 (N_3058,N_1711,N_2159);
nand U3059 (N_3059,N_1813,N_2080);
and U3060 (N_3060,N_1628,N_1930);
or U3061 (N_3061,N_2161,N_2392);
nand U3062 (N_3062,N_1992,N_2200);
nor U3063 (N_3063,N_1612,N_2177);
xor U3064 (N_3064,N_1894,N_1804);
or U3065 (N_3065,N_2352,N_2038);
xor U3066 (N_3066,N_1786,N_2180);
xnor U3067 (N_3067,N_1936,N_2301);
or U3068 (N_3068,N_2104,N_1742);
nor U3069 (N_3069,N_2125,N_1865);
nand U3070 (N_3070,N_1742,N_1834);
nor U3071 (N_3071,N_1784,N_1668);
nand U3072 (N_3072,N_1864,N_1852);
xor U3073 (N_3073,N_1676,N_1758);
xnor U3074 (N_3074,N_1730,N_2058);
nor U3075 (N_3075,N_2282,N_1656);
nand U3076 (N_3076,N_2035,N_1849);
nor U3077 (N_3077,N_2279,N_1864);
nor U3078 (N_3078,N_1887,N_2203);
and U3079 (N_3079,N_1612,N_2299);
xnor U3080 (N_3080,N_1844,N_2214);
nor U3081 (N_3081,N_2198,N_2063);
nand U3082 (N_3082,N_1808,N_1658);
xor U3083 (N_3083,N_2311,N_2365);
xor U3084 (N_3084,N_1892,N_2334);
nand U3085 (N_3085,N_1628,N_2306);
nor U3086 (N_3086,N_1630,N_2201);
xnor U3087 (N_3087,N_1986,N_2255);
and U3088 (N_3088,N_2204,N_1973);
or U3089 (N_3089,N_2161,N_1768);
xnor U3090 (N_3090,N_2120,N_1826);
nor U3091 (N_3091,N_1867,N_1730);
xnor U3092 (N_3092,N_1867,N_2102);
and U3093 (N_3093,N_1784,N_2219);
nand U3094 (N_3094,N_1966,N_1840);
nand U3095 (N_3095,N_2132,N_2032);
xor U3096 (N_3096,N_1851,N_1646);
and U3097 (N_3097,N_2332,N_1731);
nor U3098 (N_3098,N_1976,N_2365);
xor U3099 (N_3099,N_1629,N_1641);
or U3100 (N_3100,N_2232,N_1826);
nor U3101 (N_3101,N_1842,N_1941);
or U3102 (N_3102,N_1968,N_1631);
nand U3103 (N_3103,N_1768,N_2106);
and U3104 (N_3104,N_1769,N_2224);
and U3105 (N_3105,N_2346,N_2214);
nand U3106 (N_3106,N_1845,N_2186);
and U3107 (N_3107,N_2041,N_1801);
nand U3108 (N_3108,N_1781,N_2106);
or U3109 (N_3109,N_1682,N_2365);
and U3110 (N_3110,N_2199,N_1603);
nand U3111 (N_3111,N_2093,N_1627);
xor U3112 (N_3112,N_1962,N_2026);
xnor U3113 (N_3113,N_1941,N_1874);
and U3114 (N_3114,N_2377,N_2216);
or U3115 (N_3115,N_2072,N_2171);
xnor U3116 (N_3116,N_1970,N_1860);
or U3117 (N_3117,N_2191,N_2225);
nand U3118 (N_3118,N_2161,N_2357);
or U3119 (N_3119,N_1880,N_1626);
xnor U3120 (N_3120,N_1677,N_1918);
nor U3121 (N_3121,N_1674,N_1808);
xnor U3122 (N_3122,N_2142,N_1771);
xor U3123 (N_3123,N_2233,N_1856);
and U3124 (N_3124,N_2274,N_2343);
and U3125 (N_3125,N_2069,N_1735);
xnor U3126 (N_3126,N_1859,N_1705);
nor U3127 (N_3127,N_2051,N_2182);
xnor U3128 (N_3128,N_2339,N_1919);
or U3129 (N_3129,N_1688,N_2251);
xor U3130 (N_3130,N_1642,N_2266);
nor U3131 (N_3131,N_2187,N_2180);
xor U3132 (N_3132,N_1812,N_2031);
or U3133 (N_3133,N_1602,N_2220);
or U3134 (N_3134,N_2096,N_2219);
or U3135 (N_3135,N_1758,N_1806);
or U3136 (N_3136,N_1686,N_1603);
and U3137 (N_3137,N_1769,N_2238);
nor U3138 (N_3138,N_1917,N_1689);
nand U3139 (N_3139,N_2352,N_2288);
nand U3140 (N_3140,N_1861,N_1974);
xor U3141 (N_3141,N_1786,N_2273);
or U3142 (N_3142,N_1904,N_2293);
xor U3143 (N_3143,N_2273,N_2046);
or U3144 (N_3144,N_2043,N_2233);
nor U3145 (N_3145,N_2081,N_1730);
or U3146 (N_3146,N_2272,N_1734);
and U3147 (N_3147,N_1651,N_2322);
and U3148 (N_3148,N_1981,N_1600);
or U3149 (N_3149,N_1960,N_2328);
nor U3150 (N_3150,N_1748,N_1687);
nor U3151 (N_3151,N_1908,N_2292);
nor U3152 (N_3152,N_2277,N_1924);
nand U3153 (N_3153,N_2038,N_1752);
nand U3154 (N_3154,N_2274,N_2016);
nand U3155 (N_3155,N_2243,N_2258);
and U3156 (N_3156,N_1795,N_1771);
and U3157 (N_3157,N_2032,N_2093);
nor U3158 (N_3158,N_1970,N_1858);
nor U3159 (N_3159,N_1875,N_2001);
xor U3160 (N_3160,N_1892,N_1744);
nor U3161 (N_3161,N_1879,N_2259);
nor U3162 (N_3162,N_2090,N_1864);
nand U3163 (N_3163,N_2120,N_1815);
and U3164 (N_3164,N_1898,N_2102);
xor U3165 (N_3165,N_2062,N_2163);
xnor U3166 (N_3166,N_2037,N_1934);
nand U3167 (N_3167,N_2321,N_1664);
or U3168 (N_3168,N_1697,N_2325);
and U3169 (N_3169,N_2252,N_2083);
nand U3170 (N_3170,N_1914,N_2056);
or U3171 (N_3171,N_2055,N_2180);
and U3172 (N_3172,N_1935,N_1915);
nand U3173 (N_3173,N_2364,N_2145);
or U3174 (N_3174,N_2132,N_1950);
or U3175 (N_3175,N_1718,N_1940);
xnor U3176 (N_3176,N_2047,N_2204);
nor U3177 (N_3177,N_2093,N_1676);
xnor U3178 (N_3178,N_2164,N_1833);
xor U3179 (N_3179,N_1856,N_2289);
and U3180 (N_3180,N_1866,N_2339);
nor U3181 (N_3181,N_2085,N_1917);
nand U3182 (N_3182,N_1608,N_2362);
xor U3183 (N_3183,N_2232,N_1944);
or U3184 (N_3184,N_1932,N_2147);
and U3185 (N_3185,N_2360,N_2306);
or U3186 (N_3186,N_2203,N_2034);
nand U3187 (N_3187,N_1812,N_2342);
nand U3188 (N_3188,N_1785,N_1996);
nand U3189 (N_3189,N_1701,N_2318);
nor U3190 (N_3190,N_2253,N_1804);
nand U3191 (N_3191,N_2183,N_1948);
or U3192 (N_3192,N_1611,N_2394);
nor U3193 (N_3193,N_1941,N_1718);
nand U3194 (N_3194,N_2282,N_2291);
nand U3195 (N_3195,N_2309,N_2316);
or U3196 (N_3196,N_2346,N_2331);
and U3197 (N_3197,N_1838,N_1963);
or U3198 (N_3198,N_2122,N_1868);
xor U3199 (N_3199,N_1982,N_2366);
nand U3200 (N_3200,N_2461,N_2963);
nor U3201 (N_3201,N_2809,N_2422);
nor U3202 (N_3202,N_2951,N_2686);
nand U3203 (N_3203,N_2827,N_3112);
xnor U3204 (N_3204,N_2757,N_2705);
xnor U3205 (N_3205,N_2980,N_2981);
or U3206 (N_3206,N_3107,N_2846);
xnor U3207 (N_3207,N_2564,N_2822);
nor U3208 (N_3208,N_3173,N_2707);
and U3209 (N_3209,N_2685,N_2756);
xnor U3210 (N_3210,N_2887,N_2484);
and U3211 (N_3211,N_2494,N_2715);
xor U3212 (N_3212,N_2872,N_3087);
or U3213 (N_3213,N_3136,N_2433);
nand U3214 (N_3214,N_3005,N_2733);
nor U3215 (N_3215,N_2547,N_2878);
xnor U3216 (N_3216,N_3039,N_3079);
xor U3217 (N_3217,N_2505,N_2719);
and U3218 (N_3218,N_2613,N_2590);
nor U3219 (N_3219,N_2536,N_2475);
nand U3220 (N_3220,N_2879,N_3180);
xnor U3221 (N_3221,N_2896,N_2565);
xor U3222 (N_3222,N_3065,N_3046);
and U3223 (N_3223,N_2902,N_3069);
and U3224 (N_3224,N_3125,N_2845);
nor U3225 (N_3225,N_2904,N_2633);
xor U3226 (N_3226,N_3068,N_2936);
or U3227 (N_3227,N_2688,N_2413);
nor U3228 (N_3228,N_2894,N_2541);
nor U3229 (N_3229,N_2730,N_2932);
and U3230 (N_3230,N_2425,N_2670);
xnor U3231 (N_3231,N_2698,N_3137);
nand U3232 (N_3232,N_2403,N_2499);
nor U3233 (N_3233,N_2438,N_2741);
or U3234 (N_3234,N_3105,N_2824);
xnor U3235 (N_3235,N_2549,N_2501);
or U3236 (N_3236,N_2695,N_3031);
nor U3237 (N_3237,N_2857,N_2877);
and U3238 (N_3238,N_2610,N_2917);
nand U3239 (N_3239,N_2456,N_2566);
xnor U3240 (N_3240,N_2570,N_3074);
nand U3241 (N_3241,N_2407,N_2453);
nor U3242 (N_3242,N_2799,N_2411);
or U3243 (N_3243,N_2417,N_3062);
and U3244 (N_3244,N_3002,N_3148);
and U3245 (N_3245,N_2490,N_2677);
or U3246 (N_3246,N_2717,N_2623);
nor U3247 (N_3247,N_2660,N_2933);
and U3248 (N_3248,N_2989,N_2476);
nor U3249 (N_3249,N_2955,N_3055);
xor U3250 (N_3250,N_2588,N_3072);
or U3251 (N_3251,N_2840,N_2638);
nor U3252 (N_3252,N_3142,N_3108);
nand U3253 (N_3253,N_3182,N_3047);
nand U3254 (N_3254,N_2632,N_2589);
xnor U3255 (N_3255,N_3028,N_2778);
xor U3256 (N_3256,N_3004,N_3163);
xnor U3257 (N_3257,N_3167,N_2515);
and U3258 (N_3258,N_3151,N_3035);
and U3259 (N_3259,N_2574,N_3132);
nor U3260 (N_3260,N_2627,N_3126);
or U3261 (N_3261,N_3071,N_2584);
nor U3262 (N_3262,N_3038,N_2918);
nand U3263 (N_3263,N_3017,N_2777);
and U3264 (N_3264,N_2703,N_2498);
nor U3265 (N_3265,N_3129,N_2487);
or U3266 (N_3266,N_2750,N_2443);
nor U3267 (N_3267,N_2938,N_3044);
and U3268 (N_3268,N_2483,N_3048);
nand U3269 (N_3269,N_2539,N_2726);
nor U3270 (N_3270,N_2661,N_2650);
nor U3271 (N_3271,N_2713,N_3011);
nand U3272 (N_3272,N_2659,N_2924);
nand U3273 (N_3273,N_3141,N_2434);
and U3274 (N_3274,N_2897,N_2493);
and U3275 (N_3275,N_2457,N_2782);
xor U3276 (N_3276,N_2429,N_2497);
xor U3277 (N_3277,N_2943,N_3030);
xnor U3278 (N_3278,N_3159,N_2520);
nand U3279 (N_3279,N_2736,N_2546);
xnor U3280 (N_3280,N_2690,N_2751);
and U3281 (N_3281,N_2595,N_2694);
nor U3282 (N_3282,N_3152,N_3059);
or U3283 (N_3283,N_3149,N_2807);
nor U3284 (N_3284,N_2855,N_3088);
or U3285 (N_3285,N_3109,N_2854);
nor U3286 (N_3286,N_3012,N_3093);
xnor U3287 (N_3287,N_2492,N_3040);
nand U3288 (N_3288,N_2916,N_3084);
nand U3289 (N_3289,N_2525,N_2519);
xnor U3290 (N_3290,N_3155,N_2709);
or U3291 (N_3291,N_2985,N_2880);
and U3292 (N_3292,N_2728,N_2825);
nor U3293 (N_3293,N_2678,N_2727);
nor U3294 (N_3294,N_3122,N_2802);
and U3295 (N_3295,N_2965,N_2876);
nand U3296 (N_3296,N_2585,N_3172);
nor U3297 (N_3297,N_2945,N_2581);
and U3298 (N_3298,N_2642,N_2463);
and U3299 (N_3299,N_2982,N_2763);
or U3300 (N_3300,N_3123,N_2758);
nand U3301 (N_3301,N_2604,N_2785);
or U3302 (N_3302,N_3061,N_2408);
nand U3303 (N_3303,N_3086,N_3041);
nor U3304 (N_3304,N_2754,N_3058);
or U3305 (N_3305,N_2808,N_2439);
and U3306 (N_3306,N_2591,N_2423);
and U3307 (N_3307,N_2409,N_3196);
nor U3308 (N_3308,N_2962,N_2991);
and U3309 (N_3309,N_2597,N_2614);
xor U3310 (N_3310,N_2972,N_2533);
nand U3311 (N_3311,N_2668,N_2952);
nand U3312 (N_3312,N_2837,N_2772);
nand U3313 (N_3313,N_2781,N_2716);
and U3314 (N_3314,N_2414,N_2891);
nand U3315 (N_3315,N_2834,N_3094);
or U3316 (N_3316,N_2683,N_2884);
nor U3317 (N_3317,N_2853,N_2524);
nand U3318 (N_3318,N_2617,N_2998);
and U3319 (N_3319,N_2459,N_3114);
and U3320 (N_3320,N_2885,N_2959);
nor U3321 (N_3321,N_3070,N_2776);
nand U3322 (N_3322,N_3014,N_2931);
or U3323 (N_3323,N_2960,N_2559);
and U3324 (N_3324,N_2437,N_2682);
nand U3325 (N_3325,N_2544,N_2702);
nor U3326 (N_3326,N_3049,N_2615);
nand U3327 (N_3327,N_3019,N_2485);
nor U3328 (N_3328,N_3082,N_2818);
or U3329 (N_3329,N_3037,N_2852);
nand U3330 (N_3330,N_2742,N_3145);
and U3331 (N_3331,N_2919,N_2964);
and U3332 (N_3332,N_3138,N_2723);
nor U3333 (N_3333,N_2839,N_2895);
nand U3334 (N_3334,N_2491,N_2431);
xnor U3335 (N_3335,N_2789,N_3144);
or U3336 (N_3336,N_2562,N_2948);
or U3337 (N_3337,N_2947,N_2495);
xor U3338 (N_3338,N_3118,N_3081);
nor U3339 (N_3339,N_2578,N_3099);
nand U3340 (N_3340,N_2506,N_3029);
nor U3341 (N_3341,N_2983,N_2847);
nand U3342 (N_3342,N_2405,N_3063);
xnor U3343 (N_3343,N_2576,N_2503);
and U3344 (N_3344,N_2900,N_2995);
and U3345 (N_3345,N_3073,N_2710);
and U3346 (N_3346,N_3164,N_3170);
or U3347 (N_3347,N_2783,N_2869);
or U3348 (N_3348,N_2996,N_2868);
nand U3349 (N_3349,N_2416,N_2666);
nor U3350 (N_3350,N_2594,N_2669);
or U3351 (N_3351,N_2912,N_2607);
or U3352 (N_3352,N_2511,N_2611);
xor U3353 (N_3353,N_2926,N_2812);
nand U3354 (N_3354,N_2427,N_2814);
or U3355 (N_3355,N_2592,N_2734);
and U3356 (N_3356,N_2466,N_2631);
nand U3357 (N_3357,N_2974,N_3076);
nand U3358 (N_3358,N_2628,N_2725);
or U3359 (N_3359,N_3188,N_2586);
xnor U3360 (N_3360,N_2523,N_2600);
or U3361 (N_3361,N_2472,N_2937);
nand U3362 (N_3362,N_2478,N_2620);
or U3363 (N_3363,N_2568,N_2946);
nand U3364 (N_3364,N_3143,N_2532);
xor U3365 (N_3365,N_2514,N_3111);
or U3366 (N_3366,N_2823,N_3115);
xor U3367 (N_3367,N_2537,N_3190);
nand U3368 (N_3368,N_2759,N_2921);
nand U3369 (N_3369,N_3007,N_3067);
nand U3370 (N_3370,N_3127,N_2833);
and U3371 (N_3371,N_2862,N_2890);
or U3372 (N_3372,N_2583,N_3169);
nand U3373 (N_3373,N_2500,N_2909);
nor U3374 (N_3374,N_2882,N_2780);
nor U3375 (N_3375,N_2761,N_2821);
and U3376 (N_3376,N_3154,N_2521);
nor U3377 (N_3377,N_3080,N_2477);
nand U3378 (N_3378,N_2630,N_2651);
nor U3379 (N_3379,N_2779,N_2704);
nor U3380 (N_3380,N_2739,N_2898);
and U3381 (N_3381,N_3171,N_2528);
nand U3382 (N_3382,N_2410,N_2977);
and U3383 (N_3383,N_3100,N_2889);
nor U3384 (N_3384,N_2970,N_3027);
nand U3385 (N_3385,N_2722,N_2820);
or U3386 (N_3386,N_2667,N_2681);
and U3387 (N_3387,N_2442,N_3120);
nand U3388 (N_3388,N_2954,N_2700);
or U3389 (N_3389,N_2870,N_3033);
nor U3390 (N_3390,N_2606,N_2618);
or U3391 (N_3391,N_3006,N_2817);
nand U3392 (N_3392,N_2768,N_2629);
nor U3393 (N_3393,N_3195,N_2486);
xnor U3394 (N_3394,N_3090,N_2447);
or U3395 (N_3395,N_2658,N_2979);
and U3396 (N_3396,N_3153,N_2573);
nor U3397 (N_3397,N_2625,N_2556);
xor U3398 (N_3398,N_2412,N_3178);
nand U3399 (N_3399,N_2801,N_2450);
or U3400 (N_3400,N_3117,N_3022);
xnor U3401 (N_3401,N_3043,N_2957);
xnor U3402 (N_3402,N_2819,N_2811);
or U3403 (N_3403,N_3192,N_2555);
or U3404 (N_3404,N_2451,N_2563);
nor U3405 (N_3405,N_2545,N_2421);
nand U3406 (N_3406,N_2708,N_2452);
and U3407 (N_3407,N_2930,N_2458);
or U3408 (N_3408,N_2910,N_3010);
nor U3409 (N_3409,N_2550,N_3193);
and U3410 (N_3410,N_3097,N_3139);
nand U3411 (N_3411,N_3054,N_2626);
nor U3412 (N_3412,N_2637,N_2803);
and U3413 (N_3413,N_3194,N_2699);
and U3414 (N_3414,N_3051,N_3121);
and U3415 (N_3415,N_2720,N_2866);
or U3416 (N_3416,N_2567,N_2692);
nand U3417 (N_3417,N_2798,N_3134);
nor U3418 (N_3418,N_2696,N_2792);
or U3419 (N_3419,N_2496,N_2831);
and U3420 (N_3420,N_2913,N_2764);
nand U3421 (N_3421,N_2440,N_2731);
xnor U3422 (N_3422,N_2893,N_2706);
xnor U3423 (N_3423,N_2806,N_3113);
nand U3424 (N_3424,N_2529,N_2724);
nor U3425 (N_3425,N_2940,N_2969);
nor U3426 (N_3426,N_2762,N_2835);
and U3427 (N_3427,N_2883,N_2420);
and U3428 (N_3428,N_3179,N_2624);
or U3429 (N_3429,N_2616,N_2657);
nor U3430 (N_3430,N_2455,N_2797);
nand U3431 (N_3431,N_2749,N_2400);
nand U3432 (N_3432,N_2986,N_3092);
nand U3433 (N_3433,N_3198,N_3189);
and U3434 (N_3434,N_2596,N_3034);
nand U3435 (N_3435,N_3199,N_2517);
nor U3436 (N_3436,N_3021,N_2679);
nand U3437 (N_3437,N_2747,N_2471);
and U3438 (N_3438,N_3124,N_2697);
and U3439 (N_3439,N_2793,N_2791);
nor U3440 (N_3440,N_3023,N_2428);
nor U3441 (N_3441,N_2956,N_3146);
and U3442 (N_3442,N_2609,N_2784);
xor U3443 (N_3443,N_2424,N_2460);
nand U3444 (N_3444,N_2579,N_2619);
nor U3445 (N_3445,N_2843,N_2881);
nand U3446 (N_3446,N_2675,N_2988);
and U3447 (N_3447,N_2467,N_2530);
nand U3448 (N_3448,N_3119,N_2674);
nand U3449 (N_3449,N_3003,N_2480);
or U3450 (N_3450,N_2680,N_2856);
or U3451 (N_3451,N_2676,N_2445);
and U3452 (N_3452,N_2850,N_3060);
or U3453 (N_3453,N_3026,N_2771);
nor U3454 (N_3454,N_3161,N_2978);
xnor U3455 (N_3455,N_2577,N_3089);
xnor U3456 (N_3456,N_2465,N_3133);
nand U3457 (N_3457,N_2639,N_2531);
and U3458 (N_3458,N_2915,N_2552);
and U3459 (N_3459,N_2795,N_2786);
nand U3460 (N_3460,N_3095,N_2920);
nand U3461 (N_3461,N_2643,N_3103);
nand U3462 (N_3462,N_2987,N_2804);
and U3463 (N_3463,N_2929,N_2448);
nand U3464 (N_3464,N_2663,N_3128);
nor U3465 (N_3465,N_2748,N_3175);
xor U3466 (N_3466,N_2800,N_2838);
nand U3467 (N_3467,N_2548,N_2753);
xor U3468 (N_3468,N_2836,N_2419);
nor U3469 (N_3469,N_3098,N_2518);
or U3470 (N_3470,N_2415,N_2906);
nor U3471 (N_3471,N_3083,N_2640);
xor U3472 (N_3472,N_2941,N_2635);
nor U3473 (N_3473,N_2794,N_2928);
or U3474 (N_3474,N_2671,N_3183);
xor U3475 (N_3475,N_2587,N_2621);
or U3476 (N_3476,N_3130,N_3042);
xnor U3477 (N_3477,N_2554,N_3053);
nor U3478 (N_3478,N_2901,N_3187);
nand U3479 (N_3479,N_3064,N_2788);
nor U3480 (N_3480,N_2871,N_2489);
xnor U3481 (N_3481,N_2464,N_2645);
and U3482 (N_3482,N_2765,N_2907);
or U3483 (N_3483,N_3140,N_2542);
nor U3484 (N_3484,N_2968,N_2790);
nor U3485 (N_3485,N_2481,N_2861);
xnor U3486 (N_3486,N_3001,N_2867);
nor U3487 (N_3487,N_2949,N_2469);
xor U3488 (N_3488,N_2534,N_2815);
nor U3489 (N_3489,N_2436,N_2527);
xnor U3490 (N_3490,N_2770,N_2608);
and U3491 (N_3491,N_3147,N_2653);
nor U3492 (N_3492,N_2601,N_2971);
or U3493 (N_3493,N_2558,N_2976);
nand U3494 (N_3494,N_3184,N_3181);
and U3495 (N_3495,N_3102,N_2828);
xor U3496 (N_3496,N_2557,N_2551);
xnor U3497 (N_3497,N_2418,N_3050);
or U3498 (N_3498,N_2769,N_2752);
xnor U3499 (N_3499,N_2402,N_2444);
and U3500 (N_3500,N_2886,N_2430);
nor U3501 (N_3501,N_2634,N_2504);
xnor U3502 (N_3502,N_2860,N_2406);
nor U3503 (N_3503,N_2864,N_3166);
or U3504 (N_3504,N_2766,N_2598);
xor U3505 (N_3505,N_2687,N_2488);
xnor U3506 (N_3506,N_2888,N_2865);
nand U3507 (N_3507,N_2961,N_2435);
xnor U3508 (N_3508,N_2543,N_3009);
nand U3509 (N_3509,N_2923,N_2816);
xnor U3510 (N_3510,N_2644,N_2718);
nand U3511 (N_3511,N_3008,N_2662);
nor U3512 (N_3512,N_3106,N_2841);
and U3513 (N_3513,N_3186,N_2999);
xor U3514 (N_3514,N_3104,N_2569);
nand U3515 (N_3515,N_2649,N_2652);
nor U3516 (N_3516,N_2721,N_2535);
and U3517 (N_3517,N_2973,N_2605);
nand U3518 (N_3518,N_3018,N_2958);
and U3519 (N_3519,N_2911,N_3197);
nand U3520 (N_3520,N_3000,N_3036);
or U3521 (N_3521,N_2571,N_2874);
xor U3522 (N_3522,N_2648,N_2729);
xnor U3523 (N_3523,N_2966,N_3078);
nand U3524 (N_3524,N_2711,N_2851);
or U3525 (N_3525,N_2502,N_3176);
nor U3526 (N_3526,N_2844,N_3015);
and U3527 (N_3527,N_2636,N_3158);
nor U3528 (N_3528,N_3096,N_2810);
nand U3529 (N_3529,N_2482,N_3032);
xnor U3530 (N_3530,N_2673,N_3016);
xnor U3531 (N_3531,N_2787,N_3075);
xor U3532 (N_3532,N_2599,N_2401);
xor U3533 (N_3533,N_3110,N_2903);
and U3534 (N_3534,N_2832,N_3116);
nand U3535 (N_3535,N_2712,N_3165);
nand U3536 (N_3536,N_2944,N_2905);
xor U3537 (N_3537,N_3160,N_2684);
nor U3538 (N_3538,N_2942,N_2509);
or U3539 (N_3539,N_3131,N_2967);
nand U3540 (N_3540,N_2714,N_2441);
xnor U3541 (N_3541,N_2516,N_2664);
xor U3542 (N_3542,N_2701,N_2654);
or U3543 (N_3543,N_3162,N_2646);
nand U3544 (N_3544,N_2934,N_2656);
or U3545 (N_3545,N_2859,N_3077);
or U3546 (N_3546,N_2426,N_2593);
and U3547 (N_3547,N_2743,N_2849);
xnor U3548 (N_3548,N_3024,N_2953);
nor U3549 (N_3549,N_2735,N_3185);
or U3550 (N_3550,N_2908,N_2693);
nand U3551 (N_3551,N_2922,N_2826);
nand U3552 (N_3552,N_2773,N_2829);
or U3553 (N_3553,N_2939,N_3156);
nand U3554 (N_3554,N_3157,N_2522);
nor U3555 (N_3555,N_2540,N_2602);
nand U3556 (N_3556,N_2927,N_2848);
nor U3557 (N_3557,N_2473,N_2997);
and U3558 (N_3558,N_3066,N_2479);
and U3559 (N_3559,N_2892,N_2508);
nand U3560 (N_3560,N_2994,N_2914);
or U3561 (N_3561,N_2560,N_2744);
or U3562 (N_3562,N_2575,N_2432);
and U3563 (N_3563,N_2760,N_3168);
nand U3564 (N_3564,N_2984,N_2858);
nor U3565 (N_3565,N_3191,N_2992);
nor U3566 (N_3566,N_2449,N_2513);
nand U3567 (N_3567,N_2404,N_2603);
xnor U3568 (N_3568,N_2468,N_3020);
or U3569 (N_3569,N_2899,N_2538);
nor U3570 (N_3570,N_2622,N_2462);
xor U3571 (N_3571,N_2510,N_2612);
xor U3572 (N_3572,N_2474,N_3056);
nand U3573 (N_3573,N_3177,N_2842);
and U3574 (N_3574,N_2580,N_2993);
nor U3575 (N_3575,N_2805,N_2689);
nor U3576 (N_3576,N_3101,N_3013);
nand U3577 (N_3577,N_2561,N_2830);
xor U3578 (N_3578,N_2737,N_2935);
nor U3579 (N_3579,N_2507,N_2732);
and U3580 (N_3580,N_2655,N_2796);
and U3581 (N_3581,N_3174,N_2775);
xor U3582 (N_3582,N_2774,N_3057);
nand U3583 (N_3583,N_2975,N_2745);
xnor U3584 (N_3584,N_2647,N_2738);
xor U3585 (N_3585,N_3025,N_2990);
and U3586 (N_3586,N_2740,N_2691);
or U3587 (N_3587,N_3052,N_2512);
nor U3588 (N_3588,N_2526,N_2875);
xnor U3589 (N_3589,N_2925,N_2813);
nand U3590 (N_3590,N_2950,N_3135);
and U3591 (N_3591,N_2672,N_2665);
nand U3592 (N_3592,N_2446,N_2553);
and U3593 (N_3593,N_2454,N_2767);
and U3594 (N_3594,N_2582,N_2873);
and U3595 (N_3595,N_2863,N_2572);
nor U3596 (N_3596,N_3045,N_2755);
and U3597 (N_3597,N_3091,N_2746);
and U3598 (N_3598,N_3085,N_3150);
and U3599 (N_3599,N_2470,N_2641);
or U3600 (N_3600,N_2565,N_3158);
or U3601 (N_3601,N_3170,N_2809);
and U3602 (N_3602,N_2590,N_2870);
nand U3603 (N_3603,N_2749,N_2539);
or U3604 (N_3604,N_2541,N_2448);
or U3605 (N_3605,N_2674,N_2720);
nor U3606 (N_3606,N_2784,N_2693);
and U3607 (N_3607,N_3146,N_2694);
and U3608 (N_3608,N_2743,N_3147);
and U3609 (N_3609,N_2923,N_3000);
xnor U3610 (N_3610,N_3189,N_2636);
and U3611 (N_3611,N_3194,N_2895);
and U3612 (N_3612,N_2713,N_2692);
xor U3613 (N_3613,N_2968,N_2492);
xor U3614 (N_3614,N_2651,N_2501);
or U3615 (N_3615,N_2731,N_2694);
nor U3616 (N_3616,N_2874,N_3104);
xor U3617 (N_3617,N_2793,N_2403);
or U3618 (N_3618,N_2802,N_3136);
nor U3619 (N_3619,N_3056,N_2994);
and U3620 (N_3620,N_2498,N_2460);
and U3621 (N_3621,N_2737,N_2634);
nand U3622 (N_3622,N_3109,N_2888);
and U3623 (N_3623,N_2721,N_2716);
and U3624 (N_3624,N_2821,N_2922);
xnor U3625 (N_3625,N_2520,N_2411);
nand U3626 (N_3626,N_2728,N_2499);
and U3627 (N_3627,N_2548,N_2697);
or U3628 (N_3628,N_2715,N_2617);
nor U3629 (N_3629,N_2477,N_2480);
nor U3630 (N_3630,N_3014,N_2803);
or U3631 (N_3631,N_2925,N_2546);
and U3632 (N_3632,N_2987,N_2813);
or U3633 (N_3633,N_2478,N_3136);
or U3634 (N_3634,N_2544,N_2865);
nor U3635 (N_3635,N_2938,N_2982);
nand U3636 (N_3636,N_2816,N_2727);
nor U3637 (N_3637,N_3001,N_2483);
xor U3638 (N_3638,N_2703,N_2903);
nand U3639 (N_3639,N_3157,N_2621);
and U3640 (N_3640,N_3194,N_2420);
xnor U3641 (N_3641,N_2955,N_2646);
nor U3642 (N_3642,N_2889,N_3150);
xnor U3643 (N_3643,N_2952,N_3177);
nor U3644 (N_3644,N_2622,N_2620);
or U3645 (N_3645,N_3083,N_3185);
nor U3646 (N_3646,N_3115,N_3013);
nand U3647 (N_3647,N_2629,N_3064);
xor U3648 (N_3648,N_3102,N_2737);
nand U3649 (N_3649,N_3182,N_2892);
xnor U3650 (N_3650,N_2869,N_3101);
xor U3651 (N_3651,N_2961,N_2820);
nand U3652 (N_3652,N_2645,N_2791);
and U3653 (N_3653,N_2801,N_2505);
xnor U3654 (N_3654,N_2908,N_2885);
xor U3655 (N_3655,N_3127,N_2872);
or U3656 (N_3656,N_3107,N_3148);
xnor U3657 (N_3657,N_2429,N_2422);
or U3658 (N_3658,N_3163,N_2918);
nor U3659 (N_3659,N_2746,N_2655);
nor U3660 (N_3660,N_2430,N_3052);
xnor U3661 (N_3661,N_2698,N_2700);
xnor U3662 (N_3662,N_2729,N_2731);
xnor U3663 (N_3663,N_2559,N_3006);
and U3664 (N_3664,N_2958,N_2689);
nand U3665 (N_3665,N_2500,N_2533);
nor U3666 (N_3666,N_3002,N_2922);
and U3667 (N_3667,N_2693,N_2750);
xor U3668 (N_3668,N_2744,N_2561);
xnor U3669 (N_3669,N_2716,N_2950);
and U3670 (N_3670,N_2708,N_3074);
nand U3671 (N_3671,N_3118,N_2605);
and U3672 (N_3672,N_2876,N_3097);
and U3673 (N_3673,N_2913,N_2858);
xor U3674 (N_3674,N_2938,N_2451);
or U3675 (N_3675,N_2414,N_3164);
and U3676 (N_3676,N_2813,N_2404);
and U3677 (N_3677,N_2819,N_2991);
and U3678 (N_3678,N_2748,N_2761);
and U3679 (N_3679,N_3124,N_2440);
nor U3680 (N_3680,N_3102,N_3100);
xor U3681 (N_3681,N_2536,N_3156);
xnor U3682 (N_3682,N_2712,N_2785);
nand U3683 (N_3683,N_2852,N_2401);
nand U3684 (N_3684,N_3131,N_3163);
xor U3685 (N_3685,N_2694,N_2888);
nand U3686 (N_3686,N_2706,N_2862);
nand U3687 (N_3687,N_2531,N_2406);
nor U3688 (N_3688,N_3152,N_3040);
nor U3689 (N_3689,N_2410,N_3083);
and U3690 (N_3690,N_3098,N_3118);
and U3691 (N_3691,N_2960,N_2811);
nand U3692 (N_3692,N_2456,N_2821);
or U3693 (N_3693,N_2434,N_2476);
or U3694 (N_3694,N_3152,N_3132);
and U3695 (N_3695,N_2837,N_2848);
nand U3696 (N_3696,N_2823,N_2591);
or U3697 (N_3697,N_2685,N_3135);
or U3698 (N_3698,N_2668,N_3172);
nand U3699 (N_3699,N_3172,N_2539);
xor U3700 (N_3700,N_2652,N_3099);
and U3701 (N_3701,N_2951,N_3072);
nand U3702 (N_3702,N_2925,N_2467);
xor U3703 (N_3703,N_2762,N_3049);
nand U3704 (N_3704,N_2739,N_2948);
and U3705 (N_3705,N_3044,N_2942);
or U3706 (N_3706,N_2998,N_2646);
nand U3707 (N_3707,N_2407,N_2919);
or U3708 (N_3708,N_3073,N_3124);
or U3709 (N_3709,N_3192,N_3010);
xnor U3710 (N_3710,N_3183,N_2901);
or U3711 (N_3711,N_2877,N_2454);
or U3712 (N_3712,N_3021,N_3072);
nand U3713 (N_3713,N_2460,N_3008);
xnor U3714 (N_3714,N_2881,N_2604);
nor U3715 (N_3715,N_2612,N_2412);
nand U3716 (N_3716,N_3166,N_2918);
or U3717 (N_3717,N_2930,N_2688);
nand U3718 (N_3718,N_3113,N_2434);
or U3719 (N_3719,N_3199,N_2572);
nand U3720 (N_3720,N_2935,N_2497);
nand U3721 (N_3721,N_2864,N_3129);
nand U3722 (N_3722,N_2520,N_2847);
and U3723 (N_3723,N_2694,N_2947);
nor U3724 (N_3724,N_2717,N_3083);
xor U3725 (N_3725,N_2655,N_2584);
nor U3726 (N_3726,N_2531,N_2825);
and U3727 (N_3727,N_3114,N_2617);
xor U3728 (N_3728,N_2969,N_3193);
xor U3729 (N_3729,N_2762,N_3009);
or U3730 (N_3730,N_2490,N_3147);
nand U3731 (N_3731,N_3049,N_2711);
xnor U3732 (N_3732,N_2994,N_2606);
nand U3733 (N_3733,N_2460,N_2447);
and U3734 (N_3734,N_2604,N_2520);
or U3735 (N_3735,N_2513,N_2993);
nor U3736 (N_3736,N_2555,N_2937);
xnor U3737 (N_3737,N_3169,N_2771);
xnor U3738 (N_3738,N_2534,N_2743);
xnor U3739 (N_3739,N_3033,N_2901);
xor U3740 (N_3740,N_2457,N_3073);
and U3741 (N_3741,N_2622,N_3151);
and U3742 (N_3742,N_2493,N_2787);
xnor U3743 (N_3743,N_2913,N_3171);
or U3744 (N_3744,N_2844,N_2731);
and U3745 (N_3745,N_2793,N_3117);
and U3746 (N_3746,N_2675,N_3105);
nand U3747 (N_3747,N_2463,N_2935);
xnor U3748 (N_3748,N_2614,N_3000);
nor U3749 (N_3749,N_2641,N_2439);
or U3750 (N_3750,N_2538,N_2531);
and U3751 (N_3751,N_2676,N_2791);
xor U3752 (N_3752,N_2412,N_3110);
nor U3753 (N_3753,N_2835,N_2528);
nand U3754 (N_3754,N_2620,N_2433);
and U3755 (N_3755,N_2422,N_2995);
or U3756 (N_3756,N_2986,N_2690);
nor U3757 (N_3757,N_2677,N_2812);
xor U3758 (N_3758,N_2658,N_3096);
nor U3759 (N_3759,N_2958,N_2533);
nand U3760 (N_3760,N_3184,N_3032);
or U3761 (N_3761,N_2806,N_2684);
xor U3762 (N_3762,N_2518,N_3174);
nor U3763 (N_3763,N_2526,N_2432);
or U3764 (N_3764,N_2885,N_3148);
and U3765 (N_3765,N_2945,N_2516);
nand U3766 (N_3766,N_2411,N_2587);
nor U3767 (N_3767,N_2454,N_3157);
xnor U3768 (N_3768,N_2654,N_3184);
and U3769 (N_3769,N_2652,N_2735);
or U3770 (N_3770,N_2880,N_3051);
and U3771 (N_3771,N_2533,N_2438);
and U3772 (N_3772,N_2599,N_2823);
and U3773 (N_3773,N_2595,N_2597);
nand U3774 (N_3774,N_2514,N_3130);
xor U3775 (N_3775,N_3167,N_2948);
xnor U3776 (N_3776,N_2534,N_2443);
xnor U3777 (N_3777,N_2518,N_3129);
and U3778 (N_3778,N_3125,N_2781);
nand U3779 (N_3779,N_3029,N_3021);
nand U3780 (N_3780,N_2677,N_2665);
or U3781 (N_3781,N_2451,N_2507);
xor U3782 (N_3782,N_2677,N_3056);
or U3783 (N_3783,N_3107,N_2725);
or U3784 (N_3784,N_2848,N_3138);
and U3785 (N_3785,N_2978,N_3195);
or U3786 (N_3786,N_2513,N_2785);
or U3787 (N_3787,N_3078,N_3116);
xor U3788 (N_3788,N_3192,N_2400);
xor U3789 (N_3789,N_2562,N_2972);
or U3790 (N_3790,N_2947,N_3127);
xor U3791 (N_3791,N_2972,N_2677);
or U3792 (N_3792,N_3134,N_2679);
nand U3793 (N_3793,N_3049,N_3056);
xnor U3794 (N_3794,N_2406,N_2790);
xnor U3795 (N_3795,N_2452,N_2642);
nor U3796 (N_3796,N_3156,N_2550);
nor U3797 (N_3797,N_2541,N_2530);
nor U3798 (N_3798,N_3084,N_2667);
or U3799 (N_3799,N_2858,N_3119);
or U3800 (N_3800,N_2406,N_3158);
xnor U3801 (N_3801,N_2904,N_2684);
nor U3802 (N_3802,N_2987,N_2580);
nand U3803 (N_3803,N_3198,N_3150);
or U3804 (N_3804,N_2797,N_2742);
or U3805 (N_3805,N_2904,N_3195);
and U3806 (N_3806,N_2463,N_2551);
xnor U3807 (N_3807,N_2996,N_2974);
nand U3808 (N_3808,N_2910,N_3084);
nand U3809 (N_3809,N_2434,N_2537);
and U3810 (N_3810,N_3100,N_3189);
and U3811 (N_3811,N_3129,N_2996);
and U3812 (N_3812,N_3052,N_2445);
xnor U3813 (N_3813,N_2885,N_2714);
and U3814 (N_3814,N_2593,N_2548);
or U3815 (N_3815,N_2821,N_2628);
xnor U3816 (N_3816,N_2876,N_2861);
nand U3817 (N_3817,N_2742,N_2459);
nand U3818 (N_3818,N_3168,N_2744);
or U3819 (N_3819,N_3126,N_2792);
and U3820 (N_3820,N_2905,N_2577);
and U3821 (N_3821,N_2668,N_2473);
and U3822 (N_3822,N_2915,N_2425);
xnor U3823 (N_3823,N_2712,N_2814);
or U3824 (N_3824,N_2506,N_2841);
nor U3825 (N_3825,N_2565,N_2745);
nand U3826 (N_3826,N_2716,N_2786);
xnor U3827 (N_3827,N_3002,N_3063);
and U3828 (N_3828,N_2640,N_2886);
nor U3829 (N_3829,N_3120,N_2435);
xor U3830 (N_3830,N_3141,N_2444);
xnor U3831 (N_3831,N_2717,N_2605);
xnor U3832 (N_3832,N_3065,N_2934);
nand U3833 (N_3833,N_2666,N_3119);
or U3834 (N_3834,N_2610,N_2997);
nand U3835 (N_3835,N_2516,N_2599);
and U3836 (N_3836,N_3137,N_2961);
and U3837 (N_3837,N_2713,N_2940);
or U3838 (N_3838,N_2956,N_2909);
nand U3839 (N_3839,N_2735,N_2907);
and U3840 (N_3840,N_2465,N_2660);
and U3841 (N_3841,N_2638,N_3073);
xor U3842 (N_3842,N_2728,N_2447);
or U3843 (N_3843,N_2596,N_2576);
or U3844 (N_3844,N_2828,N_2994);
xnor U3845 (N_3845,N_3089,N_2966);
nor U3846 (N_3846,N_2777,N_2894);
nand U3847 (N_3847,N_2746,N_3128);
nor U3848 (N_3848,N_3195,N_2944);
and U3849 (N_3849,N_3039,N_2614);
xor U3850 (N_3850,N_2968,N_2963);
and U3851 (N_3851,N_2795,N_2567);
or U3852 (N_3852,N_3157,N_2681);
or U3853 (N_3853,N_2692,N_2849);
xnor U3854 (N_3854,N_3018,N_3171);
or U3855 (N_3855,N_2435,N_2858);
and U3856 (N_3856,N_2726,N_2674);
nor U3857 (N_3857,N_2728,N_2740);
xor U3858 (N_3858,N_2844,N_3145);
nor U3859 (N_3859,N_3181,N_2884);
nand U3860 (N_3860,N_2735,N_3195);
nor U3861 (N_3861,N_3196,N_3041);
or U3862 (N_3862,N_3139,N_2625);
nor U3863 (N_3863,N_2527,N_2720);
nor U3864 (N_3864,N_2688,N_2818);
nand U3865 (N_3865,N_2969,N_2948);
xor U3866 (N_3866,N_2808,N_2624);
xor U3867 (N_3867,N_2684,N_2697);
or U3868 (N_3868,N_2926,N_2736);
nor U3869 (N_3869,N_2513,N_2934);
nand U3870 (N_3870,N_2843,N_2811);
nand U3871 (N_3871,N_2908,N_2443);
xor U3872 (N_3872,N_2968,N_2704);
and U3873 (N_3873,N_2869,N_2419);
xnor U3874 (N_3874,N_2620,N_2470);
nand U3875 (N_3875,N_3013,N_2764);
or U3876 (N_3876,N_2870,N_2849);
xor U3877 (N_3877,N_3091,N_2834);
xor U3878 (N_3878,N_2585,N_2602);
nor U3879 (N_3879,N_3146,N_2605);
and U3880 (N_3880,N_2943,N_3122);
or U3881 (N_3881,N_3029,N_2487);
xnor U3882 (N_3882,N_3004,N_2489);
and U3883 (N_3883,N_2699,N_2933);
and U3884 (N_3884,N_2938,N_2704);
nor U3885 (N_3885,N_3087,N_2695);
xnor U3886 (N_3886,N_3042,N_2977);
or U3887 (N_3887,N_2551,N_2658);
and U3888 (N_3888,N_3148,N_2851);
or U3889 (N_3889,N_2814,N_2893);
and U3890 (N_3890,N_2994,N_2957);
xor U3891 (N_3891,N_2510,N_3044);
and U3892 (N_3892,N_2557,N_2509);
and U3893 (N_3893,N_2884,N_3075);
nand U3894 (N_3894,N_2868,N_3162);
xor U3895 (N_3895,N_2935,N_3054);
or U3896 (N_3896,N_2495,N_3167);
nor U3897 (N_3897,N_2624,N_2796);
nand U3898 (N_3898,N_3001,N_2498);
or U3899 (N_3899,N_3178,N_2687);
or U3900 (N_3900,N_2601,N_2542);
nand U3901 (N_3901,N_2580,N_2508);
or U3902 (N_3902,N_2602,N_3096);
nor U3903 (N_3903,N_2717,N_3003);
nor U3904 (N_3904,N_3105,N_2860);
nand U3905 (N_3905,N_2463,N_2977);
or U3906 (N_3906,N_2984,N_2797);
and U3907 (N_3907,N_2492,N_2635);
and U3908 (N_3908,N_2590,N_2400);
xnor U3909 (N_3909,N_3172,N_2533);
and U3910 (N_3910,N_2547,N_3097);
xnor U3911 (N_3911,N_2755,N_2935);
xnor U3912 (N_3912,N_2576,N_2654);
nor U3913 (N_3913,N_2778,N_2571);
nor U3914 (N_3914,N_2404,N_2964);
or U3915 (N_3915,N_2871,N_2484);
xor U3916 (N_3916,N_3196,N_2529);
nor U3917 (N_3917,N_2644,N_3055);
nor U3918 (N_3918,N_2711,N_3136);
xnor U3919 (N_3919,N_2849,N_2948);
nor U3920 (N_3920,N_2400,N_2821);
or U3921 (N_3921,N_2998,N_2830);
xor U3922 (N_3922,N_3065,N_2899);
nor U3923 (N_3923,N_3167,N_2980);
nand U3924 (N_3924,N_2528,N_3062);
or U3925 (N_3925,N_2861,N_2746);
nor U3926 (N_3926,N_3190,N_2834);
and U3927 (N_3927,N_2687,N_2691);
xor U3928 (N_3928,N_2503,N_2746);
nand U3929 (N_3929,N_2542,N_3067);
nand U3930 (N_3930,N_3109,N_2860);
nor U3931 (N_3931,N_3157,N_3021);
nor U3932 (N_3932,N_2489,N_2940);
or U3933 (N_3933,N_2434,N_3103);
nand U3934 (N_3934,N_2515,N_2459);
xnor U3935 (N_3935,N_2929,N_2978);
xnor U3936 (N_3936,N_2998,N_2459);
xnor U3937 (N_3937,N_2755,N_3165);
and U3938 (N_3938,N_2938,N_2657);
or U3939 (N_3939,N_2791,N_2951);
xor U3940 (N_3940,N_3165,N_2828);
xor U3941 (N_3941,N_2921,N_2419);
or U3942 (N_3942,N_3134,N_2817);
nand U3943 (N_3943,N_2765,N_2501);
nand U3944 (N_3944,N_2599,N_2781);
nand U3945 (N_3945,N_2529,N_3064);
or U3946 (N_3946,N_2544,N_3091);
nor U3947 (N_3947,N_2479,N_2998);
nand U3948 (N_3948,N_3170,N_2859);
nor U3949 (N_3949,N_2408,N_3142);
or U3950 (N_3950,N_3010,N_2560);
or U3951 (N_3951,N_2411,N_2861);
and U3952 (N_3952,N_2603,N_3184);
nand U3953 (N_3953,N_3147,N_2662);
and U3954 (N_3954,N_2749,N_2894);
or U3955 (N_3955,N_3177,N_2534);
nor U3956 (N_3956,N_2440,N_2910);
and U3957 (N_3957,N_3063,N_2952);
xnor U3958 (N_3958,N_2833,N_2563);
and U3959 (N_3959,N_2834,N_2795);
and U3960 (N_3960,N_2457,N_3099);
xor U3961 (N_3961,N_2903,N_2559);
or U3962 (N_3962,N_2679,N_2651);
or U3963 (N_3963,N_2640,N_2496);
and U3964 (N_3964,N_2450,N_2864);
and U3965 (N_3965,N_2615,N_3056);
nand U3966 (N_3966,N_2908,N_2407);
nor U3967 (N_3967,N_2656,N_2548);
and U3968 (N_3968,N_2711,N_3056);
xor U3969 (N_3969,N_3168,N_2971);
nor U3970 (N_3970,N_2901,N_3073);
nor U3971 (N_3971,N_3051,N_3013);
and U3972 (N_3972,N_2536,N_2816);
and U3973 (N_3973,N_3106,N_2875);
nor U3974 (N_3974,N_2980,N_2590);
nor U3975 (N_3975,N_2800,N_2745);
nand U3976 (N_3976,N_2945,N_2828);
xor U3977 (N_3977,N_2932,N_2801);
nand U3978 (N_3978,N_2651,N_2949);
or U3979 (N_3979,N_3030,N_3038);
nor U3980 (N_3980,N_3143,N_3189);
or U3981 (N_3981,N_2750,N_2773);
nand U3982 (N_3982,N_3172,N_2477);
and U3983 (N_3983,N_3045,N_3059);
nor U3984 (N_3984,N_2406,N_2775);
xnor U3985 (N_3985,N_2469,N_2525);
nor U3986 (N_3986,N_2899,N_2876);
xnor U3987 (N_3987,N_2715,N_3014);
or U3988 (N_3988,N_3079,N_2756);
nor U3989 (N_3989,N_2815,N_3095);
nand U3990 (N_3990,N_2489,N_2511);
xor U3991 (N_3991,N_3010,N_2476);
nor U3992 (N_3992,N_2568,N_3040);
nand U3993 (N_3993,N_2900,N_3144);
nand U3994 (N_3994,N_2866,N_2871);
nand U3995 (N_3995,N_2897,N_2504);
or U3996 (N_3996,N_3091,N_2483);
or U3997 (N_3997,N_2539,N_3082);
nand U3998 (N_3998,N_2674,N_2978);
nor U3999 (N_3999,N_3018,N_2661);
nor U4000 (N_4000,N_3424,N_3860);
nor U4001 (N_4001,N_3605,N_3897);
or U4002 (N_4002,N_3712,N_3554);
nand U4003 (N_4003,N_3524,N_3368);
nor U4004 (N_4004,N_3737,N_3866);
xor U4005 (N_4005,N_3539,N_3233);
xnor U4006 (N_4006,N_3365,N_3544);
nand U4007 (N_4007,N_3586,N_3883);
nor U4008 (N_4008,N_3732,N_3326);
xnor U4009 (N_4009,N_3954,N_3612);
or U4010 (N_4010,N_3742,N_3655);
nand U4011 (N_4011,N_3611,N_3670);
and U4012 (N_4012,N_3689,N_3425);
or U4013 (N_4013,N_3476,N_3826);
xnor U4014 (N_4014,N_3767,N_3523);
nor U4015 (N_4015,N_3288,N_3933);
and U4016 (N_4016,N_3473,N_3458);
xnor U4017 (N_4017,N_3775,N_3362);
xor U4018 (N_4018,N_3211,N_3527);
xnor U4019 (N_4019,N_3867,N_3769);
nand U4020 (N_4020,N_3295,N_3234);
nand U4021 (N_4021,N_3841,N_3237);
and U4022 (N_4022,N_3747,N_3340);
nor U4023 (N_4023,N_3555,N_3394);
nand U4024 (N_4024,N_3799,N_3694);
nand U4025 (N_4025,N_3418,N_3270);
nor U4026 (N_4026,N_3377,N_3840);
and U4027 (N_4027,N_3433,N_3502);
nand U4028 (N_4028,N_3462,N_3629);
or U4029 (N_4029,N_3852,N_3479);
nand U4030 (N_4030,N_3946,N_3552);
xor U4031 (N_4031,N_3949,N_3361);
nand U4032 (N_4032,N_3207,N_3532);
nor U4033 (N_4033,N_3378,N_3600);
nand U4034 (N_4034,N_3596,N_3864);
and U4035 (N_4035,N_3692,N_3617);
and U4036 (N_4036,N_3940,N_3318);
nor U4037 (N_4037,N_3610,N_3878);
or U4038 (N_4038,N_3263,N_3344);
and U4039 (N_4039,N_3561,N_3950);
nor U4040 (N_4040,N_3483,N_3576);
nand U4041 (N_4041,N_3464,N_3879);
or U4042 (N_4042,N_3325,N_3314);
nor U4043 (N_4043,N_3333,N_3967);
xnor U4044 (N_4044,N_3204,N_3328);
nor U4045 (N_4045,N_3764,N_3277);
or U4046 (N_4046,N_3456,N_3603);
xnor U4047 (N_4047,N_3740,N_3397);
nand U4048 (N_4048,N_3391,N_3278);
nand U4049 (N_4049,N_3616,N_3281);
or U4050 (N_4050,N_3531,N_3514);
and U4051 (N_4051,N_3836,N_3206);
and U4052 (N_4052,N_3491,N_3307);
or U4053 (N_4053,N_3265,N_3851);
nand U4054 (N_4054,N_3711,N_3256);
xor U4055 (N_4055,N_3327,N_3918);
nor U4056 (N_4056,N_3224,N_3598);
nand U4057 (N_4057,N_3208,N_3247);
xor U4058 (N_4058,N_3677,N_3948);
nand U4059 (N_4059,N_3201,N_3899);
and U4060 (N_4060,N_3488,N_3832);
nand U4061 (N_4061,N_3592,N_3734);
nand U4062 (N_4062,N_3392,N_3444);
nand U4063 (N_4063,N_3792,N_3421);
or U4064 (N_4064,N_3765,N_3871);
xnor U4065 (N_4065,N_3855,N_3470);
or U4066 (N_4066,N_3405,N_3731);
or U4067 (N_4067,N_3409,N_3713);
or U4068 (N_4068,N_3917,N_3602);
xor U4069 (N_4069,N_3570,N_3778);
and U4070 (N_4070,N_3986,N_3889);
nand U4071 (N_4071,N_3516,N_3809);
or U4072 (N_4072,N_3654,N_3931);
or U4073 (N_4073,N_3750,N_3787);
nor U4074 (N_4074,N_3912,N_3309);
or U4075 (N_4075,N_3720,N_3929);
nand U4076 (N_4076,N_3494,N_3388);
xor U4077 (N_4077,N_3960,N_3335);
xor U4078 (N_4078,N_3412,N_3703);
or U4079 (N_4079,N_3426,N_3639);
nor U4080 (N_4080,N_3536,N_3565);
or U4081 (N_4081,N_3226,N_3965);
xor U4082 (N_4082,N_3302,N_3942);
and U4083 (N_4083,N_3839,N_3818);
and U4084 (N_4084,N_3419,N_3666);
or U4085 (N_4085,N_3297,N_3952);
nand U4086 (N_4086,N_3481,N_3478);
and U4087 (N_4087,N_3266,N_3865);
nand U4088 (N_4088,N_3648,N_3888);
or U4089 (N_4089,N_3892,N_3947);
or U4090 (N_4090,N_3254,N_3550);
or U4091 (N_4091,N_3622,N_3595);
nand U4092 (N_4092,N_3390,N_3752);
nor U4093 (N_4093,N_3304,N_3557);
nand U4094 (N_4094,N_3930,N_3306);
xor U4095 (N_4095,N_3364,N_3250);
nand U4096 (N_4096,N_3275,N_3467);
or U4097 (N_4097,N_3671,N_3604);
or U4098 (N_4098,N_3759,N_3649);
nand U4099 (N_4099,N_3794,N_3238);
xor U4100 (N_4100,N_3875,N_3715);
nor U4101 (N_4101,N_3439,N_3820);
xor U4102 (N_4102,N_3902,N_3756);
nand U4103 (N_4103,N_3880,N_3553);
xnor U4104 (N_4104,N_3398,N_3493);
nor U4105 (N_4105,N_3385,N_3606);
and U4106 (N_4106,N_3722,N_3487);
and U4107 (N_4107,N_3838,N_3913);
nand U4108 (N_4108,N_3690,N_3548);
or U4109 (N_4109,N_3264,N_3406);
or U4110 (N_4110,N_3995,N_3520);
nand U4111 (N_4111,N_3200,N_3342);
nor U4112 (N_4112,N_3890,N_3618);
nor U4113 (N_4113,N_3212,N_3543);
nor U4114 (N_4114,N_3781,N_3466);
xor U4115 (N_4115,N_3279,N_3345);
or U4116 (N_4116,N_3957,N_3922);
nor U4117 (N_4117,N_3643,N_3533);
nor U4118 (N_4118,N_3475,N_3435);
nand U4119 (N_4119,N_3894,N_3222);
or U4120 (N_4120,N_3810,N_3668);
and U4121 (N_4121,N_3245,N_3859);
nand U4122 (N_4122,N_3932,N_3242);
nand U4123 (N_4123,N_3373,N_3773);
and U4124 (N_4124,N_3492,N_3216);
xnor U4125 (N_4125,N_3805,N_3384);
and U4126 (N_4126,N_3296,N_3691);
xor U4127 (N_4127,N_3978,N_3664);
nor U4128 (N_4128,N_3817,N_3945);
and U4129 (N_4129,N_3909,N_3763);
nand U4130 (N_4130,N_3785,N_3627);
or U4131 (N_4131,N_3780,N_3762);
nand U4132 (N_4132,N_3442,N_3443);
nand U4133 (N_4133,N_3468,N_3573);
or U4134 (N_4134,N_3685,N_3834);
nand U4135 (N_4135,N_3506,N_3789);
or U4136 (N_4136,N_3441,N_3635);
nor U4137 (N_4137,N_3301,N_3438);
nor U4138 (N_4138,N_3798,N_3407);
nand U4139 (N_4139,N_3546,N_3459);
or U4140 (N_4140,N_3535,N_3983);
nor U4141 (N_4141,N_3374,N_3669);
xnor U4142 (N_4142,N_3626,N_3322);
nor U4143 (N_4143,N_3590,N_3228);
xnor U4144 (N_4144,N_3526,N_3854);
nand U4145 (N_4145,N_3915,N_3601);
and U4146 (N_4146,N_3900,N_3768);
xnor U4147 (N_4147,N_3971,N_3310);
nor U4148 (N_4148,N_3678,N_3387);
nand U4149 (N_4149,N_3447,N_3958);
xnor U4150 (N_4150,N_3341,N_3988);
nor U4151 (N_4151,N_3848,N_3802);
nor U4152 (N_4152,N_3574,N_3292);
nor U4153 (N_4153,N_3943,N_3628);
or U4154 (N_4154,N_3260,N_3910);
nand U4155 (N_4155,N_3287,N_3736);
or U4156 (N_4156,N_3962,N_3972);
or U4157 (N_4157,N_3579,N_3556);
and U4158 (N_4158,N_3513,N_3793);
xor U4159 (N_4159,N_3350,N_3973);
nor U4160 (N_4160,N_3294,N_3355);
xnor U4161 (N_4161,N_3837,N_3801);
nand U4162 (N_4162,N_3684,N_3563);
or U4163 (N_4163,N_3496,N_3675);
and U4164 (N_4164,N_3934,N_3709);
or U4165 (N_4165,N_3956,N_3223);
nor U4166 (N_4166,N_3624,N_3511);
nand U4167 (N_4167,N_3991,N_3744);
xnor U4168 (N_4168,N_3504,N_3395);
and U4169 (N_4169,N_3446,N_3411);
and U4170 (N_4170,N_3477,N_3501);
or U4171 (N_4171,N_3808,N_3313);
and U4172 (N_4172,N_3597,N_3886);
and U4173 (N_4173,N_3323,N_3651);
nand U4174 (N_4174,N_3990,N_3830);
nand U4175 (N_4175,N_3937,N_3680);
nand U4176 (N_4176,N_3319,N_3779);
or U4177 (N_4177,N_3724,N_3241);
nor U4178 (N_4178,N_3755,N_3873);
xor U4179 (N_4179,N_3891,N_3833);
nand U4180 (N_4180,N_3239,N_3308);
nor U4181 (N_4181,N_3803,N_3964);
and U4182 (N_4182,N_3252,N_3620);
nor U4183 (N_4183,N_3230,N_3257);
and U4184 (N_4184,N_3415,N_3243);
xnor U4185 (N_4185,N_3303,N_3876);
and U4186 (N_4186,N_3217,N_3510);
and U4187 (N_4187,N_3427,N_3339);
xor U4188 (N_4188,N_3450,N_3369);
or U4189 (N_4189,N_3813,N_3656);
and U4190 (N_4190,N_3632,N_3227);
and U4191 (N_4191,N_3614,N_3681);
or U4192 (N_4192,N_3845,N_3367);
nor U4193 (N_4193,N_3653,N_3745);
nand U4194 (N_4194,N_3522,N_3273);
nor U4195 (N_4195,N_3753,N_3400);
nor U4196 (N_4196,N_3708,N_3885);
or U4197 (N_4197,N_3797,N_3268);
nor U4198 (N_4198,N_3977,N_3647);
and U4199 (N_4199,N_3992,N_3594);
nand U4200 (N_4200,N_3231,N_3500);
nor U4201 (N_4201,N_3938,N_3356);
nor U4202 (N_4202,N_3203,N_3568);
nand U4203 (N_4203,N_3420,N_3336);
nand U4204 (N_4204,N_3824,N_3630);
nor U4205 (N_4205,N_3976,N_3727);
nand U4206 (N_4206,N_3939,N_3508);
and U4207 (N_4207,N_3469,N_3788);
nand U4208 (N_4208,N_3645,N_3719);
or U4209 (N_4209,N_3996,N_3541);
nor U4210 (N_4210,N_3843,N_3461);
nor U4211 (N_4211,N_3695,N_3825);
nand U4212 (N_4212,N_3582,N_3782);
xor U4213 (N_4213,N_3619,N_3225);
xnor U4214 (N_4214,N_3329,N_3396);
or U4215 (N_4215,N_3291,N_3253);
and U4216 (N_4216,N_3375,N_3754);
nand U4217 (N_4217,N_3766,N_3725);
xnor U4218 (N_4218,N_3663,N_3299);
nand U4219 (N_4219,N_3961,N_3363);
or U4220 (N_4220,N_3650,N_3507);
xor U4221 (N_4221,N_3261,N_3757);
or U4222 (N_4222,N_3434,N_3906);
xnor U4223 (N_4223,N_3525,N_3585);
xor U4224 (N_4224,N_3581,N_3777);
nand U4225 (N_4225,N_3298,N_3244);
xor U4226 (N_4226,N_3998,N_3312);
nand U4227 (N_4227,N_3578,N_3638);
or U4228 (N_4228,N_3800,N_3572);
xor U4229 (N_4229,N_3821,N_3783);
xnor U4230 (N_4230,N_3259,N_3517);
nand U4231 (N_4231,N_3503,N_3267);
xor U4232 (N_4232,N_3884,N_3700);
nand U4233 (N_4233,N_3665,N_3343);
or U4234 (N_4234,N_3714,N_3537);
or U4235 (N_4235,N_3348,N_3636);
nor U4236 (N_4236,N_3562,N_3621);
nand U4237 (N_4237,N_3484,N_3402);
nor U4238 (N_4238,N_3399,N_3431);
and U4239 (N_4239,N_3428,N_3529);
xor U4240 (N_4240,N_3905,N_3571);
xnor U4241 (N_4241,N_3593,N_3401);
nand U4242 (N_4242,N_3729,N_3540);
nor U4243 (N_4243,N_3354,N_3631);
and U4244 (N_4244,N_3916,N_3380);
xor U4245 (N_4245,N_3701,N_3331);
nor U4246 (N_4246,N_3213,N_3853);
nor U4247 (N_4247,N_3869,N_3403);
nand U4248 (N_4248,N_3262,N_3480);
nor U4249 (N_4249,N_3330,N_3534);
nor U4250 (N_4250,N_3451,N_3271);
or U4251 (N_4251,N_3874,N_3795);
nand U4252 (N_4252,N_3219,N_3786);
or U4253 (N_4253,N_3707,N_3515);
xor U4254 (N_4254,N_3816,N_3413);
nor U4255 (N_4255,N_3454,N_3505);
or U4256 (N_4256,N_3584,N_3726);
xnor U4257 (N_4257,N_3613,N_3587);
nand U4258 (N_4258,N_3749,N_3386);
nand U4259 (N_4259,N_3856,N_3702);
xor U4260 (N_4260,N_3575,N_3209);
xor U4261 (N_4261,N_3283,N_3963);
or U4262 (N_4262,N_3662,N_3347);
or U4263 (N_4263,N_3993,N_3471);
nand U4264 (N_4264,N_3658,N_3615);
nor U4265 (N_4265,N_3417,N_3733);
or U4266 (N_4266,N_3440,N_3682);
and U4267 (N_4267,N_3673,N_3743);
nor U4268 (N_4268,N_3410,N_3349);
nor U4269 (N_4269,N_3735,N_3460);
xor U4270 (N_4270,N_3293,N_3968);
nand U4271 (N_4271,N_3981,N_3436);
nor U4272 (N_4272,N_3887,N_3474);
nor U4273 (N_4273,N_3358,N_3966);
nor U4274 (N_4274,N_3920,N_3704);
or U4275 (N_4275,N_3280,N_3844);
xor U4276 (N_4276,N_3337,N_3284);
xnor U4277 (N_4277,N_3577,N_3862);
and U4278 (N_4278,N_3521,N_3989);
and U4279 (N_4279,N_3235,N_3672);
and U4280 (N_4280,N_3804,N_3738);
xnor U4281 (N_4281,N_3904,N_3907);
or U4282 (N_4282,N_3580,N_3652);
xor U4283 (N_4283,N_3360,N_3538);
and U4284 (N_4284,N_3850,N_3936);
xor U4285 (N_4285,N_3895,N_3591);
nor U4286 (N_4286,N_3218,N_3370);
xor U4287 (N_4287,N_3376,N_3482);
nand U4288 (N_4288,N_3898,N_3741);
or U4289 (N_4289,N_3697,N_3559);
nand U4290 (N_4290,N_3637,N_3642);
or U4291 (N_4291,N_3389,N_3646);
or U4292 (N_4292,N_3255,N_3249);
xnor U4293 (N_4293,N_3659,N_3351);
and U4294 (N_4294,N_3974,N_3286);
and U4295 (N_4295,N_3760,N_3717);
or U4296 (N_4296,N_3776,N_3588);
and U4297 (N_4297,N_3289,N_3497);
and U4298 (N_4298,N_3359,N_3999);
nor U4299 (N_4299,N_3274,N_3625);
xor U4300 (N_4300,N_3774,N_3269);
xnor U4301 (N_4301,N_3758,N_3698);
and U4302 (N_4302,N_3790,N_3202);
xor U4303 (N_4303,N_3896,N_3317);
xor U4304 (N_4304,N_3432,N_3366);
and U4305 (N_4305,N_3644,N_3589);
xor U4306 (N_4306,N_3706,N_3485);
and U4307 (N_4307,N_3723,N_3877);
xnor U4308 (N_4308,N_3872,N_3449);
and U4309 (N_4309,N_3382,N_3679);
or U4310 (N_4310,N_3908,N_3236);
nor U4311 (N_4311,N_3205,N_3893);
nor U4312 (N_4312,N_3985,N_3282);
or U4313 (N_4313,N_3829,N_3495);
xor U4314 (N_4314,N_3530,N_3842);
xor U4315 (N_4315,N_3953,N_3372);
nor U4316 (N_4316,N_3453,N_3560);
xor U4317 (N_4317,N_3490,N_3549);
nand U4318 (N_4318,N_3919,N_3519);
or U4319 (N_4319,N_3583,N_3499);
nand U4320 (N_4320,N_3660,N_3465);
and U4321 (N_4321,N_3807,N_3558);
xor U4322 (N_4322,N_3332,N_3811);
nand U4323 (N_4323,N_3835,N_3849);
xor U4324 (N_4324,N_3846,N_3970);
or U4325 (N_4325,N_3868,N_3822);
nor U4326 (N_4326,N_3857,N_3608);
and U4327 (N_4327,N_3901,N_3831);
or U4328 (N_4328,N_3925,N_3416);
nand U4329 (N_4329,N_3545,N_3994);
nor U4330 (N_4330,N_3315,N_3667);
nor U4331 (N_4331,N_3982,N_3823);
nor U4332 (N_4332,N_3567,N_3633);
and U4333 (N_4333,N_3984,N_3847);
nor U4334 (N_4334,N_3926,N_3393);
or U4335 (N_4335,N_3599,N_3352);
and U4336 (N_4336,N_3607,N_3791);
xor U4337 (N_4337,N_3751,N_3728);
nand U4338 (N_4338,N_3861,N_3687);
xor U4339 (N_4339,N_3634,N_3955);
nand U4340 (N_4340,N_3923,N_3346);
nor U4341 (N_4341,N_3489,N_3542);
and U4342 (N_4342,N_3674,N_3547);
and U4343 (N_4343,N_3941,N_3324);
nor U4344 (N_4344,N_3408,N_3739);
and U4345 (N_4345,N_3229,N_3300);
xor U4346 (N_4346,N_3321,N_3928);
xor U4347 (N_4347,N_3214,N_3979);
nor U4348 (N_4348,N_3472,N_3240);
and U4349 (N_4349,N_3819,N_3696);
or U4350 (N_4350,N_3980,N_3371);
nor U4351 (N_4351,N_3509,N_3951);
xor U4352 (N_4352,N_3686,N_3338);
nor U4353 (N_4353,N_3641,N_3882);
nand U4354 (N_4354,N_3383,N_3320);
nor U4355 (N_4355,N_3693,N_3921);
or U4356 (N_4356,N_3870,N_3498);
xnor U4357 (N_4357,N_3858,N_3463);
nand U4358 (N_4358,N_3414,N_3718);
and U4359 (N_4359,N_3828,N_3455);
nor U4360 (N_4360,N_3448,N_3457);
nand U4361 (N_4361,N_3258,N_3609);
nor U4362 (N_4362,N_3676,N_3657);
nor U4363 (N_4363,N_3311,N_3430);
nand U4364 (N_4364,N_3987,N_3569);
or U4365 (N_4365,N_3251,N_3452);
nand U4366 (N_4366,N_3437,N_3551);
xor U4367 (N_4367,N_3944,N_3812);
and U4368 (N_4368,N_3285,N_3699);
xor U4369 (N_4369,N_3688,N_3730);
xor U4370 (N_4370,N_3975,N_3705);
nor U4371 (N_4371,N_3969,N_3305);
nor U4372 (N_4372,N_3863,N_3486);
and U4373 (N_4373,N_3221,N_3640);
and U4374 (N_4374,N_3814,N_3683);
xnor U4375 (N_4375,N_3716,N_3796);
nor U4376 (N_4376,N_3911,N_3784);
or U4377 (N_4377,N_3353,N_3512);
nand U4378 (N_4378,N_3564,N_3827);
xnor U4379 (N_4379,N_3623,N_3445);
nor U4380 (N_4380,N_3232,N_3246);
or U4381 (N_4381,N_3215,N_3220);
and U4382 (N_4382,N_3379,N_3334);
or U4383 (N_4383,N_3272,N_3959);
nor U4384 (N_4384,N_3806,N_3566);
xnor U4385 (N_4385,N_3914,N_3770);
and U4386 (N_4386,N_3290,N_3903);
or U4387 (N_4387,N_3422,N_3815);
nand U4388 (N_4388,N_3528,N_3710);
xnor U4389 (N_4389,N_3276,N_3761);
or U4390 (N_4390,N_3316,N_3661);
nor U4391 (N_4391,N_3381,N_3423);
xnor U4392 (N_4392,N_3518,N_3927);
nand U4393 (N_4393,N_3210,N_3997);
nor U4394 (N_4394,N_3357,N_3404);
or U4395 (N_4395,N_3248,N_3924);
and U4396 (N_4396,N_3746,N_3935);
nand U4397 (N_4397,N_3771,N_3772);
nor U4398 (N_4398,N_3881,N_3748);
nand U4399 (N_4399,N_3721,N_3429);
or U4400 (N_4400,N_3570,N_3667);
xor U4401 (N_4401,N_3214,N_3854);
and U4402 (N_4402,N_3866,N_3733);
xnor U4403 (N_4403,N_3644,N_3510);
nor U4404 (N_4404,N_3420,N_3559);
and U4405 (N_4405,N_3477,N_3245);
xor U4406 (N_4406,N_3400,N_3890);
nand U4407 (N_4407,N_3479,N_3639);
and U4408 (N_4408,N_3836,N_3990);
and U4409 (N_4409,N_3427,N_3633);
xnor U4410 (N_4410,N_3537,N_3457);
and U4411 (N_4411,N_3375,N_3274);
nor U4412 (N_4412,N_3628,N_3677);
nand U4413 (N_4413,N_3363,N_3722);
nand U4414 (N_4414,N_3710,N_3782);
and U4415 (N_4415,N_3801,N_3418);
or U4416 (N_4416,N_3354,N_3220);
or U4417 (N_4417,N_3792,N_3976);
or U4418 (N_4418,N_3218,N_3381);
xor U4419 (N_4419,N_3367,N_3700);
and U4420 (N_4420,N_3467,N_3600);
or U4421 (N_4421,N_3346,N_3303);
nor U4422 (N_4422,N_3267,N_3910);
and U4423 (N_4423,N_3415,N_3806);
and U4424 (N_4424,N_3779,N_3402);
xnor U4425 (N_4425,N_3867,N_3730);
xor U4426 (N_4426,N_3808,N_3733);
nand U4427 (N_4427,N_3990,N_3420);
nor U4428 (N_4428,N_3601,N_3458);
nand U4429 (N_4429,N_3687,N_3821);
nand U4430 (N_4430,N_3987,N_3422);
or U4431 (N_4431,N_3562,N_3225);
nor U4432 (N_4432,N_3965,N_3345);
nor U4433 (N_4433,N_3471,N_3394);
or U4434 (N_4434,N_3200,N_3666);
nand U4435 (N_4435,N_3638,N_3856);
nand U4436 (N_4436,N_3357,N_3381);
nor U4437 (N_4437,N_3344,N_3827);
xor U4438 (N_4438,N_3677,N_3436);
or U4439 (N_4439,N_3407,N_3952);
nor U4440 (N_4440,N_3788,N_3672);
nor U4441 (N_4441,N_3583,N_3594);
and U4442 (N_4442,N_3417,N_3671);
nand U4443 (N_4443,N_3672,N_3602);
and U4444 (N_4444,N_3361,N_3739);
or U4445 (N_4445,N_3416,N_3352);
xor U4446 (N_4446,N_3749,N_3787);
and U4447 (N_4447,N_3915,N_3233);
nor U4448 (N_4448,N_3410,N_3446);
or U4449 (N_4449,N_3611,N_3820);
xor U4450 (N_4450,N_3486,N_3224);
nand U4451 (N_4451,N_3804,N_3391);
and U4452 (N_4452,N_3495,N_3572);
xnor U4453 (N_4453,N_3517,N_3684);
nand U4454 (N_4454,N_3522,N_3500);
nor U4455 (N_4455,N_3907,N_3346);
and U4456 (N_4456,N_3925,N_3404);
and U4457 (N_4457,N_3716,N_3521);
nand U4458 (N_4458,N_3485,N_3906);
and U4459 (N_4459,N_3587,N_3856);
nand U4460 (N_4460,N_3449,N_3317);
or U4461 (N_4461,N_3858,N_3295);
nand U4462 (N_4462,N_3498,N_3218);
nand U4463 (N_4463,N_3965,N_3251);
or U4464 (N_4464,N_3626,N_3228);
nand U4465 (N_4465,N_3946,N_3884);
xnor U4466 (N_4466,N_3931,N_3680);
and U4467 (N_4467,N_3580,N_3394);
or U4468 (N_4468,N_3481,N_3442);
xnor U4469 (N_4469,N_3314,N_3666);
nor U4470 (N_4470,N_3571,N_3609);
xor U4471 (N_4471,N_3380,N_3912);
nand U4472 (N_4472,N_3986,N_3462);
or U4473 (N_4473,N_3779,N_3741);
nand U4474 (N_4474,N_3410,N_3584);
or U4475 (N_4475,N_3495,N_3304);
nor U4476 (N_4476,N_3825,N_3557);
xor U4477 (N_4477,N_3710,N_3797);
nand U4478 (N_4478,N_3332,N_3954);
nor U4479 (N_4479,N_3891,N_3294);
nor U4480 (N_4480,N_3770,N_3940);
nor U4481 (N_4481,N_3222,N_3334);
xor U4482 (N_4482,N_3809,N_3280);
or U4483 (N_4483,N_3545,N_3971);
nand U4484 (N_4484,N_3948,N_3467);
nand U4485 (N_4485,N_3715,N_3376);
or U4486 (N_4486,N_3248,N_3695);
nand U4487 (N_4487,N_3986,N_3795);
and U4488 (N_4488,N_3243,N_3585);
or U4489 (N_4489,N_3267,N_3700);
nor U4490 (N_4490,N_3718,N_3686);
or U4491 (N_4491,N_3709,N_3670);
nor U4492 (N_4492,N_3624,N_3953);
or U4493 (N_4493,N_3996,N_3612);
nand U4494 (N_4494,N_3268,N_3475);
and U4495 (N_4495,N_3215,N_3229);
nor U4496 (N_4496,N_3280,N_3533);
and U4497 (N_4497,N_3213,N_3480);
and U4498 (N_4498,N_3776,N_3644);
nand U4499 (N_4499,N_3603,N_3204);
nand U4500 (N_4500,N_3809,N_3225);
nor U4501 (N_4501,N_3990,N_3410);
nor U4502 (N_4502,N_3668,N_3798);
xnor U4503 (N_4503,N_3322,N_3349);
nor U4504 (N_4504,N_3781,N_3612);
nand U4505 (N_4505,N_3318,N_3256);
nor U4506 (N_4506,N_3283,N_3304);
and U4507 (N_4507,N_3950,N_3499);
xnor U4508 (N_4508,N_3613,N_3984);
and U4509 (N_4509,N_3710,N_3344);
xnor U4510 (N_4510,N_3669,N_3326);
nor U4511 (N_4511,N_3832,N_3569);
or U4512 (N_4512,N_3441,N_3352);
nand U4513 (N_4513,N_3834,N_3755);
nor U4514 (N_4514,N_3289,N_3604);
and U4515 (N_4515,N_3314,N_3749);
xnor U4516 (N_4516,N_3908,N_3584);
nor U4517 (N_4517,N_3618,N_3241);
xnor U4518 (N_4518,N_3847,N_3878);
nand U4519 (N_4519,N_3913,N_3438);
xor U4520 (N_4520,N_3720,N_3255);
and U4521 (N_4521,N_3480,N_3395);
and U4522 (N_4522,N_3435,N_3246);
nand U4523 (N_4523,N_3382,N_3401);
nor U4524 (N_4524,N_3261,N_3564);
and U4525 (N_4525,N_3260,N_3805);
or U4526 (N_4526,N_3440,N_3888);
nor U4527 (N_4527,N_3476,N_3913);
nor U4528 (N_4528,N_3620,N_3684);
xnor U4529 (N_4529,N_3505,N_3395);
or U4530 (N_4530,N_3631,N_3206);
nor U4531 (N_4531,N_3797,N_3318);
nand U4532 (N_4532,N_3409,N_3515);
and U4533 (N_4533,N_3310,N_3665);
or U4534 (N_4534,N_3616,N_3354);
nand U4535 (N_4535,N_3349,N_3218);
nand U4536 (N_4536,N_3389,N_3388);
and U4537 (N_4537,N_3802,N_3566);
nand U4538 (N_4538,N_3513,N_3425);
or U4539 (N_4539,N_3858,N_3457);
xnor U4540 (N_4540,N_3912,N_3940);
and U4541 (N_4541,N_3357,N_3583);
nand U4542 (N_4542,N_3735,N_3505);
nand U4543 (N_4543,N_3237,N_3940);
and U4544 (N_4544,N_3385,N_3209);
nand U4545 (N_4545,N_3302,N_3365);
nor U4546 (N_4546,N_3846,N_3266);
xor U4547 (N_4547,N_3892,N_3739);
or U4548 (N_4548,N_3753,N_3321);
nand U4549 (N_4549,N_3516,N_3264);
nor U4550 (N_4550,N_3595,N_3752);
or U4551 (N_4551,N_3898,N_3926);
xnor U4552 (N_4552,N_3941,N_3795);
xnor U4553 (N_4553,N_3638,N_3886);
xor U4554 (N_4554,N_3264,N_3949);
or U4555 (N_4555,N_3217,N_3750);
xor U4556 (N_4556,N_3969,N_3457);
nand U4557 (N_4557,N_3245,N_3660);
or U4558 (N_4558,N_3967,N_3620);
or U4559 (N_4559,N_3979,N_3825);
and U4560 (N_4560,N_3297,N_3822);
or U4561 (N_4561,N_3810,N_3797);
or U4562 (N_4562,N_3893,N_3829);
nand U4563 (N_4563,N_3583,N_3787);
xor U4564 (N_4564,N_3742,N_3401);
xnor U4565 (N_4565,N_3608,N_3970);
and U4566 (N_4566,N_3573,N_3880);
nor U4567 (N_4567,N_3690,N_3963);
nor U4568 (N_4568,N_3508,N_3490);
and U4569 (N_4569,N_3843,N_3312);
or U4570 (N_4570,N_3699,N_3550);
nor U4571 (N_4571,N_3251,N_3357);
xor U4572 (N_4572,N_3493,N_3261);
and U4573 (N_4573,N_3650,N_3289);
nor U4574 (N_4574,N_3895,N_3521);
nor U4575 (N_4575,N_3785,N_3606);
or U4576 (N_4576,N_3635,N_3778);
nor U4577 (N_4577,N_3576,N_3718);
or U4578 (N_4578,N_3564,N_3464);
nand U4579 (N_4579,N_3997,N_3900);
xor U4580 (N_4580,N_3695,N_3561);
nor U4581 (N_4581,N_3480,N_3819);
xnor U4582 (N_4582,N_3481,N_3886);
and U4583 (N_4583,N_3935,N_3872);
xnor U4584 (N_4584,N_3307,N_3439);
or U4585 (N_4585,N_3624,N_3568);
nor U4586 (N_4586,N_3684,N_3990);
nand U4587 (N_4587,N_3730,N_3871);
nor U4588 (N_4588,N_3411,N_3295);
nand U4589 (N_4589,N_3884,N_3394);
nor U4590 (N_4590,N_3432,N_3222);
or U4591 (N_4591,N_3882,N_3814);
nor U4592 (N_4592,N_3521,N_3480);
xnor U4593 (N_4593,N_3957,N_3481);
and U4594 (N_4594,N_3853,N_3617);
nand U4595 (N_4595,N_3335,N_3882);
nand U4596 (N_4596,N_3446,N_3518);
xnor U4597 (N_4597,N_3946,N_3880);
nor U4598 (N_4598,N_3276,N_3444);
xnor U4599 (N_4599,N_3543,N_3618);
nand U4600 (N_4600,N_3573,N_3522);
and U4601 (N_4601,N_3698,N_3358);
xnor U4602 (N_4602,N_3485,N_3291);
nand U4603 (N_4603,N_3994,N_3302);
nand U4604 (N_4604,N_3921,N_3725);
nand U4605 (N_4605,N_3333,N_3397);
and U4606 (N_4606,N_3992,N_3376);
nand U4607 (N_4607,N_3377,N_3734);
or U4608 (N_4608,N_3443,N_3285);
xnor U4609 (N_4609,N_3988,N_3301);
nand U4610 (N_4610,N_3343,N_3555);
nor U4611 (N_4611,N_3923,N_3644);
nand U4612 (N_4612,N_3267,N_3244);
xor U4613 (N_4613,N_3831,N_3693);
nand U4614 (N_4614,N_3945,N_3923);
xor U4615 (N_4615,N_3863,N_3801);
nand U4616 (N_4616,N_3312,N_3486);
or U4617 (N_4617,N_3984,N_3358);
nor U4618 (N_4618,N_3498,N_3932);
nand U4619 (N_4619,N_3290,N_3299);
xnor U4620 (N_4620,N_3440,N_3361);
nand U4621 (N_4621,N_3794,N_3804);
and U4622 (N_4622,N_3599,N_3547);
and U4623 (N_4623,N_3228,N_3475);
nor U4624 (N_4624,N_3598,N_3250);
nand U4625 (N_4625,N_3971,N_3873);
nor U4626 (N_4626,N_3284,N_3914);
or U4627 (N_4627,N_3962,N_3908);
nand U4628 (N_4628,N_3489,N_3906);
and U4629 (N_4629,N_3281,N_3964);
nor U4630 (N_4630,N_3293,N_3344);
nand U4631 (N_4631,N_3963,N_3491);
xnor U4632 (N_4632,N_3770,N_3889);
nand U4633 (N_4633,N_3838,N_3930);
xor U4634 (N_4634,N_3211,N_3354);
or U4635 (N_4635,N_3846,N_3967);
nand U4636 (N_4636,N_3834,N_3588);
or U4637 (N_4637,N_3506,N_3998);
or U4638 (N_4638,N_3457,N_3798);
or U4639 (N_4639,N_3731,N_3734);
nand U4640 (N_4640,N_3724,N_3226);
nor U4641 (N_4641,N_3874,N_3727);
and U4642 (N_4642,N_3539,N_3352);
nor U4643 (N_4643,N_3572,N_3692);
nor U4644 (N_4644,N_3897,N_3250);
nor U4645 (N_4645,N_3293,N_3704);
nor U4646 (N_4646,N_3617,N_3464);
xnor U4647 (N_4647,N_3948,N_3462);
nor U4648 (N_4648,N_3508,N_3538);
nor U4649 (N_4649,N_3603,N_3469);
nand U4650 (N_4650,N_3923,N_3859);
or U4651 (N_4651,N_3958,N_3852);
and U4652 (N_4652,N_3415,N_3999);
nand U4653 (N_4653,N_3401,N_3383);
and U4654 (N_4654,N_3937,N_3311);
nand U4655 (N_4655,N_3206,N_3962);
xnor U4656 (N_4656,N_3849,N_3233);
or U4657 (N_4657,N_3805,N_3208);
or U4658 (N_4658,N_3333,N_3541);
and U4659 (N_4659,N_3507,N_3403);
or U4660 (N_4660,N_3501,N_3225);
and U4661 (N_4661,N_3477,N_3386);
xor U4662 (N_4662,N_3805,N_3410);
or U4663 (N_4663,N_3475,N_3845);
or U4664 (N_4664,N_3251,N_3995);
or U4665 (N_4665,N_3661,N_3355);
nand U4666 (N_4666,N_3300,N_3381);
nor U4667 (N_4667,N_3411,N_3688);
or U4668 (N_4668,N_3800,N_3963);
nor U4669 (N_4669,N_3489,N_3881);
nor U4670 (N_4670,N_3318,N_3639);
and U4671 (N_4671,N_3623,N_3566);
xnor U4672 (N_4672,N_3837,N_3481);
xnor U4673 (N_4673,N_3381,N_3824);
nand U4674 (N_4674,N_3982,N_3931);
nor U4675 (N_4675,N_3557,N_3705);
nand U4676 (N_4676,N_3215,N_3317);
xor U4677 (N_4677,N_3973,N_3585);
nor U4678 (N_4678,N_3657,N_3800);
or U4679 (N_4679,N_3638,N_3775);
nand U4680 (N_4680,N_3351,N_3554);
nand U4681 (N_4681,N_3574,N_3433);
and U4682 (N_4682,N_3917,N_3912);
or U4683 (N_4683,N_3840,N_3905);
nand U4684 (N_4684,N_3561,N_3942);
xnor U4685 (N_4685,N_3288,N_3915);
nand U4686 (N_4686,N_3778,N_3508);
xor U4687 (N_4687,N_3751,N_3681);
nand U4688 (N_4688,N_3661,N_3703);
xor U4689 (N_4689,N_3496,N_3292);
nor U4690 (N_4690,N_3201,N_3536);
nand U4691 (N_4691,N_3383,N_3544);
or U4692 (N_4692,N_3540,N_3242);
or U4693 (N_4693,N_3285,N_3958);
nand U4694 (N_4694,N_3725,N_3660);
nor U4695 (N_4695,N_3284,N_3297);
xor U4696 (N_4696,N_3579,N_3505);
or U4697 (N_4697,N_3440,N_3749);
or U4698 (N_4698,N_3273,N_3454);
xnor U4699 (N_4699,N_3455,N_3398);
or U4700 (N_4700,N_3306,N_3414);
nor U4701 (N_4701,N_3583,N_3404);
or U4702 (N_4702,N_3777,N_3523);
nand U4703 (N_4703,N_3376,N_3208);
nor U4704 (N_4704,N_3266,N_3291);
nor U4705 (N_4705,N_3304,N_3453);
nor U4706 (N_4706,N_3534,N_3258);
or U4707 (N_4707,N_3368,N_3843);
or U4708 (N_4708,N_3583,N_3947);
nand U4709 (N_4709,N_3406,N_3631);
nand U4710 (N_4710,N_3421,N_3802);
nor U4711 (N_4711,N_3970,N_3956);
xnor U4712 (N_4712,N_3700,N_3773);
nand U4713 (N_4713,N_3444,N_3822);
nand U4714 (N_4714,N_3338,N_3493);
nor U4715 (N_4715,N_3205,N_3393);
nor U4716 (N_4716,N_3441,N_3335);
nor U4717 (N_4717,N_3899,N_3656);
nor U4718 (N_4718,N_3824,N_3551);
nand U4719 (N_4719,N_3718,N_3317);
nand U4720 (N_4720,N_3504,N_3528);
xor U4721 (N_4721,N_3333,N_3262);
and U4722 (N_4722,N_3921,N_3398);
and U4723 (N_4723,N_3868,N_3348);
or U4724 (N_4724,N_3456,N_3876);
and U4725 (N_4725,N_3338,N_3565);
or U4726 (N_4726,N_3257,N_3231);
xnor U4727 (N_4727,N_3874,N_3285);
and U4728 (N_4728,N_3896,N_3681);
and U4729 (N_4729,N_3865,N_3560);
or U4730 (N_4730,N_3891,N_3511);
nand U4731 (N_4731,N_3597,N_3466);
or U4732 (N_4732,N_3711,N_3982);
xor U4733 (N_4733,N_3804,N_3524);
nand U4734 (N_4734,N_3821,N_3705);
or U4735 (N_4735,N_3439,N_3490);
xor U4736 (N_4736,N_3670,N_3265);
and U4737 (N_4737,N_3714,N_3596);
xor U4738 (N_4738,N_3332,N_3612);
xnor U4739 (N_4739,N_3904,N_3382);
xnor U4740 (N_4740,N_3337,N_3579);
and U4741 (N_4741,N_3626,N_3315);
and U4742 (N_4742,N_3949,N_3842);
nand U4743 (N_4743,N_3627,N_3756);
or U4744 (N_4744,N_3249,N_3315);
or U4745 (N_4745,N_3884,N_3920);
nor U4746 (N_4746,N_3776,N_3839);
and U4747 (N_4747,N_3916,N_3351);
xnor U4748 (N_4748,N_3592,N_3406);
xor U4749 (N_4749,N_3996,N_3291);
nor U4750 (N_4750,N_3542,N_3845);
nand U4751 (N_4751,N_3572,N_3712);
and U4752 (N_4752,N_3322,N_3534);
and U4753 (N_4753,N_3455,N_3597);
nand U4754 (N_4754,N_3585,N_3701);
nand U4755 (N_4755,N_3586,N_3696);
and U4756 (N_4756,N_3761,N_3935);
and U4757 (N_4757,N_3211,N_3870);
and U4758 (N_4758,N_3871,N_3507);
nand U4759 (N_4759,N_3882,N_3516);
xnor U4760 (N_4760,N_3431,N_3373);
or U4761 (N_4761,N_3243,N_3760);
nand U4762 (N_4762,N_3451,N_3681);
or U4763 (N_4763,N_3500,N_3200);
nand U4764 (N_4764,N_3873,N_3991);
nor U4765 (N_4765,N_3846,N_3687);
and U4766 (N_4766,N_3326,N_3701);
xnor U4767 (N_4767,N_3692,N_3646);
nand U4768 (N_4768,N_3459,N_3469);
nor U4769 (N_4769,N_3964,N_3587);
nand U4770 (N_4770,N_3703,N_3260);
and U4771 (N_4771,N_3920,N_3558);
and U4772 (N_4772,N_3873,N_3385);
xor U4773 (N_4773,N_3889,N_3589);
or U4774 (N_4774,N_3921,N_3222);
and U4775 (N_4775,N_3588,N_3409);
nand U4776 (N_4776,N_3494,N_3890);
xnor U4777 (N_4777,N_3632,N_3248);
nor U4778 (N_4778,N_3543,N_3470);
nand U4779 (N_4779,N_3941,N_3777);
and U4780 (N_4780,N_3757,N_3966);
nor U4781 (N_4781,N_3568,N_3799);
or U4782 (N_4782,N_3971,N_3655);
nor U4783 (N_4783,N_3658,N_3616);
nor U4784 (N_4784,N_3520,N_3844);
xor U4785 (N_4785,N_3272,N_3663);
or U4786 (N_4786,N_3650,N_3399);
nand U4787 (N_4787,N_3972,N_3653);
nand U4788 (N_4788,N_3611,N_3236);
xor U4789 (N_4789,N_3491,N_3966);
and U4790 (N_4790,N_3438,N_3591);
nor U4791 (N_4791,N_3258,N_3550);
and U4792 (N_4792,N_3515,N_3499);
and U4793 (N_4793,N_3313,N_3499);
and U4794 (N_4794,N_3595,N_3406);
nor U4795 (N_4795,N_3441,N_3871);
xor U4796 (N_4796,N_3808,N_3577);
or U4797 (N_4797,N_3757,N_3531);
xor U4798 (N_4798,N_3858,N_3623);
and U4799 (N_4799,N_3553,N_3280);
nand U4800 (N_4800,N_4720,N_4516);
xnor U4801 (N_4801,N_4697,N_4433);
xor U4802 (N_4802,N_4467,N_4015);
nand U4803 (N_4803,N_4346,N_4369);
nand U4804 (N_4804,N_4021,N_4569);
and U4805 (N_4805,N_4031,N_4297);
xor U4806 (N_4806,N_4455,N_4044);
nand U4807 (N_4807,N_4544,N_4529);
xor U4808 (N_4808,N_4773,N_4396);
nor U4809 (N_4809,N_4154,N_4225);
or U4810 (N_4810,N_4246,N_4728);
and U4811 (N_4811,N_4434,N_4120);
and U4812 (N_4812,N_4014,N_4118);
nand U4813 (N_4813,N_4289,N_4703);
nand U4814 (N_4814,N_4729,N_4394);
xor U4815 (N_4815,N_4230,N_4468);
nand U4816 (N_4816,N_4579,N_4315);
xor U4817 (N_4817,N_4384,N_4349);
nor U4818 (N_4818,N_4584,N_4294);
or U4819 (N_4819,N_4058,N_4410);
or U4820 (N_4820,N_4690,N_4519);
nand U4821 (N_4821,N_4514,N_4328);
or U4822 (N_4822,N_4511,N_4020);
xnor U4823 (N_4823,N_4647,N_4064);
nand U4824 (N_4824,N_4160,N_4745);
nand U4825 (N_4825,N_4568,N_4431);
nand U4826 (N_4826,N_4252,N_4793);
and U4827 (N_4827,N_4056,N_4236);
xnor U4828 (N_4828,N_4784,N_4070);
or U4829 (N_4829,N_4596,N_4408);
or U4830 (N_4830,N_4721,N_4435);
nor U4831 (N_4831,N_4525,N_4678);
xnor U4832 (N_4832,N_4608,N_4286);
nor U4833 (N_4833,N_4597,N_4221);
xor U4834 (N_4834,N_4028,N_4622);
or U4835 (N_4835,N_4082,N_4293);
nor U4836 (N_4836,N_4701,N_4126);
nand U4837 (N_4837,N_4642,N_4344);
and U4838 (N_4838,N_4567,N_4530);
nand U4839 (N_4839,N_4095,N_4254);
xor U4840 (N_4840,N_4256,N_4442);
nor U4841 (N_4841,N_4389,N_4207);
or U4842 (N_4842,N_4366,N_4782);
nor U4843 (N_4843,N_4499,N_4444);
and U4844 (N_4844,N_4534,N_4262);
nor U4845 (N_4845,N_4418,N_4491);
nor U4846 (N_4846,N_4603,N_4423);
nor U4847 (N_4847,N_4245,N_4117);
nand U4848 (N_4848,N_4365,N_4350);
nor U4849 (N_4849,N_4779,N_4108);
nand U4850 (N_4850,N_4688,N_4576);
xor U4851 (N_4851,N_4089,N_4553);
nand U4852 (N_4852,N_4149,N_4086);
nor U4853 (N_4853,N_4589,N_4482);
nor U4854 (N_4854,N_4724,N_4247);
xnor U4855 (N_4855,N_4222,N_4096);
and U4856 (N_4856,N_4269,N_4535);
and U4857 (N_4857,N_4799,N_4422);
xnor U4858 (N_4858,N_4605,N_4224);
xnor U4859 (N_4859,N_4092,N_4476);
or U4860 (N_4860,N_4486,N_4751);
or U4861 (N_4861,N_4611,N_4138);
and U4862 (N_4862,N_4776,N_4133);
and U4863 (N_4863,N_4322,N_4065);
xor U4864 (N_4864,N_4066,N_4474);
nor U4865 (N_4865,N_4536,N_4448);
nor U4866 (N_4866,N_4746,N_4740);
and U4867 (N_4867,N_4285,N_4201);
or U4868 (N_4868,N_4123,N_4662);
nand U4869 (N_4869,N_4367,N_4053);
or U4870 (N_4870,N_4152,N_4456);
xor U4871 (N_4871,N_4683,N_4507);
or U4872 (N_4872,N_4135,N_4570);
nor U4873 (N_4873,N_4517,N_4166);
nand U4874 (N_4874,N_4428,N_4374);
nor U4875 (N_4875,N_4099,N_4227);
and U4876 (N_4876,N_4763,N_4577);
and U4877 (N_4877,N_4541,N_4758);
nand U4878 (N_4878,N_4103,N_4665);
xnor U4879 (N_4879,N_4427,N_4698);
xor U4880 (N_4880,N_4627,N_4786);
nand U4881 (N_4881,N_4337,N_4676);
xnor U4882 (N_4882,N_4318,N_4582);
nor U4883 (N_4883,N_4006,N_4079);
nor U4884 (N_4884,N_4275,N_4296);
or U4885 (N_4885,N_4426,N_4136);
xor U4886 (N_4886,N_4235,N_4736);
nor U4887 (N_4887,N_4493,N_4791);
nand U4888 (N_4888,N_4595,N_4749);
xnor U4889 (N_4889,N_4357,N_4156);
nor U4890 (N_4890,N_4393,N_4528);
nand U4891 (N_4891,N_4131,N_4324);
and U4892 (N_4892,N_4051,N_4167);
and U4893 (N_4893,N_4378,N_4756);
and U4894 (N_4894,N_4424,N_4327);
nor U4895 (N_4895,N_4764,N_4205);
xor U4896 (N_4896,N_4777,N_4109);
or U4897 (N_4897,N_4760,N_4656);
nand U4898 (N_4898,N_4008,N_4592);
xor U4899 (N_4899,N_4283,N_4446);
or U4900 (N_4900,N_4307,N_4391);
and U4901 (N_4901,N_4206,N_4667);
xnor U4902 (N_4902,N_4005,N_4795);
nand U4903 (N_4903,N_4498,N_4716);
nor U4904 (N_4904,N_4073,N_4602);
nand U4905 (N_4905,N_4364,N_4342);
nand U4906 (N_4906,N_4267,N_4069);
nor U4907 (N_4907,N_4203,N_4362);
and U4908 (N_4908,N_4604,N_4071);
and U4909 (N_4909,N_4310,N_4420);
nand U4910 (N_4910,N_4274,N_4129);
nand U4911 (N_4911,N_4626,N_4417);
nand U4912 (N_4912,N_4032,N_4072);
or U4913 (N_4913,N_4340,N_4437);
nor U4914 (N_4914,N_4657,N_4195);
or U4915 (N_4915,N_4727,N_4502);
and U4916 (N_4916,N_4062,N_4067);
xor U4917 (N_4917,N_4638,N_4292);
or U4918 (N_4918,N_4194,N_4034);
or U4919 (N_4919,N_4329,N_4587);
and U4920 (N_4920,N_4325,N_4668);
nand U4921 (N_4921,N_4334,N_4445);
nand U4922 (N_4922,N_4217,N_4359);
and U4923 (N_4923,N_4027,N_4029);
xor U4924 (N_4924,N_4231,N_4765);
or U4925 (N_4925,N_4425,N_4026);
nand U4926 (N_4926,N_4271,N_4047);
xnor U4927 (N_4927,N_4239,N_4780);
nand U4928 (N_4928,N_4343,N_4505);
or U4929 (N_4929,N_4465,N_4214);
nor U4930 (N_4930,N_4007,N_4717);
nor U4931 (N_4931,N_4093,N_4674);
xnor U4932 (N_4932,N_4709,N_4124);
or U4933 (N_4933,N_4741,N_4450);
and U4934 (N_4934,N_4770,N_4001);
nand U4935 (N_4935,N_4232,N_4515);
xor U4936 (N_4936,N_4700,N_4648);
nand U4937 (N_4937,N_4742,N_4766);
or U4938 (N_4938,N_4664,N_4218);
xor U4939 (N_4939,N_4409,N_4651);
nor U4940 (N_4940,N_4671,N_4685);
or U4941 (N_4941,N_4681,N_4375);
xnor U4942 (N_4942,N_4052,N_4303);
and U4943 (N_4943,N_4533,N_4270);
nand U4944 (N_4944,N_4261,N_4351);
nor U4945 (N_4945,N_4022,N_4625);
and U4946 (N_4946,N_4043,N_4354);
nand U4947 (N_4947,N_4219,N_4753);
nor U4948 (N_4948,N_4250,N_4299);
or U4949 (N_4949,N_4107,N_4543);
nand U4950 (N_4950,N_4600,N_4726);
xnor U4951 (N_4951,N_4237,N_4390);
or U4952 (N_4952,N_4345,N_4652);
and U4953 (N_4953,N_4240,N_4451);
and U4954 (N_4954,N_4488,N_4305);
or U4955 (N_4955,N_4102,N_4682);
xnor U4956 (N_4956,N_4041,N_4737);
or U4957 (N_4957,N_4115,N_4613);
xor U4958 (N_4958,N_4188,N_4302);
nand U4959 (N_4959,N_4150,N_4537);
or U4960 (N_4960,N_4755,N_4348);
nor U4961 (N_4961,N_4010,N_4457);
nor U4962 (N_4962,N_4615,N_4085);
nor U4963 (N_4963,N_4769,N_4513);
nor U4964 (N_4964,N_4172,N_4501);
xor U4965 (N_4965,N_4161,N_4162);
and U4966 (N_4966,N_4508,N_4171);
or U4967 (N_4967,N_4370,N_4272);
nor U4968 (N_4968,N_4460,N_4732);
and U4969 (N_4969,N_4183,N_4104);
nand U4970 (N_4970,N_4691,N_4128);
or U4971 (N_4971,N_4407,N_4125);
and U4972 (N_4972,N_4191,N_4616);
nor U4973 (N_4973,N_4278,N_4540);
nor U4974 (N_4974,N_4273,N_4168);
nand U4975 (N_4975,N_4494,N_4670);
or U4976 (N_4976,N_4238,N_4331);
or U4977 (N_4977,N_4398,N_4190);
or U4978 (N_4978,N_4101,N_4134);
nand U4979 (N_4979,N_4531,N_4735);
nor U4980 (N_4980,N_4074,N_4573);
or U4981 (N_4981,N_4288,N_4377);
or U4982 (N_4982,N_4045,N_4633);
nand U4983 (N_4983,N_4555,N_4586);
nand U4984 (N_4984,N_4105,N_4178);
or U4985 (N_4985,N_4185,N_4308);
and U4986 (N_4986,N_4719,N_4771);
nor U4987 (N_4987,N_4618,N_4241);
nand U4988 (N_4988,N_4313,N_4312);
xor U4989 (N_4989,N_4326,N_4414);
xor U4990 (N_4990,N_4556,N_4287);
or U4991 (N_4991,N_4580,N_4649);
nand U4992 (N_4992,N_4012,N_4257);
xnor U4993 (N_4993,N_4504,N_4754);
xnor U4994 (N_4994,N_4386,N_4768);
nand U4995 (N_4995,N_4042,N_4144);
xor U4996 (N_4996,N_4554,N_4419);
xor U4997 (N_4997,N_4694,N_4562);
nand U4998 (N_4998,N_4335,N_4304);
xnor U4999 (N_4999,N_4215,N_4019);
nand U5000 (N_5000,N_4202,N_4757);
nand U5001 (N_5001,N_4684,N_4588);
xor U5002 (N_5002,N_4094,N_4263);
nand U5003 (N_5003,N_4163,N_4752);
xor U5004 (N_5004,N_4487,N_4411);
or U5005 (N_5005,N_4495,N_4170);
nand U5006 (N_5006,N_4653,N_4628);
or U5007 (N_5007,N_4748,N_4148);
nor U5008 (N_5008,N_4229,N_4549);
xnor U5009 (N_5009,N_4443,N_4199);
nand U5010 (N_5010,N_4571,N_4087);
or U5011 (N_5011,N_4258,N_4100);
and U5012 (N_5012,N_4037,N_4265);
and U5013 (N_5013,N_4255,N_4209);
and U5014 (N_5014,N_4759,N_4677);
and U5015 (N_5015,N_4114,N_4228);
and U5016 (N_5016,N_4057,N_4672);
nor U5017 (N_5017,N_4298,N_4610);
nor U5018 (N_5018,N_4492,N_4281);
nor U5019 (N_5019,N_4778,N_4775);
or U5020 (N_5020,N_4518,N_4405);
xor U5021 (N_5021,N_4796,N_4524);
nor U5022 (N_5022,N_4180,N_4300);
nor U5023 (N_5023,N_4084,N_4702);
nor U5024 (N_5024,N_4211,N_4061);
and U5025 (N_5025,N_4055,N_4661);
nand U5026 (N_5026,N_4712,N_4477);
or U5027 (N_5027,N_4279,N_4459);
and U5028 (N_5028,N_4660,N_4204);
nand U5029 (N_5029,N_4248,N_4551);
nand U5030 (N_5030,N_4637,N_4030);
nand U5031 (N_5031,N_4368,N_4655);
and U5032 (N_5032,N_4243,N_4016);
and U5033 (N_5033,N_4472,N_4213);
or U5034 (N_5034,N_4506,N_4510);
xnor U5035 (N_5035,N_4738,N_4710);
xnor U5036 (N_5036,N_4548,N_4347);
or U5037 (N_5037,N_4415,N_4363);
or U5038 (N_5038,N_4695,N_4177);
or U5039 (N_5039,N_4725,N_4311);
or U5040 (N_5040,N_4761,N_4790);
and U5041 (N_5041,N_4353,N_4151);
nor U5042 (N_5042,N_4646,N_4306);
nor U5043 (N_5043,N_4621,N_4787);
xnor U5044 (N_5044,N_4438,N_4547);
nor U5045 (N_5045,N_4654,N_4747);
xor U5046 (N_5046,N_4080,N_4452);
nand U5047 (N_5047,N_4461,N_4552);
xnor U5048 (N_5048,N_4601,N_4155);
and U5049 (N_5049,N_4290,N_4339);
nand U5050 (N_5050,N_4400,N_4572);
nor U5051 (N_5051,N_4333,N_4314);
nor U5052 (N_5052,N_4762,N_4035);
nor U5053 (N_5053,N_4234,N_4489);
xnor U5054 (N_5054,N_4317,N_4282);
or U5055 (N_5055,N_4075,N_4645);
or U5056 (N_5056,N_4673,N_4500);
xnor U5057 (N_5057,N_4189,N_4119);
nor U5058 (N_5058,N_4635,N_4607);
nor U5059 (N_5059,N_4392,N_4744);
nor U5060 (N_5060,N_4223,N_4078);
xnor U5061 (N_5061,N_4193,N_4088);
and U5062 (N_5062,N_4040,N_4251);
or U5063 (N_5063,N_4192,N_4113);
xor U5064 (N_5064,N_4083,N_4539);
and U5065 (N_5065,N_4704,N_4182);
and U5066 (N_5066,N_4309,N_4046);
or U5067 (N_5067,N_4658,N_4696);
or U5068 (N_5068,N_4453,N_4382);
xor U5069 (N_5069,N_4259,N_4371);
xnor U5070 (N_5070,N_4715,N_4641);
xor U5071 (N_5071,N_4743,N_4619);
xor U5072 (N_5072,N_4212,N_4198);
nor U5073 (N_5073,N_4578,N_4112);
and U5074 (N_5074,N_4679,N_4669);
xor U5075 (N_5075,N_4301,N_4566);
or U5076 (N_5076,N_4184,N_4000);
xor U5077 (N_5077,N_4049,N_4174);
nand U5078 (N_5078,N_4785,N_4320);
nand U5079 (N_5079,N_4121,N_4464);
and U5080 (N_5080,N_4523,N_4381);
or U5081 (N_5081,N_4169,N_4323);
or U5082 (N_5082,N_4481,N_4077);
or U5083 (N_5083,N_4385,N_4629);
nand U5084 (N_5084,N_4036,N_4276);
or U5085 (N_5085,N_4797,N_4590);
xor U5086 (N_5086,N_4404,N_4666);
nand U5087 (N_5087,N_4478,N_4081);
nor U5088 (N_5088,N_4009,N_4264);
or U5089 (N_5089,N_4332,N_4557);
and U5090 (N_5090,N_4574,N_4583);
or U5091 (N_5091,N_4441,N_4479);
nor U5092 (N_5092,N_4153,N_4789);
or U5093 (N_5093,N_4004,N_4164);
nor U5094 (N_5094,N_4197,N_4527);
nand U5095 (N_5095,N_4440,N_4473);
xnor U5096 (N_5096,N_4520,N_4462);
nor U5097 (N_5097,N_4734,N_4401);
and U5098 (N_5098,N_4593,N_4122);
or U5099 (N_5099,N_4430,N_4623);
xnor U5100 (N_5100,N_4614,N_4412);
nor U5101 (N_5101,N_4559,N_4399);
xnor U5102 (N_5102,N_4249,N_4458);
nor U5103 (N_5103,N_4632,N_4447);
nand U5104 (N_5104,N_4388,N_4686);
and U5105 (N_5105,N_4565,N_4594);
or U5106 (N_5106,N_4208,N_4033);
and U5107 (N_5107,N_4220,N_4358);
or U5108 (N_5108,N_4772,N_4372);
or U5109 (N_5109,N_4352,N_4011);
nor U5110 (N_5110,N_4280,N_4620);
and U5111 (N_5111,N_4143,N_4708);
or U5112 (N_5112,N_4110,N_4512);
nand U5113 (N_5113,N_4532,N_4463);
or U5114 (N_5114,N_4675,N_4048);
xnor U5115 (N_5115,N_4050,N_4330);
and U5116 (N_5116,N_4395,N_4379);
or U5117 (N_5117,N_4175,N_4713);
nand U5118 (N_5118,N_4705,N_4127);
and U5119 (N_5119,N_4416,N_4355);
xor U5120 (N_5120,N_4630,N_4141);
nor U5121 (N_5121,N_4739,N_4397);
and U5122 (N_5122,N_4321,N_4165);
or U5123 (N_5123,N_4490,N_4116);
xor U5124 (N_5124,N_4060,N_4640);
nand U5125 (N_5125,N_4413,N_4723);
nor U5126 (N_5126,N_4360,N_4774);
nor U5127 (N_5127,N_4098,N_4781);
and U5128 (N_5128,N_4439,N_4338);
xor U5129 (N_5129,N_4023,N_4631);
xnor U5130 (N_5130,N_4609,N_4650);
nor U5131 (N_5131,N_4680,N_4159);
and U5132 (N_5132,N_4575,N_4059);
nand U5133 (N_5133,N_4585,N_4356);
or U5134 (N_5134,N_4521,N_4466);
nor U5135 (N_5135,N_4509,N_4663);
or U5136 (N_5136,N_4722,N_4454);
nand U5137 (N_5137,N_4216,N_4076);
nor U5138 (N_5138,N_4798,N_4624);
xnor U5139 (N_5139,N_4480,N_4792);
xnor U5140 (N_5140,N_4284,N_4266);
or U5141 (N_5141,N_4319,N_4699);
nor U5142 (N_5142,N_4617,N_4260);
and U5143 (N_5143,N_4106,N_4707);
and U5144 (N_5144,N_4383,N_4068);
xor U5145 (N_5145,N_4173,N_4090);
and U5146 (N_5146,N_4564,N_4475);
or U5147 (N_5147,N_4361,N_4503);
nand U5148 (N_5148,N_4538,N_4706);
and U5149 (N_5149,N_4268,N_4017);
nand U5150 (N_5150,N_4025,N_4484);
nor U5151 (N_5151,N_4130,N_4733);
or U5152 (N_5152,N_4187,N_4421);
and U5153 (N_5153,N_4469,N_4591);
and U5154 (N_5154,N_4137,N_4024);
xor U5155 (N_5155,N_4176,N_4376);
nor U5156 (N_5156,N_4471,N_4295);
nand U5157 (N_5157,N_4373,N_4750);
or U5158 (N_5158,N_4403,N_4794);
nor U5159 (N_5159,N_4380,N_4693);
and U5160 (N_5160,N_4018,N_4432);
or U5161 (N_5161,N_4429,N_4200);
nand U5162 (N_5162,N_4146,N_4643);
or U5163 (N_5163,N_4233,N_4244);
nand U5164 (N_5164,N_4226,N_4606);
xnor U5165 (N_5165,N_4242,N_4179);
nor U5166 (N_5166,N_4186,N_4711);
or U5167 (N_5167,N_4277,N_4714);
nand U5168 (N_5168,N_4145,N_4054);
and U5169 (N_5169,N_4687,N_4598);
nand U5170 (N_5170,N_4783,N_4111);
nand U5171 (N_5171,N_4718,N_4402);
nand U5172 (N_5172,N_4639,N_4788);
and U5173 (N_5173,N_4140,N_4634);
or U5174 (N_5174,N_4542,N_4387);
nor U5175 (N_5175,N_4689,N_4644);
nor U5176 (N_5176,N_4731,N_4002);
nor U5177 (N_5177,N_4210,N_4563);
nor U5178 (N_5178,N_4341,N_4406);
and U5179 (N_5179,N_4316,N_4558);
or U5180 (N_5180,N_4496,N_4063);
nor U5181 (N_5181,N_4181,N_4730);
and U5182 (N_5182,N_4139,N_4599);
nand U5183 (N_5183,N_4497,N_4485);
nand U5184 (N_5184,N_4013,N_4449);
or U5185 (N_5185,N_4091,N_4560);
nand U5186 (N_5186,N_4581,N_4038);
xor U5187 (N_5187,N_4545,N_4612);
nor U5188 (N_5188,N_4636,N_4436);
and U5189 (N_5189,N_4526,N_4158);
or U5190 (N_5190,N_4003,N_4561);
nand U5191 (N_5191,N_4132,N_4767);
nor U5192 (N_5192,N_4253,N_4522);
or U5193 (N_5193,N_4692,N_4157);
nor U5194 (N_5194,N_4336,N_4483);
xnor U5195 (N_5195,N_4550,N_4142);
xor U5196 (N_5196,N_4097,N_4147);
or U5197 (N_5197,N_4039,N_4470);
xnor U5198 (N_5198,N_4546,N_4196);
nand U5199 (N_5199,N_4291,N_4659);
or U5200 (N_5200,N_4108,N_4421);
nor U5201 (N_5201,N_4531,N_4181);
or U5202 (N_5202,N_4499,N_4147);
and U5203 (N_5203,N_4661,N_4766);
xnor U5204 (N_5204,N_4764,N_4519);
xnor U5205 (N_5205,N_4022,N_4608);
xor U5206 (N_5206,N_4459,N_4263);
nand U5207 (N_5207,N_4559,N_4687);
nand U5208 (N_5208,N_4063,N_4502);
or U5209 (N_5209,N_4784,N_4360);
xor U5210 (N_5210,N_4357,N_4089);
xnor U5211 (N_5211,N_4536,N_4433);
nor U5212 (N_5212,N_4541,N_4416);
and U5213 (N_5213,N_4173,N_4215);
or U5214 (N_5214,N_4602,N_4788);
and U5215 (N_5215,N_4583,N_4527);
or U5216 (N_5216,N_4778,N_4216);
xor U5217 (N_5217,N_4045,N_4461);
nor U5218 (N_5218,N_4700,N_4007);
and U5219 (N_5219,N_4238,N_4712);
or U5220 (N_5220,N_4336,N_4782);
xnor U5221 (N_5221,N_4540,N_4146);
nor U5222 (N_5222,N_4299,N_4428);
nor U5223 (N_5223,N_4401,N_4448);
or U5224 (N_5224,N_4214,N_4639);
xnor U5225 (N_5225,N_4140,N_4166);
or U5226 (N_5226,N_4344,N_4421);
nor U5227 (N_5227,N_4402,N_4388);
nor U5228 (N_5228,N_4352,N_4454);
xnor U5229 (N_5229,N_4290,N_4701);
or U5230 (N_5230,N_4455,N_4534);
xor U5231 (N_5231,N_4133,N_4118);
nor U5232 (N_5232,N_4307,N_4791);
nand U5233 (N_5233,N_4276,N_4649);
or U5234 (N_5234,N_4739,N_4367);
and U5235 (N_5235,N_4518,N_4014);
and U5236 (N_5236,N_4065,N_4508);
or U5237 (N_5237,N_4350,N_4011);
nand U5238 (N_5238,N_4017,N_4580);
and U5239 (N_5239,N_4771,N_4711);
or U5240 (N_5240,N_4285,N_4061);
nor U5241 (N_5241,N_4623,N_4577);
and U5242 (N_5242,N_4509,N_4474);
xor U5243 (N_5243,N_4392,N_4229);
nor U5244 (N_5244,N_4666,N_4675);
xor U5245 (N_5245,N_4695,N_4550);
nor U5246 (N_5246,N_4286,N_4776);
nor U5247 (N_5247,N_4380,N_4279);
xnor U5248 (N_5248,N_4137,N_4236);
xnor U5249 (N_5249,N_4394,N_4473);
xor U5250 (N_5250,N_4680,N_4619);
and U5251 (N_5251,N_4465,N_4569);
nor U5252 (N_5252,N_4023,N_4189);
xnor U5253 (N_5253,N_4444,N_4595);
xor U5254 (N_5254,N_4145,N_4173);
xnor U5255 (N_5255,N_4110,N_4740);
xnor U5256 (N_5256,N_4384,N_4549);
or U5257 (N_5257,N_4427,N_4458);
and U5258 (N_5258,N_4067,N_4614);
xnor U5259 (N_5259,N_4188,N_4513);
nand U5260 (N_5260,N_4718,N_4298);
nor U5261 (N_5261,N_4267,N_4390);
xnor U5262 (N_5262,N_4798,N_4616);
nand U5263 (N_5263,N_4149,N_4250);
and U5264 (N_5264,N_4122,N_4557);
nand U5265 (N_5265,N_4374,N_4474);
nor U5266 (N_5266,N_4575,N_4093);
nor U5267 (N_5267,N_4592,N_4634);
xor U5268 (N_5268,N_4326,N_4215);
nand U5269 (N_5269,N_4642,N_4397);
or U5270 (N_5270,N_4182,N_4409);
xnor U5271 (N_5271,N_4496,N_4688);
or U5272 (N_5272,N_4421,N_4624);
nor U5273 (N_5273,N_4229,N_4200);
xor U5274 (N_5274,N_4114,N_4551);
nor U5275 (N_5275,N_4065,N_4229);
or U5276 (N_5276,N_4799,N_4378);
xnor U5277 (N_5277,N_4405,N_4428);
xor U5278 (N_5278,N_4278,N_4732);
or U5279 (N_5279,N_4471,N_4179);
nand U5280 (N_5280,N_4416,N_4371);
nor U5281 (N_5281,N_4659,N_4499);
nor U5282 (N_5282,N_4263,N_4260);
or U5283 (N_5283,N_4343,N_4586);
and U5284 (N_5284,N_4456,N_4489);
and U5285 (N_5285,N_4430,N_4644);
or U5286 (N_5286,N_4469,N_4787);
nor U5287 (N_5287,N_4681,N_4031);
nand U5288 (N_5288,N_4319,N_4164);
nand U5289 (N_5289,N_4146,N_4638);
and U5290 (N_5290,N_4766,N_4424);
nand U5291 (N_5291,N_4500,N_4665);
xor U5292 (N_5292,N_4619,N_4530);
xor U5293 (N_5293,N_4595,N_4236);
xor U5294 (N_5294,N_4628,N_4159);
xnor U5295 (N_5295,N_4370,N_4337);
nand U5296 (N_5296,N_4037,N_4241);
xor U5297 (N_5297,N_4594,N_4393);
nor U5298 (N_5298,N_4707,N_4264);
or U5299 (N_5299,N_4547,N_4178);
xnor U5300 (N_5300,N_4484,N_4391);
nor U5301 (N_5301,N_4009,N_4663);
and U5302 (N_5302,N_4713,N_4675);
or U5303 (N_5303,N_4716,N_4472);
or U5304 (N_5304,N_4383,N_4268);
nand U5305 (N_5305,N_4014,N_4396);
nand U5306 (N_5306,N_4635,N_4055);
nor U5307 (N_5307,N_4436,N_4665);
or U5308 (N_5308,N_4008,N_4654);
and U5309 (N_5309,N_4446,N_4344);
or U5310 (N_5310,N_4450,N_4132);
and U5311 (N_5311,N_4689,N_4107);
nor U5312 (N_5312,N_4400,N_4763);
nand U5313 (N_5313,N_4341,N_4127);
xnor U5314 (N_5314,N_4151,N_4365);
nor U5315 (N_5315,N_4634,N_4418);
and U5316 (N_5316,N_4112,N_4610);
nand U5317 (N_5317,N_4247,N_4685);
nand U5318 (N_5318,N_4377,N_4573);
or U5319 (N_5319,N_4263,N_4340);
xnor U5320 (N_5320,N_4512,N_4352);
nor U5321 (N_5321,N_4234,N_4225);
or U5322 (N_5322,N_4528,N_4640);
or U5323 (N_5323,N_4579,N_4201);
nor U5324 (N_5324,N_4723,N_4473);
nor U5325 (N_5325,N_4024,N_4402);
and U5326 (N_5326,N_4149,N_4175);
nor U5327 (N_5327,N_4797,N_4177);
nand U5328 (N_5328,N_4721,N_4131);
xor U5329 (N_5329,N_4306,N_4563);
nor U5330 (N_5330,N_4371,N_4781);
nor U5331 (N_5331,N_4321,N_4437);
or U5332 (N_5332,N_4563,N_4353);
xnor U5333 (N_5333,N_4477,N_4633);
and U5334 (N_5334,N_4574,N_4444);
nand U5335 (N_5335,N_4314,N_4312);
or U5336 (N_5336,N_4542,N_4769);
xnor U5337 (N_5337,N_4690,N_4739);
nor U5338 (N_5338,N_4355,N_4460);
nor U5339 (N_5339,N_4445,N_4268);
nor U5340 (N_5340,N_4397,N_4775);
or U5341 (N_5341,N_4638,N_4493);
or U5342 (N_5342,N_4085,N_4469);
or U5343 (N_5343,N_4139,N_4661);
xor U5344 (N_5344,N_4164,N_4180);
and U5345 (N_5345,N_4379,N_4381);
xnor U5346 (N_5346,N_4280,N_4668);
xnor U5347 (N_5347,N_4315,N_4241);
nor U5348 (N_5348,N_4791,N_4652);
nand U5349 (N_5349,N_4279,N_4250);
nor U5350 (N_5350,N_4247,N_4293);
and U5351 (N_5351,N_4732,N_4004);
nor U5352 (N_5352,N_4307,N_4426);
xor U5353 (N_5353,N_4632,N_4072);
and U5354 (N_5354,N_4284,N_4491);
nor U5355 (N_5355,N_4447,N_4495);
or U5356 (N_5356,N_4402,N_4110);
or U5357 (N_5357,N_4386,N_4050);
or U5358 (N_5358,N_4528,N_4334);
nand U5359 (N_5359,N_4054,N_4647);
nand U5360 (N_5360,N_4140,N_4429);
and U5361 (N_5361,N_4015,N_4549);
or U5362 (N_5362,N_4761,N_4799);
nor U5363 (N_5363,N_4607,N_4428);
nor U5364 (N_5364,N_4070,N_4195);
xor U5365 (N_5365,N_4570,N_4373);
and U5366 (N_5366,N_4109,N_4613);
nand U5367 (N_5367,N_4725,N_4322);
nand U5368 (N_5368,N_4787,N_4300);
nor U5369 (N_5369,N_4566,N_4424);
nor U5370 (N_5370,N_4414,N_4126);
nand U5371 (N_5371,N_4191,N_4407);
or U5372 (N_5372,N_4668,N_4289);
nand U5373 (N_5373,N_4521,N_4248);
nor U5374 (N_5374,N_4230,N_4537);
and U5375 (N_5375,N_4178,N_4093);
xor U5376 (N_5376,N_4221,N_4525);
nand U5377 (N_5377,N_4312,N_4001);
nand U5378 (N_5378,N_4136,N_4694);
nand U5379 (N_5379,N_4230,N_4505);
nand U5380 (N_5380,N_4186,N_4406);
and U5381 (N_5381,N_4244,N_4650);
nor U5382 (N_5382,N_4297,N_4043);
and U5383 (N_5383,N_4560,N_4022);
xor U5384 (N_5384,N_4422,N_4626);
and U5385 (N_5385,N_4111,N_4487);
and U5386 (N_5386,N_4437,N_4275);
and U5387 (N_5387,N_4274,N_4199);
nand U5388 (N_5388,N_4025,N_4793);
and U5389 (N_5389,N_4046,N_4795);
or U5390 (N_5390,N_4221,N_4342);
and U5391 (N_5391,N_4303,N_4225);
nand U5392 (N_5392,N_4313,N_4467);
or U5393 (N_5393,N_4090,N_4343);
nand U5394 (N_5394,N_4355,N_4117);
nor U5395 (N_5395,N_4064,N_4128);
or U5396 (N_5396,N_4130,N_4574);
nor U5397 (N_5397,N_4649,N_4081);
xor U5398 (N_5398,N_4234,N_4418);
or U5399 (N_5399,N_4454,N_4106);
xnor U5400 (N_5400,N_4381,N_4224);
and U5401 (N_5401,N_4253,N_4129);
or U5402 (N_5402,N_4166,N_4494);
xor U5403 (N_5403,N_4586,N_4341);
nand U5404 (N_5404,N_4362,N_4548);
xnor U5405 (N_5405,N_4404,N_4125);
and U5406 (N_5406,N_4486,N_4360);
and U5407 (N_5407,N_4036,N_4514);
and U5408 (N_5408,N_4556,N_4139);
xnor U5409 (N_5409,N_4422,N_4394);
nand U5410 (N_5410,N_4319,N_4336);
or U5411 (N_5411,N_4147,N_4282);
and U5412 (N_5412,N_4290,N_4088);
or U5413 (N_5413,N_4636,N_4348);
or U5414 (N_5414,N_4213,N_4330);
and U5415 (N_5415,N_4628,N_4583);
and U5416 (N_5416,N_4126,N_4505);
nand U5417 (N_5417,N_4549,N_4684);
xnor U5418 (N_5418,N_4186,N_4404);
nor U5419 (N_5419,N_4036,N_4760);
nand U5420 (N_5420,N_4118,N_4664);
and U5421 (N_5421,N_4180,N_4002);
nand U5422 (N_5422,N_4190,N_4562);
xnor U5423 (N_5423,N_4185,N_4115);
or U5424 (N_5424,N_4378,N_4387);
xnor U5425 (N_5425,N_4620,N_4253);
nor U5426 (N_5426,N_4590,N_4483);
or U5427 (N_5427,N_4031,N_4527);
or U5428 (N_5428,N_4083,N_4622);
and U5429 (N_5429,N_4065,N_4620);
xnor U5430 (N_5430,N_4515,N_4181);
and U5431 (N_5431,N_4345,N_4193);
nor U5432 (N_5432,N_4430,N_4189);
and U5433 (N_5433,N_4003,N_4320);
nor U5434 (N_5434,N_4411,N_4722);
or U5435 (N_5435,N_4245,N_4575);
or U5436 (N_5436,N_4041,N_4726);
nand U5437 (N_5437,N_4489,N_4743);
or U5438 (N_5438,N_4332,N_4058);
nand U5439 (N_5439,N_4236,N_4083);
nand U5440 (N_5440,N_4303,N_4656);
nand U5441 (N_5441,N_4642,N_4053);
xor U5442 (N_5442,N_4554,N_4499);
nor U5443 (N_5443,N_4748,N_4458);
and U5444 (N_5444,N_4065,N_4547);
and U5445 (N_5445,N_4023,N_4005);
nand U5446 (N_5446,N_4166,N_4124);
and U5447 (N_5447,N_4437,N_4395);
nand U5448 (N_5448,N_4120,N_4504);
nor U5449 (N_5449,N_4228,N_4259);
nand U5450 (N_5450,N_4036,N_4788);
or U5451 (N_5451,N_4421,N_4573);
and U5452 (N_5452,N_4458,N_4038);
nand U5453 (N_5453,N_4372,N_4023);
or U5454 (N_5454,N_4787,N_4283);
xor U5455 (N_5455,N_4266,N_4411);
and U5456 (N_5456,N_4047,N_4150);
and U5457 (N_5457,N_4155,N_4483);
nand U5458 (N_5458,N_4114,N_4144);
nor U5459 (N_5459,N_4728,N_4639);
xnor U5460 (N_5460,N_4526,N_4447);
and U5461 (N_5461,N_4479,N_4750);
xnor U5462 (N_5462,N_4263,N_4393);
xnor U5463 (N_5463,N_4077,N_4641);
and U5464 (N_5464,N_4760,N_4663);
or U5465 (N_5465,N_4141,N_4146);
or U5466 (N_5466,N_4345,N_4249);
or U5467 (N_5467,N_4776,N_4424);
nand U5468 (N_5468,N_4150,N_4347);
and U5469 (N_5469,N_4691,N_4784);
or U5470 (N_5470,N_4197,N_4522);
xor U5471 (N_5471,N_4718,N_4777);
and U5472 (N_5472,N_4027,N_4640);
nor U5473 (N_5473,N_4786,N_4115);
nand U5474 (N_5474,N_4262,N_4734);
or U5475 (N_5475,N_4297,N_4519);
or U5476 (N_5476,N_4071,N_4180);
nand U5477 (N_5477,N_4622,N_4772);
nand U5478 (N_5478,N_4696,N_4368);
and U5479 (N_5479,N_4305,N_4567);
nand U5480 (N_5480,N_4225,N_4614);
and U5481 (N_5481,N_4679,N_4608);
or U5482 (N_5482,N_4471,N_4752);
xnor U5483 (N_5483,N_4491,N_4738);
nor U5484 (N_5484,N_4127,N_4542);
and U5485 (N_5485,N_4238,N_4494);
and U5486 (N_5486,N_4774,N_4158);
or U5487 (N_5487,N_4572,N_4069);
nand U5488 (N_5488,N_4111,N_4478);
nand U5489 (N_5489,N_4016,N_4603);
nor U5490 (N_5490,N_4238,N_4011);
and U5491 (N_5491,N_4699,N_4208);
or U5492 (N_5492,N_4657,N_4453);
nor U5493 (N_5493,N_4435,N_4340);
xor U5494 (N_5494,N_4111,N_4293);
or U5495 (N_5495,N_4018,N_4523);
xor U5496 (N_5496,N_4442,N_4075);
and U5497 (N_5497,N_4237,N_4494);
and U5498 (N_5498,N_4210,N_4120);
nand U5499 (N_5499,N_4532,N_4487);
or U5500 (N_5500,N_4656,N_4481);
nand U5501 (N_5501,N_4217,N_4068);
nor U5502 (N_5502,N_4531,N_4386);
nand U5503 (N_5503,N_4427,N_4640);
and U5504 (N_5504,N_4497,N_4566);
xnor U5505 (N_5505,N_4040,N_4199);
nand U5506 (N_5506,N_4080,N_4505);
xor U5507 (N_5507,N_4417,N_4366);
xnor U5508 (N_5508,N_4518,N_4797);
and U5509 (N_5509,N_4114,N_4542);
nor U5510 (N_5510,N_4008,N_4627);
nand U5511 (N_5511,N_4061,N_4233);
nand U5512 (N_5512,N_4595,N_4287);
nand U5513 (N_5513,N_4695,N_4324);
nand U5514 (N_5514,N_4158,N_4751);
or U5515 (N_5515,N_4413,N_4083);
or U5516 (N_5516,N_4319,N_4474);
or U5517 (N_5517,N_4397,N_4543);
or U5518 (N_5518,N_4676,N_4376);
nand U5519 (N_5519,N_4482,N_4110);
or U5520 (N_5520,N_4587,N_4340);
xnor U5521 (N_5521,N_4105,N_4132);
nor U5522 (N_5522,N_4485,N_4163);
or U5523 (N_5523,N_4116,N_4475);
nor U5524 (N_5524,N_4273,N_4530);
or U5525 (N_5525,N_4222,N_4219);
nand U5526 (N_5526,N_4422,N_4702);
nor U5527 (N_5527,N_4604,N_4241);
or U5528 (N_5528,N_4292,N_4276);
and U5529 (N_5529,N_4732,N_4055);
nor U5530 (N_5530,N_4273,N_4480);
and U5531 (N_5531,N_4704,N_4090);
and U5532 (N_5532,N_4259,N_4288);
or U5533 (N_5533,N_4209,N_4276);
and U5534 (N_5534,N_4132,N_4359);
nand U5535 (N_5535,N_4490,N_4785);
or U5536 (N_5536,N_4164,N_4158);
and U5537 (N_5537,N_4773,N_4185);
xor U5538 (N_5538,N_4197,N_4034);
nor U5539 (N_5539,N_4666,N_4465);
nor U5540 (N_5540,N_4673,N_4055);
or U5541 (N_5541,N_4349,N_4617);
xnor U5542 (N_5542,N_4426,N_4637);
xnor U5543 (N_5543,N_4118,N_4531);
nor U5544 (N_5544,N_4185,N_4542);
or U5545 (N_5545,N_4481,N_4477);
xor U5546 (N_5546,N_4703,N_4387);
nand U5547 (N_5547,N_4415,N_4707);
or U5548 (N_5548,N_4381,N_4388);
nor U5549 (N_5549,N_4781,N_4749);
xnor U5550 (N_5550,N_4537,N_4370);
and U5551 (N_5551,N_4319,N_4491);
and U5552 (N_5552,N_4721,N_4555);
and U5553 (N_5553,N_4261,N_4427);
nor U5554 (N_5554,N_4454,N_4317);
or U5555 (N_5555,N_4375,N_4736);
or U5556 (N_5556,N_4787,N_4176);
or U5557 (N_5557,N_4750,N_4351);
and U5558 (N_5558,N_4368,N_4054);
or U5559 (N_5559,N_4358,N_4342);
nor U5560 (N_5560,N_4099,N_4267);
nand U5561 (N_5561,N_4693,N_4675);
or U5562 (N_5562,N_4485,N_4696);
or U5563 (N_5563,N_4132,N_4442);
and U5564 (N_5564,N_4663,N_4205);
and U5565 (N_5565,N_4071,N_4700);
or U5566 (N_5566,N_4495,N_4367);
or U5567 (N_5567,N_4497,N_4575);
and U5568 (N_5568,N_4603,N_4167);
and U5569 (N_5569,N_4680,N_4119);
xor U5570 (N_5570,N_4753,N_4682);
nor U5571 (N_5571,N_4509,N_4396);
nor U5572 (N_5572,N_4560,N_4661);
nand U5573 (N_5573,N_4155,N_4306);
xor U5574 (N_5574,N_4410,N_4760);
or U5575 (N_5575,N_4444,N_4722);
nor U5576 (N_5576,N_4364,N_4772);
xor U5577 (N_5577,N_4541,N_4695);
nor U5578 (N_5578,N_4521,N_4049);
or U5579 (N_5579,N_4079,N_4718);
xnor U5580 (N_5580,N_4097,N_4714);
or U5581 (N_5581,N_4525,N_4392);
xor U5582 (N_5582,N_4388,N_4354);
and U5583 (N_5583,N_4000,N_4735);
and U5584 (N_5584,N_4663,N_4295);
or U5585 (N_5585,N_4030,N_4453);
and U5586 (N_5586,N_4256,N_4383);
nor U5587 (N_5587,N_4796,N_4562);
or U5588 (N_5588,N_4231,N_4595);
xnor U5589 (N_5589,N_4061,N_4406);
xor U5590 (N_5590,N_4148,N_4348);
nor U5591 (N_5591,N_4197,N_4621);
or U5592 (N_5592,N_4194,N_4443);
nor U5593 (N_5593,N_4243,N_4428);
nor U5594 (N_5594,N_4103,N_4010);
nand U5595 (N_5595,N_4633,N_4075);
nor U5596 (N_5596,N_4011,N_4393);
xnor U5597 (N_5597,N_4446,N_4242);
xor U5598 (N_5598,N_4459,N_4078);
or U5599 (N_5599,N_4716,N_4517);
and U5600 (N_5600,N_4911,N_5112);
xor U5601 (N_5601,N_5523,N_5336);
and U5602 (N_5602,N_4968,N_5207);
xor U5603 (N_5603,N_5076,N_5242);
xor U5604 (N_5604,N_4969,N_5331);
xnor U5605 (N_5605,N_5261,N_5543);
xor U5606 (N_5606,N_5103,N_5153);
xnor U5607 (N_5607,N_5577,N_4996);
or U5608 (N_5608,N_5193,N_4925);
or U5609 (N_5609,N_5503,N_5197);
nand U5610 (N_5610,N_4880,N_5075);
xnor U5611 (N_5611,N_5200,N_5254);
nor U5612 (N_5612,N_4932,N_5087);
xor U5613 (N_5613,N_5005,N_4975);
and U5614 (N_5614,N_5284,N_4833);
and U5615 (N_5615,N_5533,N_4820);
xor U5616 (N_5616,N_4887,N_5055);
nor U5617 (N_5617,N_5220,N_4971);
or U5618 (N_5618,N_5249,N_5451);
nand U5619 (N_5619,N_5157,N_5108);
or U5620 (N_5620,N_4940,N_5552);
nand U5621 (N_5621,N_5329,N_4837);
or U5622 (N_5622,N_4857,N_5561);
nor U5623 (N_5623,N_5148,N_4898);
xor U5624 (N_5624,N_5401,N_5469);
or U5625 (N_5625,N_5456,N_4965);
and U5626 (N_5626,N_5216,N_5045);
nor U5627 (N_5627,N_5212,N_5363);
and U5628 (N_5628,N_5548,N_5500);
xor U5629 (N_5629,N_5333,N_5154);
xnor U5630 (N_5630,N_5489,N_4856);
nor U5631 (N_5631,N_4816,N_5366);
nor U5632 (N_5632,N_5051,N_5074);
and U5633 (N_5633,N_5155,N_5360);
nand U5634 (N_5634,N_5210,N_5019);
nor U5635 (N_5635,N_4984,N_4990);
xnor U5636 (N_5636,N_4950,N_5495);
xnor U5637 (N_5637,N_5462,N_5537);
nand U5638 (N_5638,N_4846,N_4877);
and U5639 (N_5639,N_5166,N_5115);
or U5640 (N_5640,N_5560,N_4876);
nor U5641 (N_5641,N_4888,N_5158);
xnor U5642 (N_5642,N_5371,N_5128);
nand U5643 (N_5643,N_5341,N_5185);
nand U5644 (N_5644,N_5584,N_5117);
and U5645 (N_5645,N_5407,N_5000);
or U5646 (N_5646,N_5099,N_4946);
or U5647 (N_5647,N_5342,N_4811);
or U5648 (N_5648,N_5109,N_5189);
and U5649 (N_5649,N_4981,N_5149);
and U5650 (N_5650,N_5361,N_5289);
or U5651 (N_5651,N_5237,N_4802);
or U5652 (N_5652,N_5224,N_5301);
and U5653 (N_5653,N_5060,N_5332);
nand U5654 (N_5654,N_5250,N_5195);
xor U5655 (N_5655,N_4826,N_4914);
or U5656 (N_5656,N_5505,N_5564);
nand U5657 (N_5657,N_5356,N_5370);
nor U5658 (N_5658,N_5343,N_5377);
nor U5659 (N_5659,N_5473,N_4949);
and U5660 (N_5660,N_4976,N_5424);
and U5661 (N_5661,N_4861,N_5142);
nand U5662 (N_5662,N_4945,N_5047);
or U5663 (N_5663,N_4893,N_5082);
and U5664 (N_5664,N_4869,N_4912);
and U5665 (N_5665,N_5107,N_5399);
and U5666 (N_5666,N_5296,N_5455);
or U5667 (N_5667,N_4921,N_5288);
nor U5668 (N_5668,N_5397,N_4924);
xor U5669 (N_5669,N_5121,N_5202);
or U5670 (N_5670,N_5227,N_4852);
or U5671 (N_5671,N_5590,N_5431);
and U5672 (N_5672,N_5468,N_5429);
and U5673 (N_5673,N_4962,N_5066);
or U5674 (N_5674,N_5144,N_5597);
or U5675 (N_5675,N_5367,N_5072);
or U5676 (N_5676,N_5520,N_5433);
nand U5677 (N_5677,N_5257,N_5209);
and U5678 (N_5678,N_5172,N_5002);
or U5679 (N_5679,N_5165,N_4974);
nor U5680 (N_5680,N_4818,N_5111);
nand U5681 (N_5681,N_4875,N_5280);
nor U5682 (N_5682,N_5358,N_4844);
and U5683 (N_5683,N_4819,N_5547);
nor U5684 (N_5684,N_5252,N_5038);
nor U5685 (N_5685,N_5030,N_5541);
or U5686 (N_5686,N_4885,N_5273);
and U5687 (N_5687,N_5459,N_5521);
nand U5688 (N_5688,N_5088,N_5528);
or U5689 (N_5689,N_4872,N_4943);
nand U5690 (N_5690,N_5302,N_5232);
nor U5691 (N_5691,N_4874,N_5100);
nand U5692 (N_5692,N_4841,N_5398);
and U5693 (N_5693,N_5160,N_5594);
or U5694 (N_5694,N_5392,N_5434);
nand U5695 (N_5695,N_5225,N_5110);
or U5696 (N_5696,N_5316,N_5453);
and U5697 (N_5697,N_4867,N_4805);
xnor U5698 (N_5698,N_5326,N_4983);
xnor U5699 (N_5699,N_4855,N_5023);
or U5700 (N_5700,N_5522,N_5379);
or U5701 (N_5701,N_5294,N_5178);
nand U5702 (N_5702,N_4847,N_4982);
nand U5703 (N_5703,N_5490,N_5499);
xnor U5704 (N_5704,N_5063,N_4956);
or U5705 (N_5705,N_4989,N_4835);
and U5706 (N_5706,N_5069,N_4961);
or U5707 (N_5707,N_4892,N_5491);
xor U5708 (N_5708,N_5458,N_5132);
xnor U5709 (N_5709,N_5238,N_5098);
nand U5710 (N_5710,N_5230,N_4985);
nand U5711 (N_5711,N_5319,N_5595);
xnor U5712 (N_5712,N_5270,N_5324);
xor U5713 (N_5713,N_4955,N_5428);
or U5714 (N_5714,N_5339,N_4870);
or U5715 (N_5715,N_5576,N_5559);
or U5716 (N_5716,N_5420,N_5068);
nor U5717 (N_5717,N_5174,N_5152);
or U5718 (N_5718,N_4958,N_4938);
or U5719 (N_5719,N_5134,N_4913);
xor U5720 (N_5720,N_5347,N_5381);
xor U5721 (N_5721,N_4879,N_5496);
nand U5722 (N_5722,N_5018,N_4947);
or U5723 (N_5723,N_5192,N_5555);
xnor U5724 (N_5724,N_5592,N_5418);
nor U5725 (N_5725,N_5309,N_5081);
nand U5726 (N_5726,N_5394,N_5513);
and U5727 (N_5727,N_4941,N_5508);
xor U5728 (N_5728,N_5162,N_4840);
nor U5729 (N_5729,N_4928,N_5168);
or U5730 (N_5730,N_5359,N_5039);
and U5731 (N_5731,N_5125,N_5373);
nor U5732 (N_5732,N_5218,N_5263);
and U5733 (N_5733,N_5536,N_5461);
xor U5734 (N_5734,N_4908,N_4917);
nand U5735 (N_5735,N_5553,N_5599);
or U5736 (N_5736,N_4922,N_4882);
and U5737 (N_5737,N_5444,N_5223);
and U5738 (N_5738,N_5322,N_5408);
xnor U5739 (N_5739,N_5426,N_5268);
and U5740 (N_5740,N_5567,N_5078);
nor U5741 (N_5741,N_5372,N_5544);
nor U5742 (N_5742,N_5501,N_4829);
or U5743 (N_5743,N_5486,N_5146);
or U5744 (N_5744,N_4979,N_5147);
or U5745 (N_5745,N_4873,N_5390);
nand U5746 (N_5746,N_5485,N_5044);
nand U5747 (N_5747,N_4902,N_5291);
xor U5748 (N_5748,N_5382,N_5572);
nand U5749 (N_5749,N_5518,N_5042);
nand U5750 (N_5750,N_5565,N_5582);
and U5751 (N_5751,N_5150,N_4825);
or U5752 (N_5752,N_5163,N_5395);
xor U5753 (N_5753,N_5140,N_4814);
nand U5754 (N_5754,N_5413,N_5452);
xor U5755 (N_5755,N_5557,N_5457);
or U5756 (N_5756,N_5446,N_5182);
xnor U5757 (N_5757,N_4871,N_5101);
or U5758 (N_5758,N_4904,N_5450);
or U5759 (N_5759,N_4848,N_5277);
xnor U5760 (N_5760,N_5416,N_5568);
nand U5761 (N_5761,N_4994,N_5028);
xor U5762 (N_5762,N_4963,N_5037);
nor U5763 (N_5763,N_4959,N_5040);
and U5764 (N_5764,N_5169,N_5306);
xnor U5765 (N_5765,N_5131,N_5233);
and U5766 (N_5766,N_5205,N_5526);
or U5767 (N_5767,N_4832,N_5315);
nor U5768 (N_5768,N_4830,N_4973);
xnor U5769 (N_5769,N_5587,N_5550);
or U5770 (N_5770,N_5244,N_4986);
nor U5771 (N_5771,N_5164,N_5048);
or U5772 (N_5772,N_5012,N_5464);
nor U5773 (N_5773,N_5092,N_5506);
nand U5774 (N_5774,N_5203,N_5046);
xnor U5775 (N_5775,N_5036,N_5504);
nor U5776 (N_5776,N_5303,N_5391);
xor U5777 (N_5777,N_4894,N_5575);
or U5778 (N_5778,N_5586,N_5402);
or U5779 (N_5779,N_4839,N_4838);
xor U5780 (N_5780,N_5034,N_5542);
and U5781 (N_5781,N_5096,N_5293);
xnor U5782 (N_5782,N_4987,N_5380);
and U5783 (N_5783,N_5143,N_4891);
xor U5784 (N_5784,N_5090,N_5033);
nand U5785 (N_5785,N_5383,N_4907);
xor U5786 (N_5786,N_5267,N_5440);
xnor U5787 (N_5787,N_4850,N_5474);
nor U5788 (N_5788,N_5001,N_5449);
nand U5789 (N_5789,N_5460,N_4849);
nand U5790 (N_5790,N_5569,N_4853);
nor U5791 (N_5791,N_5472,N_5014);
xnor U5792 (N_5792,N_5351,N_4999);
or U5793 (N_5793,N_5077,N_4881);
or U5794 (N_5794,N_4886,N_5581);
and U5795 (N_5795,N_5053,N_5246);
and U5796 (N_5796,N_5409,N_4923);
xnor U5797 (N_5797,N_4851,N_5255);
or U5798 (N_5798,N_5405,N_5259);
and U5799 (N_5799,N_5320,N_5475);
nand U5800 (N_5800,N_5532,N_5260);
and U5801 (N_5801,N_5419,N_5578);
nor U5802 (N_5802,N_4890,N_5126);
nor U5803 (N_5803,N_5340,N_5421);
xor U5804 (N_5804,N_4821,N_4942);
nand U5805 (N_5805,N_4931,N_5050);
or U5806 (N_5806,N_4952,N_5512);
xor U5807 (N_5807,N_4901,N_5138);
or U5808 (N_5808,N_5171,N_5540);
nor U5809 (N_5809,N_5127,N_4903);
and U5810 (N_5810,N_5064,N_5353);
or U5811 (N_5811,N_5187,N_4823);
or U5812 (N_5812,N_5177,N_5245);
and U5813 (N_5813,N_4980,N_5007);
xnor U5814 (N_5814,N_5269,N_5062);
xor U5815 (N_5815,N_5524,N_5061);
or U5816 (N_5816,N_5129,N_5274);
nand U5817 (N_5817,N_5514,N_5251);
and U5818 (N_5818,N_4930,N_5374);
or U5819 (N_5819,N_5287,N_5105);
nor U5820 (N_5820,N_5412,N_5124);
and U5821 (N_5821,N_5190,N_4906);
nand U5822 (N_5822,N_5215,N_4831);
nor U5823 (N_5823,N_5411,N_5442);
xnor U5824 (N_5824,N_5248,N_4964);
xor U5825 (N_5825,N_5352,N_5511);
nor U5826 (N_5826,N_5235,N_5137);
nor U5827 (N_5827,N_5502,N_4910);
or U5828 (N_5828,N_5525,N_5009);
and U5829 (N_5829,N_5276,N_4883);
nor U5830 (N_5830,N_5243,N_5222);
nand U5831 (N_5831,N_5079,N_4977);
nor U5832 (N_5832,N_5275,N_5299);
nor U5833 (N_5833,N_5545,N_5551);
nand U5834 (N_5834,N_5049,N_4843);
or U5835 (N_5835,N_5441,N_5228);
xor U5836 (N_5836,N_4935,N_5015);
or U5837 (N_5837,N_5016,N_4936);
xnor U5838 (N_5838,N_5181,N_5167);
nor U5839 (N_5839,N_5297,N_5184);
xnor U5840 (N_5840,N_5029,N_5354);
and U5841 (N_5841,N_5487,N_5318);
or U5842 (N_5842,N_4951,N_5089);
or U5843 (N_5843,N_5241,N_5067);
nand U5844 (N_5844,N_5476,N_5211);
or U5845 (N_5845,N_5314,N_5151);
or U5846 (N_5846,N_5104,N_5338);
nand U5847 (N_5847,N_5396,N_4813);
and U5848 (N_5848,N_4859,N_4939);
or U5849 (N_5849,N_5334,N_5488);
xor U5850 (N_5850,N_4868,N_5546);
xnor U5851 (N_5851,N_5083,N_5482);
and U5852 (N_5852,N_4812,N_5304);
nand U5853 (N_5853,N_5425,N_5563);
and U5854 (N_5854,N_5020,N_5493);
and U5855 (N_5855,N_5427,N_4926);
and U5856 (N_5856,N_5510,N_5004);
nor U5857 (N_5857,N_5264,N_5170);
xnor U5858 (N_5858,N_5346,N_4953);
and U5859 (N_5859,N_5400,N_4834);
xnor U5860 (N_5860,N_5011,N_5364);
nand U5861 (N_5861,N_5198,N_5549);
nand U5862 (N_5862,N_5097,N_5204);
xnor U5863 (N_5863,N_5286,N_5480);
nor U5864 (N_5864,N_5355,N_5059);
nor U5865 (N_5865,N_5311,N_5466);
and U5866 (N_5866,N_5122,N_5335);
and U5867 (N_5867,N_4933,N_5133);
xor U5868 (N_5868,N_5021,N_5070);
xor U5869 (N_5869,N_5350,N_4920);
or U5870 (N_5870,N_5041,N_5369);
xnor U5871 (N_5871,N_5139,N_4864);
or U5872 (N_5872,N_4817,N_5135);
nand U5873 (N_5873,N_4858,N_5556);
and U5874 (N_5874,N_5598,N_5173);
xnor U5875 (N_5875,N_5196,N_5481);
and U5876 (N_5876,N_5305,N_5432);
nand U5877 (N_5877,N_5256,N_5345);
or U5878 (N_5878,N_5516,N_5471);
xor U5879 (N_5879,N_4916,N_4998);
xor U5880 (N_5880,N_5362,N_5136);
nand U5881 (N_5881,N_5517,N_5120);
nand U5882 (N_5882,N_5114,N_4865);
and U5883 (N_5883,N_4884,N_5337);
nand U5884 (N_5884,N_5531,N_5357);
nand U5885 (N_5885,N_5365,N_5253);
or U5886 (N_5886,N_5562,N_5217);
xnor U5887 (N_5887,N_5199,N_5239);
or U5888 (N_5888,N_5031,N_5262);
nor U5889 (N_5889,N_4957,N_5272);
xnor U5890 (N_5890,N_5093,N_5247);
nor U5891 (N_5891,N_5194,N_5116);
and U5892 (N_5892,N_5013,N_5483);
nor U5893 (N_5893,N_5465,N_5593);
nor U5894 (N_5894,N_5509,N_5386);
or U5895 (N_5895,N_4878,N_4827);
or U5896 (N_5896,N_5266,N_5539);
or U5897 (N_5897,N_5387,N_5085);
and U5898 (N_5898,N_5574,N_5388);
or U5899 (N_5899,N_5447,N_4960);
and U5900 (N_5900,N_4895,N_5571);
or U5901 (N_5901,N_4809,N_5058);
nor U5902 (N_5902,N_4948,N_5443);
or U5903 (N_5903,N_4966,N_4866);
nor U5904 (N_5904,N_5589,N_5430);
nand U5905 (N_5905,N_4970,N_5032);
nor U5906 (N_5906,N_4992,N_5348);
or U5907 (N_5907,N_4929,N_4995);
or U5908 (N_5908,N_4927,N_5484);
and U5909 (N_5909,N_5206,N_5529);
nand U5910 (N_5910,N_4919,N_5145);
or U5911 (N_5911,N_4824,N_5179);
and U5912 (N_5912,N_4808,N_5498);
or U5913 (N_5913,N_5024,N_5435);
nor U5914 (N_5914,N_4803,N_5006);
nand U5915 (N_5915,N_5438,N_4897);
and U5916 (N_5916,N_4822,N_5414);
nand U5917 (N_5917,N_5330,N_5588);
nor U5918 (N_5918,N_4810,N_5208);
nor U5919 (N_5919,N_5494,N_5519);
or U5920 (N_5920,N_5214,N_4896);
nor U5921 (N_5921,N_5393,N_4806);
nor U5922 (N_5922,N_4900,N_5384);
xor U5923 (N_5923,N_5527,N_4978);
and U5924 (N_5924,N_5043,N_5492);
nand U5925 (N_5925,N_5180,N_5156);
nand U5926 (N_5926,N_4815,N_5389);
or U5927 (N_5927,N_4807,N_5035);
nor U5928 (N_5928,N_5095,N_4905);
or U5929 (N_5929,N_5535,N_5327);
and U5930 (N_5930,N_4915,N_5213);
or U5931 (N_5931,N_5056,N_5317);
xor U5932 (N_5932,N_5478,N_5344);
nor U5933 (N_5933,N_5403,N_5295);
nand U5934 (N_5934,N_5566,N_4944);
nand U5935 (N_5935,N_5530,N_5583);
xnor U5936 (N_5936,N_5191,N_5176);
and U5937 (N_5937,N_4842,N_5313);
and U5938 (N_5938,N_4828,N_5422);
and U5939 (N_5939,N_5448,N_4997);
nor U5940 (N_5940,N_5017,N_5123);
nand U5941 (N_5941,N_5570,N_5368);
nand U5942 (N_5942,N_5071,N_5236);
nand U5943 (N_5943,N_5065,N_5376);
and U5944 (N_5944,N_5579,N_5282);
nor U5945 (N_5945,N_5008,N_5445);
or U5946 (N_5946,N_4854,N_5175);
xor U5947 (N_5947,N_5080,N_5410);
nor U5948 (N_5948,N_5406,N_4972);
nor U5949 (N_5949,N_5308,N_5054);
and U5950 (N_5950,N_5229,N_5307);
and U5951 (N_5951,N_5094,N_5188);
and U5952 (N_5952,N_4845,N_4967);
and U5953 (N_5953,N_5201,N_5477);
and U5954 (N_5954,N_5404,N_5423);
xor U5955 (N_5955,N_5310,N_5349);
nor U5956 (N_5956,N_5415,N_5321);
or U5957 (N_5957,N_5283,N_5436);
xnor U5958 (N_5958,N_5119,N_5507);
or U5959 (N_5959,N_4934,N_4863);
xnor U5960 (N_5960,N_5596,N_5554);
nor U5961 (N_5961,N_5534,N_5323);
xnor U5962 (N_5962,N_5052,N_4993);
or U5963 (N_5963,N_5285,N_4988);
nor U5964 (N_5964,N_5463,N_5221);
xnor U5965 (N_5965,N_5290,N_5219);
and U5966 (N_5966,N_5470,N_5010);
xor U5967 (N_5967,N_5159,N_4909);
and U5968 (N_5968,N_5258,N_5086);
xnor U5969 (N_5969,N_5439,N_5281);
xnor U5970 (N_5970,N_5417,N_5183);
and U5971 (N_5971,N_5106,N_5026);
nor U5972 (N_5972,N_5226,N_5585);
xnor U5973 (N_5973,N_5437,N_4889);
nand U5974 (N_5974,N_5161,N_5385);
nor U5975 (N_5975,N_5073,N_4836);
xnor U5976 (N_5976,N_5378,N_5186);
nand U5977 (N_5977,N_5467,N_5271);
and U5978 (N_5978,N_5591,N_5118);
and U5979 (N_5979,N_5141,N_5298);
or U5980 (N_5980,N_5292,N_5312);
and U5981 (N_5981,N_5454,N_4918);
nand U5982 (N_5982,N_5240,N_5375);
nor U5983 (N_5983,N_5558,N_5325);
nand U5984 (N_5984,N_4937,N_5278);
nor U5985 (N_5985,N_4899,N_5279);
xor U5986 (N_5986,N_5057,N_5497);
nand U5987 (N_5987,N_5113,N_4800);
xnor U5988 (N_5988,N_5091,N_4860);
nand U5989 (N_5989,N_5003,N_5538);
or U5990 (N_5990,N_5479,N_5022);
or U5991 (N_5991,N_5025,N_5084);
or U5992 (N_5992,N_4991,N_5328);
and U5993 (N_5993,N_5573,N_5515);
nor U5994 (N_5994,N_5300,N_5102);
nand U5995 (N_5995,N_5234,N_5265);
xnor U5996 (N_5996,N_5027,N_4801);
xor U5997 (N_5997,N_4862,N_4804);
xor U5998 (N_5998,N_4954,N_5130);
nand U5999 (N_5999,N_5231,N_5580);
or U6000 (N_6000,N_5275,N_5573);
or U6001 (N_6001,N_5196,N_5265);
or U6002 (N_6002,N_5582,N_5020);
nand U6003 (N_6003,N_4878,N_5142);
nor U6004 (N_6004,N_5472,N_5534);
and U6005 (N_6005,N_4869,N_5227);
xor U6006 (N_6006,N_5546,N_5579);
nand U6007 (N_6007,N_4907,N_5059);
or U6008 (N_6008,N_4828,N_4915);
nor U6009 (N_6009,N_5478,N_5125);
xor U6010 (N_6010,N_4941,N_5116);
nand U6011 (N_6011,N_4873,N_5158);
xnor U6012 (N_6012,N_5000,N_4914);
xor U6013 (N_6013,N_5446,N_5434);
or U6014 (N_6014,N_5261,N_4826);
nand U6015 (N_6015,N_5516,N_4864);
nand U6016 (N_6016,N_4812,N_4978);
xor U6017 (N_6017,N_4812,N_4805);
nor U6018 (N_6018,N_5212,N_4931);
nand U6019 (N_6019,N_5015,N_5353);
xor U6020 (N_6020,N_5105,N_5296);
and U6021 (N_6021,N_4874,N_5105);
and U6022 (N_6022,N_5074,N_5089);
xor U6023 (N_6023,N_5562,N_5235);
xnor U6024 (N_6024,N_4952,N_5435);
xor U6025 (N_6025,N_5020,N_5104);
xor U6026 (N_6026,N_4803,N_4886);
and U6027 (N_6027,N_5069,N_5048);
xor U6028 (N_6028,N_5152,N_4982);
and U6029 (N_6029,N_5035,N_5251);
nor U6030 (N_6030,N_5286,N_5597);
nor U6031 (N_6031,N_5113,N_5255);
or U6032 (N_6032,N_4879,N_5482);
xnor U6033 (N_6033,N_4847,N_5041);
or U6034 (N_6034,N_5134,N_5475);
nand U6035 (N_6035,N_5459,N_5077);
nor U6036 (N_6036,N_5387,N_5571);
xor U6037 (N_6037,N_5024,N_5549);
nand U6038 (N_6038,N_5224,N_5135);
or U6039 (N_6039,N_5101,N_5577);
or U6040 (N_6040,N_5094,N_4983);
xor U6041 (N_6041,N_5488,N_5593);
xnor U6042 (N_6042,N_5489,N_5494);
nand U6043 (N_6043,N_4963,N_4878);
or U6044 (N_6044,N_5086,N_5578);
xnor U6045 (N_6045,N_5586,N_5348);
nand U6046 (N_6046,N_5082,N_4871);
xnor U6047 (N_6047,N_5371,N_5303);
or U6048 (N_6048,N_5481,N_5017);
or U6049 (N_6049,N_4926,N_4868);
nand U6050 (N_6050,N_5250,N_5473);
or U6051 (N_6051,N_5261,N_5525);
or U6052 (N_6052,N_4959,N_4998);
nor U6053 (N_6053,N_5150,N_5255);
xor U6054 (N_6054,N_5196,N_5439);
xnor U6055 (N_6055,N_5315,N_5026);
or U6056 (N_6056,N_4908,N_5416);
xor U6057 (N_6057,N_5572,N_4924);
xnor U6058 (N_6058,N_5106,N_4901);
nand U6059 (N_6059,N_5191,N_5059);
and U6060 (N_6060,N_5471,N_5497);
nor U6061 (N_6061,N_4966,N_4814);
nor U6062 (N_6062,N_5229,N_5318);
or U6063 (N_6063,N_5460,N_5059);
nand U6064 (N_6064,N_5000,N_5011);
or U6065 (N_6065,N_4865,N_5179);
and U6066 (N_6066,N_5423,N_5590);
nor U6067 (N_6067,N_4807,N_5225);
nor U6068 (N_6068,N_4856,N_5345);
nand U6069 (N_6069,N_5266,N_5574);
nor U6070 (N_6070,N_5591,N_5490);
and U6071 (N_6071,N_5142,N_4880);
or U6072 (N_6072,N_5485,N_5581);
and U6073 (N_6073,N_5283,N_5301);
xnor U6074 (N_6074,N_5448,N_5424);
xor U6075 (N_6075,N_5151,N_5081);
nor U6076 (N_6076,N_4810,N_5265);
nand U6077 (N_6077,N_5152,N_4897);
nand U6078 (N_6078,N_5406,N_5039);
nand U6079 (N_6079,N_5152,N_5401);
nor U6080 (N_6080,N_4919,N_5460);
nor U6081 (N_6081,N_5270,N_4850);
and U6082 (N_6082,N_5162,N_5396);
nand U6083 (N_6083,N_4978,N_5454);
and U6084 (N_6084,N_4916,N_5593);
or U6085 (N_6085,N_5234,N_5348);
nand U6086 (N_6086,N_5534,N_5184);
nand U6087 (N_6087,N_5353,N_5343);
nor U6088 (N_6088,N_5383,N_5482);
and U6089 (N_6089,N_5258,N_4800);
xor U6090 (N_6090,N_4985,N_5033);
or U6091 (N_6091,N_5270,N_5209);
and U6092 (N_6092,N_5233,N_5182);
nand U6093 (N_6093,N_5529,N_4906);
nand U6094 (N_6094,N_5273,N_5276);
and U6095 (N_6095,N_5507,N_5471);
xor U6096 (N_6096,N_5276,N_4873);
nor U6097 (N_6097,N_5143,N_5467);
nor U6098 (N_6098,N_5543,N_5482);
or U6099 (N_6099,N_5351,N_5559);
or U6100 (N_6100,N_5319,N_5470);
or U6101 (N_6101,N_5111,N_5572);
xnor U6102 (N_6102,N_5374,N_4870);
nand U6103 (N_6103,N_5133,N_4809);
and U6104 (N_6104,N_4869,N_5425);
nor U6105 (N_6105,N_5399,N_4915);
nor U6106 (N_6106,N_5141,N_5144);
xor U6107 (N_6107,N_5410,N_5498);
or U6108 (N_6108,N_5218,N_5577);
and U6109 (N_6109,N_4856,N_5295);
nor U6110 (N_6110,N_5413,N_4847);
nor U6111 (N_6111,N_5097,N_4954);
and U6112 (N_6112,N_4922,N_5176);
or U6113 (N_6113,N_5477,N_5445);
nand U6114 (N_6114,N_4939,N_5112);
and U6115 (N_6115,N_5334,N_4987);
nand U6116 (N_6116,N_5282,N_5196);
or U6117 (N_6117,N_5318,N_5372);
and U6118 (N_6118,N_4838,N_5538);
nor U6119 (N_6119,N_5598,N_5284);
nor U6120 (N_6120,N_5283,N_5377);
nor U6121 (N_6121,N_5203,N_4908);
and U6122 (N_6122,N_4820,N_5119);
xnor U6123 (N_6123,N_5569,N_5518);
or U6124 (N_6124,N_5528,N_5390);
nor U6125 (N_6125,N_5198,N_5227);
nand U6126 (N_6126,N_5307,N_4978);
nor U6127 (N_6127,N_4874,N_5216);
or U6128 (N_6128,N_5339,N_5347);
xnor U6129 (N_6129,N_5475,N_4905);
xnor U6130 (N_6130,N_5045,N_4993);
and U6131 (N_6131,N_5292,N_4922);
or U6132 (N_6132,N_4805,N_5082);
and U6133 (N_6133,N_5056,N_5181);
xnor U6134 (N_6134,N_5340,N_5370);
or U6135 (N_6135,N_5378,N_4871);
and U6136 (N_6136,N_5151,N_4821);
nand U6137 (N_6137,N_4935,N_5387);
nand U6138 (N_6138,N_4950,N_5542);
or U6139 (N_6139,N_4901,N_5274);
nor U6140 (N_6140,N_5170,N_5488);
or U6141 (N_6141,N_4871,N_5521);
nor U6142 (N_6142,N_5262,N_5018);
xnor U6143 (N_6143,N_4964,N_5083);
or U6144 (N_6144,N_5571,N_5436);
or U6145 (N_6145,N_5176,N_5066);
nor U6146 (N_6146,N_5268,N_5269);
and U6147 (N_6147,N_5040,N_4918);
nand U6148 (N_6148,N_4979,N_5071);
nor U6149 (N_6149,N_5039,N_5192);
or U6150 (N_6150,N_5302,N_5376);
nor U6151 (N_6151,N_5596,N_5585);
nand U6152 (N_6152,N_4909,N_4829);
nand U6153 (N_6153,N_5160,N_5464);
and U6154 (N_6154,N_5358,N_5570);
xor U6155 (N_6155,N_5525,N_5501);
or U6156 (N_6156,N_5028,N_5592);
and U6157 (N_6157,N_5470,N_4985);
and U6158 (N_6158,N_5536,N_5446);
or U6159 (N_6159,N_4889,N_5070);
xor U6160 (N_6160,N_5136,N_5108);
or U6161 (N_6161,N_5240,N_5490);
nand U6162 (N_6162,N_4948,N_5237);
nand U6163 (N_6163,N_4919,N_5472);
or U6164 (N_6164,N_5291,N_5126);
and U6165 (N_6165,N_5214,N_5346);
nor U6166 (N_6166,N_5433,N_4973);
nor U6167 (N_6167,N_5003,N_4999);
nand U6168 (N_6168,N_5596,N_4993);
or U6169 (N_6169,N_5342,N_5006);
and U6170 (N_6170,N_5216,N_5526);
or U6171 (N_6171,N_4953,N_5373);
and U6172 (N_6172,N_5145,N_4886);
or U6173 (N_6173,N_5279,N_5169);
xor U6174 (N_6174,N_4806,N_5052);
nand U6175 (N_6175,N_5284,N_5549);
xor U6176 (N_6176,N_5216,N_5384);
nor U6177 (N_6177,N_5339,N_5467);
xnor U6178 (N_6178,N_5140,N_5400);
xnor U6179 (N_6179,N_5546,N_5261);
xnor U6180 (N_6180,N_4925,N_5532);
nand U6181 (N_6181,N_5396,N_5120);
nor U6182 (N_6182,N_4901,N_5301);
nor U6183 (N_6183,N_5496,N_5010);
xor U6184 (N_6184,N_5559,N_5328);
xnor U6185 (N_6185,N_5093,N_4854);
xor U6186 (N_6186,N_5099,N_5419);
nor U6187 (N_6187,N_5353,N_4961);
and U6188 (N_6188,N_5360,N_5462);
or U6189 (N_6189,N_4816,N_5034);
xnor U6190 (N_6190,N_5502,N_5414);
or U6191 (N_6191,N_4817,N_5468);
or U6192 (N_6192,N_5350,N_4879);
or U6193 (N_6193,N_4849,N_5409);
nand U6194 (N_6194,N_5424,N_5312);
and U6195 (N_6195,N_5248,N_5090);
nand U6196 (N_6196,N_5250,N_5531);
xnor U6197 (N_6197,N_5502,N_5318);
nand U6198 (N_6198,N_5380,N_5315);
nand U6199 (N_6199,N_5504,N_5021);
or U6200 (N_6200,N_5090,N_5269);
nand U6201 (N_6201,N_4911,N_5409);
and U6202 (N_6202,N_5040,N_5334);
or U6203 (N_6203,N_5117,N_5481);
nor U6204 (N_6204,N_5566,N_5595);
nor U6205 (N_6205,N_4826,N_5248);
nor U6206 (N_6206,N_5349,N_5449);
or U6207 (N_6207,N_4807,N_5451);
or U6208 (N_6208,N_5474,N_5530);
and U6209 (N_6209,N_5252,N_5478);
and U6210 (N_6210,N_5376,N_4846);
nor U6211 (N_6211,N_5051,N_5185);
xor U6212 (N_6212,N_5578,N_5249);
nor U6213 (N_6213,N_5547,N_5275);
nand U6214 (N_6214,N_5575,N_5337);
nand U6215 (N_6215,N_4924,N_5176);
or U6216 (N_6216,N_5449,N_5467);
xnor U6217 (N_6217,N_5003,N_5231);
and U6218 (N_6218,N_5051,N_5011);
nor U6219 (N_6219,N_5582,N_5270);
nand U6220 (N_6220,N_4927,N_5425);
xnor U6221 (N_6221,N_4957,N_5006);
or U6222 (N_6222,N_5436,N_5029);
nor U6223 (N_6223,N_5548,N_5082);
nor U6224 (N_6224,N_5207,N_4861);
and U6225 (N_6225,N_5154,N_4963);
nor U6226 (N_6226,N_5315,N_4968);
xnor U6227 (N_6227,N_5344,N_5418);
xnor U6228 (N_6228,N_5003,N_4905);
xor U6229 (N_6229,N_5115,N_5482);
or U6230 (N_6230,N_5140,N_4845);
xnor U6231 (N_6231,N_5070,N_5490);
nor U6232 (N_6232,N_4858,N_5338);
and U6233 (N_6233,N_5512,N_4877);
xnor U6234 (N_6234,N_5458,N_4865);
xnor U6235 (N_6235,N_5170,N_5297);
nor U6236 (N_6236,N_5113,N_5474);
nor U6237 (N_6237,N_4866,N_5422);
xnor U6238 (N_6238,N_4818,N_5562);
or U6239 (N_6239,N_4877,N_5158);
xor U6240 (N_6240,N_5530,N_5187);
xnor U6241 (N_6241,N_5271,N_5454);
or U6242 (N_6242,N_4820,N_5347);
nor U6243 (N_6243,N_5230,N_5295);
and U6244 (N_6244,N_4986,N_5584);
nor U6245 (N_6245,N_5445,N_5031);
or U6246 (N_6246,N_5006,N_4887);
and U6247 (N_6247,N_5239,N_5374);
or U6248 (N_6248,N_5598,N_5404);
nand U6249 (N_6249,N_4847,N_5591);
or U6250 (N_6250,N_4841,N_5448);
nand U6251 (N_6251,N_5522,N_5378);
or U6252 (N_6252,N_5200,N_5416);
nor U6253 (N_6253,N_5146,N_4868);
and U6254 (N_6254,N_5562,N_4977);
nand U6255 (N_6255,N_5115,N_5365);
xor U6256 (N_6256,N_5464,N_5207);
nand U6257 (N_6257,N_5047,N_5506);
xor U6258 (N_6258,N_5248,N_5117);
nor U6259 (N_6259,N_4832,N_4980);
and U6260 (N_6260,N_4987,N_5461);
and U6261 (N_6261,N_5488,N_4952);
nor U6262 (N_6262,N_5410,N_4810);
or U6263 (N_6263,N_5077,N_4960);
xor U6264 (N_6264,N_4924,N_5050);
and U6265 (N_6265,N_5114,N_5088);
xnor U6266 (N_6266,N_5361,N_5395);
and U6267 (N_6267,N_5082,N_5192);
nor U6268 (N_6268,N_4895,N_4870);
or U6269 (N_6269,N_5241,N_4811);
or U6270 (N_6270,N_5403,N_4870);
nand U6271 (N_6271,N_5477,N_4994);
nor U6272 (N_6272,N_5579,N_4805);
and U6273 (N_6273,N_5379,N_5518);
or U6274 (N_6274,N_4965,N_5224);
and U6275 (N_6275,N_5143,N_5035);
or U6276 (N_6276,N_5143,N_4881);
and U6277 (N_6277,N_5463,N_5567);
and U6278 (N_6278,N_4808,N_5182);
nand U6279 (N_6279,N_4879,N_5527);
xor U6280 (N_6280,N_5407,N_5409);
and U6281 (N_6281,N_4858,N_5195);
nand U6282 (N_6282,N_4948,N_5160);
nand U6283 (N_6283,N_5434,N_5437);
and U6284 (N_6284,N_4965,N_5060);
xnor U6285 (N_6285,N_5488,N_5137);
or U6286 (N_6286,N_5231,N_5531);
or U6287 (N_6287,N_5584,N_5051);
nor U6288 (N_6288,N_5036,N_5108);
nor U6289 (N_6289,N_4821,N_5275);
nor U6290 (N_6290,N_5136,N_4823);
nand U6291 (N_6291,N_5032,N_5175);
nor U6292 (N_6292,N_5435,N_4891);
nor U6293 (N_6293,N_5102,N_5592);
nor U6294 (N_6294,N_4865,N_4943);
or U6295 (N_6295,N_4918,N_5465);
or U6296 (N_6296,N_5295,N_5538);
and U6297 (N_6297,N_4983,N_5056);
and U6298 (N_6298,N_5229,N_4836);
nand U6299 (N_6299,N_4970,N_5280);
nor U6300 (N_6300,N_4996,N_5460);
or U6301 (N_6301,N_4830,N_5262);
or U6302 (N_6302,N_5158,N_5364);
or U6303 (N_6303,N_4834,N_5299);
xnor U6304 (N_6304,N_5090,N_5520);
and U6305 (N_6305,N_5245,N_5205);
nor U6306 (N_6306,N_4999,N_5117);
or U6307 (N_6307,N_5591,N_5305);
nor U6308 (N_6308,N_5012,N_5423);
or U6309 (N_6309,N_5291,N_5568);
nor U6310 (N_6310,N_5431,N_4800);
nand U6311 (N_6311,N_4833,N_5555);
and U6312 (N_6312,N_5418,N_4983);
and U6313 (N_6313,N_5552,N_5117);
or U6314 (N_6314,N_5530,N_5073);
or U6315 (N_6315,N_5061,N_5230);
xor U6316 (N_6316,N_4815,N_5115);
and U6317 (N_6317,N_5491,N_5201);
nor U6318 (N_6318,N_5340,N_5543);
xor U6319 (N_6319,N_5298,N_5277);
nand U6320 (N_6320,N_5276,N_5155);
nor U6321 (N_6321,N_5334,N_5111);
or U6322 (N_6322,N_4963,N_4903);
nor U6323 (N_6323,N_5431,N_5221);
nand U6324 (N_6324,N_5000,N_5164);
xor U6325 (N_6325,N_4960,N_5397);
nand U6326 (N_6326,N_5539,N_4814);
nand U6327 (N_6327,N_5036,N_5558);
and U6328 (N_6328,N_5248,N_4895);
or U6329 (N_6329,N_5584,N_5578);
nand U6330 (N_6330,N_5147,N_5012);
or U6331 (N_6331,N_5142,N_5569);
and U6332 (N_6332,N_5077,N_5393);
or U6333 (N_6333,N_5535,N_5391);
nor U6334 (N_6334,N_5368,N_5339);
xnor U6335 (N_6335,N_5134,N_5031);
xnor U6336 (N_6336,N_5594,N_5528);
or U6337 (N_6337,N_5435,N_4988);
nand U6338 (N_6338,N_5022,N_5559);
and U6339 (N_6339,N_4819,N_5146);
or U6340 (N_6340,N_5312,N_5293);
xnor U6341 (N_6341,N_5263,N_5174);
nor U6342 (N_6342,N_4985,N_5010);
or U6343 (N_6343,N_4985,N_5541);
nor U6344 (N_6344,N_5235,N_5127);
or U6345 (N_6345,N_4826,N_5175);
and U6346 (N_6346,N_5108,N_5188);
xor U6347 (N_6347,N_5381,N_4998);
or U6348 (N_6348,N_5331,N_5452);
xnor U6349 (N_6349,N_4987,N_4943);
nor U6350 (N_6350,N_5441,N_5080);
or U6351 (N_6351,N_5265,N_4929);
nand U6352 (N_6352,N_5100,N_4875);
nor U6353 (N_6353,N_5384,N_5567);
nor U6354 (N_6354,N_4802,N_4958);
nor U6355 (N_6355,N_5513,N_4989);
and U6356 (N_6356,N_5367,N_5532);
nand U6357 (N_6357,N_4994,N_5588);
nor U6358 (N_6358,N_4922,N_5156);
nand U6359 (N_6359,N_4840,N_5399);
nand U6360 (N_6360,N_5209,N_5504);
nor U6361 (N_6361,N_4804,N_5335);
nand U6362 (N_6362,N_5000,N_4920);
and U6363 (N_6363,N_5138,N_5171);
nand U6364 (N_6364,N_5249,N_5001);
and U6365 (N_6365,N_5579,N_5364);
or U6366 (N_6366,N_5157,N_5572);
xor U6367 (N_6367,N_4966,N_5054);
or U6368 (N_6368,N_5072,N_5244);
xnor U6369 (N_6369,N_5202,N_5323);
nand U6370 (N_6370,N_5146,N_4807);
xnor U6371 (N_6371,N_5479,N_5486);
xor U6372 (N_6372,N_5351,N_4868);
xor U6373 (N_6373,N_5371,N_5360);
nor U6374 (N_6374,N_5338,N_5391);
nand U6375 (N_6375,N_5289,N_5533);
and U6376 (N_6376,N_5315,N_5163);
nand U6377 (N_6377,N_4856,N_5442);
and U6378 (N_6378,N_5446,N_5567);
nor U6379 (N_6379,N_4819,N_4918);
nor U6380 (N_6380,N_5412,N_5561);
and U6381 (N_6381,N_4848,N_5409);
or U6382 (N_6382,N_5434,N_5429);
nor U6383 (N_6383,N_5390,N_5475);
or U6384 (N_6384,N_5191,N_5290);
nand U6385 (N_6385,N_5081,N_5412);
nand U6386 (N_6386,N_5316,N_4986);
and U6387 (N_6387,N_5078,N_4865);
nand U6388 (N_6388,N_4820,N_5567);
or U6389 (N_6389,N_5385,N_5292);
xnor U6390 (N_6390,N_5402,N_5027);
or U6391 (N_6391,N_5057,N_4880);
nor U6392 (N_6392,N_5131,N_4850);
and U6393 (N_6393,N_5369,N_4941);
nand U6394 (N_6394,N_5363,N_5064);
nand U6395 (N_6395,N_5194,N_5262);
nand U6396 (N_6396,N_5005,N_4915);
nand U6397 (N_6397,N_5127,N_5301);
xor U6398 (N_6398,N_5552,N_5427);
and U6399 (N_6399,N_5104,N_5206);
xor U6400 (N_6400,N_5909,N_6223);
nor U6401 (N_6401,N_6043,N_6385);
or U6402 (N_6402,N_5654,N_5904);
nand U6403 (N_6403,N_5686,N_6330);
nor U6404 (N_6404,N_6205,N_5605);
and U6405 (N_6405,N_6143,N_5976);
nand U6406 (N_6406,N_6389,N_6125);
nand U6407 (N_6407,N_5847,N_5691);
nor U6408 (N_6408,N_6329,N_5939);
and U6409 (N_6409,N_5756,N_6068);
nand U6410 (N_6410,N_6147,N_5794);
or U6411 (N_6411,N_5834,N_5688);
nor U6412 (N_6412,N_5879,N_5713);
and U6413 (N_6413,N_5946,N_6221);
or U6414 (N_6414,N_5937,N_6238);
and U6415 (N_6415,N_5769,N_6104);
xnor U6416 (N_6416,N_6088,N_5817);
and U6417 (N_6417,N_5626,N_5839);
xnor U6418 (N_6418,N_6006,N_6346);
xor U6419 (N_6419,N_6055,N_5902);
xor U6420 (N_6420,N_6155,N_5696);
nor U6421 (N_6421,N_5803,N_5938);
nor U6422 (N_6422,N_5742,N_5670);
and U6423 (N_6423,N_5884,N_6067);
nor U6424 (N_6424,N_5918,N_5759);
nor U6425 (N_6425,N_5727,N_5699);
or U6426 (N_6426,N_5666,N_5674);
xor U6427 (N_6427,N_5960,N_6153);
nor U6428 (N_6428,N_6278,N_6197);
xnor U6429 (N_6429,N_6102,N_6179);
xnor U6430 (N_6430,N_5963,N_5747);
nand U6431 (N_6431,N_5640,N_6076);
nor U6432 (N_6432,N_6216,N_5914);
and U6433 (N_6433,N_5734,N_5876);
xor U6434 (N_6434,N_6158,N_6367);
nor U6435 (N_6435,N_5702,N_5889);
nor U6436 (N_6436,N_6062,N_6256);
nor U6437 (N_6437,N_5882,N_5796);
nor U6438 (N_6438,N_6239,N_5956);
nand U6439 (N_6439,N_5706,N_5786);
or U6440 (N_6440,N_5764,N_5888);
and U6441 (N_6441,N_5779,N_5931);
nand U6442 (N_6442,N_6119,N_6274);
xor U6443 (N_6443,N_5651,N_5892);
nor U6444 (N_6444,N_5875,N_5693);
and U6445 (N_6445,N_6266,N_6378);
nor U6446 (N_6446,N_6218,N_6314);
nand U6447 (N_6447,N_6350,N_5646);
or U6448 (N_6448,N_5784,N_6328);
or U6449 (N_6449,N_5830,N_5788);
or U6450 (N_6450,N_6032,N_6142);
or U6451 (N_6451,N_5715,N_5912);
nand U6452 (N_6452,N_5631,N_6152);
nand U6453 (N_6453,N_6165,N_5653);
nor U6454 (N_6454,N_6276,N_6210);
or U6455 (N_6455,N_5851,N_6263);
nor U6456 (N_6456,N_5837,N_6016);
nand U6457 (N_6457,N_5991,N_5676);
or U6458 (N_6458,N_5695,N_6353);
or U6459 (N_6459,N_5947,N_5869);
xor U6460 (N_6460,N_6325,N_6261);
nor U6461 (N_6461,N_5744,N_5896);
or U6462 (N_6462,N_6253,N_5637);
nand U6463 (N_6463,N_6192,N_6316);
nor U6464 (N_6464,N_5999,N_5872);
or U6465 (N_6465,N_5878,N_5733);
or U6466 (N_6466,N_6277,N_6307);
nand U6467 (N_6467,N_5964,N_6168);
and U6468 (N_6468,N_6213,N_5671);
nand U6469 (N_6469,N_6196,N_6004);
or U6470 (N_6470,N_6294,N_6324);
or U6471 (N_6471,N_6392,N_6275);
nand U6472 (N_6472,N_5968,N_6061);
nor U6473 (N_6473,N_5883,N_6198);
and U6474 (N_6474,N_6014,N_6347);
and U6475 (N_6475,N_5980,N_5940);
nand U6476 (N_6476,N_6206,N_6241);
nand U6477 (N_6477,N_5636,N_6387);
nand U6478 (N_6478,N_6090,N_6260);
and U6479 (N_6479,N_6011,N_6010);
nand U6480 (N_6480,N_5746,N_5682);
or U6481 (N_6481,N_6030,N_6345);
nor U6482 (N_6482,N_5880,N_5773);
xor U6483 (N_6483,N_6078,N_6111);
and U6484 (N_6484,N_5607,N_5738);
nor U6485 (N_6485,N_5903,N_5885);
and U6486 (N_6486,N_5762,N_5655);
xor U6487 (N_6487,N_6255,N_6121);
nor U6488 (N_6488,N_5948,N_6342);
nand U6489 (N_6489,N_5729,N_6137);
nor U6490 (N_6490,N_5859,N_6243);
xnor U6491 (N_6491,N_6200,N_5719);
nand U6492 (N_6492,N_6313,N_5728);
nand U6493 (N_6493,N_6398,N_5850);
nand U6494 (N_6494,N_6273,N_6020);
or U6495 (N_6495,N_6097,N_6052);
or U6496 (N_6496,N_5819,N_5955);
nor U6497 (N_6497,N_6122,N_5805);
xor U6498 (N_6498,N_5966,N_5987);
xor U6499 (N_6499,N_6133,N_6240);
nor U6500 (N_6500,N_6064,N_5697);
xnor U6501 (N_6501,N_5934,N_6291);
nor U6502 (N_6502,N_5632,N_5775);
and U6503 (N_6503,N_6336,N_6351);
and U6504 (N_6504,N_6355,N_5967);
and U6505 (N_6505,N_6149,N_6364);
and U6506 (N_6506,N_5743,N_6303);
or U6507 (N_6507,N_5766,N_6250);
and U6508 (N_6508,N_6323,N_5887);
nand U6509 (N_6509,N_5898,N_6359);
and U6510 (N_6510,N_6322,N_5615);
and U6511 (N_6511,N_6176,N_5996);
or U6512 (N_6512,N_6047,N_5618);
or U6513 (N_6513,N_5985,N_6219);
and U6514 (N_6514,N_6368,N_5721);
nand U6515 (N_6515,N_6194,N_6396);
xor U6516 (N_6516,N_6005,N_6201);
nand U6517 (N_6517,N_5957,N_5608);
nor U6518 (N_6518,N_5926,N_5848);
and U6519 (N_6519,N_6018,N_5649);
nand U6520 (N_6520,N_5737,N_5951);
and U6521 (N_6521,N_6365,N_6229);
and U6522 (N_6522,N_5714,N_6031);
xnor U6523 (N_6523,N_5652,N_5907);
nand U6524 (N_6524,N_6344,N_5970);
and U6525 (N_6525,N_6093,N_5731);
xnor U6526 (N_6526,N_6366,N_6017);
xnor U6527 (N_6527,N_5795,N_5983);
nand U6528 (N_6528,N_5771,N_6115);
and U6529 (N_6529,N_6204,N_5611);
or U6530 (N_6530,N_5755,N_6002);
xor U6531 (N_6531,N_5823,N_5690);
xor U6532 (N_6532,N_5809,N_6375);
or U6533 (N_6533,N_6383,N_6272);
nor U6534 (N_6534,N_6098,N_5910);
and U6535 (N_6535,N_5920,N_5675);
nor U6536 (N_6536,N_5992,N_5712);
and U6537 (N_6537,N_6227,N_6001);
and U6538 (N_6538,N_5776,N_5614);
xor U6539 (N_6539,N_6025,N_6315);
nor U6540 (N_6540,N_5613,N_6167);
nand U6541 (N_6541,N_5831,N_6299);
or U6542 (N_6542,N_6056,N_5698);
nor U6543 (N_6543,N_5790,N_6038);
nand U6544 (N_6544,N_6070,N_5833);
xnor U6545 (N_6545,N_6354,N_5827);
and U6546 (N_6546,N_5886,N_6117);
or U6547 (N_6547,N_6144,N_6222);
and U6548 (N_6548,N_5804,N_5659);
or U6549 (N_6549,N_5933,N_5711);
or U6550 (N_6550,N_6259,N_6042);
xor U6551 (N_6551,N_5873,N_6084);
nand U6552 (N_6552,N_6129,N_6304);
and U6553 (N_6553,N_5893,N_6252);
and U6554 (N_6554,N_6019,N_5890);
nor U6555 (N_6555,N_6360,N_6071);
xnor U6556 (N_6556,N_6040,N_5864);
or U6557 (N_6557,N_5801,N_6258);
nand U6558 (N_6558,N_5656,N_6361);
nor U6559 (N_6559,N_6271,N_6159);
nor U6560 (N_6560,N_6319,N_6357);
nor U6561 (N_6561,N_6349,N_5768);
nand U6562 (N_6562,N_6333,N_6321);
or U6563 (N_6563,N_6109,N_5797);
nand U6564 (N_6564,N_5720,N_6053);
nand U6565 (N_6565,N_5821,N_6292);
nor U6566 (N_6566,N_5984,N_5602);
nand U6567 (N_6567,N_6251,N_6188);
nand U6568 (N_6568,N_5612,N_6298);
nor U6569 (N_6569,N_6235,N_6136);
nand U6570 (N_6570,N_6135,N_6236);
xnor U6571 (N_6571,N_5802,N_5757);
xor U6572 (N_6572,N_6191,N_6376);
or U6573 (N_6573,N_6095,N_5783);
nand U6574 (N_6574,N_5681,N_5772);
nor U6575 (N_6575,N_5667,N_6352);
nor U6576 (N_6576,N_5927,N_5924);
and U6577 (N_6577,N_5761,N_6334);
nand U6578 (N_6578,N_6094,N_6037);
xnor U6579 (N_6579,N_6063,N_5741);
nand U6580 (N_6580,N_5945,N_5891);
nand U6581 (N_6581,N_6085,N_5818);
or U6582 (N_6582,N_5978,N_6060);
xor U6583 (N_6583,N_6295,N_5622);
nand U6584 (N_6584,N_5730,N_5854);
nor U6585 (N_6585,N_5662,N_6369);
or U6586 (N_6586,N_6270,N_5680);
nor U6587 (N_6587,N_5658,N_6289);
nand U6588 (N_6588,N_6287,N_5913);
nor U6589 (N_6589,N_6058,N_6190);
nor U6590 (N_6590,N_6300,N_6332);
xnor U6591 (N_6591,N_6215,N_6145);
nor U6592 (N_6592,N_6171,N_5716);
xnor U6593 (N_6593,N_5603,N_6081);
or U6594 (N_6594,N_5844,N_6110);
and U6595 (N_6595,N_5616,N_6099);
xnor U6596 (N_6596,N_6343,N_5645);
or U6597 (N_6597,N_5723,N_6246);
xor U6598 (N_6598,N_6281,N_6399);
and U6599 (N_6599,N_6169,N_5717);
xnor U6600 (N_6600,N_6123,N_6247);
nand U6601 (N_6601,N_5989,N_6262);
nor U6602 (N_6602,N_6083,N_5861);
and U6603 (N_6603,N_6077,N_6086);
or U6604 (N_6604,N_6202,N_5917);
nor U6605 (N_6605,N_6000,N_5857);
nand U6606 (N_6606,N_5677,N_5650);
nor U6607 (N_6607,N_5816,N_6214);
nor U6608 (N_6608,N_5647,N_5994);
and U6609 (N_6609,N_5973,N_5829);
nor U6610 (N_6610,N_6107,N_6013);
or U6611 (N_6611,N_5758,N_6373);
and U6612 (N_6612,N_6338,N_5694);
nand U6613 (N_6613,N_6379,N_6029);
and U6614 (N_6614,N_6148,N_6103);
xor U6615 (N_6615,N_5791,N_5689);
nor U6616 (N_6616,N_5881,N_5942);
nor U6617 (N_6617,N_5787,N_5824);
or U6618 (N_6618,N_5672,N_5822);
xor U6619 (N_6619,N_5634,N_6157);
nor U6620 (N_6620,N_6301,N_5799);
nand U6621 (N_6621,N_6126,N_5894);
nor U6622 (N_6622,N_6065,N_5877);
nand U6623 (N_6623,N_5661,N_5641);
or U6624 (N_6624,N_5778,N_5700);
nor U6625 (N_6625,N_6134,N_5644);
xnor U6626 (N_6626,N_6154,N_6249);
or U6627 (N_6627,N_5812,N_5986);
nor U6628 (N_6628,N_6230,N_5606);
nor U6629 (N_6629,N_5793,N_5722);
xor U6630 (N_6630,N_5840,N_5789);
nor U6631 (N_6631,N_5754,N_5745);
xor U6632 (N_6632,N_6268,N_6184);
xnor U6633 (N_6633,N_5604,N_5905);
and U6634 (N_6634,N_6377,N_6187);
nor U6635 (N_6635,N_5624,N_6228);
nor U6636 (N_6636,N_5687,N_5908);
and U6637 (N_6637,N_5814,N_6138);
nand U6638 (N_6638,N_6339,N_6226);
xor U6639 (N_6639,N_5977,N_6370);
and U6640 (N_6640,N_6131,N_5638);
or U6641 (N_6641,N_5961,N_6008);
and U6642 (N_6642,N_6069,N_6362);
xnor U6643 (N_6643,N_6381,N_6384);
and U6644 (N_6644,N_5750,N_5988);
and U6645 (N_6645,N_6181,N_6244);
or U6646 (N_6646,N_5665,N_5943);
xor U6647 (N_6647,N_5995,N_5916);
or U6648 (N_6648,N_5765,N_6035);
nor U6649 (N_6649,N_6170,N_6356);
nand U6650 (N_6650,N_6028,N_5954);
nand U6651 (N_6651,N_6189,N_6174);
and U6652 (N_6652,N_6124,N_6391);
nand U6653 (N_6653,N_5770,N_6279);
nand U6654 (N_6654,N_5684,N_6348);
nor U6655 (N_6655,N_6089,N_6073);
or U6656 (N_6656,N_6305,N_6096);
and U6657 (N_6657,N_6269,N_5867);
and U6658 (N_6658,N_5609,N_6156);
or U6659 (N_6659,N_5621,N_5748);
nand U6660 (N_6660,N_6224,N_5838);
and U6661 (N_6661,N_5969,N_6130);
nand U6662 (N_6662,N_5932,N_5863);
and U6663 (N_6663,N_6337,N_5664);
xor U6664 (N_6664,N_5941,N_5753);
nand U6665 (N_6665,N_6150,N_5899);
nand U6666 (N_6666,N_5625,N_6380);
xor U6667 (N_6667,N_6265,N_6340);
nor U6668 (N_6668,N_6212,N_6393);
nor U6669 (N_6669,N_5856,N_6091);
nor U6670 (N_6670,N_6310,N_5993);
or U6671 (N_6671,N_5897,N_5981);
nand U6672 (N_6672,N_6066,N_6033);
and U6673 (N_6673,N_5953,N_5990);
and U6674 (N_6674,N_5707,N_6326);
and U6675 (N_6675,N_6286,N_6185);
nand U6676 (N_6676,N_6302,N_6049);
xor U6677 (N_6677,N_5925,N_6007);
and U6678 (N_6678,N_5668,N_6282);
or U6679 (N_6679,N_6397,N_6208);
xor U6680 (N_6680,N_5813,N_5781);
and U6681 (N_6681,N_5623,N_6160);
xor U6682 (N_6682,N_5669,N_6290);
or U6683 (N_6683,N_6163,N_5846);
and U6684 (N_6684,N_5726,N_6080);
nor U6685 (N_6685,N_6003,N_5635);
nand U6686 (N_6686,N_5922,N_6161);
nand U6687 (N_6687,N_5928,N_6220);
xnor U6688 (N_6688,N_5852,N_6386);
nand U6689 (N_6689,N_6127,N_5835);
and U6690 (N_6690,N_6059,N_5923);
nand U6691 (N_6691,N_6092,N_6039);
nand U6692 (N_6692,N_5901,N_6105);
nand U6693 (N_6693,N_5806,N_5868);
nand U6694 (N_6694,N_6394,N_6172);
or U6695 (N_6695,N_6363,N_5958);
and U6696 (N_6696,N_5836,N_5703);
nand U6697 (N_6697,N_5643,N_6317);
or U6698 (N_6698,N_5739,N_5617);
and U6699 (N_6699,N_6232,N_6183);
nor U6700 (N_6700,N_5627,N_5639);
or U6701 (N_6701,N_6318,N_6164);
nand U6702 (N_6702,N_6254,N_5815);
nand U6703 (N_6703,N_6045,N_6335);
nor U6704 (N_6704,N_6054,N_5629);
nor U6705 (N_6705,N_5732,N_5620);
xor U6706 (N_6706,N_5842,N_6118);
nor U6707 (N_6707,N_6358,N_5701);
nor U6708 (N_6708,N_6108,N_5683);
and U6709 (N_6709,N_6320,N_6044);
nand U6710 (N_6710,N_6036,N_6285);
and U6711 (N_6711,N_6233,N_5704);
nor U6712 (N_6712,N_6022,N_5709);
xnor U6713 (N_6713,N_6341,N_5808);
nor U6714 (N_6714,N_5705,N_5843);
nor U6715 (N_6715,N_5785,N_5870);
nor U6716 (N_6716,N_5792,N_6371);
and U6717 (N_6717,N_5915,N_6225);
nand U6718 (N_6718,N_6141,N_6331);
and U6719 (N_6719,N_6217,N_5900);
and U6720 (N_6720,N_5935,N_5962);
or U6721 (N_6721,N_6057,N_6177);
or U6722 (N_6722,N_6199,N_5865);
and U6723 (N_6723,N_6106,N_5777);
xor U6724 (N_6724,N_5736,N_6182);
xnor U6725 (N_6725,N_6113,N_6151);
and U6726 (N_6726,N_6048,N_5630);
and U6727 (N_6727,N_6186,N_5692);
xnor U6728 (N_6728,N_6026,N_6041);
nand U6729 (N_6729,N_6390,N_5965);
nand U6730 (N_6730,N_5642,N_5735);
and U6731 (N_6731,N_5774,N_5798);
or U6732 (N_6732,N_6372,N_5853);
and U6733 (N_6733,N_5921,N_6234);
nor U6734 (N_6734,N_6231,N_6293);
nand U6735 (N_6735,N_5972,N_5807);
nand U6736 (N_6736,N_6051,N_6034);
and U6737 (N_6737,N_6024,N_6101);
nand U6738 (N_6738,N_5944,N_5858);
nor U6739 (N_6739,N_5751,N_5826);
and U6740 (N_6740,N_6312,N_6211);
or U6741 (N_6741,N_6072,N_5782);
xnor U6742 (N_6742,N_6308,N_6178);
nand U6743 (N_6743,N_5959,N_6112);
nor U6744 (N_6744,N_5708,N_5660);
and U6745 (N_6745,N_5998,N_6023);
nand U6746 (N_6746,N_6245,N_5979);
xor U6747 (N_6747,N_6203,N_6237);
nand U6748 (N_6748,N_5906,N_5895);
nand U6749 (N_6749,N_5862,N_5749);
or U6750 (N_6750,N_6114,N_5845);
xor U6751 (N_6751,N_5855,N_5930);
and U6752 (N_6752,N_5860,N_5619);
and U6753 (N_6753,N_5982,N_5911);
nand U6754 (N_6754,N_5820,N_5828);
xor U6755 (N_6755,N_6140,N_6327);
nor U6756 (N_6756,N_5811,N_5936);
and U6757 (N_6757,N_5633,N_6082);
nor U6758 (N_6758,N_5950,N_6284);
or U6759 (N_6759,N_6009,N_6382);
nand U6760 (N_6760,N_5825,N_6046);
nor U6761 (N_6761,N_5600,N_6207);
nand U6762 (N_6762,N_6388,N_5685);
xnor U6763 (N_6763,N_5832,N_5678);
xnor U6764 (N_6764,N_6395,N_5780);
xnor U6765 (N_6765,N_6175,N_6100);
or U6766 (N_6766,N_5952,N_5874);
or U6767 (N_6767,N_6146,N_5610);
nor U6768 (N_6768,N_6050,N_6374);
xnor U6769 (N_6769,N_6257,N_6075);
xnor U6770 (N_6770,N_6079,N_5810);
nand U6771 (N_6771,N_6162,N_5725);
nand U6772 (N_6772,N_5710,N_5628);
and U6773 (N_6773,N_5919,N_6074);
xor U6774 (N_6774,N_5974,N_6087);
or U6775 (N_6775,N_5718,N_6132);
and U6776 (N_6776,N_5663,N_6021);
nor U6777 (N_6777,N_5997,N_5601);
xnor U6778 (N_6778,N_6296,N_5724);
or U6779 (N_6779,N_6128,N_6193);
nor U6780 (N_6780,N_6166,N_6264);
and U6781 (N_6781,N_5648,N_6195);
nor U6782 (N_6782,N_5767,N_6173);
and U6783 (N_6783,N_5871,N_6242);
and U6784 (N_6784,N_6288,N_6209);
xnor U6785 (N_6785,N_6180,N_6120);
nand U6786 (N_6786,N_6139,N_6297);
nor U6787 (N_6787,N_5841,N_5760);
xnor U6788 (N_6788,N_6027,N_5929);
and U6789 (N_6789,N_6116,N_6280);
nor U6790 (N_6790,N_6311,N_5971);
xor U6791 (N_6791,N_6015,N_5657);
xnor U6792 (N_6792,N_5679,N_6012);
or U6793 (N_6793,N_5752,N_5740);
and U6794 (N_6794,N_6283,N_6267);
and U6795 (N_6795,N_6248,N_6309);
nand U6796 (N_6796,N_6306,N_5763);
or U6797 (N_6797,N_5849,N_5673);
xnor U6798 (N_6798,N_5866,N_5975);
xor U6799 (N_6799,N_5949,N_5800);
nand U6800 (N_6800,N_5952,N_5777);
nand U6801 (N_6801,N_6289,N_5646);
xnor U6802 (N_6802,N_5624,N_6350);
and U6803 (N_6803,N_5920,N_6252);
nand U6804 (N_6804,N_5610,N_5609);
nor U6805 (N_6805,N_5763,N_6276);
or U6806 (N_6806,N_5955,N_6304);
or U6807 (N_6807,N_5862,N_5806);
and U6808 (N_6808,N_5679,N_6317);
nand U6809 (N_6809,N_6262,N_5732);
or U6810 (N_6810,N_5728,N_6049);
and U6811 (N_6811,N_5690,N_5858);
or U6812 (N_6812,N_5658,N_5908);
and U6813 (N_6813,N_6268,N_5924);
and U6814 (N_6814,N_6327,N_5795);
and U6815 (N_6815,N_6296,N_6219);
nand U6816 (N_6816,N_6235,N_6353);
nand U6817 (N_6817,N_6011,N_6083);
or U6818 (N_6818,N_6150,N_6261);
nand U6819 (N_6819,N_5718,N_6087);
xnor U6820 (N_6820,N_6346,N_5770);
nor U6821 (N_6821,N_6065,N_5621);
or U6822 (N_6822,N_5715,N_6255);
nor U6823 (N_6823,N_6195,N_5679);
nor U6824 (N_6824,N_5916,N_5681);
nand U6825 (N_6825,N_6365,N_6094);
or U6826 (N_6826,N_6057,N_6132);
or U6827 (N_6827,N_5887,N_5682);
nor U6828 (N_6828,N_5845,N_5906);
and U6829 (N_6829,N_5878,N_5938);
nor U6830 (N_6830,N_5855,N_6372);
nand U6831 (N_6831,N_5720,N_6337);
xnor U6832 (N_6832,N_5780,N_5740);
nand U6833 (N_6833,N_6139,N_5967);
and U6834 (N_6834,N_6262,N_6202);
and U6835 (N_6835,N_6132,N_6036);
or U6836 (N_6836,N_6005,N_5904);
xor U6837 (N_6837,N_5713,N_6392);
nand U6838 (N_6838,N_6125,N_5996);
nand U6839 (N_6839,N_5689,N_5701);
xor U6840 (N_6840,N_5911,N_6045);
nand U6841 (N_6841,N_5760,N_6320);
xor U6842 (N_6842,N_6097,N_5902);
or U6843 (N_6843,N_6079,N_6069);
xor U6844 (N_6844,N_6279,N_6015);
and U6845 (N_6845,N_5766,N_6242);
nor U6846 (N_6846,N_6235,N_6289);
and U6847 (N_6847,N_6198,N_6386);
xor U6848 (N_6848,N_6167,N_5760);
xor U6849 (N_6849,N_5906,N_5805);
nor U6850 (N_6850,N_5634,N_6075);
and U6851 (N_6851,N_5696,N_5663);
nor U6852 (N_6852,N_5608,N_6201);
and U6853 (N_6853,N_6035,N_5893);
and U6854 (N_6854,N_5648,N_5618);
and U6855 (N_6855,N_5659,N_6343);
and U6856 (N_6856,N_5912,N_5816);
or U6857 (N_6857,N_6181,N_6153);
or U6858 (N_6858,N_5948,N_5709);
or U6859 (N_6859,N_5780,N_6361);
and U6860 (N_6860,N_6343,N_6151);
and U6861 (N_6861,N_6262,N_5833);
nand U6862 (N_6862,N_6011,N_6280);
and U6863 (N_6863,N_5870,N_6376);
and U6864 (N_6864,N_5976,N_5873);
nor U6865 (N_6865,N_6073,N_5807);
and U6866 (N_6866,N_5785,N_5828);
nor U6867 (N_6867,N_6006,N_6030);
nor U6868 (N_6868,N_5884,N_6089);
nand U6869 (N_6869,N_5723,N_6176);
or U6870 (N_6870,N_5647,N_6309);
or U6871 (N_6871,N_5654,N_5726);
nand U6872 (N_6872,N_5692,N_5649);
nand U6873 (N_6873,N_5878,N_5896);
nor U6874 (N_6874,N_6274,N_5853);
xnor U6875 (N_6875,N_5878,N_6148);
xnor U6876 (N_6876,N_6082,N_6131);
nand U6877 (N_6877,N_6086,N_5700);
nor U6878 (N_6878,N_5678,N_5777);
nor U6879 (N_6879,N_5866,N_6347);
and U6880 (N_6880,N_5729,N_6281);
and U6881 (N_6881,N_6372,N_5876);
and U6882 (N_6882,N_5923,N_6197);
and U6883 (N_6883,N_6158,N_6192);
or U6884 (N_6884,N_6031,N_6323);
xor U6885 (N_6885,N_6367,N_5983);
or U6886 (N_6886,N_6320,N_5866);
and U6887 (N_6887,N_5899,N_6199);
and U6888 (N_6888,N_6265,N_5820);
nor U6889 (N_6889,N_5775,N_5620);
nor U6890 (N_6890,N_5786,N_5616);
nand U6891 (N_6891,N_6106,N_5623);
nand U6892 (N_6892,N_5668,N_6330);
or U6893 (N_6893,N_5785,N_5862);
or U6894 (N_6894,N_6178,N_5709);
xor U6895 (N_6895,N_6188,N_5815);
and U6896 (N_6896,N_5776,N_5727);
and U6897 (N_6897,N_5689,N_6338);
xor U6898 (N_6898,N_6151,N_6298);
or U6899 (N_6899,N_5863,N_6234);
nor U6900 (N_6900,N_6283,N_5689);
or U6901 (N_6901,N_5889,N_6346);
nor U6902 (N_6902,N_6297,N_6002);
and U6903 (N_6903,N_5963,N_5741);
nor U6904 (N_6904,N_6295,N_5862);
or U6905 (N_6905,N_6026,N_6218);
nor U6906 (N_6906,N_5973,N_6345);
xor U6907 (N_6907,N_6234,N_6272);
or U6908 (N_6908,N_5772,N_6353);
or U6909 (N_6909,N_5917,N_6365);
nor U6910 (N_6910,N_5617,N_6319);
or U6911 (N_6911,N_6219,N_5746);
nand U6912 (N_6912,N_5999,N_6243);
or U6913 (N_6913,N_6386,N_5806);
nand U6914 (N_6914,N_5656,N_5652);
xor U6915 (N_6915,N_5736,N_6067);
and U6916 (N_6916,N_6171,N_6383);
nand U6917 (N_6917,N_6161,N_6032);
nor U6918 (N_6918,N_5996,N_6309);
or U6919 (N_6919,N_6198,N_5982);
or U6920 (N_6920,N_5984,N_5753);
or U6921 (N_6921,N_6283,N_5992);
and U6922 (N_6922,N_6387,N_5940);
and U6923 (N_6923,N_6277,N_5903);
nand U6924 (N_6924,N_6239,N_6108);
and U6925 (N_6925,N_6323,N_6126);
or U6926 (N_6926,N_5799,N_6037);
or U6927 (N_6927,N_5882,N_5947);
nand U6928 (N_6928,N_6025,N_5968);
nor U6929 (N_6929,N_5800,N_6319);
xor U6930 (N_6930,N_6210,N_6377);
and U6931 (N_6931,N_5628,N_6224);
and U6932 (N_6932,N_6110,N_5708);
nand U6933 (N_6933,N_5732,N_5683);
nand U6934 (N_6934,N_6366,N_5601);
xor U6935 (N_6935,N_6084,N_6120);
nor U6936 (N_6936,N_6247,N_6155);
nor U6937 (N_6937,N_5798,N_5900);
nand U6938 (N_6938,N_5951,N_6274);
xor U6939 (N_6939,N_6000,N_6391);
nand U6940 (N_6940,N_6087,N_6330);
nor U6941 (N_6941,N_6051,N_5847);
nor U6942 (N_6942,N_5866,N_5939);
or U6943 (N_6943,N_6095,N_6298);
nor U6944 (N_6944,N_6391,N_6247);
or U6945 (N_6945,N_5865,N_6117);
nand U6946 (N_6946,N_6085,N_6035);
nor U6947 (N_6947,N_5968,N_6050);
and U6948 (N_6948,N_6149,N_6045);
and U6949 (N_6949,N_5980,N_6206);
nor U6950 (N_6950,N_5705,N_5865);
xor U6951 (N_6951,N_6383,N_6199);
or U6952 (N_6952,N_6099,N_5663);
xor U6953 (N_6953,N_6370,N_6353);
nand U6954 (N_6954,N_5830,N_6280);
and U6955 (N_6955,N_5721,N_5602);
xnor U6956 (N_6956,N_5893,N_6324);
xor U6957 (N_6957,N_6190,N_6132);
nor U6958 (N_6958,N_6352,N_6022);
nand U6959 (N_6959,N_6380,N_5953);
or U6960 (N_6960,N_6036,N_6388);
nand U6961 (N_6961,N_6134,N_5936);
xor U6962 (N_6962,N_6378,N_5876);
and U6963 (N_6963,N_5792,N_6271);
nor U6964 (N_6964,N_6235,N_5620);
nand U6965 (N_6965,N_5648,N_6024);
xnor U6966 (N_6966,N_6290,N_5875);
or U6967 (N_6967,N_5779,N_5628);
nor U6968 (N_6968,N_5986,N_6339);
xor U6969 (N_6969,N_6135,N_6109);
xor U6970 (N_6970,N_6169,N_5879);
and U6971 (N_6971,N_6067,N_6095);
nand U6972 (N_6972,N_6296,N_5934);
nand U6973 (N_6973,N_6376,N_6331);
or U6974 (N_6974,N_6282,N_5999);
nor U6975 (N_6975,N_5949,N_5753);
and U6976 (N_6976,N_5873,N_5930);
nand U6977 (N_6977,N_6281,N_5828);
xnor U6978 (N_6978,N_5766,N_5750);
nor U6979 (N_6979,N_5940,N_5754);
nor U6980 (N_6980,N_5616,N_6363);
nor U6981 (N_6981,N_6103,N_6287);
xnor U6982 (N_6982,N_5964,N_5746);
nand U6983 (N_6983,N_5710,N_6172);
or U6984 (N_6984,N_5800,N_6190);
or U6985 (N_6985,N_6368,N_6031);
nor U6986 (N_6986,N_6222,N_6170);
nor U6987 (N_6987,N_6227,N_5970);
and U6988 (N_6988,N_5615,N_6017);
nand U6989 (N_6989,N_6001,N_6157);
xor U6990 (N_6990,N_5835,N_6398);
and U6991 (N_6991,N_6284,N_5611);
nand U6992 (N_6992,N_6242,N_6189);
and U6993 (N_6993,N_6115,N_5892);
nor U6994 (N_6994,N_6325,N_5823);
nand U6995 (N_6995,N_6232,N_5615);
and U6996 (N_6996,N_6211,N_5926);
nor U6997 (N_6997,N_5974,N_6240);
xnor U6998 (N_6998,N_5788,N_5670);
and U6999 (N_6999,N_5755,N_6302);
xor U7000 (N_7000,N_6332,N_5724);
or U7001 (N_7001,N_5614,N_5951);
xnor U7002 (N_7002,N_5825,N_5753);
or U7003 (N_7003,N_5856,N_6348);
and U7004 (N_7004,N_6326,N_5801);
xor U7005 (N_7005,N_5998,N_6320);
xor U7006 (N_7006,N_5789,N_6055);
xnor U7007 (N_7007,N_6114,N_6302);
nor U7008 (N_7008,N_5633,N_6330);
nor U7009 (N_7009,N_6365,N_6283);
nor U7010 (N_7010,N_6292,N_5894);
xnor U7011 (N_7011,N_5967,N_5766);
and U7012 (N_7012,N_5626,N_5826);
and U7013 (N_7013,N_5957,N_5660);
nor U7014 (N_7014,N_6359,N_6155);
and U7015 (N_7015,N_5988,N_6297);
nor U7016 (N_7016,N_6007,N_6312);
or U7017 (N_7017,N_5753,N_5804);
xor U7018 (N_7018,N_5901,N_5684);
and U7019 (N_7019,N_6255,N_5954);
nand U7020 (N_7020,N_5968,N_5874);
or U7021 (N_7021,N_6062,N_5980);
and U7022 (N_7022,N_6150,N_5783);
nand U7023 (N_7023,N_6225,N_6390);
xor U7024 (N_7024,N_6174,N_5695);
xnor U7025 (N_7025,N_6321,N_5631);
or U7026 (N_7026,N_6387,N_6230);
and U7027 (N_7027,N_6024,N_6273);
and U7028 (N_7028,N_5758,N_5882);
nand U7029 (N_7029,N_6009,N_6248);
xnor U7030 (N_7030,N_6112,N_5901);
nand U7031 (N_7031,N_6157,N_6350);
or U7032 (N_7032,N_5688,N_6029);
nand U7033 (N_7033,N_6074,N_5633);
and U7034 (N_7034,N_5653,N_5640);
nand U7035 (N_7035,N_5883,N_5639);
and U7036 (N_7036,N_6240,N_5613);
and U7037 (N_7037,N_6342,N_5841);
nor U7038 (N_7038,N_6389,N_6110);
or U7039 (N_7039,N_6190,N_5665);
xnor U7040 (N_7040,N_5718,N_6097);
nor U7041 (N_7041,N_6294,N_6131);
or U7042 (N_7042,N_6251,N_5918);
nand U7043 (N_7043,N_6186,N_6322);
and U7044 (N_7044,N_6373,N_5648);
and U7045 (N_7045,N_5610,N_5677);
nor U7046 (N_7046,N_5662,N_5639);
xor U7047 (N_7047,N_6331,N_5917);
xnor U7048 (N_7048,N_5912,N_5883);
xnor U7049 (N_7049,N_6233,N_6089);
or U7050 (N_7050,N_5938,N_6238);
nand U7051 (N_7051,N_6333,N_5848);
nor U7052 (N_7052,N_6146,N_6206);
or U7053 (N_7053,N_6164,N_5893);
xnor U7054 (N_7054,N_6365,N_6384);
or U7055 (N_7055,N_5975,N_6009);
and U7056 (N_7056,N_6318,N_6131);
xnor U7057 (N_7057,N_6289,N_6081);
xor U7058 (N_7058,N_6347,N_5780);
nand U7059 (N_7059,N_6150,N_5718);
nand U7060 (N_7060,N_5780,N_6309);
and U7061 (N_7061,N_6121,N_6296);
xor U7062 (N_7062,N_5970,N_6369);
xor U7063 (N_7063,N_6047,N_5839);
nand U7064 (N_7064,N_6047,N_5937);
nor U7065 (N_7065,N_6366,N_5990);
and U7066 (N_7066,N_6208,N_5756);
nor U7067 (N_7067,N_5991,N_5879);
or U7068 (N_7068,N_6005,N_5745);
xor U7069 (N_7069,N_6297,N_5834);
and U7070 (N_7070,N_5892,N_6177);
and U7071 (N_7071,N_6195,N_6280);
nor U7072 (N_7072,N_6079,N_6111);
xnor U7073 (N_7073,N_6058,N_6353);
and U7074 (N_7074,N_5930,N_5935);
nor U7075 (N_7075,N_5800,N_6230);
nor U7076 (N_7076,N_5672,N_6180);
nand U7077 (N_7077,N_6132,N_5654);
nand U7078 (N_7078,N_6292,N_6124);
nand U7079 (N_7079,N_6335,N_6331);
xnor U7080 (N_7080,N_6355,N_5731);
or U7081 (N_7081,N_6362,N_5760);
and U7082 (N_7082,N_6268,N_5629);
xnor U7083 (N_7083,N_5950,N_6232);
nand U7084 (N_7084,N_6007,N_5781);
and U7085 (N_7085,N_6147,N_5984);
nor U7086 (N_7086,N_5949,N_5786);
or U7087 (N_7087,N_5678,N_5602);
xor U7088 (N_7088,N_5789,N_6389);
or U7089 (N_7089,N_6221,N_5739);
and U7090 (N_7090,N_6105,N_6097);
and U7091 (N_7091,N_6372,N_6215);
or U7092 (N_7092,N_5877,N_5810);
nor U7093 (N_7093,N_6184,N_6395);
or U7094 (N_7094,N_6340,N_5843);
or U7095 (N_7095,N_6368,N_6331);
and U7096 (N_7096,N_6212,N_6122);
nor U7097 (N_7097,N_6085,N_5961);
or U7098 (N_7098,N_5821,N_6393);
or U7099 (N_7099,N_6024,N_5809);
nand U7100 (N_7100,N_6332,N_5709);
nor U7101 (N_7101,N_6248,N_5780);
xor U7102 (N_7102,N_5713,N_6324);
and U7103 (N_7103,N_5948,N_6193);
nand U7104 (N_7104,N_6297,N_6005);
or U7105 (N_7105,N_6013,N_5925);
or U7106 (N_7106,N_6315,N_6155);
or U7107 (N_7107,N_6324,N_6061);
and U7108 (N_7108,N_5617,N_6261);
and U7109 (N_7109,N_5739,N_5686);
and U7110 (N_7110,N_5629,N_5980);
and U7111 (N_7111,N_5811,N_6131);
and U7112 (N_7112,N_5874,N_5634);
nand U7113 (N_7113,N_6028,N_6225);
nor U7114 (N_7114,N_6007,N_5818);
nand U7115 (N_7115,N_6169,N_6190);
and U7116 (N_7116,N_5645,N_5925);
xor U7117 (N_7117,N_6263,N_5818);
or U7118 (N_7118,N_5746,N_5752);
and U7119 (N_7119,N_6255,N_6071);
and U7120 (N_7120,N_5896,N_6024);
and U7121 (N_7121,N_5706,N_5944);
nand U7122 (N_7122,N_6257,N_5832);
and U7123 (N_7123,N_6307,N_5792);
xor U7124 (N_7124,N_5749,N_6288);
xor U7125 (N_7125,N_6196,N_5966);
xnor U7126 (N_7126,N_6215,N_6266);
and U7127 (N_7127,N_5946,N_5744);
nand U7128 (N_7128,N_6375,N_6395);
nor U7129 (N_7129,N_6054,N_6193);
xnor U7130 (N_7130,N_6294,N_6353);
xor U7131 (N_7131,N_5743,N_6361);
or U7132 (N_7132,N_6234,N_6390);
xnor U7133 (N_7133,N_5974,N_6235);
nor U7134 (N_7134,N_5914,N_6276);
and U7135 (N_7135,N_5731,N_5964);
or U7136 (N_7136,N_5978,N_5724);
or U7137 (N_7137,N_6218,N_6295);
nor U7138 (N_7138,N_6251,N_6128);
xnor U7139 (N_7139,N_5656,N_5985);
nand U7140 (N_7140,N_5735,N_5893);
xnor U7141 (N_7141,N_5810,N_6066);
and U7142 (N_7142,N_5633,N_6087);
or U7143 (N_7143,N_5774,N_5878);
nand U7144 (N_7144,N_6274,N_6258);
or U7145 (N_7145,N_5989,N_5972);
xor U7146 (N_7146,N_5848,N_6332);
nor U7147 (N_7147,N_6112,N_6038);
or U7148 (N_7148,N_5729,N_5735);
or U7149 (N_7149,N_5937,N_5769);
nand U7150 (N_7150,N_5622,N_6196);
nand U7151 (N_7151,N_5757,N_6038);
or U7152 (N_7152,N_6261,N_5940);
xnor U7153 (N_7153,N_5680,N_6175);
nand U7154 (N_7154,N_5833,N_6390);
or U7155 (N_7155,N_5941,N_5990);
nor U7156 (N_7156,N_6067,N_6005);
nor U7157 (N_7157,N_6300,N_6114);
or U7158 (N_7158,N_6374,N_6380);
or U7159 (N_7159,N_5947,N_5900);
or U7160 (N_7160,N_6050,N_6328);
and U7161 (N_7161,N_5660,N_5738);
xor U7162 (N_7162,N_6086,N_6161);
or U7163 (N_7163,N_5873,N_5818);
xor U7164 (N_7164,N_6031,N_6115);
and U7165 (N_7165,N_5686,N_6164);
or U7166 (N_7166,N_6283,N_6031);
nand U7167 (N_7167,N_5807,N_6152);
or U7168 (N_7168,N_6255,N_5686);
xor U7169 (N_7169,N_5850,N_6306);
and U7170 (N_7170,N_5780,N_6322);
or U7171 (N_7171,N_5974,N_5679);
xor U7172 (N_7172,N_5640,N_6377);
and U7173 (N_7173,N_6322,N_6063);
nand U7174 (N_7174,N_6152,N_5876);
nor U7175 (N_7175,N_6167,N_5853);
xor U7176 (N_7176,N_5754,N_6001);
or U7177 (N_7177,N_6385,N_5670);
and U7178 (N_7178,N_5638,N_5798);
nor U7179 (N_7179,N_6091,N_5794);
xnor U7180 (N_7180,N_5624,N_5805);
nor U7181 (N_7181,N_6082,N_6257);
xor U7182 (N_7182,N_6016,N_5914);
nand U7183 (N_7183,N_5691,N_5651);
or U7184 (N_7184,N_6192,N_6324);
or U7185 (N_7185,N_5966,N_6002);
nand U7186 (N_7186,N_5941,N_5667);
or U7187 (N_7187,N_5879,N_5685);
nor U7188 (N_7188,N_5685,N_6202);
and U7189 (N_7189,N_6292,N_6011);
and U7190 (N_7190,N_5837,N_6000);
xor U7191 (N_7191,N_6022,N_5956);
nor U7192 (N_7192,N_5836,N_6298);
or U7193 (N_7193,N_6322,N_6128);
nand U7194 (N_7194,N_5990,N_5727);
xor U7195 (N_7195,N_6051,N_5971);
or U7196 (N_7196,N_5683,N_6300);
or U7197 (N_7197,N_6043,N_5698);
nor U7198 (N_7198,N_6093,N_6379);
nor U7199 (N_7199,N_5798,N_6209);
nor U7200 (N_7200,N_6689,N_6530);
or U7201 (N_7201,N_7114,N_6639);
nor U7202 (N_7202,N_6946,N_6407);
nor U7203 (N_7203,N_6536,N_6429);
or U7204 (N_7204,N_6507,N_6494);
xor U7205 (N_7205,N_6665,N_6666);
nor U7206 (N_7206,N_6551,N_6858);
nand U7207 (N_7207,N_6515,N_6539);
xnor U7208 (N_7208,N_7050,N_6955);
nand U7209 (N_7209,N_6403,N_6546);
and U7210 (N_7210,N_6445,N_6766);
nand U7211 (N_7211,N_6464,N_7074);
and U7212 (N_7212,N_6710,N_6805);
nor U7213 (N_7213,N_7036,N_6757);
or U7214 (N_7214,N_6457,N_7132);
or U7215 (N_7215,N_6756,N_7080);
xor U7216 (N_7216,N_7161,N_6960);
nor U7217 (N_7217,N_6884,N_6453);
xnor U7218 (N_7218,N_6609,N_6888);
nor U7219 (N_7219,N_6881,N_6613);
nand U7220 (N_7220,N_7109,N_6486);
nor U7221 (N_7221,N_6942,N_7154);
or U7222 (N_7222,N_6557,N_6779);
nor U7223 (N_7223,N_7006,N_6706);
xor U7224 (N_7224,N_6840,N_6599);
xnor U7225 (N_7225,N_6619,N_6450);
nor U7226 (N_7226,N_6852,N_6480);
nand U7227 (N_7227,N_6508,N_6413);
xnor U7228 (N_7228,N_6424,N_6459);
or U7229 (N_7229,N_6427,N_6820);
xor U7230 (N_7230,N_7060,N_6969);
nor U7231 (N_7231,N_6502,N_6650);
and U7232 (N_7232,N_6673,N_6719);
nand U7233 (N_7233,N_6487,N_6535);
nor U7234 (N_7234,N_6987,N_7140);
xor U7235 (N_7235,N_6700,N_7082);
and U7236 (N_7236,N_7097,N_6493);
or U7237 (N_7237,N_6560,N_6793);
or U7238 (N_7238,N_6895,N_6642);
nor U7239 (N_7239,N_6923,N_6981);
or U7240 (N_7240,N_6477,N_6596);
xnor U7241 (N_7241,N_6688,N_6498);
or U7242 (N_7242,N_7093,N_6762);
nor U7243 (N_7243,N_6683,N_6777);
or U7244 (N_7244,N_7033,N_6815);
and U7245 (N_7245,N_6782,N_7106);
or U7246 (N_7246,N_7111,N_6824);
nor U7247 (N_7247,N_6721,N_7027);
and U7248 (N_7248,N_6918,N_6564);
nor U7249 (N_7249,N_6513,N_6423);
nand U7250 (N_7250,N_6913,N_7178);
xor U7251 (N_7251,N_6412,N_6811);
or U7252 (N_7252,N_7049,N_6677);
nor U7253 (N_7253,N_6476,N_6416);
xor U7254 (N_7254,N_6890,N_6853);
and U7255 (N_7255,N_6543,N_6602);
nand U7256 (N_7256,N_6587,N_6966);
nand U7257 (N_7257,N_6442,N_7020);
or U7258 (N_7258,N_6621,N_6780);
nand U7259 (N_7259,N_7069,N_6695);
or U7260 (N_7260,N_7090,N_7122);
xor U7261 (N_7261,N_6556,N_6626);
xnor U7262 (N_7262,N_6875,N_6474);
or U7263 (N_7263,N_6746,N_6522);
nor U7264 (N_7264,N_6750,N_7126);
or U7265 (N_7265,N_6951,N_6723);
xnor U7266 (N_7266,N_6934,N_6916);
nand U7267 (N_7267,N_6774,N_6735);
and U7268 (N_7268,N_7046,N_6646);
nor U7269 (N_7269,N_6702,N_6404);
xor U7270 (N_7270,N_6839,N_6426);
or U7271 (N_7271,N_6465,N_6542);
nor U7272 (N_7272,N_7192,N_6973);
xnor U7273 (N_7273,N_7019,N_6940);
nor U7274 (N_7274,N_6889,N_7177);
nor U7275 (N_7275,N_6899,N_7068);
or U7276 (N_7276,N_6819,N_7117);
nand U7277 (N_7277,N_7149,N_6926);
or U7278 (N_7278,N_7040,N_7044);
nand U7279 (N_7279,N_6958,N_7175);
nor U7280 (N_7280,N_6860,N_6791);
xnor U7281 (N_7281,N_7061,N_6527);
xnor U7282 (N_7282,N_7143,N_7145);
and U7283 (N_7283,N_7130,N_7001);
nor U7284 (N_7284,N_7197,N_6990);
nand U7285 (N_7285,N_6849,N_6526);
or U7286 (N_7286,N_7063,N_7039);
or U7287 (N_7287,N_6767,N_6991);
or U7288 (N_7288,N_6730,N_6797);
and U7289 (N_7289,N_7008,N_7113);
nor U7290 (N_7290,N_6441,N_6796);
nand U7291 (N_7291,N_6533,N_6680);
xnor U7292 (N_7292,N_6927,N_6548);
and U7293 (N_7293,N_6428,N_6577);
nor U7294 (N_7294,N_7081,N_7042);
or U7295 (N_7295,N_6961,N_6864);
or U7296 (N_7296,N_6994,N_6885);
or U7297 (N_7297,N_6794,N_6947);
nand U7298 (N_7298,N_6967,N_6489);
nand U7299 (N_7299,N_6630,N_6469);
or U7300 (N_7300,N_6622,N_6595);
xnor U7301 (N_7301,N_7142,N_7084);
nor U7302 (N_7302,N_6669,N_6816);
or U7303 (N_7303,N_6826,N_6488);
nor U7304 (N_7304,N_6549,N_6582);
and U7305 (N_7305,N_6971,N_6709);
and U7306 (N_7306,N_6830,N_6759);
or U7307 (N_7307,N_6785,N_6886);
nor U7308 (N_7308,N_6541,N_6733);
nand U7309 (N_7309,N_6635,N_6936);
or U7310 (N_7310,N_7191,N_6985);
nand U7311 (N_7311,N_6804,N_6753);
nor U7312 (N_7312,N_7184,N_7155);
xnor U7313 (N_7313,N_6847,N_6623);
or U7314 (N_7314,N_6789,N_7195);
or U7315 (N_7315,N_7171,N_7102);
or U7316 (N_7316,N_6662,N_6932);
nand U7317 (N_7317,N_6657,N_6887);
and U7318 (N_7318,N_6908,N_6633);
nand U7319 (N_7319,N_7123,N_7173);
nor U7320 (N_7320,N_6846,N_6484);
nor U7321 (N_7321,N_6438,N_6935);
xor U7322 (N_7322,N_6965,N_7116);
and U7323 (N_7323,N_6589,N_6712);
or U7324 (N_7324,N_6612,N_6503);
and U7325 (N_7325,N_6795,N_7104);
xnor U7326 (N_7326,N_7165,N_7013);
nor U7327 (N_7327,N_6892,N_7185);
nand U7328 (N_7328,N_6628,N_7089);
nand U7329 (N_7329,N_6871,N_7190);
nand U7330 (N_7330,N_6866,N_6655);
or U7331 (N_7331,N_7196,N_6863);
nor U7332 (N_7332,N_6415,N_6620);
or U7333 (N_7333,N_6638,N_6959);
nand U7334 (N_7334,N_6974,N_6996);
and U7335 (N_7335,N_6798,N_7048);
xnor U7336 (N_7336,N_7189,N_6829);
or U7337 (N_7337,N_7032,N_7099);
xnor U7338 (N_7338,N_6500,N_6763);
and U7339 (N_7339,N_6781,N_6914);
and U7340 (N_7340,N_6550,N_6714);
nand U7341 (N_7341,N_6808,N_6525);
or U7342 (N_7342,N_6993,N_6873);
and U7343 (N_7343,N_6732,N_6983);
nand U7344 (N_7344,N_7086,N_6768);
or U7345 (N_7345,N_6904,N_6933);
nand U7346 (N_7346,N_6571,N_6705);
nand U7347 (N_7347,N_6406,N_7139);
nor U7348 (N_7348,N_7057,N_6722);
nand U7349 (N_7349,N_7166,N_6569);
xnor U7350 (N_7350,N_6401,N_6769);
xnor U7351 (N_7351,N_6809,N_6760);
nand U7352 (N_7352,N_6472,N_6580);
and U7353 (N_7353,N_7101,N_6828);
nor U7354 (N_7354,N_7121,N_7026);
nor U7355 (N_7355,N_6685,N_6775);
and U7356 (N_7356,N_6982,N_7129);
nor U7357 (N_7357,N_6636,N_7159);
nor U7358 (N_7358,N_7172,N_6470);
nand U7359 (N_7359,N_7125,N_7188);
and U7360 (N_7360,N_7124,N_7078);
or U7361 (N_7361,N_6510,N_6456);
or U7362 (N_7362,N_6772,N_7127);
or U7363 (N_7363,N_6497,N_6707);
or U7364 (N_7364,N_6574,N_7062);
nand U7365 (N_7365,N_6962,N_6418);
nor U7366 (N_7366,N_6739,N_6893);
xnor U7367 (N_7367,N_7029,N_6856);
or U7368 (N_7368,N_6976,N_6562);
nand U7369 (N_7369,N_6745,N_6431);
or U7370 (N_7370,N_7077,N_6499);
nand U7371 (N_7371,N_7164,N_7193);
xnor U7372 (N_7372,N_6443,N_6479);
xnor U7373 (N_7373,N_6854,N_7181);
and U7374 (N_7374,N_7131,N_7056);
and U7375 (N_7375,N_7054,N_6701);
nor U7376 (N_7376,N_6614,N_6693);
or U7377 (N_7377,N_6440,N_6667);
xnor U7378 (N_7378,N_7141,N_7169);
nand U7379 (N_7379,N_6468,N_6572);
nor U7380 (N_7380,N_7180,N_6868);
nor U7381 (N_7381,N_6656,N_7176);
nor U7382 (N_7382,N_7085,N_6696);
and U7383 (N_7383,N_6601,N_6736);
nand U7384 (N_7384,N_6411,N_6570);
nor U7385 (N_7385,N_6616,N_6925);
and U7386 (N_7386,N_6678,N_6711);
or U7387 (N_7387,N_6979,N_6617);
and U7388 (N_7388,N_6867,N_6862);
xnor U7389 (N_7389,N_6605,N_7105);
and U7390 (N_7390,N_6608,N_6783);
and U7391 (N_7391,N_7035,N_6409);
nand U7392 (N_7392,N_6728,N_6747);
nand U7393 (N_7393,N_7138,N_6697);
or U7394 (N_7394,N_7134,N_7043);
nor U7395 (N_7395,N_6910,N_6752);
xor U7396 (N_7396,N_6716,N_6740);
and U7397 (N_7397,N_6851,N_6674);
and U7398 (N_7398,N_7004,N_6975);
nand U7399 (N_7399,N_6640,N_6603);
xor U7400 (N_7400,N_7094,N_6691);
and U7401 (N_7401,N_7148,N_6654);
and U7402 (N_7402,N_6754,N_6578);
nand U7403 (N_7403,N_6482,N_6842);
or U7404 (N_7404,N_7010,N_6417);
nand U7405 (N_7405,N_6818,N_6988);
nor U7406 (N_7406,N_6490,N_6911);
xor U7407 (N_7407,N_6773,N_6540);
and U7408 (N_7408,N_6585,N_6724);
nand U7409 (N_7409,N_6604,N_6405);
and U7410 (N_7410,N_6668,N_6806);
nor U7411 (N_7411,N_6496,N_6637);
and U7412 (N_7412,N_6624,N_6749);
or U7413 (N_7413,N_7016,N_6672);
nor U7414 (N_7414,N_6410,N_6447);
nand U7415 (N_7415,N_6518,N_7073);
nor U7416 (N_7416,N_6670,N_7014);
nor U7417 (N_7417,N_6523,N_6565);
nor U7418 (N_7418,N_6717,N_7199);
and U7419 (N_7419,N_6869,N_6992);
and U7420 (N_7420,N_6963,N_6491);
or U7421 (N_7421,N_6896,N_7064);
xor U7422 (N_7422,N_7112,N_7153);
and U7423 (N_7423,N_6586,N_6653);
or U7424 (N_7424,N_6634,N_7087);
or U7425 (N_7425,N_6425,N_6687);
nand U7426 (N_7426,N_6454,N_6611);
or U7427 (N_7427,N_6776,N_6742);
and U7428 (N_7428,N_6843,N_6627);
and U7429 (N_7429,N_6787,N_7133);
or U7430 (N_7430,N_6434,N_6520);
or U7431 (N_7431,N_6692,N_6400);
nor U7432 (N_7432,N_7168,N_6583);
and U7433 (N_7433,N_6592,N_6483);
nor U7434 (N_7434,N_6827,N_6597);
nor U7435 (N_7435,N_6610,N_7058);
or U7436 (N_7436,N_6986,N_7152);
xor U7437 (N_7437,N_6978,N_7002);
nand U7438 (N_7438,N_6699,N_6641);
and U7439 (N_7439,N_6836,N_6439);
or U7440 (N_7440,N_7051,N_7187);
nand U7441 (N_7441,N_6770,N_6831);
nor U7442 (N_7442,N_7047,N_7136);
or U7443 (N_7443,N_7071,N_7135);
and U7444 (N_7444,N_6584,N_6694);
nand U7445 (N_7445,N_6481,N_6519);
nor U7446 (N_7446,N_6949,N_6652);
or U7447 (N_7447,N_6765,N_7198);
and U7448 (N_7448,N_6944,N_6492);
or U7449 (N_7449,N_6743,N_6984);
and U7450 (N_7450,N_6531,N_6938);
xor U7451 (N_7451,N_6715,N_7118);
or U7452 (N_7452,N_6485,N_6581);
and U7453 (N_7453,N_6600,N_7182);
nand U7454 (N_7454,N_6919,N_6865);
nor U7455 (N_7455,N_6807,N_6544);
nor U7456 (N_7456,N_6822,N_6857);
nor U7457 (N_7457,N_6408,N_6738);
and U7458 (N_7458,N_6941,N_6803);
and U7459 (N_7459,N_6894,N_7146);
nor U7460 (N_7460,N_6729,N_6686);
xnor U7461 (N_7461,N_7076,N_6467);
xor U7462 (N_7462,N_7151,N_6575);
nor U7463 (N_7463,N_7167,N_6660);
and U7464 (N_7464,N_6861,N_7179);
and U7465 (N_7465,N_6924,N_7018);
nor U7466 (N_7466,N_6931,N_6997);
or U7467 (N_7467,N_6552,N_6566);
or U7468 (N_7468,N_6594,N_6471);
or U7469 (N_7469,N_6877,N_7000);
nand U7470 (N_7470,N_6436,N_6505);
or U7471 (N_7471,N_7059,N_6506);
and U7472 (N_7472,N_6900,N_7137);
xnor U7473 (N_7473,N_6661,N_7023);
or U7474 (N_7474,N_7003,N_6547);
or U7475 (N_7475,N_6573,N_6648);
or U7476 (N_7476,N_7045,N_6989);
nor U7477 (N_7477,N_7194,N_6649);
nor U7478 (N_7478,N_7092,N_6524);
and U7479 (N_7479,N_6598,N_6664);
and U7480 (N_7480,N_6446,N_6554);
nand U7481 (N_7481,N_6907,N_6511);
nor U7482 (N_7482,N_6943,N_6870);
xnor U7483 (N_7483,N_6948,N_6629);
and U7484 (N_7484,N_6658,N_6802);
or U7485 (N_7485,N_7186,N_7066);
nor U7486 (N_7486,N_7147,N_6891);
xor U7487 (N_7487,N_7021,N_6837);
xnor U7488 (N_7488,N_6731,N_6844);
xor U7489 (N_7489,N_6880,N_6521);
and U7490 (N_7490,N_7156,N_7028);
nor U7491 (N_7491,N_6593,N_6473);
nand U7492 (N_7492,N_6420,N_6449);
xor U7493 (N_7493,N_7024,N_6579);
xnor U7494 (N_7494,N_6751,N_6957);
nand U7495 (N_7495,N_6625,N_7055);
nand U7496 (N_7496,N_6901,N_6906);
or U7497 (N_7497,N_6495,N_6461);
or U7498 (N_7498,N_6872,N_6537);
nand U7499 (N_7499,N_6437,N_6455);
or U7500 (N_7500,N_7005,N_7065);
nor U7501 (N_7501,N_7144,N_7012);
nand U7502 (N_7502,N_6433,N_6466);
xnor U7503 (N_7503,N_6703,N_6823);
and U7504 (N_7504,N_6771,N_6509);
or U7505 (N_7505,N_6671,N_6972);
and U7506 (N_7506,N_6812,N_6929);
nand U7507 (N_7507,N_6720,N_7157);
or U7508 (N_7508,N_6644,N_6953);
or U7509 (N_7509,N_6834,N_6778);
or U7510 (N_7510,N_7072,N_6708);
and U7511 (N_7511,N_7070,N_6528);
or U7512 (N_7512,N_7041,N_7037);
and U7513 (N_7513,N_6792,N_6725);
and U7514 (N_7514,N_6555,N_7053);
xor U7515 (N_7515,N_6419,N_6448);
xnor U7516 (N_7516,N_6645,N_6930);
or U7517 (N_7517,N_6801,N_6463);
or U7518 (N_7518,N_6761,N_6713);
or U7519 (N_7519,N_7038,N_6748);
or U7520 (N_7520,N_6444,N_6813);
and U7521 (N_7521,N_6859,N_7017);
and U7522 (N_7522,N_6838,N_6451);
nor U7523 (N_7523,N_6841,N_6647);
nor U7524 (N_7524,N_6920,N_6952);
xor U7525 (N_7525,N_6800,N_7022);
nand U7526 (N_7526,N_6675,N_7128);
nor U7527 (N_7527,N_6939,N_6897);
nor U7528 (N_7528,N_6538,N_6999);
or U7529 (N_7529,N_6903,N_7083);
nand U7530 (N_7530,N_6741,N_6825);
and U7531 (N_7531,N_6727,N_6788);
nor U7532 (N_7532,N_6898,N_7079);
xnor U7533 (N_7533,N_6790,N_6902);
xor U7534 (N_7534,N_6917,N_6452);
and U7535 (N_7535,N_6590,N_6529);
nor U7536 (N_7536,N_6845,N_6921);
or U7537 (N_7537,N_7075,N_6977);
nor U7538 (N_7538,N_6882,N_6651);
nor U7539 (N_7539,N_6821,N_6964);
and U7540 (N_7540,N_7031,N_6682);
nand U7541 (N_7541,N_6567,N_6501);
or U7542 (N_7542,N_6876,N_6734);
or U7543 (N_7543,N_7025,N_6832);
and U7544 (N_7544,N_6737,N_7011);
and U7545 (N_7545,N_7119,N_6517);
or U7546 (N_7546,N_6937,N_6970);
nand U7547 (N_7547,N_6786,N_7160);
nor U7548 (N_7548,N_6618,N_7158);
nand U7549 (N_7549,N_6718,N_6588);
nand U7550 (N_7550,N_6534,N_6690);
or U7551 (N_7551,N_6478,N_7052);
nand U7552 (N_7552,N_6460,N_7067);
nand U7553 (N_7553,N_7103,N_7034);
nand U7554 (N_7554,N_6784,N_6606);
or U7555 (N_7555,N_6659,N_6817);
or U7556 (N_7556,N_6475,N_6950);
xnor U7557 (N_7557,N_7150,N_6545);
nand U7558 (N_7558,N_6512,N_6855);
xnor U7559 (N_7559,N_7030,N_6912);
nand U7560 (N_7560,N_6421,N_6402);
nand U7561 (N_7561,N_7120,N_6995);
nor U7562 (N_7562,N_6504,N_6631);
and U7563 (N_7563,N_6532,N_7183);
nor U7564 (N_7564,N_6615,N_7007);
or U7565 (N_7565,N_6435,N_6833);
nand U7566 (N_7566,N_6432,N_6848);
nor U7567 (N_7567,N_7100,N_6643);
and U7568 (N_7568,N_6883,N_7091);
xnor U7569 (N_7569,N_7174,N_6799);
or U7570 (N_7570,N_7162,N_6663);
nor U7571 (N_7571,N_6878,N_6905);
or U7572 (N_7572,N_7110,N_6956);
or U7573 (N_7573,N_6922,N_6698);
nor U7574 (N_7574,N_6563,N_7096);
and U7575 (N_7575,N_6909,N_6558);
nor U7576 (N_7576,N_7088,N_6850);
or U7577 (N_7577,N_6559,N_7115);
and U7578 (N_7578,N_6764,N_6755);
xor U7579 (N_7579,N_6998,N_6561);
or U7580 (N_7580,N_7108,N_6568);
nand U7581 (N_7581,N_6514,N_6430);
nor U7582 (N_7582,N_7163,N_6726);
and U7583 (N_7583,N_6945,N_6810);
nand U7584 (N_7584,N_6458,N_6553);
nand U7585 (N_7585,N_6576,N_7095);
nand U7586 (N_7586,N_6422,N_6758);
and U7587 (N_7587,N_7098,N_6835);
nand U7588 (N_7588,N_6632,N_6968);
xor U7589 (N_7589,N_6462,N_6414);
nand U7590 (N_7590,N_6915,N_6681);
nor U7591 (N_7591,N_7107,N_7009);
and U7592 (N_7592,N_7015,N_6684);
xnor U7593 (N_7593,N_6874,N_6879);
or U7594 (N_7594,N_6954,N_6928);
or U7595 (N_7595,N_6607,N_6516);
xor U7596 (N_7596,N_6814,N_6591);
xor U7597 (N_7597,N_6744,N_6676);
nand U7598 (N_7598,N_6679,N_6980);
nor U7599 (N_7599,N_6704,N_7170);
xnor U7600 (N_7600,N_6633,N_6497);
or U7601 (N_7601,N_6695,N_7138);
and U7602 (N_7602,N_6434,N_6804);
nor U7603 (N_7603,N_6721,N_7086);
nand U7604 (N_7604,N_6791,N_6812);
nand U7605 (N_7605,N_6482,N_6692);
or U7606 (N_7606,N_6564,N_6430);
or U7607 (N_7607,N_6864,N_6725);
nor U7608 (N_7608,N_7104,N_6967);
nand U7609 (N_7609,N_6656,N_6615);
nor U7610 (N_7610,N_6551,N_6411);
nand U7611 (N_7611,N_6683,N_6782);
or U7612 (N_7612,N_7136,N_7034);
or U7613 (N_7613,N_6505,N_7116);
or U7614 (N_7614,N_6951,N_6546);
xor U7615 (N_7615,N_7092,N_6558);
xor U7616 (N_7616,N_6715,N_6748);
nor U7617 (N_7617,N_6578,N_7152);
nor U7618 (N_7618,N_6557,N_7019);
nor U7619 (N_7619,N_6430,N_6954);
nor U7620 (N_7620,N_6761,N_6843);
nor U7621 (N_7621,N_6757,N_6571);
nand U7622 (N_7622,N_6929,N_7019);
xor U7623 (N_7623,N_6670,N_7021);
xor U7624 (N_7624,N_6856,N_7025);
nand U7625 (N_7625,N_7103,N_6601);
nor U7626 (N_7626,N_6987,N_6448);
and U7627 (N_7627,N_6928,N_7157);
nor U7628 (N_7628,N_6611,N_7010);
and U7629 (N_7629,N_6721,N_6983);
or U7630 (N_7630,N_7064,N_6976);
xor U7631 (N_7631,N_6728,N_7059);
and U7632 (N_7632,N_6567,N_6523);
nand U7633 (N_7633,N_6735,N_6575);
nor U7634 (N_7634,N_6916,N_6823);
nor U7635 (N_7635,N_7102,N_7076);
nor U7636 (N_7636,N_6869,N_6802);
and U7637 (N_7637,N_7055,N_6524);
nand U7638 (N_7638,N_6958,N_6481);
nor U7639 (N_7639,N_6795,N_6742);
nor U7640 (N_7640,N_6526,N_6554);
xor U7641 (N_7641,N_7095,N_6665);
xor U7642 (N_7642,N_6809,N_6549);
xor U7643 (N_7643,N_7068,N_7107);
or U7644 (N_7644,N_6722,N_6509);
nor U7645 (N_7645,N_6723,N_6760);
and U7646 (N_7646,N_6721,N_6684);
nand U7647 (N_7647,N_6768,N_6821);
nand U7648 (N_7648,N_6627,N_7154);
and U7649 (N_7649,N_6513,N_6983);
nand U7650 (N_7650,N_7153,N_6977);
and U7651 (N_7651,N_6741,N_6727);
nand U7652 (N_7652,N_7071,N_6828);
nand U7653 (N_7653,N_7124,N_6841);
and U7654 (N_7654,N_6582,N_6863);
nand U7655 (N_7655,N_6572,N_7109);
and U7656 (N_7656,N_6655,N_6463);
xnor U7657 (N_7657,N_6412,N_6692);
xor U7658 (N_7658,N_7062,N_6477);
nor U7659 (N_7659,N_6921,N_6674);
nor U7660 (N_7660,N_7105,N_7039);
or U7661 (N_7661,N_6815,N_6826);
xnor U7662 (N_7662,N_7000,N_7156);
nor U7663 (N_7663,N_6894,N_7160);
nor U7664 (N_7664,N_6788,N_6591);
nor U7665 (N_7665,N_7191,N_7113);
nor U7666 (N_7666,N_7099,N_6511);
and U7667 (N_7667,N_6581,N_6402);
nor U7668 (N_7668,N_6486,N_6606);
nor U7669 (N_7669,N_6545,N_6899);
nand U7670 (N_7670,N_6977,N_6793);
xnor U7671 (N_7671,N_6503,N_6934);
xnor U7672 (N_7672,N_6631,N_6467);
and U7673 (N_7673,N_6637,N_6452);
xnor U7674 (N_7674,N_6829,N_6952);
nand U7675 (N_7675,N_6609,N_7091);
nand U7676 (N_7676,N_6527,N_6732);
and U7677 (N_7677,N_7189,N_6779);
nor U7678 (N_7678,N_6549,N_6908);
and U7679 (N_7679,N_6464,N_6726);
nor U7680 (N_7680,N_7194,N_6812);
xor U7681 (N_7681,N_7083,N_6704);
xor U7682 (N_7682,N_6855,N_6858);
or U7683 (N_7683,N_6892,N_6877);
or U7684 (N_7684,N_6417,N_6514);
xor U7685 (N_7685,N_6550,N_6745);
or U7686 (N_7686,N_6982,N_6690);
and U7687 (N_7687,N_6885,N_6453);
nor U7688 (N_7688,N_6633,N_6907);
or U7689 (N_7689,N_6486,N_6616);
or U7690 (N_7690,N_6796,N_6817);
and U7691 (N_7691,N_6409,N_6745);
nand U7692 (N_7692,N_7144,N_6917);
nor U7693 (N_7693,N_6721,N_6549);
nand U7694 (N_7694,N_6749,N_7085);
xnor U7695 (N_7695,N_6882,N_6603);
and U7696 (N_7696,N_6896,N_6426);
nor U7697 (N_7697,N_6496,N_6536);
nand U7698 (N_7698,N_6688,N_6961);
nor U7699 (N_7699,N_7032,N_6775);
nor U7700 (N_7700,N_6445,N_6507);
and U7701 (N_7701,N_6675,N_6431);
nor U7702 (N_7702,N_6415,N_6991);
or U7703 (N_7703,N_6565,N_6659);
or U7704 (N_7704,N_7124,N_6597);
nor U7705 (N_7705,N_6492,N_6528);
nand U7706 (N_7706,N_6958,N_6944);
and U7707 (N_7707,N_6669,N_6731);
xor U7708 (N_7708,N_6715,N_7134);
and U7709 (N_7709,N_7178,N_6852);
nor U7710 (N_7710,N_6651,N_6789);
and U7711 (N_7711,N_7138,N_6637);
and U7712 (N_7712,N_6929,N_6993);
and U7713 (N_7713,N_6861,N_6669);
nor U7714 (N_7714,N_7119,N_6701);
nor U7715 (N_7715,N_6815,N_6606);
nor U7716 (N_7716,N_6668,N_6962);
and U7717 (N_7717,N_6492,N_7058);
or U7718 (N_7718,N_6890,N_6858);
nor U7719 (N_7719,N_6527,N_6865);
or U7720 (N_7720,N_6555,N_7000);
nand U7721 (N_7721,N_6791,N_6856);
nor U7722 (N_7722,N_6682,N_7081);
nand U7723 (N_7723,N_6650,N_7122);
nor U7724 (N_7724,N_6673,N_7083);
or U7725 (N_7725,N_7049,N_6556);
nand U7726 (N_7726,N_6702,N_6808);
nand U7727 (N_7727,N_6822,N_6495);
and U7728 (N_7728,N_6605,N_6439);
xor U7729 (N_7729,N_6680,N_6844);
and U7730 (N_7730,N_6931,N_6595);
or U7731 (N_7731,N_6532,N_6793);
or U7732 (N_7732,N_6919,N_6836);
xnor U7733 (N_7733,N_7065,N_6922);
and U7734 (N_7734,N_6458,N_6867);
and U7735 (N_7735,N_6653,N_7001);
xnor U7736 (N_7736,N_6938,N_7085);
and U7737 (N_7737,N_6682,N_6914);
nor U7738 (N_7738,N_7179,N_6754);
nand U7739 (N_7739,N_6514,N_6891);
nand U7740 (N_7740,N_6964,N_6619);
xnor U7741 (N_7741,N_7056,N_6475);
xnor U7742 (N_7742,N_6878,N_6966);
nor U7743 (N_7743,N_7009,N_6535);
nand U7744 (N_7744,N_7190,N_6783);
and U7745 (N_7745,N_7037,N_6401);
nand U7746 (N_7746,N_6567,N_6725);
xor U7747 (N_7747,N_6542,N_6610);
nor U7748 (N_7748,N_6973,N_7060);
or U7749 (N_7749,N_6919,N_6573);
xor U7750 (N_7750,N_6484,N_6607);
nand U7751 (N_7751,N_6803,N_6842);
nor U7752 (N_7752,N_6463,N_6612);
xor U7753 (N_7753,N_6430,N_6708);
xnor U7754 (N_7754,N_6778,N_6730);
or U7755 (N_7755,N_7175,N_6746);
nand U7756 (N_7756,N_6861,N_6993);
nand U7757 (N_7757,N_7045,N_6976);
nor U7758 (N_7758,N_6796,N_6942);
nor U7759 (N_7759,N_6748,N_7116);
nand U7760 (N_7760,N_7080,N_6515);
and U7761 (N_7761,N_6461,N_6824);
xnor U7762 (N_7762,N_6802,N_6940);
nor U7763 (N_7763,N_7199,N_6720);
and U7764 (N_7764,N_7073,N_7096);
nor U7765 (N_7765,N_6739,N_7168);
or U7766 (N_7766,N_6869,N_6714);
nand U7767 (N_7767,N_6864,N_6887);
nor U7768 (N_7768,N_7071,N_6432);
nor U7769 (N_7769,N_6743,N_6988);
and U7770 (N_7770,N_6649,N_7021);
xnor U7771 (N_7771,N_7003,N_6903);
or U7772 (N_7772,N_6693,N_7107);
or U7773 (N_7773,N_7138,N_6780);
and U7774 (N_7774,N_6626,N_6766);
and U7775 (N_7775,N_6721,N_6994);
nor U7776 (N_7776,N_6700,N_6617);
nor U7777 (N_7777,N_6509,N_6700);
nor U7778 (N_7778,N_7094,N_7108);
nor U7779 (N_7779,N_6517,N_6433);
nor U7780 (N_7780,N_6932,N_6635);
or U7781 (N_7781,N_6973,N_6673);
and U7782 (N_7782,N_7133,N_6658);
or U7783 (N_7783,N_6514,N_6455);
nor U7784 (N_7784,N_7066,N_7016);
nand U7785 (N_7785,N_6868,N_7117);
or U7786 (N_7786,N_6474,N_6905);
or U7787 (N_7787,N_6609,N_7093);
nor U7788 (N_7788,N_7186,N_6895);
nand U7789 (N_7789,N_7131,N_6903);
xnor U7790 (N_7790,N_6546,N_6786);
xnor U7791 (N_7791,N_6605,N_6908);
nand U7792 (N_7792,N_6925,N_7049);
xnor U7793 (N_7793,N_7098,N_6690);
nand U7794 (N_7794,N_7017,N_6642);
xnor U7795 (N_7795,N_6963,N_6821);
or U7796 (N_7796,N_6569,N_6764);
nor U7797 (N_7797,N_6964,N_6483);
nor U7798 (N_7798,N_6950,N_6980);
or U7799 (N_7799,N_7165,N_6407);
and U7800 (N_7800,N_7188,N_7185);
nand U7801 (N_7801,N_6806,N_6852);
nor U7802 (N_7802,N_6741,N_6565);
nor U7803 (N_7803,N_6684,N_6577);
nand U7804 (N_7804,N_6579,N_6660);
or U7805 (N_7805,N_7113,N_6974);
and U7806 (N_7806,N_6615,N_6911);
and U7807 (N_7807,N_6673,N_6600);
xor U7808 (N_7808,N_6792,N_6843);
or U7809 (N_7809,N_6649,N_6576);
or U7810 (N_7810,N_6462,N_6851);
nor U7811 (N_7811,N_6851,N_6642);
xnor U7812 (N_7812,N_6905,N_7188);
and U7813 (N_7813,N_6968,N_6563);
xor U7814 (N_7814,N_6552,N_6888);
xnor U7815 (N_7815,N_7068,N_6483);
nor U7816 (N_7816,N_6875,N_7178);
nand U7817 (N_7817,N_7073,N_7023);
nand U7818 (N_7818,N_6753,N_6509);
or U7819 (N_7819,N_6749,N_6471);
nor U7820 (N_7820,N_7135,N_6402);
or U7821 (N_7821,N_6820,N_7031);
nor U7822 (N_7822,N_7073,N_7063);
nor U7823 (N_7823,N_6481,N_6796);
or U7824 (N_7824,N_6863,N_7073);
xor U7825 (N_7825,N_6522,N_6684);
nand U7826 (N_7826,N_6954,N_6579);
nand U7827 (N_7827,N_6748,N_6581);
and U7828 (N_7828,N_6848,N_6844);
and U7829 (N_7829,N_7128,N_6532);
or U7830 (N_7830,N_6977,N_6887);
xor U7831 (N_7831,N_6708,N_6583);
nor U7832 (N_7832,N_7054,N_7140);
or U7833 (N_7833,N_6807,N_6442);
or U7834 (N_7834,N_6910,N_7117);
or U7835 (N_7835,N_6531,N_6629);
nand U7836 (N_7836,N_6597,N_7103);
and U7837 (N_7837,N_7095,N_7080);
and U7838 (N_7838,N_6916,N_6895);
or U7839 (N_7839,N_6994,N_6525);
nor U7840 (N_7840,N_6855,N_6659);
and U7841 (N_7841,N_6945,N_7104);
xnor U7842 (N_7842,N_6517,N_6877);
nor U7843 (N_7843,N_7164,N_7108);
and U7844 (N_7844,N_6711,N_7165);
or U7845 (N_7845,N_6862,N_6551);
xnor U7846 (N_7846,N_6427,N_6910);
and U7847 (N_7847,N_7156,N_7008);
and U7848 (N_7848,N_6413,N_6493);
and U7849 (N_7849,N_6684,N_6647);
xnor U7850 (N_7850,N_6822,N_6513);
xor U7851 (N_7851,N_7001,N_6930);
nand U7852 (N_7852,N_7069,N_6794);
nor U7853 (N_7853,N_6860,N_6426);
xor U7854 (N_7854,N_6574,N_7109);
or U7855 (N_7855,N_6677,N_7051);
nand U7856 (N_7856,N_7103,N_6750);
nand U7857 (N_7857,N_7049,N_7185);
and U7858 (N_7858,N_7055,N_6651);
nor U7859 (N_7859,N_6454,N_6460);
and U7860 (N_7860,N_6948,N_6989);
nor U7861 (N_7861,N_6473,N_7051);
nor U7862 (N_7862,N_7118,N_6796);
xnor U7863 (N_7863,N_6450,N_6777);
nor U7864 (N_7864,N_6566,N_7064);
nand U7865 (N_7865,N_6455,N_6874);
or U7866 (N_7866,N_6863,N_6818);
nand U7867 (N_7867,N_6742,N_6606);
xnor U7868 (N_7868,N_6818,N_6789);
or U7869 (N_7869,N_6925,N_6538);
nor U7870 (N_7870,N_7018,N_6896);
nand U7871 (N_7871,N_6930,N_7177);
or U7872 (N_7872,N_6510,N_6812);
nor U7873 (N_7873,N_6888,N_6817);
nor U7874 (N_7874,N_6704,N_6803);
nor U7875 (N_7875,N_6865,N_6905);
or U7876 (N_7876,N_6480,N_6547);
nor U7877 (N_7877,N_6561,N_6569);
nor U7878 (N_7878,N_6997,N_7042);
and U7879 (N_7879,N_6834,N_6633);
nor U7880 (N_7880,N_7100,N_7108);
xnor U7881 (N_7881,N_7084,N_6559);
or U7882 (N_7882,N_6706,N_7103);
and U7883 (N_7883,N_7122,N_6486);
nor U7884 (N_7884,N_6965,N_7087);
nand U7885 (N_7885,N_6577,N_6820);
xnor U7886 (N_7886,N_6961,N_6777);
or U7887 (N_7887,N_6872,N_7135);
nand U7888 (N_7888,N_7170,N_6430);
nor U7889 (N_7889,N_7033,N_6811);
nand U7890 (N_7890,N_6498,N_7016);
nor U7891 (N_7891,N_6807,N_6618);
nor U7892 (N_7892,N_6923,N_7175);
nor U7893 (N_7893,N_6769,N_7118);
or U7894 (N_7894,N_6724,N_6755);
nand U7895 (N_7895,N_7113,N_6458);
xnor U7896 (N_7896,N_6795,N_6685);
and U7897 (N_7897,N_7141,N_6557);
or U7898 (N_7898,N_6515,N_6720);
or U7899 (N_7899,N_6949,N_7184);
nand U7900 (N_7900,N_6721,N_6579);
xor U7901 (N_7901,N_6532,N_7006);
nand U7902 (N_7902,N_6967,N_6520);
xor U7903 (N_7903,N_6418,N_6800);
nand U7904 (N_7904,N_6773,N_7134);
nand U7905 (N_7905,N_7177,N_6601);
or U7906 (N_7906,N_6406,N_6832);
or U7907 (N_7907,N_6936,N_7143);
or U7908 (N_7908,N_7086,N_6764);
or U7909 (N_7909,N_6618,N_6899);
and U7910 (N_7910,N_7044,N_6841);
or U7911 (N_7911,N_6853,N_6525);
nor U7912 (N_7912,N_6677,N_6807);
nand U7913 (N_7913,N_6405,N_6987);
nor U7914 (N_7914,N_6657,N_6411);
or U7915 (N_7915,N_6486,N_7001);
nor U7916 (N_7916,N_6802,N_6925);
nor U7917 (N_7917,N_6606,N_6633);
and U7918 (N_7918,N_6928,N_6880);
nand U7919 (N_7919,N_6762,N_6804);
xnor U7920 (N_7920,N_6556,N_6734);
nor U7921 (N_7921,N_6526,N_6941);
and U7922 (N_7922,N_7131,N_7163);
and U7923 (N_7923,N_6455,N_7113);
nor U7924 (N_7924,N_7001,N_7190);
and U7925 (N_7925,N_6633,N_6677);
nor U7926 (N_7926,N_6698,N_6416);
nand U7927 (N_7927,N_7103,N_7029);
xnor U7928 (N_7928,N_6703,N_7087);
or U7929 (N_7929,N_6535,N_6437);
nor U7930 (N_7930,N_6476,N_6607);
xnor U7931 (N_7931,N_6788,N_7000);
and U7932 (N_7932,N_7144,N_6730);
nor U7933 (N_7933,N_6546,N_6587);
or U7934 (N_7934,N_6640,N_7059);
nor U7935 (N_7935,N_7165,N_6948);
and U7936 (N_7936,N_7054,N_6790);
and U7937 (N_7937,N_6600,N_6537);
nand U7938 (N_7938,N_6520,N_6635);
nor U7939 (N_7939,N_6604,N_6807);
nand U7940 (N_7940,N_7065,N_7157);
or U7941 (N_7941,N_6612,N_6507);
xnor U7942 (N_7942,N_6728,N_6464);
xnor U7943 (N_7943,N_6839,N_6505);
xor U7944 (N_7944,N_7071,N_6995);
or U7945 (N_7945,N_6646,N_6801);
nand U7946 (N_7946,N_6611,N_6643);
xnor U7947 (N_7947,N_6714,N_7094);
or U7948 (N_7948,N_6642,N_6622);
nor U7949 (N_7949,N_7031,N_6821);
xnor U7950 (N_7950,N_7002,N_6542);
nand U7951 (N_7951,N_6436,N_6991);
nand U7952 (N_7952,N_6998,N_6543);
nor U7953 (N_7953,N_6475,N_7110);
nand U7954 (N_7954,N_6568,N_6841);
xnor U7955 (N_7955,N_6487,N_7015);
nor U7956 (N_7956,N_6810,N_6553);
nand U7957 (N_7957,N_7195,N_6980);
and U7958 (N_7958,N_7062,N_6489);
or U7959 (N_7959,N_6441,N_7121);
nor U7960 (N_7960,N_6548,N_7199);
nand U7961 (N_7961,N_6790,N_6748);
and U7962 (N_7962,N_6725,N_7049);
and U7963 (N_7963,N_6461,N_7126);
and U7964 (N_7964,N_7103,N_6572);
nand U7965 (N_7965,N_6757,N_7171);
xor U7966 (N_7966,N_6912,N_7136);
xor U7967 (N_7967,N_6406,N_6823);
nand U7968 (N_7968,N_6860,N_7150);
xor U7969 (N_7969,N_6986,N_6987);
nand U7970 (N_7970,N_7046,N_6572);
or U7971 (N_7971,N_6768,N_6482);
or U7972 (N_7972,N_6602,N_6476);
xor U7973 (N_7973,N_7177,N_7034);
xor U7974 (N_7974,N_6712,N_6426);
or U7975 (N_7975,N_7091,N_6683);
nand U7976 (N_7976,N_6815,N_6767);
and U7977 (N_7977,N_6634,N_6870);
nand U7978 (N_7978,N_7187,N_7117);
xnor U7979 (N_7979,N_7114,N_6873);
or U7980 (N_7980,N_6622,N_6938);
and U7981 (N_7981,N_6951,N_7086);
or U7982 (N_7982,N_6790,N_6885);
and U7983 (N_7983,N_6619,N_7006);
nand U7984 (N_7984,N_7038,N_6461);
and U7985 (N_7985,N_6690,N_6417);
or U7986 (N_7986,N_6890,N_7086);
nand U7987 (N_7987,N_6433,N_7138);
xor U7988 (N_7988,N_7122,N_7190);
and U7989 (N_7989,N_6407,N_6897);
and U7990 (N_7990,N_6863,N_6629);
nor U7991 (N_7991,N_6846,N_7078);
nand U7992 (N_7992,N_6432,N_6641);
or U7993 (N_7993,N_6544,N_6573);
nor U7994 (N_7994,N_6834,N_6484);
and U7995 (N_7995,N_6824,N_6740);
or U7996 (N_7996,N_6546,N_6868);
xnor U7997 (N_7997,N_6809,N_6868);
nor U7998 (N_7998,N_6947,N_6764);
or U7999 (N_7999,N_6739,N_7199);
nor U8000 (N_8000,N_7734,N_7366);
xor U8001 (N_8001,N_7392,N_7990);
and U8002 (N_8002,N_7808,N_7283);
nor U8003 (N_8003,N_7668,N_7715);
nand U8004 (N_8004,N_7699,N_7867);
nand U8005 (N_8005,N_7304,N_7434);
nor U8006 (N_8006,N_7839,N_7653);
and U8007 (N_8007,N_7978,N_7625);
and U8008 (N_8008,N_7953,N_7816);
or U8009 (N_8009,N_7402,N_7705);
and U8010 (N_8010,N_7235,N_7834);
xor U8011 (N_8011,N_7977,N_7988);
and U8012 (N_8012,N_7963,N_7841);
xnor U8013 (N_8013,N_7894,N_7923);
or U8014 (N_8014,N_7400,N_7346);
xor U8015 (N_8015,N_7640,N_7900);
and U8016 (N_8016,N_7524,N_7437);
nand U8017 (N_8017,N_7499,N_7296);
nand U8018 (N_8018,N_7754,N_7258);
or U8019 (N_8019,N_7790,N_7908);
xor U8020 (N_8020,N_7377,N_7695);
and U8021 (N_8021,N_7770,N_7445);
nor U8022 (N_8022,N_7692,N_7512);
xnor U8023 (N_8023,N_7814,N_7472);
xor U8024 (N_8024,N_7347,N_7343);
or U8025 (N_8025,N_7441,N_7473);
nand U8026 (N_8026,N_7788,N_7540);
or U8027 (N_8027,N_7865,N_7233);
or U8028 (N_8028,N_7658,N_7855);
nor U8029 (N_8029,N_7305,N_7667);
nand U8030 (N_8030,N_7356,N_7644);
nor U8031 (N_8031,N_7419,N_7778);
or U8032 (N_8032,N_7310,N_7306);
nand U8033 (N_8033,N_7757,N_7338);
and U8034 (N_8034,N_7767,N_7902);
and U8035 (N_8035,N_7966,N_7874);
xor U8036 (N_8036,N_7301,N_7538);
nand U8037 (N_8037,N_7421,N_7341);
xor U8038 (N_8038,N_7753,N_7284);
and U8039 (N_8039,N_7394,N_7243);
nand U8040 (N_8040,N_7641,N_7286);
nand U8041 (N_8041,N_7871,N_7917);
nand U8042 (N_8042,N_7761,N_7643);
nand U8043 (N_8043,N_7315,N_7417);
nor U8044 (N_8044,N_7504,N_7592);
xnor U8045 (N_8045,N_7317,N_7401);
nor U8046 (N_8046,N_7440,N_7630);
or U8047 (N_8047,N_7520,N_7460);
or U8048 (N_8048,N_7257,N_7833);
nor U8049 (N_8049,N_7222,N_7427);
xnor U8050 (N_8050,N_7242,N_7911);
or U8051 (N_8051,N_7555,N_7797);
or U8052 (N_8052,N_7464,N_7262);
and U8053 (N_8053,N_7961,N_7799);
nand U8054 (N_8054,N_7649,N_7677);
nand U8055 (N_8055,N_7873,N_7951);
xor U8056 (N_8056,N_7380,N_7551);
nand U8057 (N_8057,N_7432,N_7830);
nand U8058 (N_8058,N_7636,N_7395);
xnor U8059 (N_8059,N_7360,N_7719);
and U8060 (N_8060,N_7603,N_7971);
nand U8061 (N_8061,N_7599,N_7929);
xnor U8062 (N_8062,N_7954,N_7948);
and U8063 (N_8063,N_7756,N_7452);
xnor U8064 (N_8064,N_7375,N_7435);
or U8065 (N_8065,N_7960,N_7528);
and U8066 (N_8066,N_7789,N_7736);
nor U8067 (N_8067,N_7541,N_7981);
xor U8068 (N_8068,N_7796,N_7527);
nor U8069 (N_8069,N_7918,N_7406);
nand U8070 (N_8070,N_7983,N_7864);
or U8071 (N_8071,N_7311,N_7626);
xnor U8072 (N_8072,N_7950,N_7623);
or U8073 (N_8073,N_7570,N_7422);
nand U8074 (N_8074,N_7241,N_7609);
or U8075 (N_8075,N_7484,N_7991);
nor U8076 (N_8076,N_7281,N_7606);
xor U8077 (N_8077,N_7675,N_7821);
or U8078 (N_8078,N_7348,N_7312);
nor U8079 (N_8079,N_7506,N_7491);
or U8080 (N_8080,N_7822,N_7568);
nand U8081 (N_8081,N_7280,N_7457);
nand U8082 (N_8082,N_7259,N_7666);
or U8083 (N_8083,N_7605,N_7308);
and U8084 (N_8084,N_7218,N_7938);
and U8085 (N_8085,N_7396,N_7854);
nand U8086 (N_8086,N_7439,N_7863);
nor U8087 (N_8087,N_7480,N_7278);
xor U8088 (N_8088,N_7836,N_7279);
nor U8089 (N_8089,N_7654,N_7333);
and U8090 (N_8090,N_7783,N_7591);
and U8091 (N_8091,N_7344,N_7706);
and U8092 (N_8092,N_7998,N_7800);
xnor U8093 (N_8093,N_7709,N_7361);
nand U8094 (N_8094,N_7391,N_7933);
and U8095 (N_8095,N_7536,N_7525);
xnor U8096 (N_8096,N_7203,N_7274);
xor U8097 (N_8097,N_7443,N_7271);
nand U8098 (N_8098,N_7967,N_7268);
and U8099 (N_8099,N_7420,N_7733);
or U8100 (N_8100,N_7828,N_7980);
nor U8101 (N_8101,N_7937,N_7487);
nor U8102 (N_8102,N_7263,N_7412);
nand U8103 (N_8103,N_7206,N_7632);
and U8104 (N_8104,N_7759,N_7393);
xnor U8105 (N_8105,N_7915,N_7261);
or U8106 (N_8106,N_7604,N_7972);
xor U8107 (N_8107,N_7357,N_7297);
and U8108 (N_8108,N_7342,N_7737);
nor U8109 (N_8109,N_7426,N_7547);
or U8110 (N_8110,N_7999,N_7248);
and U8111 (N_8111,N_7680,N_7982);
xor U8112 (N_8112,N_7866,N_7897);
nand U8113 (N_8113,N_7881,N_7328);
or U8114 (N_8114,N_7817,N_7334);
xnor U8115 (N_8115,N_7912,N_7215);
or U8116 (N_8116,N_7728,N_7648);
and U8117 (N_8117,N_7228,N_7246);
or U8118 (N_8118,N_7404,N_7812);
xnor U8119 (N_8119,N_7968,N_7493);
nand U8120 (N_8120,N_7852,N_7708);
or U8121 (N_8121,N_7878,N_7887);
or U8122 (N_8122,N_7721,N_7616);
xnor U8123 (N_8123,N_7735,N_7781);
xnor U8124 (N_8124,N_7384,N_7220);
or U8125 (N_8125,N_7505,N_7634);
and U8126 (N_8126,N_7752,N_7921);
or U8127 (N_8127,N_7236,N_7353);
or U8128 (N_8128,N_7478,N_7217);
or U8129 (N_8129,N_7823,N_7408);
xnor U8130 (N_8130,N_7230,N_7582);
nor U8131 (N_8131,N_7850,N_7762);
nand U8132 (N_8132,N_7859,N_7806);
nor U8133 (N_8133,N_7594,N_7679);
or U8134 (N_8134,N_7544,N_7463);
or U8135 (N_8135,N_7738,N_7523);
or U8136 (N_8136,N_7612,N_7827);
and U8137 (N_8137,N_7300,N_7503);
or U8138 (N_8138,N_7820,N_7664);
nor U8139 (N_8139,N_7613,N_7492);
nand U8140 (N_8140,N_7952,N_7891);
xnor U8141 (N_8141,N_7496,N_7819);
xnor U8142 (N_8142,N_7904,N_7932);
nor U8143 (N_8143,N_7226,N_7451);
nand U8144 (N_8144,N_7232,N_7683);
nor U8145 (N_8145,N_7860,N_7847);
and U8146 (N_8146,N_7554,N_7913);
or U8147 (N_8147,N_7454,N_7558);
nand U8148 (N_8148,N_7798,N_7602);
nor U8149 (N_8149,N_7947,N_7483);
and U8150 (N_8150,N_7793,N_7979);
nand U8151 (N_8151,N_7619,N_7382);
or U8152 (N_8152,N_7890,N_7646);
and U8153 (N_8153,N_7772,N_7862);
xor U8154 (N_8154,N_7655,N_7424);
or U8155 (N_8155,N_7571,N_7211);
xor U8156 (N_8156,N_7651,N_7893);
nor U8157 (N_8157,N_7269,N_7748);
xor U8158 (N_8158,N_7906,N_7689);
xor U8159 (N_8159,N_7247,N_7231);
xor U8160 (N_8160,N_7690,N_7760);
and U8161 (N_8161,N_7920,N_7946);
xnor U8162 (N_8162,N_7251,N_7326);
nand U8163 (N_8163,N_7224,N_7880);
xnor U8164 (N_8164,N_7813,N_7562);
or U8165 (N_8165,N_7374,N_7488);
or U8166 (N_8166,N_7892,N_7962);
and U8167 (N_8167,N_7320,N_7291);
nor U8168 (N_8168,N_7239,N_7702);
xnor U8169 (N_8169,N_7707,N_7794);
xnor U8170 (N_8170,N_7586,N_7475);
and U8171 (N_8171,N_7621,N_7701);
xnor U8172 (N_8172,N_7955,N_7332);
or U8173 (N_8173,N_7389,N_7691);
xnor U8174 (N_8174,N_7294,N_7786);
nor U8175 (N_8175,N_7513,N_7238);
and U8176 (N_8176,N_7515,N_7886);
nand U8177 (N_8177,N_7992,N_7957);
nor U8178 (N_8178,N_7227,N_7337);
nor U8179 (N_8179,N_7614,N_7383);
xor U8180 (N_8180,N_7245,N_7455);
nor U8181 (N_8181,N_7944,N_7372);
xor U8182 (N_8182,N_7745,N_7548);
and U8183 (N_8183,N_7959,N_7943);
xnor U8184 (N_8184,N_7498,N_7635);
and U8185 (N_8185,N_7670,N_7267);
or U8186 (N_8186,N_7674,N_7712);
nor U8187 (N_8187,N_7608,N_7497);
nor U8188 (N_8188,N_7747,N_7717);
xnor U8189 (N_8189,N_7316,N_7809);
nand U8190 (N_8190,N_7755,N_7359);
nand U8191 (N_8191,N_7939,N_7637);
xnor U8192 (N_8192,N_7610,N_7696);
and U8193 (N_8193,N_7832,N_7293);
nand U8194 (N_8194,N_7598,N_7381);
xor U8195 (N_8195,N_7656,N_7622);
nor U8196 (N_8196,N_7928,N_7995);
nand U8197 (N_8197,N_7266,N_7430);
nor U8198 (N_8198,N_7660,N_7723);
or U8199 (N_8199,N_7704,N_7367);
and U8200 (N_8200,N_7924,N_7510);
or U8201 (N_8201,N_7214,N_7456);
nand U8202 (N_8202,N_7295,N_7787);
or U8203 (N_8203,N_7405,N_7556);
nand U8204 (N_8204,N_7414,N_7397);
nor U8205 (N_8205,N_7249,N_7576);
and U8206 (N_8206,N_7225,N_7672);
nor U8207 (N_8207,N_7601,N_7889);
nand U8208 (N_8208,N_7386,N_7898);
and U8209 (N_8209,N_7627,N_7546);
and U8210 (N_8210,N_7750,N_7662);
nor U8211 (N_8211,N_7438,N_7428);
or U8212 (N_8212,N_7565,N_7254);
or U8213 (N_8213,N_7910,N_7740);
nor U8214 (N_8214,N_7535,N_7985);
or U8215 (N_8215,N_7204,N_7354);
and U8216 (N_8216,N_7250,N_7645);
or U8217 (N_8217,N_7407,N_7801);
nand U8218 (N_8218,N_7774,N_7669);
nor U8219 (N_8219,N_7916,N_7638);
nand U8220 (N_8220,N_7824,N_7355);
or U8221 (N_8221,N_7849,N_7673);
nand U8222 (N_8222,N_7792,N_7327);
and U8223 (N_8223,N_7577,N_7415);
or U8224 (N_8224,N_7872,N_7588);
nand U8225 (N_8225,N_7829,N_7469);
and U8226 (N_8226,N_7468,N_7618);
nor U8227 (N_8227,N_7791,N_7726);
xnor U8228 (N_8228,N_7256,N_7216);
nand U8229 (N_8229,N_7663,N_7746);
xor U8230 (N_8230,N_7322,N_7964);
xor U8231 (N_8231,N_7986,N_7563);
nand U8232 (N_8232,N_7732,N_7495);
nand U8233 (N_8233,N_7202,N_7209);
nor U8234 (N_8234,N_7803,N_7779);
xor U8235 (N_8235,N_7201,N_7615);
or U8236 (N_8236,N_7516,N_7869);
xnor U8237 (N_8237,N_7378,N_7825);
nor U8238 (N_8238,N_7771,N_7578);
or U8239 (N_8239,N_7518,N_7743);
xnor U8240 (N_8240,N_7277,N_7620);
and U8241 (N_8241,N_7240,N_7633);
or U8242 (N_8242,N_7365,N_7494);
nand U8243 (N_8243,N_7210,N_7773);
and U8244 (N_8244,N_7909,N_7661);
xnor U8245 (N_8245,N_7449,N_7471);
and U8246 (N_8246,N_7583,N_7965);
xnor U8247 (N_8247,N_7530,N_7290);
and U8248 (N_8248,N_7330,N_7739);
xnor U8249 (N_8249,N_7436,N_7351);
and U8250 (N_8250,N_7936,N_7877);
xnor U8251 (N_8251,N_7587,N_7511);
nor U8252 (N_8252,N_7935,N_7521);
or U8253 (N_8253,N_7289,N_7370);
or U8254 (N_8254,N_7818,N_7581);
and U8255 (N_8255,N_7403,N_7973);
xor U8256 (N_8256,N_7318,N_7987);
nor U8257 (N_8257,N_7907,N_7223);
nand U8258 (N_8258,N_7329,N_7508);
and U8259 (N_8259,N_7758,N_7940);
or U8260 (N_8260,N_7490,N_7539);
nand U8261 (N_8261,N_7369,N_7273);
nor U8262 (N_8262,N_7462,N_7727);
nor U8263 (N_8263,N_7303,N_7479);
nor U8264 (N_8264,N_7458,N_7398);
nand U8265 (N_8265,N_7597,N_7914);
nand U8266 (N_8266,N_7519,N_7693);
nand U8267 (N_8267,N_7785,N_7567);
xnor U8268 (N_8268,N_7489,N_7288);
or U8269 (N_8269,N_7688,N_7345);
and U8270 (N_8270,N_7835,N_7742);
xnor U8271 (N_8271,N_7461,N_7362);
nand U8272 (N_8272,N_7718,N_7879);
and U8273 (N_8273,N_7275,N_7975);
and U8274 (N_8274,N_7264,N_7888);
nand U8275 (N_8275,N_7244,N_7444);
or U8276 (N_8276,N_7569,N_7659);
nor U8277 (N_8277,N_7298,N_7840);
nor U8278 (N_8278,N_7467,N_7481);
nand U8279 (N_8279,N_7861,N_7331);
or U8280 (N_8280,N_7376,N_7844);
xor U8281 (N_8281,N_7219,N_7585);
nand U8282 (N_8282,N_7945,N_7260);
nand U8283 (N_8283,N_7368,N_7363);
nand U8284 (N_8284,N_7642,N_7207);
or U8285 (N_8285,N_7205,N_7676);
nor U8286 (N_8286,N_7416,N_7399);
nor U8287 (N_8287,N_7212,N_7650);
nor U8288 (N_8288,N_7722,N_7501);
nor U8289 (N_8289,N_7710,N_7390);
nand U8290 (N_8290,N_7514,N_7270);
nand U8291 (N_8291,N_7697,N_7553);
nand U8292 (N_8292,N_7926,N_7552);
nand U8293 (N_8293,N_7564,N_7678);
and U8294 (N_8294,N_7784,N_7804);
or U8295 (N_8295,N_7931,N_7253);
or U8296 (N_8296,N_7611,N_7507);
or U8297 (N_8297,N_7352,N_7993);
nor U8298 (N_8298,N_7956,N_7371);
and U8299 (N_8299,N_7542,N_7319);
xor U8300 (N_8300,N_7580,N_7875);
or U8301 (N_8301,N_7573,N_7805);
nand U8302 (N_8302,N_7927,N_7379);
or U8303 (N_8303,N_7321,N_7766);
nor U8304 (N_8304,N_7550,N_7868);
nand U8305 (N_8305,N_7922,N_7325);
xor U8306 (N_8306,N_7252,N_7777);
or U8307 (N_8307,N_7453,N_7532);
nor U8308 (N_8308,N_7851,N_7600);
nor U8309 (N_8309,N_7561,N_7431);
and U8310 (N_8310,N_7533,N_7486);
or U8311 (N_8311,N_7845,N_7930);
or U8312 (N_8312,N_7896,N_7373);
or U8313 (N_8313,N_7470,N_7589);
nand U8314 (N_8314,N_7448,N_7831);
xor U8315 (N_8315,N_7639,N_7885);
nand U8316 (N_8316,N_7815,N_7350);
xor U8317 (N_8317,N_7684,N_7903);
nand U8318 (N_8318,N_7846,N_7485);
nor U8319 (N_8319,N_7826,N_7703);
and U8320 (N_8320,N_7276,N_7749);
or U8321 (N_8321,N_7631,N_7423);
xor U8322 (N_8322,N_7730,N_7731);
xor U8323 (N_8323,N_7358,N_7299);
xor U8324 (N_8324,N_7687,N_7543);
xor U8325 (N_8325,N_7477,N_7526);
and U8326 (N_8326,N_7744,N_7853);
xnor U8327 (N_8327,N_7895,N_7324);
and U8328 (N_8328,N_7335,N_7593);
nor U8329 (N_8329,N_7714,N_7617);
xor U8330 (N_8330,N_7200,N_7810);
xnor U8331 (N_8331,N_7969,N_7919);
nand U8332 (N_8332,N_7883,N_7694);
and U8333 (N_8333,N_7837,N_7681);
xor U8334 (N_8334,N_7566,N_7517);
nor U8335 (N_8335,N_7811,N_7459);
and U8336 (N_8336,N_7628,N_7925);
nand U8337 (N_8337,N_7349,N_7265);
nor U8338 (N_8338,N_7465,N_7557);
and U8339 (N_8339,N_7843,N_7870);
nor U8340 (N_8340,N_7221,N_7997);
and U8341 (N_8341,N_7857,N_7385);
and U8342 (N_8342,N_7234,N_7309);
and U8343 (N_8343,N_7858,N_7958);
and U8344 (N_8344,N_7652,N_7237);
xnor U8345 (N_8345,N_7775,N_7575);
and U8346 (N_8346,N_7522,N_7531);
and U8347 (N_8347,N_7842,N_7229);
nor U8348 (N_8348,N_7549,N_7629);
or U8349 (N_8349,N_7725,N_7970);
or U8350 (N_8350,N_7899,N_7765);
xor U8351 (N_8351,N_7624,N_7884);
or U8352 (N_8352,N_7905,N_7534);
xnor U8353 (N_8353,N_7769,N_7856);
nand U8354 (N_8354,N_7560,N_7647);
nor U8355 (N_8355,N_7387,N_7942);
nand U8356 (N_8356,N_7314,N_7579);
xnor U8357 (N_8357,N_7720,N_7807);
xnor U8358 (N_8358,N_7429,N_7848);
or U8359 (N_8359,N_7764,N_7433);
nand U8360 (N_8360,N_7751,N_7388);
xnor U8361 (N_8361,N_7994,N_7574);
xor U8362 (N_8362,N_7776,N_7559);
nor U8363 (N_8363,N_7364,N_7292);
xnor U8364 (N_8364,N_7302,N_7442);
nor U8365 (N_8365,N_7411,N_7313);
nand U8366 (N_8366,N_7716,N_7795);
or U8367 (N_8367,N_7802,N_7782);
xnor U8368 (N_8368,N_7336,N_7425);
or U8369 (N_8369,N_7949,N_7272);
and U8370 (N_8370,N_7671,N_7711);
nand U8371 (N_8371,N_7323,N_7208);
xor U8372 (N_8372,N_7450,N_7713);
nor U8373 (N_8373,N_7665,N_7529);
or U8374 (N_8374,N_7876,N_7339);
nand U8375 (N_8375,N_7595,N_7882);
or U8376 (N_8376,N_7698,N_7989);
or U8377 (N_8377,N_7213,N_7941);
and U8378 (N_8378,N_7976,N_7741);
nand U8379 (N_8379,N_7340,N_7418);
nor U8380 (N_8380,N_7768,N_7545);
or U8381 (N_8381,N_7763,N_7413);
and U8382 (N_8382,N_7285,N_7596);
nand U8383 (N_8383,N_7287,N_7502);
nor U8384 (N_8384,N_7474,N_7476);
xor U8385 (N_8385,N_7686,N_7409);
nor U8386 (N_8386,N_7590,N_7282);
nor U8387 (N_8387,N_7307,N_7974);
xor U8388 (N_8388,N_7509,N_7700);
or U8389 (N_8389,N_7901,N_7500);
and U8390 (N_8390,N_7572,N_7447);
or U8391 (N_8391,N_7446,N_7838);
xor U8392 (N_8392,N_7984,N_7607);
or U8393 (N_8393,N_7729,N_7682);
nor U8394 (N_8394,N_7482,N_7780);
or U8395 (N_8395,N_7996,N_7584);
and U8396 (N_8396,N_7724,N_7410);
nand U8397 (N_8397,N_7934,N_7657);
or U8398 (N_8398,N_7685,N_7255);
or U8399 (N_8399,N_7537,N_7466);
and U8400 (N_8400,N_7762,N_7947);
and U8401 (N_8401,N_7407,N_7469);
xor U8402 (N_8402,N_7941,N_7272);
nor U8403 (N_8403,N_7497,N_7282);
xor U8404 (N_8404,N_7356,N_7296);
xor U8405 (N_8405,N_7381,N_7641);
or U8406 (N_8406,N_7923,N_7985);
or U8407 (N_8407,N_7734,N_7284);
or U8408 (N_8408,N_7454,N_7957);
nor U8409 (N_8409,N_7979,N_7422);
and U8410 (N_8410,N_7306,N_7215);
or U8411 (N_8411,N_7440,N_7679);
xnor U8412 (N_8412,N_7889,N_7575);
and U8413 (N_8413,N_7561,N_7995);
nand U8414 (N_8414,N_7843,N_7284);
nor U8415 (N_8415,N_7658,N_7669);
nor U8416 (N_8416,N_7924,N_7821);
and U8417 (N_8417,N_7947,N_7914);
nand U8418 (N_8418,N_7362,N_7962);
xor U8419 (N_8419,N_7569,N_7263);
and U8420 (N_8420,N_7416,N_7508);
nor U8421 (N_8421,N_7861,N_7580);
and U8422 (N_8422,N_7774,N_7999);
or U8423 (N_8423,N_7359,N_7783);
xor U8424 (N_8424,N_7301,N_7559);
and U8425 (N_8425,N_7721,N_7969);
nor U8426 (N_8426,N_7568,N_7972);
xnor U8427 (N_8427,N_7632,N_7532);
or U8428 (N_8428,N_7563,N_7387);
nor U8429 (N_8429,N_7674,N_7660);
or U8430 (N_8430,N_7316,N_7903);
nor U8431 (N_8431,N_7799,N_7795);
nand U8432 (N_8432,N_7923,N_7346);
or U8433 (N_8433,N_7727,N_7686);
or U8434 (N_8434,N_7986,N_7700);
xnor U8435 (N_8435,N_7560,N_7976);
nor U8436 (N_8436,N_7651,N_7544);
nor U8437 (N_8437,N_7488,N_7257);
nor U8438 (N_8438,N_7519,N_7711);
or U8439 (N_8439,N_7329,N_7778);
or U8440 (N_8440,N_7599,N_7354);
and U8441 (N_8441,N_7938,N_7912);
xnor U8442 (N_8442,N_7380,N_7753);
or U8443 (N_8443,N_7530,N_7963);
and U8444 (N_8444,N_7996,N_7404);
and U8445 (N_8445,N_7317,N_7588);
and U8446 (N_8446,N_7864,N_7552);
and U8447 (N_8447,N_7979,N_7503);
nand U8448 (N_8448,N_7366,N_7867);
nor U8449 (N_8449,N_7361,N_7498);
or U8450 (N_8450,N_7472,N_7641);
or U8451 (N_8451,N_7528,N_7999);
nand U8452 (N_8452,N_7229,N_7273);
and U8453 (N_8453,N_7254,N_7850);
nor U8454 (N_8454,N_7722,N_7675);
xor U8455 (N_8455,N_7255,N_7718);
nor U8456 (N_8456,N_7544,N_7693);
nor U8457 (N_8457,N_7871,N_7718);
or U8458 (N_8458,N_7705,N_7458);
nand U8459 (N_8459,N_7598,N_7328);
nand U8460 (N_8460,N_7383,N_7686);
and U8461 (N_8461,N_7360,N_7840);
nor U8462 (N_8462,N_7895,N_7265);
xor U8463 (N_8463,N_7386,N_7401);
and U8464 (N_8464,N_7755,N_7355);
nor U8465 (N_8465,N_7966,N_7601);
and U8466 (N_8466,N_7925,N_7411);
xor U8467 (N_8467,N_7509,N_7237);
and U8468 (N_8468,N_7964,N_7705);
or U8469 (N_8469,N_7710,N_7204);
nand U8470 (N_8470,N_7894,N_7333);
nor U8471 (N_8471,N_7803,N_7584);
nand U8472 (N_8472,N_7494,N_7304);
nor U8473 (N_8473,N_7945,N_7517);
nand U8474 (N_8474,N_7753,N_7646);
nor U8475 (N_8475,N_7494,N_7712);
and U8476 (N_8476,N_7681,N_7534);
nand U8477 (N_8477,N_7337,N_7852);
xnor U8478 (N_8478,N_7311,N_7918);
nor U8479 (N_8479,N_7652,N_7472);
and U8480 (N_8480,N_7729,N_7782);
or U8481 (N_8481,N_7333,N_7411);
or U8482 (N_8482,N_7736,N_7816);
and U8483 (N_8483,N_7522,N_7258);
xor U8484 (N_8484,N_7965,N_7285);
and U8485 (N_8485,N_7734,N_7969);
and U8486 (N_8486,N_7476,N_7829);
xnor U8487 (N_8487,N_7528,N_7273);
xor U8488 (N_8488,N_7654,N_7667);
and U8489 (N_8489,N_7291,N_7549);
nand U8490 (N_8490,N_7716,N_7227);
xnor U8491 (N_8491,N_7448,N_7384);
nor U8492 (N_8492,N_7818,N_7560);
and U8493 (N_8493,N_7750,N_7705);
or U8494 (N_8494,N_7996,N_7646);
or U8495 (N_8495,N_7982,N_7791);
nor U8496 (N_8496,N_7933,N_7860);
nand U8497 (N_8497,N_7582,N_7604);
and U8498 (N_8498,N_7913,N_7579);
nor U8499 (N_8499,N_7955,N_7918);
xnor U8500 (N_8500,N_7922,N_7951);
nor U8501 (N_8501,N_7462,N_7525);
xor U8502 (N_8502,N_7401,N_7374);
nand U8503 (N_8503,N_7378,N_7345);
and U8504 (N_8504,N_7470,N_7549);
nand U8505 (N_8505,N_7235,N_7511);
or U8506 (N_8506,N_7597,N_7550);
and U8507 (N_8507,N_7785,N_7740);
nand U8508 (N_8508,N_7851,N_7860);
or U8509 (N_8509,N_7772,N_7259);
or U8510 (N_8510,N_7229,N_7775);
nand U8511 (N_8511,N_7473,N_7839);
and U8512 (N_8512,N_7216,N_7491);
xnor U8513 (N_8513,N_7658,N_7245);
xnor U8514 (N_8514,N_7674,N_7966);
nor U8515 (N_8515,N_7393,N_7491);
nor U8516 (N_8516,N_7397,N_7437);
nor U8517 (N_8517,N_7867,N_7631);
xor U8518 (N_8518,N_7765,N_7692);
or U8519 (N_8519,N_7745,N_7860);
and U8520 (N_8520,N_7787,N_7373);
and U8521 (N_8521,N_7267,N_7532);
or U8522 (N_8522,N_7317,N_7394);
and U8523 (N_8523,N_7816,N_7415);
or U8524 (N_8524,N_7930,N_7340);
and U8525 (N_8525,N_7630,N_7791);
nand U8526 (N_8526,N_7586,N_7661);
nor U8527 (N_8527,N_7988,N_7529);
or U8528 (N_8528,N_7768,N_7628);
and U8529 (N_8529,N_7233,N_7361);
xnor U8530 (N_8530,N_7907,N_7702);
or U8531 (N_8531,N_7741,N_7386);
nand U8532 (N_8532,N_7323,N_7355);
xnor U8533 (N_8533,N_7683,N_7542);
xor U8534 (N_8534,N_7761,N_7833);
nand U8535 (N_8535,N_7557,N_7259);
and U8536 (N_8536,N_7955,N_7200);
xnor U8537 (N_8537,N_7479,N_7801);
nand U8538 (N_8538,N_7870,N_7448);
xor U8539 (N_8539,N_7292,N_7506);
nor U8540 (N_8540,N_7327,N_7682);
and U8541 (N_8541,N_7367,N_7569);
nand U8542 (N_8542,N_7572,N_7873);
or U8543 (N_8543,N_7722,N_7984);
nor U8544 (N_8544,N_7280,N_7963);
xor U8545 (N_8545,N_7432,N_7904);
nand U8546 (N_8546,N_7934,N_7841);
nand U8547 (N_8547,N_7904,N_7347);
or U8548 (N_8548,N_7370,N_7839);
xnor U8549 (N_8549,N_7490,N_7853);
nand U8550 (N_8550,N_7274,N_7709);
nor U8551 (N_8551,N_7539,N_7419);
nand U8552 (N_8552,N_7503,N_7974);
and U8553 (N_8553,N_7689,N_7992);
nor U8554 (N_8554,N_7923,N_7445);
and U8555 (N_8555,N_7818,N_7450);
nor U8556 (N_8556,N_7402,N_7740);
or U8557 (N_8557,N_7660,N_7938);
and U8558 (N_8558,N_7231,N_7523);
and U8559 (N_8559,N_7474,N_7879);
nand U8560 (N_8560,N_7816,N_7212);
nand U8561 (N_8561,N_7866,N_7936);
or U8562 (N_8562,N_7897,N_7208);
and U8563 (N_8563,N_7835,N_7962);
nor U8564 (N_8564,N_7670,N_7425);
nor U8565 (N_8565,N_7293,N_7236);
and U8566 (N_8566,N_7697,N_7812);
nand U8567 (N_8567,N_7599,N_7230);
or U8568 (N_8568,N_7912,N_7654);
xnor U8569 (N_8569,N_7276,N_7543);
and U8570 (N_8570,N_7859,N_7406);
nand U8571 (N_8571,N_7793,N_7635);
xnor U8572 (N_8572,N_7237,N_7508);
nand U8573 (N_8573,N_7955,N_7251);
nor U8574 (N_8574,N_7725,N_7948);
nand U8575 (N_8575,N_7778,N_7650);
xor U8576 (N_8576,N_7403,N_7588);
and U8577 (N_8577,N_7921,N_7604);
nor U8578 (N_8578,N_7225,N_7821);
or U8579 (N_8579,N_7416,N_7582);
xnor U8580 (N_8580,N_7779,N_7334);
or U8581 (N_8581,N_7524,N_7473);
or U8582 (N_8582,N_7283,N_7964);
nor U8583 (N_8583,N_7347,N_7262);
or U8584 (N_8584,N_7205,N_7886);
xnor U8585 (N_8585,N_7664,N_7379);
or U8586 (N_8586,N_7470,N_7397);
and U8587 (N_8587,N_7400,N_7233);
xnor U8588 (N_8588,N_7248,N_7807);
nand U8589 (N_8589,N_7710,N_7860);
or U8590 (N_8590,N_7504,N_7875);
xnor U8591 (N_8591,N_7206,N_7333);
and U8592 (N_8592,N_7723,N_7866);
and U8593 (N_8593,N_7232,N_7406);
or U8594 (N_8594,N_7706,N_7909);
nand U8595 (N_8595,N_7517,N_7948);
nor U8596 (N_8596,N_7770,N_7987);
nor U8597 (N_8597,N_7341,N_7460);
nor U8598 (N_8598,N_7875,N_7959);
nand U8599 (N_8599,N_7244,N_7701);
nor U8600 (N_8600,N_7443,N_7749);
and U8601 (N_8601,N_7638,N_7665);
or U8602 (N_8602,N_7268,N_7801);
or U8603 (N_8603,N_7286,N_7332);
nand U8604 (N_8604,N_7287,N_7689);
or U8605 (N_8605,N_7511,N_7353);
and U8606 (N_8606,N_7534,N_7887);
xnor U8607 (N_8607,N_7976,N_7289);
nand U8608 (N_8608,N_7456,N_7927);
or U8609 (N_8609,N_7861,N_7863);
xor U8610 (N_8610,N_7755,N_7982);
and U8611 (N_8611,N_7767,N_7730);
or U8612 (N_8612,N_7711,N_7672);
xnor U8613 (N_8613,N_7625,N_7844);
nor U8614 (N_8614,N_7283,N_7797);
or U8615 (N_8615,N_7363,N_7220);
nor U8616 (N_8616,N_7803,N_7660);
or U8617 (N_8617,N_7409,N_7358);
or U8618 (N_8618,N_7423,N_7976);
and U8619 (N_8619,N_7486,N_7407);
nand U8620 (N_8620,N_7408,N_7723);
nor U8621 (N_8621,N_7839,N_7577);
xor U8622 (N_8622,N_7382,N_7715);
or U8623 (N_8623,N_7255,N_7941);
nor U8624 (N_8624,N_7445,N_7962);
nand U8625 (N_8625,N_7346,N_7720);
and U8626 (N_8626,N_7748,N_7268);
xnor U8627 (N_8627,N_7670,N_7269);
and U8628 (N_8628,N_7726,N_7557);
and U8629 (N_8629,N_7427,N_7209);
nand U8630 (N_8630,N_7815,N_7297);
xor U8631 (N_8631,N_7380,N_7377);
and U8632 (N_8632,N_7973,N_7337);
xor U8633 (N_8633,N_7672,N_7215);
or U8634 (N_8634,N_7513,N_7977);
and U8635 (N_8635,N_7800,N_7380);
nor U8636 (N_8636,N_7841,N_7311);
nand U8637 (N_8637,N_7958,N_7510);
or U8638 (N_8638,N_7440,N_7978);
or U8639 (N_8639,N_7608,N_7623);
nand U8640 (N_8640,N_7431,N_7361);
nand U8641 (N_8641,N_7396,N_7489);
or U8642 (N_8642,N_7316,N_7547);
xnor U8643 (N_8643,N_7889,N_7325);
nor U8644 (N_8644,N_7789,N_7365);
nor U8645 (N_8645,N_7439,N_7614);
nand U8646 (N_8646,N_7744,N_7500);
nand U8647 (N_8647,N_7854,N_7323);
or U8648 (N_8648,N_7635,N_7929);
nor U8649 (N_8649,N_7510,N_7436);
xor U8650 (N_8650,N_7349,N_7443);
nor U8651 (N_8651,N_7917,N_7529);
nor U8652 (N_8652,N_7373,N_7224);
nor U8653 (N_8653,N_7389,N_7512);
or U8654 (N_8654,N_7703,N_7730);
nand U8655 (N_8655,N_7441,N_7488);
nor U8656 (N_8656,N_7641,N_7916);
and U8657 (N_8657,N_7673,N_7649);
xor U8658 (N_8658,N_7841,N_7799);
or U8659 (N_8659,N_7618,N_7421);
nor U8660 (N_8660,N_7948,N_7593);
xnor U8661 (N_8661,N_7650,N_7528);
xor U8662 (N_8662,N_7986,N_7917);
nand U8663 (N_8663,N_7445,N_7540);
nand U8664 (N_8664,N_7513,N_7930);
or U8665 (N_8665,N_7455,N_7374);
and U8666 (N_8666,N_7412,N_7358);
nor U8667 (N_8667,N_7424,N_7469);
nor U8668 (N_8668,N_7425,N_7834);
xor U8669 (N_8669,N_7315,N_7536);
xor U8670 (N_8670,N_7275,N_7467);
and U8671 (N_8671,N_7260,N_7858);
and U8672 (N_8672,N_7459,N_7431);
nor U8673 (N_8673,N_7554,N_7873);
and U8674 (N_8674,N_7246,N_7726);
or U8675 (N_8675,N_7846,N_7362);
xnor U8676 (N_8676,N_7755,N_7932);
xnor U8677 (N_8677,N_7819,N_7206);
nand U8678 (N_8678,N_7711,N_7465);
nor U8679 (N_8679,N_7689,N_7621);
xnor U8680 (N_8680,N_7368,N_7312);
xor U8681 (N_8681,N_7403,N_7714);
nor U8682 (N_8682,N_7921,N_7712);
and U8683 (N_8683,N_7514,N_7437);
or U8684 (N_8684,N_7247,N_7496);
and U8685 (N_8685,N_7697,N_7369);
nand U8686 (N_8686,N_7659,N_7930);
nand U8687 (N_8687,N_7472,N_7232);
nand U8688 (N_8688,N_7370,N_7909);
nor U8689 (N_8689,N_7806,N_7926);
xor U8690 (N_8690,N_7570,N_7253);
xnor U8691 (N_8691,N_7210,N_7220);
or U8692 (N_8692,N_7556,N_7800);
and U8693 (N_8693,N_7915,N_7384);
nor U8694 (N_8694,N_7903,N_7907);
nand U8695 (N_8695,N_7500,N_7342);
xor U8696 (N_8696,N_7596,N_7278);
xor U8697 (N_8697,N_7935,N_7220);
nor U8698 (N_8698,N_7806,N_7234);
or U8699 (N_8699,N_7394,N_7486);
and U8700 (N_8700,N_7215,N_7783);
nand U8701 (N_8701,N_7875,N_7920);
nand U8702 (N_8702,N_7728,N_7639);
nand U8703 (N_8703,N_7858,N_7495);
or U8704 (N_8704,N_7442,N_7848);
and U8705 (N_8705,N_7312,N_7715);
xor U8706 (N_8706,N_7748,N_7530);
nor U8707 (N_8707,N_7404,N_7516);
or U8708 (N_8708,N_7351,N_7768);
nor U8709 (N_8709,N_7253,N_7482);
and U8710 (N_8710,N_7232,N_7342);
and U8711 (N_8711,N_7859,N_7385);
xor U8712 (N_8712,N_7785,N_7696);
xor U8713 (N_8713,N_7830,N_7237);
xnor U8714 (N_8714,N_7771,N_7734);
or U8715 (N_8715,N_7739,N_7979);
nor U8716 (N_8716,N_7639,N_7674);
and U8717 (N_8717,N_7751,N_7930);
or U8718 (N_8718,N_7384,N_7614);
nor U8719 (N_8719,N_7952,N_7900);
and U8720 (N_8720,N_7748,N_7891);
nor U8721 (N_8721,N_7448,N_7985);
nand U8722 (N_8722,N_7786,N_7617);
or U8723 (N_8723,N_7223,N_7871);
xnor U8724 (N_8724,N_7416,N_7242);
xnor U8725 (N_8725,N_7223,N_7873);
xnor U8726 (N_8726,N_7869,N_7497);
nand U8727 (N_8727,N_7385,N_7866);
nand U8728 (N_8728,N_7812,N_7480);
nor U8729 (N_8729,N_7287,N_7249);
nor U8730 (N_8730,N_7712,N_7860);
xor U8731 (N_8731,N_7854,N_7940);
nor U8732 (N_8732,N_7575,N_7309);
nor U8733 (N_8733,N_7441,N_7912);
and U8734 (N_8734,N_7889,N_7879);
or U8735 (N_8735,N_7735,N_7464);
nor U8736 (N_8736,N_7530,N_7670);
or U8737 (N_8737,N_7230,N_7220);
or U8738 (N_8738,N_7341,N_7470);
nor U8739 (N_8739,N_7522,N_7490);
xnor U8740 (N_8740,N_7980,N_7734);
xnor U8741 (N_8741,N_7931,N_7233);
or U8742 (N_8742,N_7739,N_7501);
or U8743 (N_8743,N_7637,N_7215);
and U8744 (N_8744,N_7471,N_7654);
and U8745 (N_8745,N_7739,N_7900);
nand U8746 (N_8746,N_7496,N_7861);
and U8747 (N_8747,N_7876,N_7471);
or U8748 (N_8748,N_7902,N_7892);
or U8749 (N_8749,N_7832,N_7358);
xnor U8750 (N_8750,N_7949,N_7602);
or U8751 (N_8751,N_7243,N_7746);
nor U8752 (N_8752,N_7388,N_7213);
nand U8753 (N_8753,N_7733,N_7829);
nand U8754 (N_8754,N_7814,N_7907);
or U8755 (N_8755,N_7799,N_7894);
and U8756 (N_8756,N_7791,N_7764);
and U8757 (N_8757,N_7864,N_7459);
and U8758 (N_8758,N_7716,N_7329);
or U8759 (N_8759,N_7820,N_7712);
and U8760 (N_8760,N_7601,N_7278);
nor U8761 (N_8761,N_7780,N_7720);
nand U8762 (N_8762,N_7720,N_7799);
nand U8763 (N_8763,N_7603,N_7810);
xnor U8764 (N_8764,N_7360,N_7758);
xor U8765 (N_8765,N_7356,N_7387);
nand U8766 (N_8766,N_7271,N_7779);
xnor U8767 (N_8767,N_7866,N_7988);
xor U8768 (N_8768,N_7294,N_7209);
nand U8769 (N_8769,N_7389,N_7510);
or U8770 (N_8770,N_7229,N_7795);
nand U8771 (N_8771,N_7668,N_7956);
nor U8772 (N_8772,N_7647,N_7428);
xor U8773 (N_8773,N_7259,N_7526);
xnor U8774 (N_8774,N_7264,N_7209);
or U8775 (N_8775,N_7631,N_7730);
nand U8776 (N_8776,N_7830,N_7911);
or U8777 (N_8777,N_7219,N_7218);
nor U8778 (N_8778,N_7624,N_7941);
nand U8779 (N_8779,N_7780,N_7893);
or U8780 (N_8780,N_7763,N_7254);
or U8781 (N_8781,N_7945,N_7820);
or U8782 (N_8782,N_7578,N_7427);
and U8783 (N_8783,N_7585,N_7368);
nor U8784 (N_8784,N_7239,N_7976);
nand U8785 (N_8785,N_7369,N_7536);
nand U8786 (N_8786,N_7478,N_7975);
xnor U8787 (N_8787,N_7493,N_7259);
nand U8788 (N_8788,N_7968,N_7649);
and U8789 (N_8789,N_7465,N_7879);
xor U8790 (N_8790,N_7474,N_7817);
or U8791 (N_8791,N_7695,N_7256);
and U8792 (N_8792,N_7324,N_7440);
xnor U8793 (N_8793,N_7718,N_7914);
or U8794 (N_8794,N_7787,N_7298);
xnor U8795 (N_8795,N_7729,N_7740);
xor U8796 (N_8796,N_7233,N_7822);
or U8797 (N_8797,N_7891,N_7348);
nor U8798 (N_8798,N_7212,N_7526);
nand U8799 (N_8799,N_7670,N_7706);
or U8800 (N_8800,N_8182,N_8699);
nand U8801 (N_8801,N_8291,N_8202);
and U8802 (N_8802,N_8424,N_8485);
or U8803 (N_8803,N_8562,N_8788);
nand U8804 (N_8804,N_8635,N_8393);
xnor U8805 (N_8805,N_8010,N_8784);
or U8806 (N_8806,N_8041,N_8461);
nor U8807 (N_8807,N_8483,N_8370);
nor U8808 (N_8808,N_8326,N_8675);
and U8809 (N_8809,N_8630,N_8772);
or U8810 (N_8810,N_8312,N_8789);
or U8811 (N_8811,N_8498,N_8445);
xnor U8812 (N_8812,N_8356,N_8217);
and U8813 (N_8813,N_8048,N_8354);
or U8814 (N_8814,N_8503,N_8529);
and U8815 (N_8815,N_8062,N_8589);
and U8816 (N_8816,N_8741,N_8147);
and U8817 (N_8817,N_8344,N_8053);
and U8818 (N_8818,N_8223,N_8543);
nor U8819 (N_8819,N_8558,N_8614);
and U8820 (N_8820,N_8272,N_8081);
or U8821 (N_8821,N_8690,N_8317);
xor U8822 (N_8822,N_8594,N_8135);
nor U8823 (N_8823,N_8071,N_8436);
or U8824 (N_8824,N_8311,N_8346);
and U8825 (N_8825,N_8547,N_8186);
nor U8826 (N_8826,N_8411,N_8045);
nand U8827 (N_8827,N_8094,N_8238);
nor U8828 (N_8828,N_8753,N_8103);
and U8829 (N_8829,N_8585,N_8571);
nand U8830 (N_8830,N_8545,N_8012);
nand U8831 (N_8831,N_8099,N_8752);
nor U8832 (N_8832,N_8262,N_8438);
or U8833 (N_8833,N_8277,N_8179);
nand U8834 (N_8834,N_8781,N_8671);
nor U8835 (N_8835,N_8225,N_8009);
nand U8836 (N_8836,N_8063,N_8456);
and U8837 (N_8837,N_8639,N_8085);
or U8838 (N_8838,N_8260,N_8764);
or U8839 (N_8839,N_8112,N_8361);
nand U8840 (N_8840,N_8601,N_8122);
and U8841 (N_8841,N_8603,N_8318);
xor U8842 (N_8842,N_8373,N_8597);
nor U8843 (N_8843,N_8372,N_8013);
xnor U8844 (N_8844,N_8153,N_8345);
nand U8845 (N_8845,N_8723,N_8609);
and U8846 (N_8846,N_8522,N_8139);
nand U8847 (N_8847,N_8487,N_8284);
or U8848 (N_8848,N_8049,N_8582);
xnor U8849 (N_8849,N_8204,N_8641);
and U8850 (N_8850,N_8495,N_8005);
or U8851 (N_8851,N_8568,N_8499);
nand U8852 (N_8852,N_8758,N_8777);
or U8853 (N_8853,N_8766,N_8165);
xor U8854 (N_8854,N_8124,N_8590);
and U8855 (N_8855,N_8246,N_8618);
nand U8856 (N_8856,N_8377,N_8211);
or U8857 (N_8857,N_8338,N_8565);
or U8858 (N_8858,N_8251,N_8156);
xnor U8859 (N_8859,N_8263,N_8504);
or U8860 (N_8860,N_8793,N_8267);
and U8861 (N_8861,N_8158,N_8666);
xor U8862 (N_8862,N_8588,N_8092);
nor U8863 (N_8863,N_8196,N_8799);
nand U8864 (N_8864,N_8610,N_8314);
nand U8865 (N_8865,N_8019,N_8660);
or U8866 (N_8866,N_8198,N_8683);
or U8867 (N_8867,N_8736,N_8070);
or U8868 (N_8868,N_8608,N_8001);
nand U8869 (N_8869,N_8043,N_8442);
xnor U8870 (N_8870,N_8125,N_8060);
xnor U8871 (N_8871,N_8496,N_8554);
nand U8872 (N_8872,N_8705,N_8360);
nand U8873 (N_8873,N_8400,N_8686);
nor U8874 (N_8874,N_8680,N_8340);
nand U8875 (N_8875,N_8231,N_8336);
xor U8876 (N_8876,N_8180,N_8261);
nor U8877 (N_8877,N_8020,N_8624);
xnor U8878 (N_8878,N_8364,N_8188);
and U8879 (N_8879,N_8380,N_8634);
nor U8880 (N_8880,N_8247,N_8044);
nor U8881 (N_8881,N_8693,N_8331);
nand U8882 (N_8882,N_8700,N_8655);
or U8883 (N_8883,N_8038,N_8566);
xor U8884 (N_8884,N_8516,N_8484);
xnor U8885 (N_8885,N_8378,N_8287);
nor U8886 (N_8886,N_8304,N_8408);
xor U8887 (N_8887,N_8144,N_8502);
nand U8888 (N_8888,N_8110,N_8451);
or U8889 (N_8889,N_8226,N_8711);
nand U8890 (N_8890,N_8220,N_8232);
nor U8891 (N_8891,N_8082,N_8093);
or U8892 (N_8892,N_8111,N_8123);
and U8893 (N_8893,N_8518,N_8584);
and U8894 (N_8894,N_8510,N_8425);
or U8895 (N_8895,N_8383,N_8459);
nor U8896 (N_8896,N_8678,N_8138);
nand U8897 (N_8897,N_8187,N_8177);
nor U8898 (N_8898,N_8195,N_8573);
nand U8899 (N_8899,N_8754,N_8358);
and U8900 (N_8900,N_8074,N_8391);
or U8901 (N_8901,N_8493,N_8620);
nand U8902 (N_8902,N_8170,N_8507);
or U8903 (N_8903,N_8371,N_8473);
nand U8904 (N_8904,N_8339,N_8537);
nand U8905 (N_8905,N_8406,N_8482);
nor U8906 (N_8906,N_8292,N_8611);
and U8907 (N_8907,N_8595,N_8677);
or U8908 (N_8908,N_8076,N_8409);
or U8909 (N_8909,N_8778,N_8270);
xor U8910 (N_8910,N_8337,N_8037);
xor U8911 (N_8911,N_8768,N_8593);
xnor U8912 (N_8912,N_8527,N_8604);
xor U8913 (N_8913,N_8613,N_8649);
and U8914 (N_8914,N_8404,N_8720);
or U8915 (N_8915,N_8707,N_8780);
nand U8916 (N_8916,N_8249,N_8519);
and U8917 (N_8917,N_8034,N_8405);
nor U8918 (N_8918,N_8018,N_8556);
xor U8919 (N_8919,N_8167,N_8745);
or U8920 (N_8920,N_8040,N_8176);
nor U8921 (N_8921,N_8143,N_8388);
or U8922 (N_8922,N_8435,N_8694);
or U8923 (N_8923,N_8441,N_8230);
nand U8924 (N_8924,N_8448,N_8418);
nand U8925 (N_8925,N_8329,N_8695);
xor U8926 (N_8926,N_8779,N_8760);
xor U8927 (N_8927,N_8283,N_8587);
nand U8928 (N_8928,N_8255,N_8450);
or U8929 (N_8929,N_8228,N_8455);
or U8930 (N_8930,N_8015,N_8648);
or U8931 (N_8931,N_8559,N_8434);
nand U8932 (N_8932,N_8327,N_8363);
nor U8933 (N_8933,N_8084,N_8150);
or U8934 (N_8934,N_8280,N_8157);
and U8935 (N_8935,N_8245,N_8574);
xnor U8936 (N_8936,N_8091,N_8126);
nand U8937 (N_8937,N_8658,N_8214);
nor U8938 (N_8938,N_8352,N_8673);
xnor U8939 (N_8939,N_8264,N_8059);
nand U8940 (N_8940,N_8108,N_8464);
nand U8941 (N_8941,N_8302,N_8715);
nor U8942 (N_8942,N_8762,N_8517);
nand U8943 (N_8943,N_8315,N_8178);
and U8944 (N_8944,N_8029,N_8365);
nor U8945 (N_8945,N_8446,N_8310);
nor U8946 (N_8946,N_8600,N_8787);
nor U8947 (N_8947,N_8007,N_8119);
and U8948 (N_8948,N_8643,N_8419);
nor U8949 (N_8949,N_8576,N_8353);
nor U8950 (N_8950,N_8794,N_8426);
and U8951 (N_8951,N_8164,N_8319);
and U8952 (N_8952,N_8166,N_8728);
xor U8953 (N_8953,N_8115,N_8541);
nand U8954 (N_8954,N_8689,N_8306);
nand U8955 (N_8955,N_8382,N_8374);
and U8956 (N_8956,N_8146,N_8531);
and U8957 (N_8957,N_8117,N_8324);
nor U8958 (N_8958,N_8325,N_8549);
or U8959 (N_8959,N_8023,N_8189);
nand U8960 (N_8960,N_8797,N_8569);
nand U8961 (N_8961,N_8055,N_8343);
and U8962 (N_8962,N_8077,N_8172);
nor U8963 (N_8963,N_8369,N_8664);
nor U8964 (N_8964,N_8348,N_8309);
nand U8965 (N_8965,N_8751,N_8767);
and U8966 (N_8966,N_8016,N_8756);
or U8967 (N_8967,N_8490,N_8056);
nor U8968 (N_8968,N_8417,N_8663);
nand U8969 (N_8969,N_8497,N_8002);
nor U8970 (N_8970,N_8069,N_8470);
nand U8971 (N_8971,N_8730,N_8242);
nand U8972 (N_8972,N_8386,N_8021);
nor U8973 (N_8973,N_8719,N_8513);
or U8974 (N_8974,N_8116,N_8357);
nand U8975 (N_8975,N_8640,N_8712);
nor U8976 (N_8976,N_8474,N_8581);
or U8977 (N_8977,N_8349,N_8632);
or U8978 (N_8978,N_8181,N_8617);
nand U8979 (N_8979,N_8792,N_8253);
nand U8980 (N_8980,N_8027,N_8668);
nand U8981 (N_8981,N_8506,N_8453);
nand U8982 (N_8982,N_8185,N_8625);
or U8983 (N_8983,N_8390,N_8252);
nor U8984 (N_8984,N_8449,N_8145);
nand U8985 (N_8985,N_8533,N_8335);
nand U8986 (N_8986,N_8042,N_8203);
nand U8987 (N_8987,N_8500,N_8136);
or U8988 (N_8988,N_8224,N_8615);
nand U8989 (N_8989,N_8539,N_8121);
nor U8990 (N_8990,N_8362,N_8621);
and U8991 (N_8991,N_8248,N_8175);
or U8992 (N_8992,N_8278,N_8681);
and U8993 (N_8993,N_8258,N_8279);
xnor U8994 (N_8994,N_8114,N_8704);
and U8995 (N_8995,N_8536,N_8701);
nand U8996 (N_8996,N_8684,N_8207);
or U8997 (N_8997,N_8414,N_8530);
or U8998 (N_8998,N_8551,N_8472);
xnor U8999 (N_8999,N_8266,N_8216);
and U9000 (N_9000,N_8141,N_8739);
xnor U9001 (N_9001,N_8465,N_8692);
nor U9002 (N_9002,N_8674,N_8259);
or U9003 (N_9003,N_8421,N_8078);
nor U9004 (N_9004,N_8046,N_8706);
nand U9005 (N_9005,N_8783,N_8330);
or U9006 (N_9006,N_8650,N_8697);
and U9007 (N_9007,N_8651,N_8403);
or U9008 (N_9008,N_8733,N_8612);
nand U9009 (N_9009,N_8740,N_8729);
or U9010 (N_9010,N_8665,N_8222);
and U9011 (N_9011,N_8713,N_8384);
xnor U9012 (N_9012,N_8402,N_8477);
nand U9013 (N_9013,N_8127,N_8734);
or U9014 (N_9014,N_8645,N_8570);
or U9015 (N_9015,N_8737,N_8328);
xor U9016 (N_9016,N_8169,N_8320);
or U9017 (N_9017,N_8047,N_8460);
and U9018 (N_9018,N_8749,N_8299);
xor U9019 (N_9019,N_8440,N_8798);
or U9020 (N_9020,N_8423,N_8437);
nand U9021 (N_9021,N_8535,N_8061);
nor U9022 (N_9022,N_8457,N_8239);
and U9023 (N_9023,N_8416,N_8233);
xor U9024 (N_9024,N_8396,N_8322);
nand U9025 (N_9025,N_8183,N_8308);
xnor U9026 (N_9026,N_8068,N_8432);
or U9027 (N_9027,N_8725,N_8033);
xor U9028 (N_9028,N_8087,N_8162);
and U9029 (N_9029,N_8785,N_8347);
or U9030 (N_9030,N_8035,N_8572);
nor U9031 (N_9031,N_8716,N_8489);
xnor U9032 (N_9032,N_8596,N_8269);
and U9033 (N_9033,N_8301,N_8759);
xor U9034 (N_9034,N_8702,N_8036);
and U9035 (N_9035,N_8546,N_8237);
xor U9036 (N_9036,N_8721,N_8795);
and U9037 (N_9037,N_8622,N_8151);
nand U9038 (N_9038,N_8726,N_8469);
and U9039 (N_9039,N_8774,N_8244);
or U9040 (N_9040,N_8101,N_8190);
and U9041 (N_9041,N_8750,N_8698);
nor U9042 (N_9042,N_8782,N_8392);
or U9043 (N_9043,N_8105,N_8652);
nand U9044 (N_9044,N_8095,N_8148);
nor U9045 (N_9045,N_8168,N_8109);
xor U9046 (N_9046,N_8508,N_8086);
or U9047 (N_9047,N_8636,N_8064);
or U9048 (N_9048,N_8275,N_8366);
nor U9049 (N_9049,N_8107,N_8466);
xnor U9050 (N_9050,N_8526,N_8647);
and U9051 (N_9051,N_8462,N_8332);
xnor U9052 (N_9052,N_8379,N_8028);
nor U9053 (N_9053,N_8544,N_8209);
or U9054 (N_9054,N_8717,N_8375);
and U9055 (N_9055,N_8542,N_8149);
xnor U9056 (N_9056,N_8219,N_8118);
and U9057 (N_9057,N_8367,N_8385);
nor U9058 (N_9058,N_8557,N_8747);
or U9059 (N_9059,N_8765,N_8140);
nand U9060 (N_9060,N_8297,N_8427);
and U9061 (N_9061,N_8454,N_8743);
or U9062 (N_9062,N_8598,N_8083);
nor U9063 (N_9063,N_8057,N_8644);
and U9064 (N_9064,N_8213,N_8234);
and U9065 (N_9065,N_8528,N_8065);
and U9066 (N_9066,N_8268,N_8467);
xnor U9067 (N_9067,N_8488,N_8241);
or U9068 (N_9068,N_8578,N_8004);
nor U9069 (N_9069,N_8205,N_8642);
nor U9070 (N_9070,N_8184,N_8293);
nand U9071 (N_9071,N_8236,N_8724);
or U9072 (N_9072,N_8271,N_8192);
and U9073 (N_9073,N_8703,N_8577);
or U9074 (N_9074,N_8676,N_8415);
nand U9075 (N_9075,N_8017,N_8654);
or U9076 (N_9076,N_8512,N_8659);
nand U9077 (N_9077,N_8025,N_8351);
and U9078 (N_9078,N_8710,N_8088);
nor U9079 (N_9079,N_8090,N_8395);
nand U9080 (N_9080,N_8532,N_8341);
or U9081 (N_9081,N_8394,N_8381);
or U9082 (N_9082,N_8265,N_8605);
and U9083 (N_9083,N_8133,N_8286);
nand U9084 (N_9084,N_8452,N_8334);
xor U9085 (N_9085,N_8769,N_8709);
nor U9086 (N_9086,N_8429,N_8511);
and U9087 (N_9087,N_8727,N_8113);
xor U9088 (N_9088,N_8128,N_8491);
xnor U9089 (N_9089,N_8662,N_8250);
or U9090 (N_9090,N_8152,N_8746);
nor U9091 (N_9091,N_8669,N_8431);
xnor U9092 (N_9092,N_8321,N_8579);
nor U9093 (N_9093,N_8410,N_8206);
nor U9094 (N_9094,N_8355,N_8682);
and U9095 (N_9095,N_8407,N_8359);
nor U9096 (N_9096,N_8627,N_8524);
xnor U9097 (N_9097,N_8420,N_8691);
or U9098 (N_9098,N_8300,N_8106);
nor U9099 (N_9099,N_8763,N_8790);
nor U9100 (N_9100,N_8137,N_8097);
nand U9101 (N_9101,N_8742,N_8398);
nand U9102 (N_9102,N_8240,N_8458);
nand U9103 (N_9103,N_8548,N_8439);
or U9104 (N_9104,N_8560,N_8591);
or U9105 (N_9105,N_8468,N_8633);
and U9106 (N_9106,N_8030,N_8534);
nand U9107 (N_9107,N_8313,N_8290);
or U9108 (N_9108,N_8494,N_8350);
or U9109 (N_9109,N_8586,N_8142);
nand U9110 (N_9110,N_8521,N_8066);
nand U9111 (N_9111,N_8563,N_8098);
xor U9112 (N_9112,N_8102,N_8744);
nand U9113 (N_9113,N_8776,N_8104);
nand U9114 (N_9114,N_8479,N_8303);
nor U9115 (N_9115,N_8285,N_8024);
and U9116 (N_9116,N_8443,N_8227);
or U9117 (N_9117,N_8032,N_8134);
nand U9118 (N_9118,N_8638,N_8679);
and U9119 (N_9119,N_8342,N_8773);
and U9120 (N_9120,N_8646,N_8525);
and U9121 (N_9121,N_8444,N_8592);
or U9122 (N_9122,N_8583,N_8289);
or U9123 (N_9123,N_8550,N_8413);
xor U9124 (N_9124,N_8052,N_8555);
or U9125 (N_9125,N_8771,N_8738);
nor U9126 (N_9126,N_8256,N_8637);
and U9127 (N_9127,N_8626,N_8039);
or U9128 (N_9128,N_8770,N_8486);
and U9129 (N_9129,N_8463,N_8218);
nor U9130 (N_9130,N_8003,N_8079);
nand U9131 (N_9131,N_8687,N_8599);
or U9132 (N_9132,N_8412,N_8051);
or U9133 (N_9133,N_8796,N_8401);
or U9134 (N_9134,N_8159,N_8096);
or U9135 (N_9135,N_8130,N_8201);
nor U9136 (N_9136,N_8672,N_8008);
nor U9137 (N_9137,N_8171,N_8476);
xnor U9138 (N_9138,N_8564,N_8561);
nand U9139 (N_9139,N_8430,N_8161);
nand U9140 (N_9140,N_8212,N_8235);
xor U9141 (N_9141,N_8131,N_8080);
xor U9142 (N_9142,N_8154,N_8616);
or U9143 (N_9143,N_8791,N_8670);
nand U9144 (N_9144,N_8389,N_8520);
xor U9145 (N_9145,N_8656,N_8215);
or U9146 (N_9146,N_8732,N_8775);
and U9147 (N_9147,N_8174,N_8075);
nor U9148 (N_9148,N_8688,N_8387);
or U9149 (N_9149,N_8433,N_8100);
nand U9150 (N_9150,N_8786,N_8399);
nor U9151 (N_9151,N_8607,N_8072);
nor U9152 (N_9152,N_8282,N_8155);
nor U9153 (N_9153,N_8631,N_8514);
nand U9154 (N_9154,N_8054,N_8653);
and U9155 (N_9155,N_8050,N_8197);
xnor U9156 (N_9156,N_8480,N_8022);
nand U9157 (N_9157,N_8580,N_8492);
and U9158 (N_9158,N_8011,N_8718);
xnor U9159 (N_9159,N_8481,N_8619);
and U9160 (N_9160,N_8333,N_8058);
and U9161 (N_9161,N_8567,N_8714);
nor U9162 (N_9162,N_8229,N_8553);
xnor U9163 (N_9163,N_8296,N_8295);
and U9164 (N_9164,N_8120,N_8200);
or U9165 (N_9165,N_8523,N_8173);
or U9166 (N_9166,N_8509,N_8602);
nor U9167 (N_9167,N_8208,N_8210);
nand U9168 (N_9168,N_8129,N_8505);
nor U9169 (N_9169,N_8722,N_8163);
and U9170 (N_9170,N_8428,N_8273);
nand U9171 (N_9171,N_8376,N_8628);
and U9172 (N_9172,N_8657,N_8132);
and U9173 (N_9173,N_8755,N_8294);
nand U9174 (N_9174,N_8191,N_8257);
or U9175 (N_9175,N_8014,N_8667);
nand U9176 (N_9176,N_8288,N_8538);
xor U9177 (N_9177,N_8515,N_8623);
xor U9178 (N_9178,N_8276,N_8447);
and U9179 (N_9179,N_8606,N_8397);
nand U9180 (N_9180,N_8708,N_8194);
xor U9181 (N_9181,N_8006,N_8748);
nand U9182 (N_9182,N_8031,N_8629);
and U9183 (N_9183,N_8073,N_8478);
nand U9184 (N_9184,N_8575,N_8026);
nor U9185 (N_9185,N_8552,N_8274);
nand U9186 (N_9186,N_8471,N_8368);
nor U9187 (N_9187,N_8254,N_8316);
nand U9188 (N_9188,N_8160,N_8757);
xnor U9189 (N_9189,N_8305,N_8323);
xor U9190 (N_9190,N_8735,N_8193);
nand U9191 (N_9191,N_8000,N_8089);
nand U9192 (N_9192,N_8307,N_8243);
or U9193 (N_9193,N_8761,N_8298);
and U9194 (N_9194,N_8540,N_8501);
nand U9195 (N_9195,N_8281,N_8067);
xor U9196 (N_9196,N_8422,N_8199);
xnor U9197 (N_9197,N_8221,N_8731);
nor U9198 (N_9198,N_8475,N_8685);
nand U9199 (N_9199,N_8696,N_8661);
xnor U9200 (N_9200,N_8598,N_8305);
xnor U9201 (N_9201,N_8494,N_8396);
nor U9202 (N_9202,N_8302,N_8168);
xnor U9203 (N_9203,N_8796,N_8005);
or U9204 (N_9204,N_8677,N_8644);
nor U9205 (N_9205,N_8260,N_8274);
xor U9206 (N_9206,N_8609,N_8720);
or U9207 (N_9207,N_8227,N_8150);
and U9208 (N_9208,N_8092,N_8073);
and U9209 (N_9209,N_8765,N_8745);
nor U9210 (N_9210,N_8744,N_8482);
nor U9211 (N_9211,N_8454,N_8655);
nor U9212 (N_9212,N_8733,N_8378);
nor U9213 (N_9213,N_8080,N_8013);
xor U9214 (N_9214,N_8528,N_8767);
xor U9215 (N_9215,N_8213,N_8255);
nand U9216 (N_9216,N_8505,N_8246);
nor U9217 (N_9217,N_8496,N_8648);
nor U9218 (N_9218,N_8443,N_8451);
xor U9219 (N_9219,N_8115,N_8221);
xnor U9220 (N_9220,N_8766,N_8087);
xor U9221 (N_9221,N_8765,N_8479);
nor U9222 (N_9222,N_8482,N_8694);
nor U9223 (N_9223,N_8692,N_8559);
nand U9224 (N_9224,N_8717,N_8492);
and U9225 (N_9225,N_8772,N_8411);
nor U9226 (N_9226,N_8252,N_8482);
or U9227 (N_9227,N_8417,N_8636);
and U9228 (N_9228,N_8473,N_8362);
nand U9229 (N_9229,N_8129,N_8458);
and U9230 (N_9230,N_8294,N_8290);
or U9231 (N_9231,N_8551,N_8241);
and U9232 (N_9232,N_8287,N_8666);
nand U9233 (N_9233,N_8641,N_8168);
xnor U9234 (N_9234,N_8641,N_8165);
nor U9235 (N_9235,N_8591,N_8182);
nand U9236 (N_9236,N_8274,N_8039);
or U9237 (N_9237,N_8498,N_8722);
nand U9238 (N_9238,N_8320,N_8474);
xor U9239 (N_9239,N_8258,N_8452);
nor U9240 (N_9240,N_8572,N_8566);
or U9241 (N_9241,N_8742,N_8696);
xor U9242 (N_9242,N_8654,N_8179);
or U9243 (N_9243,N_8254,N_8069);
or U9244 (N_9244,N_8274,N_8116);
xnor U9245 (N_9245,N_8042,N_8538);
nand U9246 (N_9246,N_8011,N_8504);
and U9247 (N_9247,N_8717,N_8793);
and U9248 (N_9248,N_8646,N_8780);
nand U9249 (N_9249,N_8522,N_8055);
or U9250 (N_9250,N_8682,N_8594);
nand U9251 (N_9251,N_8318,N_8105);
xor U9252 (N_9252,N_8770,N_8028);
and U9253 (N_9253,N_8096,N_8576);
xor U9254 (N_9254,N_8374,N_8336);
or U9255 (N_9255,N_8783,N_8643);
nand U9256 (N_9256,N_8246,N_8758);
and U9257 (N_9257,N_8774,N_8383);
or U9258 (N_9258,N_8689,N_8081);
and U9259 (N_9259,N_8167,N_8544);
or U9260 (N_9260,N_8553,N_8282);
xor U9261 (N_9261,N_8037,N_8738);
nor U9262 (N_9262,N_8241,N_8793);
nor U9263 (N_9263,N_8075,N_8412);
nor U9264 (N_9264,N_8195,N_8155);
and U9265 (N_9265,N_8624,N_8348);
nand U9266 (N_9266,N_8029,N_8509);
nor U9267 (N_9267,N_8566,N_8164);
xnor U9268 (N_9268,N_8581,N_8413);
xor U9269 (N_9269,N_8353,N_8796);
or U9270 (N_9270,N_8682,N_8579);
nor U9271 (N_9271,N_8383,N_8757);
xnor U9272 (N_9272,N_8408,N_8543);
nor U9273 (N_9273,N_8002,N_8395);
or U9274 (N_9274,N_8444,N_8624);
nand U9275 (N_9275,N_8707,N_8729);
or U9276 (N_9276,N_8600,N_8022);
nor U9277 (N_9277,N_8583,N_8190);
xor U9278 (N_9278,N_8653,N_8019);
or U9279 (N_9279,N_8009,N_8067);
and U9280 (N_9280,N_8487,N_8273);
xnor U9281 (N_9281,N_8082,N_8004);
and U9282 (N_9282,N_8260,N_8468);
nor U9283 (N_9283,N_8601,N_8328);
and U9284 (N_9284,N_8503,N_8630);
xor U9285 (N_9285,N_8369,N_8046);
nand U9286 (N_9286,N_8488,N_8028);
nor U9287 (N_9287,N_8268,N_8534);
xnor U9288 (N_9288,N_8569,N_8580);
and U9289 (N_9289,N_8635,N_8384);
or U9290 (N_9290,N_8761,N_8287);
or U9291 (N_9291,N_8641,N_8327);
xnor U9292 (N_9292,N_8293,N_8116);
and U9293 (N_9293,N_8446,N_8444);
nor U9294 (N_9294,N_8452,N_8594);
nand U9295 (N_9295,N_8267,N_8781);
and U9296 (N_9296,N_8439,N_8423);
nand U9297 (N_9297,N_8035,N_8778);
nor U9298 (N_9298,N_8524,N_8403);
and U9299 (N_9299,N_8099,N_8421);
nor U9300 (N_9300,N_8267,N_8743);
xnor U9301 (N_9301,N_8236,N_8122);
nand U9302 (N_9302,N_8129,N_8170);
or U9303 (N_9303,N_8713,N_8548);
xnor U9304 (N_9304,N_8005,N_8271);
and U9305 (N_9305,N_8071,N_8313);
nor U9306 (N_9306,N_8289,N_8481);
and U9307 (N_9307,N_8190,N_8246);
nand U9308 (N_9308,N_8098,N_8539);
nor U9309 (N_9309,N_8230,N_8280);
and U9310 (N_9310,N_8631,N_8119);
xor U9311 (N_9311,N_8155,N_8268);
xnor U9312 (N_9312,N_8587,N_8017);
and U9313 (N_9313,N_8173,N_8392);
and U9314 (N_9314,N_8177,N_8693);
nand U9315 (N_9315,N_8370,N_8782);
and U9316 (N_9316,N_8634,N_8301);
or U9317 (N_9317,N_8711,N_8408);
xnor U9318 (N_9318,N_8664,N_8207);
nand U9319 (N_9319,N_8776,N_8784);
nor U9320 (N_9320,N_8131,N_8501);
xor U9321 (N_9321,N_8420,N_8154);
nor U9322 (N_9322,N_8516,N_8532);
nand U9323 (N_9323,N_8521,N_8260);
or U9324 (N_9324,N_8738,N_8490);
or U9325 (N_9325,N_8027,N_8682);
nand U9326 (N_9326,N_8512,N_8776);
xnor U9327 (N_9327,N_8399,N_8159);
nand U9328 (N_9328,N_8786,N_8357);
or U9329 (N_9329,N_8543,N_8681);
or U9330 (N_9330,N_8203,N_8564);
or U9331 (N_9331,N_8117,N_8430);
nand U9332 (N_9332,N_8474,N_8076);
nand U9333 (N_9333,N_8089,N_8440);
nor U9334 (N_9334,N_8433,N_8740);
and U9335 (N_9335,N_8430,N_8597);
or U9336 (N_9336,N_8462,N_8529);
or U9337 (N_9337,N_8146,N_8087);
nor U9338 (N_9338,N_8122,N_8256);
nor U9339 (N_9339,N_8170,N_8728);
nand U9340 (N_9340,N_8762,N_8774);
and U9341 (N_9341,N_8273,N_8443);
nand U9342 (N_9342,N_8024,N_8646);
and U9343 (N_9343,N_8283,N_8655);
or U9344 (N_9344,N_8715,N_8137);
nor U9345 (N_9345,N_8532,N_8489);
and U9346 (N_9346,N_8074,N_8315);
or U9347 (N_9347,N_8251,N_8231);
xnor U9348 (N_9348,N_8434,N_8490);
nor U9349 (N_9349,N_8170,N_8174);
nand U9350 (N_9350,N_8233,N_8364);
xor U9351 (N_9351,N_8573,N_8596);
and U9352 (N_9352,N_8789,N_8596);
or U9353 (N_9353,N_8419,N_8586);
and U9354 (N_9354,N_8640,N_8760);
or U9355 (N_9355,N_8407,N_8778);
or U9356 (N_9356,N_8290,N_8352);
xnor U9357 (N_9357,N_8157,N_8547);
nand U9358 (N_9358,N_8353,N_8384);
nand U9359 (N_9359,N_8370,N_8564);
and U9360 (N_9360,N_8310,N_8706);
xnor U9361 (N_9361,N_8558,N_8036);
xor U9362 (N_9362,N_8735,N_8620);
xnor U9363 (N_9363,N_8167,N_8647);
xnor U9364 (N_9364,N_8442,N_8762);
and U9365 (N_9365,N_8022,N_8770);
or U9366 (N_9366,N_8300,N_8701);
or U9367 (N_9367,N_8456,N_8412);
or U9368 (N_9368,N_8157,N_8689);
xor U9369 (N_9369,N_8222,N_8346);
xnor U9370 (N_9370,N_8422,N_8260);
nand U9371 (N_9371,N_8349,N_8586);
nor U9372 (N_9372,N_8140,N_8697);
or U9373 (N_9373,N_8691,N_8032);
nand U9374 (N_9374,N_8447,N_8430);
xor U9375 (N_9375,N_8708,N_8091);
nor U9376 (N_9376,N_8041,N_8170);
and U9377 (N_9377,N_8087,N_8702);
xnor U9378 (N_9378,N_8215,N_8062);
nand U9379 (N_9379,N_8214,N_8231);
nor U9380 (N_9380,N_8655,N_8172);
or U9381 (N_9381,N_8373,N_8181);
or U9382 (N_9382,N_8509,N_8122);
xnor U9383 (N_9383,N_8114,N_8448);
or U9384 (N_9384,N_8322,N_8274);
and U9385 (N_9385,N_8317,N_8658);
nand U9386 (N_9386,N_8173,N_8053);
or U9387 (N_9387,N_8397,N_8415);
and U9388 (N_9388,N_8201,N_8194);
xnor U9389 (N_9389,N_8081,N_8459);
nor U9390 (N_9390,N_8049,N_8520);
or U9391 (N_9391,N_8217,N_8563);
and U9392 (N_9392,N_8117,N_8638);
or U9393 (N_9393,N_8298,N_8665);
and U9394 (N_9394,N_8002,N_8256);
and U9395 (N_9395,N_8079,N_8125);
xor U9396 (N_9396,N_8493,N_8223);
nor U9397 (N_9397,N_8515,N_8060);
xnor U9398 (N_9398,N_8280,N_8650);
or U9399 (N_9399,N_8469,N_8032);
and U9400 (N_9400,N_8162,N_8478);
nor U9401 (N_9401,N_8627,N_8635);
xnor U9402 (N_9402,N_8146,N_8611);
and U9403 (N_9403,N_8723,N_8732);
or U9404 (N_9404,N_8388,N_8169);
xnor U9405 (N_9405,N_8352,N_8634);
and U9406 (N_9406,N_8029,N_8254);
nand U9407 (N_9407,N_8593,N_8648);
nor U9408 (N_9408,N_8600,N_8127);
nor U9409 (N_9409,N_8695,N_8619);
and U9410 (N_9410,N_8154,N_8407);
xor U9411 (N_9411,N_8537,N_8497);
and U9412 (N_9412,N_8535,N_8166);
and U9413 (N_9413,N_8036,N_8226);
and U9414 (N_9414,N_8787,N_8105);
nand U9415 (N_9415,N_8041,N_8121);
and U9416 (N_9416,N_8445,N_8682);
xnor U9417 (N_9417,N_8148,N_8370);
and U9418 (N_9418,N_8242,N_8659);
nor U9419 (N_9419,N_8515,N_8760);
nand U9420 (N_9420,N_8764,N_8119);
and U9421 (N_9421,N_8751,N_8026);
and U9422 (N_9422,N_8213,N_8034);
and U9423 (N_9423,N_8623,N_8777);
xor U9424 (N_9424,N_8084,N_8144);
nor U9425 (N_9425,N_8550,N_8768);
xnor U9426 (N_9426,N_8056,N_8788);
and U9427 (N_9427,N_8540,N_8244);
xor U9428 (N_9428,N_8503,N_8265);
xnor U9429 (N_9429,N_8776,N_8627);
xnor U9430 (N_9430,N_8408,N_8075);
and U9431 (N_9431,N_8569,N_8558);
xor U9432 (N_9432,N_8626,N_8629);
nor U9433 (N_9433,N_8031,N_8667);
or U9434 (N_9434,N_8091,N_8401);
xnor U9435 (N_9435,N_8704,N_8084);
xor U9436 (N_9436,N_8458,N_8545);
nand U9437 (N_9437,N_8233,N_8081);
nand U9438 (N_9438,N_8044,N_8280);
or U9439 (N_9439,N_8268,N_8232);
and U9440 (N_9440,N_8357,N_8492);
and U9441 (N_9441,N_8193,N_8183);
or U9442 (N_9442,N_8424,N_8116);
xor U9443 (N_9443,N_8437,N_8570);
or U9444 (N_9444,N_8384,N_8620);
xor U9445 (N_9445,N_8638,N_8674);
nor U9446 (N_9446,N_8349,N_8300);
and U9447 (N_9447,N_8753,N_8691);
nor U9448 (N_9448,N_8777,N_8011);
xnor U9449 (N_9449,N_8096,N_8179);
nand U9450 (N_9450,N_8315,N_8551);
xnor U9451 (N_9451,N_8689,N_8587);
and U9452 (N_9452,N_8665,N_8542);
nor U9453 (N_9453,N_8583,N_8346);
or U9454 (N_9454,N_8383,N_8533);
and U9455 (N_9455,N_8179,N_8330);
xor U9456 (N_9456,N_8169,N_8194);
and U9457 (N_9457,N_8439,N_8520);
xnor U9458 (N_9458,N_8436,N_8737);
xor U9459 (N_9459,N_8195,N_8268);
or U9460 (N_9460,N_8105,N_8093);
xor U9461 (N_9461,N_8627,N_8261);
nor U9462 (N_9462,N_8691,N_8292);
or U9463 (N_9463,N_8093,N_8362);
or U9464 (N_9464,N_8058,N_8747);
nand U9465 (N_9465,N_8534,N_8636);
and U9466 (N_9466,N_8583,N_8572);
xnor U9467 (N_9467,N_8448,N_8084);
and U9468 (N_9468,N_8789,N_8636);
and U9469 (N_9469,N_8358,N_8772);
nor U9470 (N_9470,N_8025,N_8193);
xnor U9471 (N_9471,N_8056,N_8102);
or U9472 (N_9472,N_8402,N_8354);
and U9473 (N_9473,N_8167,N_8698);
nor U9474 (N_9474,N_8417,N_8635);
nand U9475 (N_9475,N_8282,N_8111);
and U9476 (N_9476,N_8785,N_8729);
nand U9477 (N_9477,N_8034,N_8323);
nor U9478 (N_9478,N_8740,N_8107);
xor U9479 (N_9479,N_8736,N_8429);
nor U9480 (N_9480,N_8380,N_8639);
xor U9481 (N_9481,N_8595,N_8151);
or U9482 (N_9482,N_8528,N_8042);
nand U9483 (N_9483,N_8724,N_8383);
xnor U9484 (N_9484,N_8508,N_8200);
nand U9485 (N_9485,N_8536,N_8563);
nor U9486 (N_9486,N_8741,N_8590);
and U9487 (N_9487,N_8540,N_8424);
and U9488 (N_9488,N_8406,N_8613);
and U9489 (N_9489,N_8073,N_8766);
or U9490 (N_9490,N_8360,N_8058);
or U9491 (N_9491,N_8385,N_8455);
nor U9492 (N_9492,N_8122,N_8314);
nand U9493 (N_9493,N_8614,N_8511);
nand U9494 (N_9494,N_8661,N_8764);
or U9495 (N_9495,N_8319,N_8156);
nand U9496 (N_9496,N_8099,N_8529);
or U9497 (N_9497,N_8431,N_8799);
nor U9498 (N_9498,N_8018,N_8340);
xnor U9499 (N_9499,N_8605,N_8176);
xor U9500 (N_9500,N_8213,N_8662);
and U9501 (N_9501,N_8628,N_8737);
xnor U9502 (N_9502,N_8260,N_8065);
xnor U9503 (N_9503,N_8765,N_8519);
and U9504 (N_9504,N_8635,N_8729);
nand U9505 (N_9505,N_8725,N_8040);
and U9506 (N_9506,N_8042,N_8378);
nor U9507 (N_9507,N_8151,N_8662);
and U9508 (N_9508,N_8695,N_8420);
nand U9509 (N_9509,N_8146,N_8401);
nand U9510 (N_9510,N_8748,N_8310);
and U9511 (N_9511,N_8026,N_8346);
and U9512 (N_9512,N_8319,N_8392);
or U9513 (N_9513,N_8528,N_8591);
nand U9514 (N_9514,N_8529,N_8239);
or U9515 (N_9515,N_8147,N_8788);
xnor U9516 (N_9516,N_8231,N_8786);
xor U9517 (N_9517,N_8463,N_8291);
nand U9518 (N_9518,N_8794,N_8721);
nor U9519 (N_9519,N_8165,N_8657);
xor U9520 (N_9520,N_8109,N_8487);
nand U9521 (N_9521,N_8487,N_8560);
nor U9522 (N_9522,N_8040,N_8518);
nand U9523 (N_9523,N_8703,N_8304);
nand U9524 (N_9524,N_8458,N_8792);
and U9525 (N_9525,N_8285,N_8761);
nor U9526 (N_9526,N_8184,N_8060);
xnor U9527 (N_9527,N_8588,N_8286);
nand U9528 (N_9528,N_8039,N_8371);
nor U9529 (N_9529,N_8215,N_8144);
and U9530 (N_9530,N_8157,N_8137);
nand U9531 (N_9531,N_8653,N_8098);
xnor U9532 (N_9532,N_8733,N_8530);
nor U9533 (N_9533,N_8744,N_8020);
nand U9534 (N_9534,N_8455,N_8552);
nand U9535 (N_9535,N_8384,N_8765);
or U9536 (N_9536,N_8222,N_8495);
xnor U9537 (N_9537,N_8581,N_8273);
nor U9538 (N_9538,N_8664,N_8167);
and U9539 (N_9539,N_8170,N_8648);
or U9540 (N_9540,N_8369,N_8465);
or U9541 (N_9541,N_8667,N_8117);
nand U9542 (N_9542,N_8048,N_8756);
nand U9543 (N_9543,N_8694,N_8692);
or U9544 (N_9544,N_8337,N_8229);
and U9545 (N_9545,N_8688,N_8460);
or U9546 (N_9546,N_8537,N_8456);
nor U9547 (N_9547,N_8402,N_8790);
xor U9548 (N_9548,N_8340,N_8584);
xnor U9549 (N_9549,N_8031,N_8307);
or U9550 (N_9550,N_8418,N_8158);
and U9551 (N_9551,N_8485,N_8586);
and U9552 (N_9552,N_8629,N_8458);
nand U9553 (N_9553,N_8724,N_8281);
nand U9554 (N_9554,N_8491,N_8681);
or U9555 (N_9555,N_8715,N_8072);
or U9556 (N_9556,N_8158,N_8076);
and U9557 (N_9557,N_8574,N_8181);
nand U9558 (N_9558,N_8179,N_8338);
or U9559 (N_9559,N_8796,N_8325);
nor U9560 (N_9560,N_8072,N_8361);
and U9561 (N_9561,N_8114,N_8208);
xor U9562 (N_9562,N_8078,N_8282);
nand U9563 (N_9563,N_8602,N_8450);
xor U9564 (N_9564,N_8531,N_8726);
xor U9565 (N_9565,N_8267,N_8792);
nor U9566 (N_9566,N_8713,N_8365);
xor U9567 (N_9567,N_8592,N_8562);
or U9568 (N_9568,N_8531,N_8600);
or U9569 (N_9569,N_8436,N_8249);
nand U9570 (N_9570,N_8556,N_8032);
xor U9571 (N_9571,N_8599,N_8406);
nor U9572 (N_9572,N_8207,N_8308);
nand U9573 (N_9573,N_8200,N_8647);
xnor U9574 (N_9574,N_8616,N_8209);
xor U9575 (N_9575,N_8325,N_8162);
and U9576 (N_9576,N_8586,N_8136);
xor U9577 (N_9577,N_8407,N_8423);
and U9578 (N_9578,N_8118,N_8379);
or U9579 (N_9579,N_8050,N_8796);
nand U9580 (N_9580,N_8292,N_8594);
nand U9581 (N_9581,N_8415,N_8209);
xnor U9582 (N_9582,N_8222,N_8010);
nand U9583 (N_9583,N_8268,N_8293);
nand U9584 (N_9584,N_8441,N_8132);
nor U9585 (N_9585,N_8297,N_8464);
xor U9586 (N_9586,N_8594,N_8344);
nor U9587 (N_9587,N_8322,N_8705);
xnor U9588 (N_9588,N_8642,N_8410);
xor U9589 (N_9589,N_8142,N_8186);
nand U9590 (N_9590,N_8095,N_8431);
xnor U9591 (N_9591,N_8249,N_8199);
nand U9592 (N_9592,N_8497,N_8368);
nor U9593 (N_9593,N_8192,N_8358);
xnor U9594 (N_9594,N_8590,N_8329);
nand U9595 (N_9595,N_8542,N_8588);
nand U9596 (N_9596,N_8310,N_8618);
and U9597 (N_9597,N_8676,N_8681);
xor U9598 (N_9598,N_8443,N_8542);
and U9599 (N_9599,N_8652,N_8558);
and U9600 (N_9600,N_9435,N_9144);
and U9601 (N_9601,N_8944,N_9349);
or U9602 (N_9602,N_9269,N_9221);
xor U9603 (N_9603,N_9500,N_9576);
and U9604 (N_9604,N_9208,N_8840);
nor U9605 (N_9605,N_9263,N_9053);
xor U9606 (N_9606,N_8909,N_9499);
or U9607 (N_9607,N_9241,N_9385);
xnor U9608 (N_9608,N_8984,N_9292);
and U9609 (N_9609,N_8947,N_9235);
xor U9610 (N_9610,N_9219,N_9578);
nor U9611 (N_9611,N_8910,N_9534);
or U9612 (N_9612,N_8849,N_8807);
or U9613 (N_9613,N_9587,N_9255);
nand U9614 (N_9614,N_9492,N_9428);
nor U9615 (N_9615,N_9001,N_9038);
xor U9616 (N_9616,N_9481,N_9515);
nor U9617 (N_9617,N_8899,N_9400);
nand U9618 (N_9618,N_8986,N_9555);
nor U9619 (N_9619,N_8813,N_9368);
nand U9620 (N_9620,N_9225,N_9384);
nand U9621 (N_9621,N_8943,N_8878);
nor U9622 (N_9622,N_9175,N_9130);
nor U9623 (N_9623,N_9011,N_9065);
or U9624 (N_9624,N_9405,N_8903);
nand U9625 (N_9625,N_9547,N_9033);
nor U9626 (N_9626,N_8806,N_9083);
or U9627 (N_9627,N_8845,N_9094);
nor U9628 (N_9628,N_9423,N_9062);
or U9629 (N_9629,N_9229,N_8847);
xnor U9630 (N_9630,N_9098,N_9359);
xnor U9631 (N_9631,N_9202,N_8988);
or U9632 (N_9632,N_9569,N_9309);
nor U9633 (N_9633,N_9126,N_9556);
and U9634 (N_9634,N_9333,N_9074);
nand U9635 (N_9635,N_9592,N_9138);
or U9636 (N_9636,N_8974,N_9482);
xnor U9637 (N_9637,N_9203,N_9174);
nor U9638 (N_9638,N_9531,N_9467);
and U9639 (N_9639,N_9490,N_8859);
xor U9640 (N_9640,N_9566,N_8976);
nand U9641 (N_9641,N_8851,N_9119);
xor U9642 (N_9642,N_9581,N_9313);
nand U9643 (N_9643,N_8980,N_8825);
xnor U9644 (N_9644,N_9565,N_9013);
nand U9645 (N_9645,N_9117,N_9502);
xnor U9646 (N_9646,N_9245,N_9549);
nand U9647 (N_9647,N_9442,N_8837);
nor U9648 (N_9648,N_9382,N_9527);
xnor U9649 (N_9649,N_8844,N_9319);
and U9650 (N_9650,N_8804,N_9217);
or U9651 (N_9651,N_9304,N_9373);
and U9652 (N_9652,N_9476,N_9586);
xor U9653 (N_9653,N_9332,N_9045);
xor U9654 (N_9654,N_9437,N_9051);
xnor U9655 (N_9655,N_9529,N_8811);
or U9656 (N_9656,N_9338,N_9157);
and U9657 (N_9657,N_9517,N_9550);
nor U9658 (N_9658,N_9109,N_9439);
xnor U9659 (N_9659,N_8870,N_9068);
xnor U9660 (N_9660,N_9369,N_9206);
nor U9661 (N_9661,N_8956,N_9543);
or U9662 (N_9662,N_9243,N_9315);
or U9663 (N_9663,N_9411,N_8889);
and U9664 (N_9664,N_9343,N_9105);
nor U9665 (N_9665,N_9034,N_9451);
nand U9666 (N_9666,N_9047,N_8805);
nand U9667 (N_9667,N_8820,N_9140);
nand U9668 (N_9668,N_9182,N_9307);
xnor U9669 (N_9669,N_9345,N_8936);
or U9670 (N_9670,N_9133,N_9267);
or U9671 (N_9671,N_9177,N_9380);
and U9672 (N_9672,N_8992,N_9378);
and U9673 (N_9673,N_9113,N_9060);
and U9674 (N_9674,N_9372,N_9455);
and U9675 (N_9675,N_8816,N_9535);
xor U9676 (N_9676,N_9357,N_9223);
nor U9677 (N_9677,N_8955,N_8832);
xnor U9678 (N_9678,N_9468,N_8921);
xnor U9679 (N_9679,N_8856,N_9327);
and U9680 (N_9680,N_9185,N_9471);
nor U9681 (N_9681,N_9295,N_9399);
xor U9682 (N_9682,N_9107,N_9247);
nor U9683 (N_9683,N_9453,N_9434);
xor U9684 (N_9684,N_9252,N_9344);
nor U9685 (N_9685,N_9134,N_8989);
nor U9686 (N_9686,N_9342,N_8959);
xnor U9687 (N_9687,N_9169,N_9323);
xor U9688 (N_9688,N_9283,N_8914);
xor U9689 (N_9689,N_9523,N_9008);
or U9690 (N_9690,N_9339,N_9422);
nand U9691 (N_9691,N_9386,N_9337);
nor U9692 (N_9692,N_9293,N_9306);
nor U9693 (N_9693,N_9579,N_9242);
or U9694 (N_9694,N_9533,N_9127);
nor U9695 (N_9695,N_8835,N_9154);
nor U9696 (N_9696,N_9539,N_8919);
nor U9697 (N_9697,N_8808,N_9312);
nand U9698 (N_9698,N_8862,N_9196);
xor U9699 (N_9699,N_9377,N_9446);
nand U9700 (N_9700,N_9262,N_8884);
and U9701 (N_9701,N_8841,N_9512);
or U9702 (N_9702,N_9186,N_9457);
nor U9703 (N_9703,N_8977,N_9049);
nor U9704 (N_9704,N_8890,N_9387);
xnor U9705 (N_9705,N_9155,N_9014);
nor U9706 (N_9706,N_9591,N_9129);
and U9707 (N_9707,N_8897,N_9559);
and U9708 (N_9708,N_9142,N_8821);
or U9709 (N_9709,N_9228,N_8915);
xnor U9710 (N_9710,N_8817,N_9006);
nand U9711 (N_9711,N_9264,N_8949);
nand U9712 (N_9712,N_9370,N_9136);
xnor U9713 (N_9713,N_9361,N_9141);
xnor U9714 (N_9714,N_9341,N_9234);
or U9715 (N_9715,N_9156,N_9398);
or U9716 (N_9716,N_9061,N_9139);
or U9717 (N_9717,N_9058,N_9272);
or U9718 (N_9718,N_9284,N_9183);
and U9719 (N_9719,N_9076,N_9198);
xnor U9720 (N_9720,N_8886,N_9145);
and U9721 (N_9721,N_9082,N_9450);
nor U9722 (N_9722,N_9078,N_9022);
nand U9723 (N_9723,N_9239,N_8892);
xnor U9724 (N_9724,N_8961,N_9021);
or U9725 (N_9725,N_9322,N_9355);
xnor U9726 (N_9726,N_9427,N_9577);
xnor U9727 (N_9727,N_8833,N_9005);
xnor U9728 (N_9728,N_9407,N_8998);
nor U9729 (N_9729,N_9394,N_9392);
nand U9730 (N_9730,N_9420,N_9470);
nor U9731 (N_9731,N_8920,N_9300);
nand U9732 (N_9732,N_8819,N_9390);
xor U9733 (N_9733,N_9280,N_9176);
nand U9734 (N_9734,N_9410,N_9258);
nor U9735 (N_9735,N_9436,N_9019);
and U9736 (N_9736,N_9506,N_9404);
nand U9737 (N_9737,N_9458,N_9230);
nor U9738 (N_9738,N_8829,N_9135);
xnor U9739 (N_9739,N_9417,N_8993);
or U9740 (N_9740,N_9393,N_9366);
nand U9741 (N_9741,N_9275,N_8893);
nor U9742 (N_9742,N_8957,N_8881);
or U9743 (N_9743,N_9189,N_8995);
nor U9744 (N_9744,N_9044,N_9236);
xor U9745 (N_9745,N_9023,N_9371);
and U9746 (N_9746,N_9055,N_9201);
nand U9747 (N_9747,N_9474,N_9429);
nand U9748 (N_9748,N_9112,N_9486);
nor U9749 (N_9749,N_9016,N_9305);
and U9750 (N_9750,N_8948,N_9032);
xor U9751 (N_9751,N_8963,N_9071);
or U9752 (N_9752,N_9268,N_9519);
xor U9753 (N_9753,N_8966,N_9584);
or U9754 (N_9754,N_9571,N_9415);
and U9755 (N_9755,N_9311,N_9360);
and U9756 (N_9756,N_9121,N_9334);
xnor U9757 (N_9757,N_9353,N_9180);
xor U9758 (N_9758,N_9583,N_9096);
and U9759 (N_9759,N_9103,N_9416);
and U9760 (N_9760,N_9246,N_8945);
nand U9761 (N_9761,N_8838,N_9012);
nand U9762 (N_9762,N_9197,N_9087);
nor U9763 (N_9763,N_8962,N_9250);
xor U9764 (N_9764,N_9102,N_9381);
nand U9765 (N_9765,N_9321,N_9421);
and U9766 (N_9766,N_9483,N_9518);
and U9767 (N_9767,N_9414,N_9495);
and U9768 (N_9768,N_9020,N_9494);
and U9769 (N_9769,N_9088,N_9317);
and U9770 (N_9770,N_9256,N_9541);
nand U9771 (N_9771,N_9340,N_9302);
nand U9772 (N_9772,N_8885,N_9279);
nand U9773 (N_9773,N_9009,N_9588);
and U9774 (N_9774,N_8991,N_9084);
nand U9775 (N_9775,N_9589,N_9454);
and U9776 (N_9776,N_9158,N_9278);
nor U9777 (N_9777,N_8887,N_9194);
and U9778 (N_9778,N_9290,N_9259);
and U9779 (N_9779,N_9173,N_9025);
or U9780 (N_9780,N_8818,N_9188);
or U9781 (N_9781,N_9568,N_9150);
xnor U9782 (N_9782,N_8934,N_9310);
and U9783 (N_9783,N_9063,N_8952);
or U9784 (N_9784,N_9191,N_9426);
or U9785 (N_9785,N_9090,N_9123);
nand U9786 (N_9786,N_9465,N_9159);
or U9787 (N_9787,N_9558,N_9299);
xnor U9788 (N_9788,N_8834,N_9433);
or U9789 (N_9789,N_9479,N_9298);
nor U9790 (N_9790,N_9402,N_9276);
nor U9791 (N_9791,N_9137,N_9570);
and U9792 (N_9792,N_9200,N_9513);
nor U9793 (N_9793,N_9171,N_9473);
nor U9794 (N_9794,N_9524,N_8891);
nand U9795 (N_9795,N_9598,N_9383);
or U9796 (N_9796,N_8800,N_8932);
nand U9797 (N_9797,N_8905,N_8894);
nor U9798 (N_9798,N_9120,N_9215);
nand U9799 (N_9799,N_9017,N_9296);
nor U9800 (N_9800,N_9093,N_8941);
xor U9801 (N_9801,N_9525,N_9408);
and U9802 (N_9802,N_8990,N_8940);
and U9803 (N_9803,N_8871,N_9358);
or U9804 (N_9804,N_9240,N_9035);
xnor U9805 (N_9805,N_8860,N_9132);
nand U9806 (N_9806,N_9362,N_9147);
nor U9807 (N_9807,N_9000,N_9031);
and U9808 (N_9808,N_9395,N_8868);
or U9809 (N_9809,N_9595,N_9554);
and U9810 (N_9810,N_9516,N_9503);
nor U9811 (N_9811,N_9287,N_9075);
or U9812 (N_9812,N_9431,N_8843);
and U9813 (N_9813,N_9324,N_9079);
and U9814 (N_9814,N_9462,N_8926);
or U9815 (N_9815,N_9346,N_9057);
or U9816 (N_9816,N_9222,N_9026);
nor U9817 (N_9817,N_8827,N_8857);
and U9818 (N_9818,N_9128,N_9209);
xor U9819 (N_9819,N_9104,N_8950);
nor U9820 (N_9820,N_8918,N_9118);
or U9821 (N_9821,N_8923,N_9046);
nand U9822 (N_9822,N_9593,N_9029);
or U9823 (N_9823,N_9507,N_8848);
nand U9824 (N_9824,N_9514,N_9597);
and U9825 (N_9825,N_8971,N_9248);
nor U9826 (N_9826,N_9281,N_9505);
or U9827 (N_9827,N_8907,N_9452);
nand U9828 (N_9828,N_9314,N_9548);
xor U9829 (N_9829,N_9214,N_9210);
nor U9830 (N_9830,N_9095,N_9489);
or U9831 (N_9831,N_8965,N_9178);
xnor U9832 (N_9832,N_9294,N_9067);
or U9833 (N_9833,N_8826,N_8802);
or U9834 (N_9834,N_9449,N_9412);
nor U9835 (N_9835,N_9594,N_9545);
or U9836 (N_9836,N_8994,N_9073);
nand U9837 (N_9837,N_9496,N_8902);
nand U9838 (N_9838,N_9165,N_9551);
nor U9839 (N_9839,N_8815,N_9184);
nor U9840 (N_9840,N_9010,N_9537);
nand U9841 (N_9841,N_9086,N_9389);
nand U9842 (N_9842,N_9430,N_9152);
and U9843 (N_9843,N_8876,N_8982);
and U9844 (N_9844,N_8896,N_9160);
and U9845 (N_9845,N_9270,N_8865);
nand U9846 (N_9846,N_9085,N_9316);
nand U9847 (N_9847,N_9397,N_8901);
nor U9848 (N_9848,N_9237,N_8978);
xnor U9849 (N_9849,N_9573,N_8972);
nor U9850 (N_9850,N_9375,N_9528);
nand U9851 (N_9851,N_8812,N_9520);
or U9852 (N_9852,N_8969,N_9596);
nand U9853 (N_9853,N_8852,N_9056);
and U9854 (N_9854,N_9567,N_9491);
or U9855 (N_9855,N_9125,N_9081);
or U9856 (N_9856,N_9042,N_8850);
nor U9857 (N_9857,N_9461,N_9050);
and U9858 (N_9858,N_9116,N_9167);
nor U9859 (N_9859,N_9401,N_9204);
nand U9860 (N_9860,N_8929,N_9273);
and U9861 (N_9861,N_9418,N_8908);
nor U9862 (N_9862,N_9227,N_9224);
nor U9863 (N_9863,N_9469,N_9580);
or U9864 (N_9864,N_8983,N_9388);
and U9865 (N_9865,N_9575,N_8916);
xor U9866 (N_9866,N_9018,N_9254);
nor U9867 (N_9867,N_9153,N_9146);
xnor U9868 (N_9868,N_9376,N_9560);
xor U9869 (N_9869,N_9493,N_8861);
nor U9870 (N_9870,N_8911,N_8999);
xnor U9871 (N_9871,N_8822,N_9466);
nor U9872 (N_9872,N_8904,N_9277);
nand U9873 (N_9873,N_9069,N_9162);
and U9874 (N_9874,N_8864,N_8900);
xor U9875 (N_9875,N_9599,N_9552);
xor U9876 (N_9876,N_9498,N_9027);
nand U9877 (N_9877,N_9522,N_8906);
xnor U9878 (N_9878,N_9266,N_9037);
and U9879 (N_9879,N_9562,N_9265);
nand U9880 (N_9880,N_9168,N_8973);
nor U9881 (N_9881,N_9301,N_9124);
or U9882 (N_9882,N_9438,N_8985);
nand U9883 (N_9883,N_9488,N_9211);
and U9884 (N_9884,N_9274,N_9582);
xnor U9885 (N_9885,N_8964,N_9257);
and U9886 (N_9886,N_9335,N_9179);
or U9887 (N_9887,N_9546,N_9557);
and U9888 (N_9888,N_9511,N_9424);
nand U9889 (N_9889,N_9540,N_9080);
nand U9890 (N_9890,N_9330,N_9553);
nor U9891 (N_9891,N_9015,N_8975);
or U9892 (N_9892,N_9478,N_8928);
xor U9893 (N_9893,N_8839,N_9477);
and U9894 (N_9894,N_8855,N_9028);
or U9895 (N_9895,N_9114,N_9318);
and U9896 (N_9896,N_9475,N_9059);
and U9897 (N_9897,N_9480,N_8867);
or U9898 (N_9898,N_9444,N_8853);
nor U9899 (N_9899,N_8938,N_8831);
xnor U9900 (N_9900,N_8927,N_9286);
nor U9901 (N_9901,N_9181,N_9365);
or U9902 (N_9902,N_8951,N_8933);
or U9903 (N_9903,N_8960,N_8968);
or U9904 (N_9904,N_9066,N_9585);
nor U9905 (N_9905,N_8967,N_9232);
nor U9906 (N_9906,N_9391,N_8924);
or U9907 (N_9907,N_8823,N_9226);
or U9908 (N_9908,N_9111,N_9413);
or U9909 (N_9909,N_8895,N_9149);
nand U9910 (N_9910,N_8937,N_9356);
or U9911 (N_9911,N_9070,N_9199);
and U9912 (N_9912,N_9289,N_8930);
nand U9913 (N_9913,N_9110,N_8953);
and U9914 (N_9914,N_8883,N_9521);
xnor U9915 (N_9915,N_9205,N_8879);
xnor U9916 (N_9916,N_9396,N_8996);
nor U9917 (N_9917,N_9538,N_9350);
xor U9918 (N_9918,N_9419,N_9445);
and U9919 (N_9919,N_9352,N_9106);
nor U9920 (N_9920,N_9406,N_8875);
nor U9921 (N_9921,N_8809,N_9542);
nand U9922 (N_9922,N_9097,N_9367);
and U9923 (N_9923,N_9054,N_9456);
nand U9924 (N_9924,N_9572,N_9320);
or U9925 (N_9925,N_9212,N_9448);
and U9926 (N_9926,N_9064,N_9003);
nand U9927 (N_9927,N_9260,N_9143);
and U9928 (N_9928,N_8869,N_9271);
xor U9929 (N_9929,N_8877,N_8874);
and U9930 (N_9930,N_8958,N_9099);
nor U9931 (N_9931,N_9509,N_9348);
or U9932 (N_9932,N_8880,N_9041);
nand U9933 (N_9933,N_9460,N_9484);
nor U9934 (N_9934,N_9002,N_9331);
or U9935 (N_9935,N_9363,N_9220);
and U9936 (N_9936,N_9115,N_8931);
or U9937 (N_9937,N_9308,N_9039);
or U9938 (N_9938,N_8846,N_9485);
xnor U9939 (N_9939,N_8946,N_9024);
nand U9940 (N_9940,N_9164,N_8814);
or U9941 (N_9941,N_9432,N_9303);
and U9942 (N_9942,N_9563,N_9166);
nor U9943 (N_9943,N_8801,N_9440);
xor U9944 (N_9944,N_9036,N_8935);
and U9945 (N_9945,N_8939,N_8970);
nand U9946 (N_9946,N_9092,N_8898);
or U9947 (N_9947,N_9233,N_9508);
or U9948 (N_9948,N_9195,N_9148);
and U9949 (N_9949,N_9285,N_8858);
xor U9950 (N_9950,N_8888,N_9443);
nand U9951 (N_9951,N_9379,N_8828);
and U9952 (N_9952,N_9472,N_9336);
and U9953 (N_9953,N_8942,N_9213);
nor U9954 (N_9954,N_9249,N_9077);
nand U9955 (N_9955,N_9192,N_8912);
xnor U9956 (N_9956,N_8917,N_9325);
nor U9957 (N_9957,N_9091,N_8913);
nor U9958 (N_9958,N_9030,N_9532);
or U9959 (N_9959,N_9590,N_9218);
and U9960 (N_9960,N_9328,N_9347);
nor U9961 (N_9961,N_9122,N_9374);
nand U9962 (N_9962,N_9463,N_9244);
xor U9963 (N_9963,N_9251,N_8979);
nand U9964 (N_9964,N_9464,N_9329);
and U9965 (N_9965,N_9530,N_9409);
nor U9966 (N_9966,N_9040,N_9238);
nand U9967 (N_9967,N_9487,N_8836);
nor U9968 (N_9968,N_9151,N_9193);
nand U9969 (N_9969,N_8997,N_9497);
nor U9970 (N_9970,N_9288,N_9564);
nand U9971 (N_9971,N_9403,N_9172);
or U9972 (N_9972,N_9536,N_9501);
nand U9973 (N_9973,N_9544,N_9574);
nor U9974 (N_9974,N_8854,N_8803);
and U9975 (N_9975,N_9131,N_9170);
xor U9976 (N_9976,N_9089,N_8882);
xor U9977 (N_9977,N_8873,N_9425);
nand U9978 (N_9978,N_9108,N_8824);
nor U9979 (N_9979,N_9447,N_9510);
nor U9980 (N_9980,N_8863,N_9326);
nand U9981 (N_9981,N_9207,N_8981);
nor U9982 (N_9982,N_9282,N_9187);
xnor U9983 (N_9983,N_9004,N_9504);
or U9984 (N_9984,N_9100,N_9297);
nor U9985 (N_9985,N_9048,N_9354);
xor U9986 (N_9986,N_8842,N_8922);
and U9987 (N_9987,N_9291,N_9526);
xnor U9988 (N_9988,N_9459,N_8987);
or U9989 (N_9989,N_9231,N_9052);
nand U9990 (N_9990,N_9163,N_9364);
nor U9991 (N_9991,N_9261,N_9561);
and U9992 (N_9992,N_9190,N_8866);
xor U9993 (N_9993,N_9043,N_9101);
nor U9994 (N_9994,N_8872,N_8830);
or U9995 (N_9995,N_8954,N_8810);
nand U9996 (N_9996,N_9441,N_9253);
nor U9997 (N_9997,N_8925,N_9216);
xnor U9998 (N_9998,N_9007,N_9072);
or U9999 (N_9999,N_9351,N_9161);
and U10000 (N_10000,N_9187,N_9019);
nor U10001 (N_10001,N_9360,N_9319);
xnor U10002 (N_10002,N_9109,N_9518);
xnor U10003 (N_10003,N_9256,N_9041);
and U10004 (N_10004,N_9206,N_8813);
xor U10005 (N_10005,N_9323,N_8948);
nor U10006 (N_10006,N_9486,N_8950);
and U10007 (N_10007,N_9127,N_9201);
and U10008 (N_10008,N_9577,N_9021);
nand U10009 (N_10009,N_9180,N_8816);
and U10010 (N_10010,N_9113,N_8922);
xnor U10011 (N_10011,N_9281,N_8866);
or U10012 (N_10012,N_9481,N_9446);
nand U10013 (N_10013,N_9411,N_9478);
nor U10014 (N_10014,N_9006,N_8960);
nand U10015 (N_10015,N_9560,N_8808);
nand U10016 (N_10016,N_9355,N_9523);
xnor U10017 (N_10017,N_9354,N_8854);
or U10018 (N_10018,N_9380,N_9445);
nand U10019 (N_10019,N_8945,N_8967);
or U10020 (N_10020,N_9015,N_9448);
xnor U10021 (N_10021,N_9106,N_9166);
and U10022 (N_10022,N_9397,N_9542);
nand U10023 (N_10023,N_9491,N_9569);
and U10024 (N_10024,N_9426,N_8912);
and U10025 (N_10025,N_9230,N_9348);
xor U10026 (N_10026,N_9093,N_9134);
xnor U10027 (N_10027,N_9048,N_9138);
and U10028 (N_10028,N_9581,N_9382);
nor U10029 (N_10029,N_9033,N_8854);
nand U10030 (N_10030,N_9371,N_9357);
nor U10031 (N_10031,N_9588,N_8934);
or U10032 (N_10032,N_9467,N_9481);
nand U10033 (N_10033,N_9111,N_9298);
nand U10034 (N_10034,N_9064,N_8853);
xor U10035 (N_10035,N_8802,N_9521);
nand U10036 (N_10036,N_9519,N_9296);
or U10037 (N_10037,N_9310,N_9489);
nand U10038 (N_10038,N_9377,N_8965);
and U10039 (N_10039,N_8921,N_8962);
nor U10040 (N_10040,N_9144,N_9041);
or U10041 (N_10041,N_9487,N_9216);
and U10042 (N_10042,N_9545,N_9420);
and U10043 (N_10043,N_9555,N_9584);
or U10044 (N_10044,N_9294,N_9115);
nand U10045 (N_10045,N_9298,N_9537);
nor U10046 (N_10046,N_9433,N_9361);
nor U10047 (N_10047,N_8808,N_8801);
or U10048 (N_10048,N_9060,N_8958);
nor U10049 (N_10049,N_9486,N_9577);
nor U10050 (N_10050,N_8914,N_9295);
nand U10051 (N_10051,N_9529,N_8970);
nand U10052 (N_10052,N_8992,N_8895);
xor U10053 (N_10053,N_9131,N_9453);
or U10054 (N_10054,N_9539,N_9301);
nor U10055 (N_10055,N_8864,N_8877);
nor U10056 (N_10056,N_9595,N_9179);
nor U10057 (N_10057,N_8950,N_8998);
or U10058 (N_10058,N_8847,N_9578);
or U10059 (N_10059,N_9212,N_8915);
nor U10060 (N_10060,N_8849,N_9410);
nor U10061 (N_10061,N_9096,N_8888);
or U10062 (N_10062,N_8958,N_9332);
nor U10063 (N_10063,N_9492,N_9324);
or U10064 (N_10064,N_9434,N_9489);
xor U10065 (N_10065,N_8971,N_9463);
and U10066 (N_10066,N_9006,N_9482);
xnor U10067 (N_10067,N_8945,N_9449);
nor U10068 (N_10068,N_9356,N_9554);
xor U10069 (N_10069,N_9086,N_9065);
or U10070 (N_10070,N_9052,N_9024);
nor U10071 (N_10071,N_9461,N_9144);
nor U10072 (N_10072,N_9435,N_9167);
nand U10073 (N_10073,N_8852,N_9258);
or U10074 (N_10074,N_9571,N_9005);
and U10075 (N_10075,N_9348,N_9362);
nor U10076 (N_10076,N_8915,N_9084);
nand U10077 (N_10077,N_9286,N_9358);
nor U10078 (N_10078,N_8920,N_9211);
xnor U10079 (N_10079,N_8936,N_9164);
and U10080 (N_10080,N_9168,N_9217);
xor U10081 (N_10081,N_9283,N_9054);
nor U10082 (N_10082,N_9429,N_9294);
or U10083 (N_10083,N_9391,N_8907);
nand U10084 (N_10084,N_9423,N_8874);
xor U10085 (N_10085,N_9345,N_9036);
or U10086 (N_10086,N_9070,N_9205);
xor U10087 (N_10087,N_9589,N_9010);
and U10088 (N_10088,N_9200,N_9546);
nand U10089 (N_10089,N_9192,N_8889);
or U10090 (N_10090,N_8891,N_9473);
nor U10091 (N_10091,N_9356,N_9544);
xor U10092 (N_10092,N_9478,N_8805);
nand U10093 (N_10093,N_9281,N_9159);
xnor U10094 (N_10094,N_9016,N_9236);
nor U10095 (N_10095,N_9012,N_8873);
or U10096 (N_10096,N_8820,N_9132);
nand U10097 (N_10097,N_9008,N_9439);
nor U10098 (N_10098,N_9308,N_9001);
or U10099 (N_10099,N_9407,N_9189);
xnor U10100 (N_10100,N_8801,N_9547);
nor U10101 (N_10101,N_8954,N_9325);
nand U10102 (N_10102,N_9414,N_9470);
or U10103 (N_10103,N_8800,N_9238);
and U10104 (N_10104,N_9457,N_8895);
nor U10105 (N_10105,N_8848,N_8847);
xnor U10106 (N_10106,N_9320,N_9231);
and U10107 (N_10107,N_9121,N_9257);
and U10108 (N_10108,N_8913,N_9301);
or U10109 (N_10109,N_9578,N_8935);
and U10110 (N_10110,N_8879,N_9365);
nor U10111 (N_10111,N_9096,N_9068);
or U10112 (N_10112,N_9297,N_8818);
nor U10113 (N_10113,N_8958,N_9246);
nor U10114 (N_10114,N_9138,N_9198);
xor U10115 (N_10115,N_9441,N_9169);
nand U10116 (N_10116,N_9038,N_9386);
nor U10117 (N_10117,N_9233,N_9457);
nand U10118 (N_10118,N_9423,N_9232);
nor U10119 (N_10119,N_8828,N_9154);
xnor U10120 (N_10120,N_9229,N_9441);
xor U10121 (N_10121,N_8872,N_8996);
nor U10122 (N_10122,N_8812,N_9385);
nand U10123 (N_10123,N_9280,N_8912);
xnor U10124 (N_10124,N_9473,N_9370);
nand U10125 (N_10125,N_9546,N_8992);
or U10126 (N_10126,N_8965,N_9057);
and U10127 (N_10127,N_8832,N_8929);
and U10128 (N_10128,N_8846,N_9273);
xor U10129 (N_10129,N_9332,N_9433);
and U10130 (N_10130,N_8808,N_9388);
nand U10131 (N_10131,N_9442,N_8859);
nand U10132 (N_10132,N_9102,N_9524);
and U10133 (N_10133,N_9525,N_9307);
nand U10134 (N_10134,N_8937,N_9276);
or U10135 (N_10135,N_8845,N_9028);
nand U10136 (N_10136,N_9034,N_9018);
and U10137 (N_10137,N_9126,N_9031);
nand U10138 (N_10138,N_8822,N_9315);
nor U10139 (N_10139,N_8927,N_9127);
nor U10140 (N_10140,N_9422,N_9463);
nor U10141 (N_10141,N_9399,N_9002);
or U10142 (N_10142,N_9301,N_9556);
and U10143 (N_10143,N_9131,N_8930);
nor U10144 (N_10144,N_9532,N_9035);
nand U10145 (N_10145,N_8871,N_9591);
or U10146 (N_10146,N_9330,N_9567);
and U10147 (N_10147,N_9418,N_9332);
nor U10148 (N_10148,N_9422,N_8931);
and U10149 (N_10149,N_9056,N_9515);
xor U10150 (N_10150,N_9136,N_8972);
nor U10151 (N_10151,N_8947,N_9291);
xor U10152 (N_10152,N_8873,N_9398);
and U10153 (N_10153,N_8875,N_9483);
xnor U10154 (N_10154,N_9395,N_9518);
nand U10155 (N_10155,N_9253,N_9384);
or U10156 (N_10156,N_9384,N_9226);
and U10157 (N_10157,N_8995,N_9561);
xor U10158 (N_10158,N_9252,N_9059);
nand U10159 (N_10159,N_8815,N_9325);
and U10160 (N_10160,N_8840,N_8917);
xnor U10161 (N_10161,N_9210,N_9487);
nor U10162 (N_10162,N_9515,N_9554);
xor U10163 (N_10163,N_9327,N_9551);
or U10164 (N_10164,N_9451,N_8946);
and U10165 (N_10165,N_9548,N_9572);
nor U10166 (N_10166,N_9560,N_8974);
nor U10167 (N_10167,N_9390,N_9207);
and U10168 (N_10168,N_9036,N_9534);
xnor U10169 (N_10169,N_9084,N_9539);
or U10170 (N_10170,N_9452,N_9423);
xor U10171 (N_10171,N_8850,N_9184);
and U10172 (N_10172,N_9064,N_9364);
nand U10173 (N_10173,N_9574,N_9298);
and U10174 (N_10174,N_8946,N_9566);
xor U10175 (N_10175,N_9586,N_9048);
nand U10176 (N_10176,N_9497,N_8946);
and U10177 (N_10177,N_8925,N_9083);
and U10178 (N_10178,N_9578,N_9161);
or U10179 (N_10179,N_9133,N_8904);
xnor U10180 (N_10180,N_9292,N_9341);
or U10181 (N_10181,N_9114,N_8957);
nand U10182 (N_10182,N_8962,N_8907);
nor U10183 (N_10183,N_9129,N_9393);
and U10184 (N_10184,N_8901,N_9180);
and U10185 (N_10185,N_9538,N_9205);
or U10186 (N_10186,N_9206,N_9046);
nand U10187 (N_10187,N_9007,N_9298);
nand U10188 (N_10188,N_9057,N_9270);
nand U10189 (N_10189,N_8919,N_9113);
nor U10190 (N_10190,N_9580,N_9014);
nor U10191 (N_10191,N_8881,N_8822);
xnor U10192 (N_10192,N_9124,N_9023);
or U10193 (N_10193,N_9011,N_9003);
and U10194 (N_10194,N_8942,N_9196);
xnor U10195 (N_10195,N_9144,N_9540);
or U10196 (N_10196,N_9342,N_8841);
and U10197 (N_10197,N_8880,N_8997);
xnor U10198 (N_10198,N_9234,N_9189);
and U10199 (N_10199,N_9391,N_9305);
nand U10200 (N_10200,N_9234,N_9084);
xnor U10201 (N_10201,N_9294,N_9235);
or U10202 (N_10202,N_8859,N_9026);
and U10203 (N_10203,N_9179,N_8924);
and U10204 (N_10204,N_9016,N_8834);
nand U10205 (N_10205,N_9224,N_8816);
or U10206 (N_10206,N_9386,N_9140);
nand U10207 (N_10207,N_8882,N_9066);
and U10208 (N_10208,N_9422,N_9228);
and U10209 (N_10209,N_9437,N_9271);
nand U10210 (N_10210,N_9219,N_9359);
nand U10211 (N_10211,N_9024,N_9090);
nor U10212 (N_10212,N_9115,N_8900);
or U10213 (N_10213,N_9304,N_9325);
or U10214 (N_10214,N_9179,N_8956);
xor U10215 (N_10215,N_9182,N_9330);
and U10216 (N_10216,N_9572,N_9508);
nor U10217 (N_10217,N_9117,N_8938);
or U10218 (N_10218,N_9341,N_9515);
and U10219 (N_10219,N_9040,N_9120);
xnor U10220 (N_10220,N_8804,N_8808);
xor U10221 (N_10221,N_8856,N_8945);
or U10222 (N_10222,N_8800,N_9043);
and U10223 (N_10223,N_8811,N_9503);
nand U10224 (N_10224,N_9467,N_9410);
xnor U10225 (N_10225,N_8920,N_9038);
nor U10226 (N_10226,N_8902,N_9122);
or U10227 (N_10227,N_9259,N_9090);
or U10228 (N_10228,N_8990,N_9578);
or U10229 (N_10229,N_8978,N_9330);
and U10230 (N_10230,N_8842,N_9138);
xor U10231 (N_10231,N_9293,N_8914);
nor U10232 (N_10232,N_9454,N_9599);
nor U10233 (N_10233,N_9275,N_9190);
or U10234 (N_10234,N_9372,N_9341);
nand U10235 (N_10235,N_9449,N_9336);
nor U10236 (N_10236,N_8823,N_8931);
nor U10237 (N_10237,N_9012,N_9153);
nand U10238 (N_10238,N_9050,N_9339);
xnor U10239 (N_10239,N_9045,N_9589);
xor U10240 (N_10240,N_8805,N_8883);
or U10241 (N_10241,N_9441,N_9092);
or U10242 (N_10242,N_9204,N_9042);
or U10243 (N_10243,N_9317,N_9593);
nand U10244 (N_10244,N_9316,N_9066);
and U10245 (N_10245,N_9101,N_9077);
or U10246 (N_10246,N_9169,N_9211);
or U10247 (N_10247,N_8853,N_9148);
and U10248 (N_10248,N_8931,N_9376);
nand U10249 (N_10249,N_9490,N_8845);
xor U10250 (N_10250,N_9274,N_9532);
nand U10251 (N_10251,N_9463,N_9065);
nand U10252 (N_10252,N_8887,N_8897);
nor U10253 (N_10253,N_9057,N_8894);
xor U10254 (N_10254,N_8810,N_8997);
or U10255 (N_10255,N_9306,N_9213);
xor U10256 (N_10256,N_8923,N_9528);
xnor U10257 (N_10257,N_9374,N_9483);
and U10258 (N_10258,N_9554,N_9120);
xnor U10259 (N_10259,N_8814,N_9270);
nand U10260 (N_10260,N_9129,N_9394);
xnor U10261 (N_10261,N_8998,N_8914);
nand U10262 (N_10262,N_9561,N_9207);
or U10263 (N_10263,N_8882,N_9341);
or U10264 (N_10264,N_9423,N_8894);
and U10265 (N_10265,N_9098,N_9512);
and U10266 (N_10266,N_9086,N_9208);
or U10267 (N_10267,N_8938,N_9036);
nor U10268 (N_10268,N_9564,N_9186);
or U10269 (N_10269,N_9165,N_8831);
or U10270 (N_10270,N_9195,N_9307);
nor U10271 (N_10271,N_9511,N_9582);
and U10272 (N_10272,N_9596,N_9436);
or U10273 (N_10273,N_9210,N_9021);
or U10274 (N_10274,N_9534,N_8805);
xor U10275 (N_10275,N_9327,N_9421);
nor U10276 (N_10276,N_9330,N_8996);
xor U10277 (N_10277,N_9367,N_9027);
nor U10278 (N_10278,N_8951,N_9525);
nand U10279 (N_10279,N_9037,N_9407);
and U10280 (N_10280,N_9420,N_9366);
xnor U10281 (N_10281,N_9247,N_8932);
nor U10282 (N_10282,N_9310,N_9294);
or U10283 (N_10283,N_9141,N_9429);
nor U10284 (N_10284,N_9191,N_9092);
nand U10285 (N_10285,N_9402,N_9520);
nand U10286 (N_10286,N_9088,N_8809);
and U10287 (N_10287,N_8881,N_9013);
nor U10288 (N_10288,N_9427,N_9251);
xor U10289 (N_10289,N_9233,N_9308);
nand U10290 (N_10290,N_9089,N_9353);
or U10291 (N_10291,N_8881,N_8925);
or U10292 (N_10292,N_9505,N_8984);
and U10293 (N_10293,N_9203,N_9530);
xnor U10294 (N_10294,N_9499,N_9424);
xnor U10295 (N_10295,N_8845,N_9361);
or U10296 (N_10296,N_8984,N_9581);
nand U10297 (N_10297,N_9228,N_8837);
nand U10298 (N_10298,N_8848,N_9240);
nor U10299 (N_10299,N_8843,N_9126);
and U10300 (N_10300,N_9111,N_9183);
and U10301 (N_10301,N_9473,N_9049);
nor U10302 (N_10302,N_8853,N_9035);
and U10303 (N_10303,N_9599,N_8979);
nor U10304 (N_10304,N_9380,N_8996);
xor U10305 (N_10305,N_9072,N_9205);
or U10306 (N_10306,N_9450,N_8813);
nor U10307 (N_10307,N_9256,N_9225);
xor U10308 (N_10308,N_9360,N_9329);
xor U10309 (N_10309,N_9527,N_8900);
nand U10310 (N_10310,N_9312,N_9362);
or U10311 (N_10311,N_9223,N_9519);
and U10312 (N_10312,N_8801,N_9279);
nand U10313 (N_10313,N_9245,N_9422);
nor U10314 (N_10314,N_8965,N_9245);
and U10315 (N_10315,N_8918,N_9524);
nor U10316 (N_10316,N_8801,N_8965);
nor U10317 (N_10317,N_9439,N_9137);
xor U10318 (N_10318,N_9484,N_9128);
or U10319 (N_10319,N_9418,N_9486);
and U10320 (N_10320,N_9005,N_9457);
or U10321 (N_10321,N_9243,N_8883);
or U10322 (N_10322,N_9320,N_8990);
xor U10323 (N_10323,N_9251,N_9159);
or U10324 (N_10324,N_9038,N_9448);
xnor U10325 (N_10325,N_9328,N_8986);
nor U10326 (N_10326,N_9161,N_9589);
and U10327 (N_10327,N_9239,N_8954);
nor U10328 (N_10328,N_9145,N_8843);
nor U10329 (N_10329,N_8909,N_9406);
or U10330 (N_10330,N_9497,N_9439);
nand U10331 (N_10331,N_9018,N_9514);
or U10332 (N_10332,N_9594,N_9186);
and U10333 (N_10333,N_9378,N_9185);
and U10334 (N_10334,N_8906,N_9030);
nand U10335 (N_10335,N_9168,N_9112);
or U10336 (N_10336,N_9518,N_8856);
nand U10337 (N_10337,N_9011,N_9108);
xnor U10338 (N_10338,N_8978,N_9393);
or U10339 (N_10339,N_9579,N_8945);
and U10340 (N_10340,N_8854,N_8851);
and U10341 (N_10341,N_8833,N_8865);
nor U10342 (N_10342,N_9421,N_9514);
and U10343 (N_10343,N_9061,N_8978);
and U10344 (N_10344,N_9299,N_9184);
nor U10345 (N_10345,N_9423,N_9321);
or U10346 (N_10346,N_9051,N_9184);
xnor U10347 (N_10347,N_9405,N_9410);
nand U10348 (N_10348,N_8867,N_9187);
or U10349 (N_10349,N_8847,N_8882);
and U10350 (N_10350,N_8886,N_9022);
nor U10351 (N_10351,N_9292,N_9547);
nand U10352 (N_10352,N_8813,N_9417);
nor U10353 (N_10353,N_9141,N_9240);
nand U10354 (N_10354,N_9336,N_8931);
or U10355 (N_10355,N_9527,N_9057);
nand U10356 (N_10356,N_9186,N_9539);
and U10357 (N_10357,N_9574,N_9306);
or U10358 (N_10358,N_9010,N_8836);
xor U10359 (N_10359,N_8856,N_9139);
xnor U10360 (N_10360,N_9570,N_8800);
xor U10361 (N_10361,N_8965,N_9092);
or U10362 (N_10362,N_9197,N_8996);
or U10363 (N_10363,N_8973,N_9310);
or U10364 (N_10364,N_9157,N_9145);
and U10365 (N_10365,N_9315,N_9591);
nor U10366 (N_10366,N_8822,N_9422);
nand U10367 (N_10367,N_9561,N_9182);
and U10368 (N_10368,N_8950,N_9181);
and U10369 (N_10369,N_9214,N_9255);
and U10370 (N_10370,N_9489,N_9029);
or U10371 (N_10371,N_8845,N_9120);
xnor U10372 (N_10372,N_8877,N_9310);
nand U10373 (N_10373,N_9489,N_9283);
xnor U10374 (N_10374,N_9422,N_9117);
nand U10375 (N_10375,N_9199,N_8808);
and U10376 (N_10376,N_9555,N_9553);
and U10377 (N_10377,N_8928,N_9434);
and U10378 (N_10378,N_9102,N_9021);
nand U10379 (N_10379,N_9531,N_9182);
and U10380 (N_10380,N_9314,N_9192);
and U10381 (N_10381,N_8897,N_9500);
nor U10382 (N_10382,N_9311,N_9397);
xnor U10383 (N_10383,N_9268,N_9491);
xnor U10384 (N_10384,N_9262,N_8897);
or U10385 (N_10385,N_9307,N_9598);
nand U10386 (N_10386,N_9259,N_9214);
nor U10387 (N_10387,N_9518,N_9359);
or U10388 (N_10388,N_9232,N_9128);
and U10389 (N_10389,N_9192,N_9466);
or U10390 (N_10390,N_9488,N_9252);
nor U10391 (N_10391,N_9307,N_9260);
and U10392 (N_10392,N_8809,N_9248);
nor U10393 (N_10393,N_9302,N_8822);
nand U10394 (N_10394,N_9562,N_8904);
nor U10395 (N_10395,N_9506,N_9387);
or U10396 (N_10396,N_9076,N_8888);
nor U10397 (N_10397,N_9336,N_8958);
nor U10398 (N_10398,N_9326,N_9308);
and U10399 (N_10399,N_9279,N_9231);
nor U10400 (N_10400,N_9726,N_9844);
xor U10401 (N_10401,N_10061,N_9890);
and U10402 (N_10402,N_9697,N_10044);
and U10403 (N_10403,N_10183,N_9757);
and U10404 (N_10404,N_10031,N_10361);
xor U10405 (N_10405,N_9995,N_10166);
nor U10406 (N_10406,N_10220,N_10060);
and U10407 (N_10407,N_10265,N_9771);
or U10408 (N_10408,N_9603,N_9668);
or U10409 (N_10409,N_9893,N_10051);
nor U10410 (N_10410,N_10316,N_10058);
and U10411 (N_10411,N_10357,N_10034);
xnor U10412 (N_10412,N_9946,N_10287);
nand U10413 (N_10413,N_10279,N_10395);
nand U10414 (N_10414,N_9799,N_9795);
xnor U10415 (N_10415,N_9972,N_10340);
or U10416 (N_10416,N_10241,N_10134);
nand U10417 (N_10417,N_10016,N_10330);
and U10418 (N_10418,N_10144,N_10017);
nor U10419 (N_10419,N_10238,N_10207);
nand U10420 (N_10420,N_10264,N_10121);
or U10421 (N_10421,N_10151,N_9933);
nor U10422 (N_10422,N_10211,N_9666);
xor U10423 (N_10423,N_9631,N_10004);
and U10424 (N_10424,N_9876,N_9754);
xnor U10425 (N_10425,N_9822,N_9874);
nor U10426 (N_10426,N_9971,N_9883);
nor U10427 (N_10427,N_9963,N_9887);
and U10428 (N_10428,N_9645,N_10109);
nand U10429 (N_10429,N_9635,N_10026);
nand U10430 (N_10430,N_10071,N_9787);
nand U10431 (N_10431,N_10366,N_10378);
or U10432 (N_10432,N_10164,N_10067);
or U10433 (N_10433,N_9922,N_10070);
and U10434 (N_10434,N_9889,N_10393);
or U10435 (N_10435,N_9658,N_10075);
nor U10436 (N_10436,N_9780,N_9602);
nand U10437 (N_10437,N_10035,N_9770);
nand U10438 (N_10438,N_9669,N_9652);
or U10439 (N_10439,N_10065,N_10305);
or U10440 (N_10440,N_9953,N_10343);
xnor U10441 (N_10441,N_10028,N_9834);
xor U10442 (N_10442,N_10115,N_10310);
nand U10443 (N_10443,N_10322,N_10375);
or U10444 (N_10444,N_10222,N_9829);
nor U10445 (N_10445,N_9722,N_9760);
nor U10446 (N_10446,N_9994,N_10302);
xor U10447 (N_10447,N_9777,N_10005);
xnor U10448 (N_10448,N_10193,N_9847);
and U10449 (N_10449,N_9840,N_9960);
and U10450 (N_10450,N_9665,N_9688);
and U10451 (N_10451,N_9931,N_9858);
and U10452 (N_10452,N_10253,N_10087);
xor U10453 (N_10453,N_10092,N_9607);
xnor U10454 (N_10454,N_10176,N_9794);
nand U10455 (N_10455,N_10221,N_10122);
or U10456 (N_10456,N_10381,N_9713);
nand U10457 (N_10457,N_9888,N_10328);
and U10458 (N_10458,N_10125,N_9627);
xor U10459 (N_10459,N_9681,N_10081);
and U10460 (N_10460,N_9848,N_10289);
nand U10461 (N_10461,N_10332,N_10131);
and U10462 (N_10462,N_9618,N_9756);
xor U10463 (N_10463,N_10040,N_10311);
xnor U10464 (N_10464,N_9914,N_9800);
xnor U10465 (N_10465,N_10068,N_10059);
xnor U10466 (N_10466,N_10387,N_9601);
xor U10467 (N_10467,N_9701,N_9997);
xor U10468 (N_10468,N_10304,N_9685);
or U10469 (N_10469,N_9879,N_10203);
or U10470 (N_10470,N_9869,N_9814);
nor U10471 (N_10471,N_10111,N_10249);
xnor U10472 (N_10472,N_9942,N_10020);
nand U10473 (N_10473,N_9984,N_10064);
or U10474 (N_10474,N_10329,N_10209);
or U10475 (N_10475,N_9608,N_9789);
nor U10476 (N_10476,N_9740,N_10275);
xor U10477 (N_10477,N_10094,N_10186);
nand U10478 (N_10478,N_9943,N_9611);
nor U10479 (N_10479,N_10192,N_9988);
nand U10480 (N_10480,N_10072,N_10055);
xnor U10481 (N_10481,N_9657,N_10210);
nor U10482 (N_10482,N_9958,N_10032);
and U10483 (N_10483,N_10356,N_10339);
xor U10484 (N_10484,N_10139,N_10175);
or U10485 (N_10485,N_10224,N_10350);
xor U10486 (N_10486,N_10285,N_10128);
and U10487 (N_10487,N_9624,N_10376);
xor U10488 (N_10488,N_10011,N_10297);
and U10489 (N_10489,N_10205,N_9775);
nand U10490 (N_10490,N_10358,N_9612);
nand U10491 (N_10491,N_9664,N_9656);
and U10492 (N_10492,N_10147,N_9716);
or U10493 (N_10493,N_9815,N_10392);
xor U10494 (N_10494,N_9845,N_10283);
xor U10495 (N_10495,N_10202,N_9849);
nor U10496 (N_10496,N_10337,N_10286);
or U10497 (N_10497,N_9980,N_9918);
or U10498 (N_10498,N_9955,N_9621);
xor U10499 (N_10499,N_10012,N_9764);
xor U10500 (N_10500,N_9965,N_9606);
nor U10501 (N_10501,N_9751,N_10114);
or U10502 (N_10502,N_9974,N_9680);
nor U10503 (N_10503,N_9916,N_10019);
or U10504 (N_10504,N_10138,N_9605);
and U10505 (N_10505,N_10078,N_10007);
nand U10506 (N_10506,N_10320,N_10113);
nor U10507 (N_10507,N_9709,N_9894);
nor U10508 (N_10508,N_9675,N_9674);
or U10509 (N_10509,N_10132,N_10288);
or U10510 (N_10510,N_10083,N_9630);
nor U10511 (N_10511,N_10149,N_9617);
nor U10512 (N_10512,N_10097,N_9850);
nor U10513 (N_10513,N_10386,N_9644);
xor U10514 (N_10514,N_9626,N_10326);
and U10515 (N_10515,N_10015,N_9620);
and U10516 (N_10516,N_9982,N_10243);
nor U10517 (N_10517,N_10152,N_9654);
xor U10518 (N_10518,N_9998,N_9604);
xor U10519 (N_10519,N_9826,N_9673);
nor U10520 (N_10520,N_10272,N_10277);
xor U10521 (N_10521,N_9801,N_10187);
xor U10522 (N_10522,N_10232,N_10331);
nor U10523 (N_10523,N_9791,N_9905);
xnor U10524 (N_10524,N_9853,N_10008);
nor U10525 (N_10525,N_9941,N_10291);
xor U10526 (N_10526,N_9719,N_9952);
nand U10527 (N_10527,N_10391,N_10295);
nand U10528 (N_10528,N_10140,N_10276);
or U10529 (N_10529,N_9843,N_9745);
nor U10530 (N_10530,N_10353,N_9919);
nor U10531 (N_10531,N_10030,N_9839);
nand U10532 (N_10532,N_10240,N_9903);
or U10533 (N_10533,N_10333,N_9846);
or U10534 (N_10534,N_9975,N_10174);
nand U10535 (N_10535,N_10117,N_10052);
and U10536 (N_10536,N_9891,N_10023);
and U10537 (N_10537,N_9742,N_9906);
xnor U10538 (N_10538,N_10244,N_9950);
and U10539 (N_10539,N_9809,N_10258);
nor U10540 (N_10540,N_9802,N_10315);
nand U10541 (N_10541,N_10143,N_9643);
xnor U10542 (N_10542,N_9937,N_9727);
and U10543 (N_10543,N_10398,N_10270);
or U10544 (N_10544,N_9730,N_10198);
or U10545 (N_10545,N_10274,N_9655);
nor U10546 (N_10546,N_10158,N_10190);
or U10547 (N_10547,N_9686,N_10348);
xnor U10548 (N_10548,N_9856,N_10206);
xor U10549 (N_10549,N_9939,N_9900);
nand U10550 (N_10550,N_9739,N_9703);
nand U10551 (N_10551,N_9786,N_9798);
or U10552 (N_10552,N_9706,N_10233);
nor U10553 (N_10553,N_9734,N_10397);
or U10554 (N_10554,N_9712,N_9661);
nand U10555 (N_10555,N_9699,N_10370);
or U10556 (N_10556,N_10043,N_10334);
xnor U10557 (N_10557,N_10062,N_9841);
nor U10558 (N_10558,N_10084,N_9671);
or U10559 (N_10559,N_9738,N_9784);
xor U10560 (N_10560,N_9792,N_10146);
xor U10561 (N_10561,N_10009,N_10273);
or U10562 (N_10562,N_10119,N_9825);
or U10563 (N_10563,N_10167,N_10185);
nor U10564 (N_10564,N_9819,N_10150);
nor U10565 (N_10565,N_9733,N_10069);
xnor U10566 (N_10566,N_9614,N_10335);
or U10567 (N_10567,N_10089,N_10112);
xnor U10568 (N_10568,N_9763,N_10250);
nor U10569 (N_10569,N_9749,N_10318);
nor U10570 (N_10570,N_10215,N_10262);
xor U10571 (N_10571,N_9913,N_10372);
nand U10572 (N_10572,N_9736,N_9684);
nor U10573 (N_10573,N_9930,N_9855);
xnor U10574 (N_10574,N_10216,N_10110);
nor U10575 (N_10575,N_10255,N_10229);
nor U10576 (N_10576,N_9877,N_10266);
and U10577 (N_10577,N_10252,N_10338);
nor U10578 (N_10578,N_9857,N_10045);
and U10579 (N_10579,N_10362,N_10168);
nor U10580 (N_10580,N_9993,N_10312);
nand U10581 (N_10581,N_9642,N_10047);
xor U10582 (N_10582,N_10126,N_9728);
and U10583 (N_10583,N_9715,N_9670);
and U10584 (N_10584,N_9693,N_9724);
xor U10585 (N_10585,N_9947,N_10292);
and U10586 (N_10586,N_10018,N_10300);
or U10587 (N_10587,N_9964,N_9723);
and U10588 (N_10588,N_10095,N_9662);
or U10589 (N_10589,N_9638,N_9619);
or U10590 (N_10590,N_10345,N_10050);
or U10591 (N_10591,N_9774,N_9705);
or U10592 (N_10592,N_9827,N_10321);
and U10593 (N_10593,N_9884,N_9861);
nor U10594 (N_10594,N_9732,N_10135);
xor U10595 (N_10595,N_9651,N_9954);
nor U10596 (N_10596,N_9695,N_9737);
nand U10597 (N_10597,N_9636,N_10161);
nor U10598 (N_10598,N_10317,N_9910);
and U10599 (N_10599,N_9842,N_10389);
and U10600 (N_10600,N_9779,N_10169);
nor U10601 (N_10601,N_9629,N_10002);
nand U10602 (N_10602,N_10296,N_9793);
or U10603 (N_10603,N_10054,N_9925);
xor U10604 (N_10604,N_9623,N_10208);
nor U10605 (N_10605,N_9875,N_10088);
or U10606 (N_10606,N_9710,N_9927);
and U10607 (N_10607,N_10063,N_9783);
xnor U10608 (N_10608,N_9961,N_9862);
and U10609 (N_10609,N_9899,N_10256);
nor U10610 (N_10610,N_10336,N_9907);
or U10611 (N_10611,N_10120,N_10194);
nor U10612 (N_10612,N_10271,N_9871);
or U10613 (N_10613,N_10245,N_10165);
xor U10614 (N_10614,N_9672,N_10171);
nor U10615 (N_10615,N_9731,N_9909);
xnor U10616 (N_10616,N_10073,N_9648);
and U10617 (N_10617,N_10025,N_9812);
xor U10618 (N_10618,N_9968,N_10036);
nor U10619 (N_10619,N_9824,N_10246);
and U10620 (N_10620,N_9864,N_10077);
nor U10621 (N_10621,N_10363,N_10079);
xor U10622 (N_10622,N_10013,N_9897);
and U10623 (N_10623,N_9985,N_10090);
nor U10624 (N_10624,N_9790,N_10239);
or U10625 (N_10625,N_9837,N_10298);
xor U10626 (N_10626,N_9667,N_9967);
and U10627 (N_10627,N_9639,N_10057);
xor U10628 (N_10628,N_10319,N_9957);
or U10629 (N_10629,N_9772,N_10041);
or U10630 (N_10630,N_9797,N_9711);
xnor U10631 (N_10631,N_9778,N_10260);
or U10632 (N_10632,N_10267,N_10293);
xor U10633 (N_10633,N_9996,N_10153);
nor U10634 (N_10634,N_9677,N_9687);
nand U10635 (N_10635,N_9935,N_9981);
xor U10636 (N_10636,N_9870,N_10136);
xor U10637 (N_10637,N_10006,N_10268);
nor U10638 (N_10638,N_9649,N_9908);
nand U10639 (N_10639,N_10309,N_10029);
nand U10640 (N_10640,N_10248,N_10306);
nor U10641 (N_10641,N_10308,N_9989);
nand U10642 (N_10642,N_10213,N_9915);
or U10643 (N_10643,N_9718,N_10099);
nand U10644 (N_10644,N_9748,N_9944);
and U10645 (N_10645,N_9729,N_10235);
or U10646 (N_10646,N_10226,N_10066);
and U10647 (N_10647,N_10261,N_9945);
and U10648 (N_10648,N_10145,N_9702);
or U10649 (N_10649,N_9881,N_9938);
or U10650 (N_10650,N_10301,N_10385);
nand U10651 (N_10651,N_10303,N_10038);
and U10652 (N_10652,N_10352,N_10214);
xor U10653 (N_10653,N_9896,N_10281);
and U10654 (N_10654,N_9708,N_10101);
or U10655 (N_10655,N_10076,N_9924);
and U10656 (N_10656,N_10242,N_10096);
and U10657 (N_10657,N_9676,N_9951);
or U10658 (N_10658,N_9832,N_9948);
nand U10659 (N_10659,N_9867,N_10182);
and U10660 (N_10660,N_10173,N_9753);
and U10661 (N_10661,N_9836,N_10074);
nor U10662 (N_10662,N_9929,N_9868);
nand U10663 (N_10663,N_9973,N_9911);
nand U10664 (N_10664,N_9926,N_10347);
and U10665 (N_10665,N_9650,N_9970);
xor U10666 (N_10666,N_9634,N_10129);
nor U10667 (N_10667,N_9610,N_9936);
nand U10668 (N_10668,N_9878,N_9901);
nor U10669 (N_10669,N_10103,N_9892);
and U10670 (N_10670,N_10373,N_9885);
xor U10671 (N_10671,N_10197,N_10124);
xnor U10672 (N_10672,N_9762,N_10325);
or U10673 (N_10673,N_10284,N_9803);
or U10674 (N_10674,N_9692,N_10098);
and U10675 (N_10675,N_10037,N_10227);
nor U10676 (N_10676,N_10195,N_10091);
or U10677 (N_10677,N_10369,N_10360);
nand U10678 (N_10678,N_9743,N_9761);
xor U10679 (N_10679,N_10162,N_10106);
or U10680 (N_10680,N_10278,N_10177);
nand U10681 (N_10681,N_9808,N_9851);
nand U10682 (N_10682,N_10027,N_9758);
and U10683 (N_10683,N_10141,N_9863);
nor U10684 (N_10684,N_10048,N_10382);
and U10685 (N_10685,N_9859,N_9766);
or U10686 (N_10686,N_10156,N_10307);
nand U10687 (N_10687,N_9720,N_10003);
or U10688 (N_10688,N_9741,N_10104);
and U10689 (N_10689,N_10394,N_10396);
nor U10690 (N_10690,N_9902,N_9852);
xor U10691 (N_10691,N_10217,N_9904);
xor U10692 (N_10692,N_10148,N_9959);
nor U10693 (N_10693,N_9796,N_10200);
nand U10694 (N_10694,N_9752,N_9746);
nand U10695 (N_10695,N_10223,N_10269);
or U10696 (N_10696,N_9805,N_9725);
and U10697 (N_10697,N_10383,N_10123);
nor U10698 (N_10698,N_9917,N_9804);
nand U10699 (N_10699,N_10105,N_9707);
nand U10700 (N_10700,N_9700,N_10102);
nand U10701 (N_10701,N_9785,N_9759);
xor U10702 (N_10702,N_9691,N_10093);
and U10703 (N_10703,N_10364,N_9714);
or U10704 (N_10704,N_9912,N_10001);
or U10705 (N_10705,N_10251,N_10323);
or U10706 (N_10706,N_10201,N_9632);
xnor U10707 (N_10707,N_10294,N_9781);
xor U10708 (N_10708,N_9653,N_9646);
xnor U10709 (N_10709,N_9637,N_10230);
and U10710 (N_10710,N_10263,N_10024);
xnor U10711 (N_10711,N_9765,N_9979);
and U10712 (N_10712,N_10231,N_10184);
or U10713 (N_10713,N_9949,N_9788);
nand U10714 (N_10714,N_10170,N_9811);
xnor U10715 (N_10715,N_10142,N_9696);
and U10716 (N_10716,N_9818,N_10181);
nand U10717 (N_10717,N_10033,N_9895);
or U10718 (N_10718,N_9923,N_10355);
xnor U10719 (N_10719,N_10313,N_10327);
xor U10720 (N_10720,N_9622,N_9721);
nand U10721 (N_10721,N_9983,N_9640);
nand U10722 (N_10722,N_10046,N_10080);
xnor U10723 (N_10723,N_9999,N_10049);
and U10724 (N_10724,N_9747,N_10344);
or U10725 (N_10725,N_9616,N_10172);
nand U10726 (N_10726,N_9921,N_10179);
nand U10727 (N_10727,N_9704,N_10365);
nor U10728 (N_10728,N_9625,N_10259);
nand U10729 (N_10729,N_9820,N_10154);
nand U10730 (N_10730,N_9821,N_9698);
or U10731 (N_10731,N_10237,N_9609);
or U10732 (N_10732,N_10022,N_9830);
and U10733 (N_10733,N_9633,N_10159);
nor U10734 (N_10734,N_10053,N_10218);
xor U10735 (N_10735,N_10042,N_9831);
and U10736 (N_10736,N_9735,N_9860);
xor U10737 (N_10737,N_9962,N_10351);
nor U10738 (N_10738,N_10368,N_10257);
or U10739 (N_10739,N_10133,N_9928);
and U10740 (N_10740,N_10086,N_10204);
and U10741 (N_10741,N_9613,N_9810);
nor U10742 (N_10742,N_10130,N_9689);
nor U10743 (N_10743,N_10010,N_10082);
and U10744 (N_10744,N_10349,N_10212);
xnor U10745 (N_10745,N_10299,N_9806);
or U10746 (N_10746,N_10388,N_9750);
or U10747 (N_10747,N_10228,N_10390);
nor U10748 (N_10748,N_10236,N_10155);
or U10749 (N_10749,N_10191,N_9882);
xnor U10750 (N_10750,N_9717,N_9978);
nand U10751 (N_10751,N_9682,N_9773);
xor U10752 (N_10752,N_9854,N_10346);
and U10753 (N_10753,N_10280,N_10225);
and U10754 (N_10754,N_10085,N_10371);
xor U10755 (N_10755,N_9986,N_9873);
nand U10756 (N_10756,N_9615,N_10107);
and U10757 (N_10757,N_10374,N_9828);
and U10758 (N_10758,N_9966,N_10189);
nand U10759 (N_10759,N_10157,N_10160);
nor U10760 (N_10760,N_9823,N_10354);
and U10761 (N_10761,N_9990,N_9659);
xor U10762 (N_10762,N_10359,N_10116);
nand U10763 (N_10763,N_9683,N_9641);
nor U10764 (N_10764,N_10247,N_10056);
nor U10765 (N_10765,N_9865,N_9898);
nor U10766 (N_10766,N_9663,N_9768);
and U10767 (N_10767,N_10163,N_10367);
xnor U10768 (N_10768,N_10282,N_9647);
nor U10769 (N_10769,N_10254,N_9880);
xnor U10770 (N_10770,N_10290,N_9690);
and U10771 (N_10771,N_10380,N_9987);
or U10772 (N_10772,N_9694,N_9934);
xnor U10773 (N_10773,N_10324,N_9816);
or U10774 (N_10774,N_9817,N_9782);
or U10775 (N_10775,N_9660,N_10384);
xor U10776 (N_10776,N_9769,N_9833);
nor U10777 (N_10777,N_9992,N_10342);
or U10778 (N_10778,N_10234,N_10108);
or U10779 (N_10779,N_9969,N_9866);
nor U10780 (N_10780,N_9976,N_10180);
nor U10781 (N_10781,N_9835,N_10377);
or U10782 (N_10782,N_10021,N_10100);
xor U10783 (N_10783,N_9600,N_9744);
xor U10784 (N_10784,N_9886,N_10127);
xnor U10785 (N_10785,N_10314,N_10137);
and U10786 (N_10786,N_9678,N_10014);
and U10787 (N_10787,N_10399,N_9872);
and U10788 (N_10788,N_10219,N_10196);
and U10789 (N_10789,N_9838,N_9755);
xnor U10790 (N_10790,N_9813,N_9807);
nor U10791 (N_10791,N_10039,N_9991);
xnor U10792 (N_10792,N_10188,N_10199);
or U10793 (N_10793,N_10118,N_9679);
nand U10794 (N_10794,N_10341,N_9776);
nor U10795 (N_10795,N_10379,N_9767);
nor U10796 (N_10796,N_10000,N_9977);
nand U10797 (N_10797,N_9628,N_9940);
nor U10798 (N_10798,N_9920,N_9932);
or U10799 (N_10799,N_10178,N_9956);
and U10800 (N_10800,N_9649,N_9928);
nor U10801 (N_10801,N_9613,N_9886);
or U10802 (N_10802,N_10271,N_10096);
nor U10803 (N_10803,N_10009,N_9865);
or U10804 (N_10804,N_9715,N_10246);
nand U10805 (N_10805,N_10093,N_10199);
or U10806 (N_10806,N_10090,N_10159);
nand U10807 (N_10807,N_9808,N_10327);
nand U10808 (N_10808,N_10068,N_10170);
xor U10809 (N_10809,N_9866,N_10001);
and U10810 (N_10810,N_9822,N_10028);
and U10811 (N_10811,N_9694,N_10010);
and U10812 (N_10812,N_10135,N_10386);
xnor U10813 (N_10813,N_9961,N_9754);
xnor U10814 (N_10814,N_9609,N_10175);
xor U10815 (N_10815,N_9769,N_9805);
nor U10816 (N_10816,N_10251,N_9887);
nor U10817 (N_10817,N_9941,N_9998);
and U10818 (N_10818,N_10334,N_9621);
xnor U10819 (N_10819,N_9749,N_9867);
or U10820 (N_10820,N_9744,N_10072);
or U10821 (N_10821,N_10101,N_9748);
or U10822 (N_10822,N_10076,N_9850);
and U10823 (N_10823,N_9988,N_10352);
nor U10824 (N_10824,N_9838,N_9742);
nor U10825 (N_10825,N_10093,N_10261);
and U10826 (N_10826,N_10124,N_10234);
xor U10827 (N_10827,N_10004,N_10276);
xnor U10828 (N_10828,N_10201,N_9841);
and U10829 (N_10829,N_10268,N_9943);
nor U10830 (N_10830,N_9818,N_9819);
nor U10831 (N_10831,N_10000,N_9718);
xor U10832 (N_10832,N_9884,N_9978);
or U10833 (N_10833,N_10275,N_9720);
xnor U10834 (N_10834,N_9890,N_10119);
nor U10835 (N_10835,N_10074,N_9796);
nand U10836 (N_10836,N_10133,N_10191);
xor U10837 (N_10837,N_9829,N_9605);
xor U10838 (N_10838,N_9656,N_9787);
nor U10839 (N_10839,N_9614,N_9782);
xor U10840 (N_10840,N_10394,N_9904);
nand U10841 (N_10841,N_9690,N_10144);
xor U10842 (N_10842,N_9880,N_9954);
nand U10843 (N_10843,N_9696,N_10078);
nor U10844 (N_10844,N_9618,N_10121);
xnor U10845 (N_10845,N_10146,N_10307);
nand U10846 (N_10846,N_9871,N_9659);
nor U10847 (N_10847,N_10022,N_10375);
or U10848 (N_10848,N_10034,N_9624);
nor U10849 (N_10849,N_10327,N_9681);
xnor U10850 (N_10850,N_9777,N_9657);
xnor U10851 (N_10851,N_10017,N_9899);
xor U10852 (N_10852,N_9802,N_9764);
nand U10853 (N_10853,N_10287,N_10168);
nor U10854 (N_10854,N_10268,N_9909);
nand U10855 (N_10855,N_9951,N_9698);
nor U10856 (N_10856,N_10110,N_9808);
or U10857 (N_10857,N_10308,N_10214);
xor U10858 (N_10858,N_10015,N_9842);
nand U10859 (N_10859,N_9947,N_10002);
or U10860 (N_10860,N_9929,N_10248);
xor U10861 (N_10861,N_9630,N_10138);
and U10862 (N_10862,N_9850,N_10193);
or U10863 (N_10863,N_10087,N_9944);
and U10864 (N_10864,N_9935,N_10324);
nand U10865 (N_10865,N_9737,N_10025);
and U10866 (N_10866,N_10294,N_10265);
and U10867 (N_10867,N_9978,N_9800);
nand U10868 (N_10868,N_10168,N_10363);
nor U10869 (N_10869,N_9749,N_10217);
and U10870 (N_10870,N_10286,N_10398);
nor U10871 (N_10871,N_9941,N_10100);
and U10872 (N_10872,N_9701,N_9717);
nand U10873 (N_10873,N_9856,N_9653);
nor U10874 (N_10874,N_9641,N_9668);
and U10875 (N_10875,N_10264,N_9898);
nor U10876 (N_10876,N_10294,N_9696);
xor U10877 (N_10877,N_10307,N_9677);
and U10878 (N_10878,N_9779,N_10221);
or U10879 (N_10879,N_10240,N_10199);
and U10880 (N_10880,N_9752,N_10231);
nand U10881 (N_10881,N_9882,N_9701);
nand U10882 (N_10882,N_9606,N_9784);
nor U10883 (N_10883,N_10166,N_10151);
xnor U10884 (N_10884,N_9713,N_9936);
and U10885 (N_10885,N_10375,N_9925);
nand U10886 (N_10886,N_9918,N_10343);
and U10887 (N_10887,N_10051,N_10184);
xor U10888 (N_10888,N_10153,N_9986);
and U10889 (N_10889,N_10079,N_10156);
and U10890 (N_10890,N_10079,N_9825);
nor U10891 (N_10891,N_9664,N_9741);
xnor U10892 (N_10892,N_10156,N_9689);
and U10893 (N_10893,N_10205,N_10256);
nand U10894 (N_10894,N_9958,N_10354);
nor U10895 (N_10895,N_10291,N_9908);
and U10896 (N_10896,N_10264,N_9702);
nand U10897 (N_10897,N_9620,N_9617);
or U10898 (N_10898,N_9987,N_10387);
xor U10899 (N_10899,N_9705,N_9863);
nor U10900 (N_10900,N_9971,N_9814);
nor U10901 (N_10901,N_9723,N_10364);
or U10902 (N_10902,N_10372,N_9988);
and U10903 (N_10903,N_9687,N_10093);
and U10904 (N_10904,N_10251,N_10219);
nor U10905 (N_10905,N_10369,N_10103);
and U10906 (N_10906,N_9922,N_9755);
xor U10907 (N_10907,N_9621,N_10143);
nor U10908 (N_10908,N_9805,N_9798);
or U10909 (N_10909,N_9840,N_10351);
nor U10910 (N_10910,N_10092,N_10108);
xor U10911 (N_10911,N_10286,N_9722);
nand U10912 (N_10912,N_10168,N_9879);
and U10913 (N_10913,N_9932,N_9735);
nand U10914 (N_10914,N_10213,N_10010);
nor U10915 (N_10915,N_9958,N_10296);
or U10916 (N_10916,N_10195,N_9771);
nor U10917 (N_10917,N_9793,N_10259);
nand U10918 (N_10918,N_10227,N_10362);
and U10919 (N_10919,N_10190,N_10343);
nor U10920 (N_10920,N_9872,N_9769);
nor U10921 (N_10921,N_9898,N_9715);
or U10922 (N_10922,N_9616,N_9867);
or U10923 (N_10923,N_10318,N_9743);
or U10924 (N_10924,N_9669,N_9918);
nand U10925 (N_10925,N_10132,N_9901);
nor U10926 (N_10926,N_9684,N_10276);
nor U10927 (N_10927,N_9657,N_10039);
nand U10928 (N_10928,N_10172,N_10137);
and U10929 (N_10929,N_10395,N_10076);
nor U10930 (N_10930,N_9801,N_9815);
or U10931 (N_10931,N_9816,N_10210);
nor U10932 (N_10932,N_10343,N_10302);
nand U10933 (N_10933,N_9822,N_10256);
xor U10934 (N_10934,N_10230,N_10196);
nor U10935 (N_10935,N_9810,N_9666);
nand U10936 (N_10936,N_10386,N_9651);
nor U10937 (N_10937,N_10094,N_10056);
or U10938 (N_10938,N_10277,N_9946);
or U10939 (N_10939,N_9925,N_10267);
and U10940 (N_10940,N_10307,N_9856);
nor U10941 (N_10941,N_10138,N_10128);
xnor U10942 (N_10942,N_9688,N_10105);
nor U10943 (N_10943,N_9753,N_10200);
or U10944 (N_10944,N_9984,N_9665);
and U10945 (N_10945,N_9892,N_9925);
or U10946 (N_10946,N_10018,N_10060);
or U10947 (N_10947,N_10173,N_10067);
xnor U10948 (N_10948,N_10341,N_10313);
and U10949 (N_10949,N_9877,N_9923);
xnor U10950 (N_10950,N_10057,N_10381);
or U10951 (N_10951,N_10343,N_9790);
and U10952 (N_10952,N_9807,N_9769);
xnor U10953 (N_10953,N_9892,N_9641);
or U10954 (N_10954,N_10005,N_9738);
and U10955 (N_10955,N_9768,N_10010);
or U10956 (N_10956,N_10114,N_9804);
and U10957 (N_10957,N_10258,N_10053);
nor U10958 (N_10958,N_9966,N_10018);
nand U10959 (N_10959,N_9954,N_10095);
or U10960 (N_10960,N_9715,N_9611);
xor U10961 (N_10961,N_10352,N_10050);
nor U10962 (N_10962,N_10030,N_9996);
or U10963 (N_10963,N_10163,N_9627);
nor U10964 (N_10964,N_9933,N_9629);
nor U10965 (N_10965,N_10073,N_10104);
and U10966 (N_10966,N_9967,N_10239);
nor U10967 (N_10967,N_9894,N_9865);
xor U10968 (N_10968,N_9861,N_9818);
and U10969 (N_10969,N_10119,N_9659);
nand U10970 (N_10970,N_10193,N_9838);
xnor U10971 (N_10971,N_9725,N_9625);
and U10972 (N_10972,N_10207,N_10220);
nor U10973 (N_10973,N_9772,N_10149);
or U10974 (N_10974,N_10357,N_10061);
nor U10975 (N_10975,N_10085,N_9912);
xnor U10976 (N_10976,N_9812,N_10218);
xnor U10977 (N_10977,N_10369,N_9627);
nor U10978 (N_10978,N_9903,N_9843);
xor U10979 (N_10979,N_10306,N_9658);
xor U10980 (N_10980,N_10248,N_9678);
nor U10981 (N_10981,N_10179,N_9816);
xnor U10982 (N_10982,N_10007,N_9974);
and U10983 (N_10983,N_9626,N_10040);
xnor U10984 (N_10984,N_10041,N_9611);
nand U10985 (N_10985,N_9941,N_9615);
nand U10986 (N_10986,N_10147,N_10157);
or U10987 (N_10987,N_9736,N_10324);
nand U10988 (N_10988,N_9910,N_10397);
or U10989 (N_10989,N_10257,N_9665);
or U10990 (N_10990,N_9620,N_9811);
and U10991 (N_10991,N_9715,N_9929);
and U10992 (N_10992,N_10205,N_9827);
and U10993 (N_10993,N_10240,N_10073);
or U10994 (N_10994,N_9820,N_9699);
nand U10995 (N_10995,N_10332,N_9900);
and U10996 (N_10996,N_10252,N_9920);
or U10997 (N_10997,N_10127,N_9998);
nand U10998 (N_10998,N_9764,N_10069);
or U10999 (N_10999,N_10117,N_9970);
xnor U11000 (N_11000,N_9773,N_9808);
or U11001 (N_11001,N_9755,N_10035);
nor U11002 (N_11002,N_10120,N_9810);
xor U11003 (N_11003,N_9841,N_9977);
nor U11004 (N_11004,N_9973,N_9778);
nand U11005 (N_11005,N_10055,N_9882);
or U11006 (N_11006,N_10207,N_10146);
and U11007 (N_11007,N_9795,N_9902);
nor U11008 (N_11008,N_10073,N_10009);
and U11009 (N_11009,N_9733,N_10018);
nor U11010 (N_11010,N_10198,N_9746);
or U11011 (N_11011,N_10315,N_9906);
nor U11012 (N_11012,N_9773,N_9832);
nand U11013 (N_11013,N_9822,N_10017);
or U11014 (N_11014,N_10196,N_10264);
or U11015 (N_11015,N_10327,N_10003);
nand U11016 (N_11016,N_9652,N_10318);
nand U11017 (N_11017,N_9758,N_9989);
xor U11018 (N_11018,N_10160,N_9733);
xnor U11019 (N_11019,N_9707,N_9621);
and U11020 (N_11020,N_10052,N_10136);
nand U11021 (N_11021,N_10057,N_10317);
or U11022 (N_11022,N_10059,N_10049);
and U11023 (N_11023,N_10205,N_10031);
nand U11024 (N_11024,N_10180,N_9654);
nand U11025 (N_11025,N_9892,N_9844);
nand U11026 (N_11026,N_9799,N_9964);
nand U11027 (N_11027,N_9900,N_9804);
or U11028 (N_11028,N_9713,N_9808);
or U11029 (N_11029,N_10387,N_9609);
or U11030 (N_11030,N_10232,N_10204);
nor U11031 (N_11031,N_9703,N_10227);
and U11032 (N_11032,N_10337,N_10001);
and U11033 (N_11033,N_10090,N_10092);
nand U11034 (N_11034,N_9954,N_10149);
and U11035 (N_11035,N_9871,N_9693);
and U11036 (N_11036,N_10024,N_10223);
xnor U11037 (N_11037,N_10208,N_9652);
nor U11038 (N_11038,N_9939,N_10100);
xnor U11039 (N_11039,N_10126,N_9833);
xor U11040 (N_11040,N_10361,N_10320);
and U11041 (N_11041,N_10182,N_10136);
nand U11042 (N_11042,N_10243,N_9910);
nand U11043 (N_11043,N_10293,N_10089);
nor U11044 (N_11044,N_9671,N_10271);
xor U11045 (N_11045,N_9664,N_9644);
or U11046 (N_11046,N_9974,N_10300);
or U11047 (N_11047,N_10072,N_9978);
nor U11048 (N_11048,N_10201,N_9877);
xor U11049 (N_11049,N_9647,N_10201);
and U11050 (N_11050,N_10040,N_10144);
nor U11051 (N_11051,N_10265,N_9811);
and U11052 (N_11052,N_9640,N_10145);
or U11053 (N_11053,N_10099,N_9724);
xor U11054 (N_11054,N_9967,N_10048);
and U11055 (N_11055,N_10134,N_10311);
xnor U11056 (N_11056,N_9818,N_10064);
and U11057 (N_11057,N_10025,N_10055);
or U11058 (N_11058,N_10336,N_10248);
nor U11059 (N_11059,N_9907,N_9988);
nor U11060 (N_11060,N_9698,N_9652);
and U11061 (N_11061,N_9713,N_10043);
nor U11062 (N_11062,N_9735,N_9630);
and U11063 (N_11063,N_9972,N_10185);
or U11064 (N_11064,N_10037,N_9900);
nand U11065 (N_11065,N_10295,N_10038);
or U11066 (N_11066,N_10227,N_10018);
and U11067 (N_11067,N_10067,N_9846);
xnor U11068 (N_11068,N_9796,N_10369);
and U11069 (N_11069,N_10018,N_10242);
nor U11070 (N_11070,N_10005,N_9857);
xnor U11071 (N_11071,N_9711,N_9839);
nand U11072 (N_11072,N_10023,N_9788);
and U11073 (N_11073,N_9973,N_9621);
nor U11074 (N_11074,N_9864,N_10099);
xnor U11075 (N_11075,N_9831,N_10113);
nand U11076 (N_11076,N_9992,N_9742);
nor U11077 (N_11077,N_10062,N_9679);
or U11078 (N_11078,N_10113,N_10007);
and U11079 (N_11079,N_9660,N_10242);
or U11080 (N_11080,N_10357,N_9826);
xnor U11081 (N_11081,N_10058,N_9663);
xnor U11082 (N_11082,N_9682,N_9813);
and U11083 (N_11083,N_10230,N_9666);
nand U11084 (N_11084,N_9830,N_9854);
and U11085 (N_11085,N_9781,N_9844);
xor U11086 (N_11086,N_9698,N_10391);
or U11087 (N_11087,N_9832,N_9930);
xnor U11088 (N_11088,N_9984,N_10114);
or U11089 (N_11089,N_9794,N_10000);
and U11090 (N_11090,N_10083,N_10347);
or U11091 (N_11091,N_10274,N_9848);
xnor U11092 (N_11092,N_10391,N_9723);
xor U11093 (N_11093,N_9748,N_9922);
nor U11094 (N_11094,N_10381,N_10025);
and U11095 (N_11095,N_10280,N_10333);
nor U11096 (N_11096,N_9916,N_9881);
or U11097 (N_11097,N_9619,N_10076);
or U11098 (N_11098,N_9717,N_9665);
nand U11099 (N_11099,N_10094,N_10269);
xnor U11100 (N_11100,N_10210,N_10323);
nor U11101 (N_11101,N_9961,N_9948);
or U11102 (N_11102,N_9605,N_9697);
nor U11103 (N_11103,N_9980,N_10217);
xor U11104 (N_11104,N_9634,N_10363);
or U11105 (N_11105,N_10020,N_10138);
and U11106 (N_11106,N_10017,N_9950);
or U11107 (N_11107,N_10034,N_9998);
xor U11108 (N_11108,N_9961,N_10042);
nor U11109 (N_11109,N_10335,N_9692);
or U11110 (N_11110,N_10226,N_10231);
xnor U11111 (N_11111,N_10201,N_10393);
and U11112 (N_11112,N_9782,N_10023);
nor U11113 (N_11113,N_10274,N_9889);
or U11114 (N_11114,N_10210,N_9811);
nand U11115 (N_11115,N_10316,N_9749);
nand U11116 (N_11116,N_9615,N_9783);
and U11117 (N_11117,N_9643,N_9930);
xnor U11118 (N_11118,N_10379,N_9635);
or U11119 (N_11119,N_10283,N_9858);
nand U11120 (N_11120,N_10282,N_10207);
and U11121 (N_11121,N_9690,N_10165);
nor U11122 (N_11122,N_9811,N_10087);
and U11123 (N_11123,N_9954,N_10052);
nor U11124 (N_11124,N_9901,N_10346);
nand U11125 (N_11125,N_9780,N_9826);
nand U11126 (N_11126,N_9641,N_10277);
xor U11127 (N_11127,N_10092,N_9826);
or U11128 (N_11128,N_10070,N_10334);
xor U11129 (N_11129,N_10354,N_10136);
nand U11130 (N_11130,N_9894,N_10076);
and U11131 (N_11131,N_10074,N_9966);
nand U11132 (N_11132,N_10144,N_9988);
and U11133 (N_11133,N_10277,N_9724);
xor U11134 (N_11134,N_10373,N_10101);
nor U11135 (N_11135,N_9607,N_9708);
xor U11136 (N_11136,N_10135,N_10203);
xor U11137 (N_11137,N_10139,N_9930);
nand U11138 (N_11138,N_10136,N_10226);
nand U11139 (N_11139,N_9704,N_9746);
nand U11140 (N_11140,N_9736,N_9766);
nor U11141 (N_11141,N_10084,N_10108);
nand U11142 (N_11142,N_10382,N_9762);
xor U11143 (N_11143,N_10341,N_9766);
xnor U11144 (N_11144,N_10361,N_9743);
nand U11145 (N_11145,N_10322,N_10278);
nor U11146 (N_11146,N_10130,N_9669);
or U11147 (N_11147,N_9849,N_10192);
xor U11148 (N_11148,N_10278,N_9997);
nor U11149 (N_11149,N_9693,N_10139);
xnor U11150 (N_11150,N_9815,N_9831);
or U11151 (N_11151,N_10213,N_9868);
nor U11152 (N_11152,N_9788,N_9974);
and U11153 (N_11153,N_10312,N_9722);
or U11154 (N_11154,N_9852,N_9894);
nor U11155 (N_11155,N_9650,N_10120);
nor U11156 (N_11156,N_9930,N_9875);
or U11157 (N_11157,N_9722,N_9877);
nand U11158 (N_11158,N_9750,N_10355);
or U11159 (N_11159,N_9693,N_10355);
nor U11160 (N_11160,N_9980,N_10315);
and U11161 (N_11161,N_9722,N_10333);
nor U11162 (N_11162,N_9625,N_9972);
nor U11163 (N_11163,N_10102,N_9982);
and U11164 (N_11164,N_9897,N_9806);
or U11165 (N_11165,N_9889,N_9969);
and U11166 (N_11166,N_9823,N_10290);
xnor U11167 (N_11167,N_10062,N_10195);
nor U11168 (N_11168,N_10256,N_10088);
xor U11169 (N_11169,N_9613,N_9865);
nor U11170 (N_11170,N_10331,N_10287);
and U11171 (N_11171,N_10305,N_10260);
nor U11172 (N_11172,N_10015,N_9945);
or U11173 (N_11173,N_9625,N_10064);
xnor U11174 (N_11174,N_9647,N_9947);
nand U11175 (N_11175,N_9729,N_9902);
and U11176 (N_11176,N_9636,N_9870);
nand U11177 (N_11177,N_9839,N_10379);
nand U11178 (N_11178,N_10108,N_10383);
or U11179 (N_11179,N_10037,N_10377);
nor U11180 (N_11180,N_10001,N_10397);
or U11181 (N_11181,N_9671,N_10071);
nor U11182 (N_11182,N_10322,N_10088);
or U11183 (N_11183,N_10095,N_10065);
nand U11184 (N_11184,N_9714,N_9764);
nand U11185 (N_11185,N_10080,N_9999);
nor U11186 (N_11186,N_10296,N_9609);
xnor U11187 (N_11187,N_10326,N_10036);
nand U11188 (N_11188,N_10369,N_10005);
nor U11189 (N_11189,N_9787,N_10142);
or U11190 (N_11190,N_10278,N_10266);
nand U11191 (N_11191,N_10051,N_10379);
or U11192 (N_11192,N_10342,N_10208);
nor U11193 (N_11193,N_9970,N_9765);
nand U11194 (N_11194,N_9990,N_9877);
or U11195 (N_11195,N_9989,N_10102);
or U11196 (N_11196,N_10108,N_10176);
or U11197 (N_11197,N_10210,N_10262);
and U11198 (N_11198,N_10168,N_9828);
nand U11199 (N_11199,N_9992,N_9893);
and U11200 (N_11200,N_10739,N_10666);
nand U11201 (N_11201,N_10876,N_10866);
or U11202 (N_11202,N_11183,N_10759);
nand U11203 (N_11203,N_10492,N_10547);
xor U11204 (N_11204,N_10663,N_10472);
and U11205 (N_11205,N_11105,N_10653);
nor U11206 (N_11206,N_10977,N_10921);
or U11207 (N_11207,N_10792,N_10804);
nor U11208 (N_11208,N_10627,N_10545);
nor U11209 (N_11209,N_10907,N_10974);
or U11210 (N_11210,N_11109,N_10461);
xor U11211 (N_11211,N_11083,N_10701);
nor U11212 (N_11212,N_11057,N_11143);
nand U11213 (N_11213,N_10903,N_10772);
nor U11214 (N_11214,N_10563,N_11156);
xor U11215 (N_11215,N_11119,N_10401);
xnor U11216 (N_11216,N_10507,N_11079);
xnor U11217 (N_11217,N_10508,N_11001);
and U11218 (N_11218,N_10665,N_10433);
xnor U11219 (N_11219,N_11164,N_10931);
xnor U11220 (N_11220,N_11014,N_10798);
nand U11221 (N_11221,N_10549,N_10402);
or U11222 (N_11222,N_10744,N_10721);
nand U11223 (N_11223,N_11080,N_10446);
xor U11224 (N_11224,N_10523,N_10832);
or U11225 (N_11225,N_10825,N_10843);
xnor U11226 (N_11226,N_10990,N_10583);
xor U11227 (N_11227,N_10518,N_11177);
nand U11228 (N_11228,N_10453,N_10889);
or U11229 (N_11229,N_11029,N_10766);
and U11230 (N_11230,N_10521,N_10513);
nand U11231 (N_11231,N_10970,N_10934);
xnor U11232 (N_11232,N_10953,N_10748);
nor U11233 (N_11233,N_10763,N_10509);
nor U11234 (N_11234,N_11131,N_10878);
nor U11235 (N_11235,N_11019,N_10578);
nor U11236 (N_11236,N_10629,N_10593);
nand U11237 (N_11237,N_10613,N_10923);
xor U11238 (N_11238,N_10860,N_10617);
or U11239 (N_11239,N_10947,N_10598);
or U11240 (N_11240,N_10719,N_10528);
nor U11241 (N_11241,N_10691,N_11166);
nor U11242 (N_11242,N_11043,N_10846);
or U11243 (N_11243,N_10768,N_10526);
nor U11244 (N_11244,N_10609,N_11161);
or U11245 (N_11245,N_10722,N_10800);
or U11246 (N_11246,N_10992,N_10415);
nor U11247 (N_11247,N_10801,N_10979);
or U11248 (N_11248,N_10638,N_11005);
nor U11249 (N_11249,N_10877,N_11142);
and U11250 (N_11250,N_10569,N_10794);
or U11251 (N_11251,N_10536,N_10863);
and U11252 (N_11252,N_10475,N_10795);
nor U11253 (N_11253,N_10943,N_10965);
and U11254 (N_11254,N_11189,N_10912);
xor U11255 (N_11255,N_11162,N_10410);
or U11256 (N_11256,N_10491,N_10532);
nand U11257 (N_11257,N_11123,N_10892);
or U11258 (N_11258,N_10867,N_11058);
or U11259 (N_11259,N_11072,N_10944);
or U11260 (N_11260,N_10793,N_10622);
nor U11261 (N_11261,N_10505,N_10407);
nand U11262 (N_11262,N_10625,N_11037);
or U11263 (N_11263,N_10933,N_10618);
xnor U11264 (N_11264,N_10548,N_10477);
and U11265 (N_11265,N_10811,N_11113);
and U11266 (N_11266,N_10418,N_10836);
or U11267 (N_11267,N_10585,N_10676);
and U11268 (N_11268,N_10993,N_10678);
and U11269 (N_11269,N_10888,N_10727);
nand U11270 (N_11270,N_11153,N_10850);
nor U11271 (N_11271,N_10459,N_10753);
nor U11272 (N_11272,N_10680,N_10777);
nor U11273 (N_11273,N_10499,N_10738);
and U11274 (N_11274,N_10731,N_10637);
nand U11275 (N_11275,N_10802,N_10538);
xor U11276 (N_11276,N_10874,N_10660);
or U11277 (N_11277,N_10964,N_10790);
nand U11278 (N_11278,N_10774,N_11071);
or U11279 (N_11279,N_11016,N_10529);
xnor U11280 (N_11280,N_11170,N_11084);
xor U11281 (N_11281,N_10769,N_10754);
and U11282 (N_11282,N_11158,N_10899);
xor U11283 (N_11283,N_11042,N_10403);
nand U11284 (N_11284,N_11012,N_11063);
and U11285 (N_11285,N_10434,N_11068);
or U11286 (N_11286,N_10833,N_10568);
xor U11287 (N_11287,N_10565,N_10514);
xor U11288 (N_11288,N_11052,N_10670);
and U11289 (N_11289,N_11046,N_11098);
nor U11290 (N_11290,N_10460,N_10881);
nand U11291 (N_11291,N_11074,N_10740);
or U11292 (N_11292,N_10552,N_10695);
or U11293 (N_11293,N_11184,N_10601);
or U11294 (N_11294,N_10983,N_11127);
xnor U11295 (N_11295,N_11062,N_10517);
nand U11296 (N_11296,N_10996,N_11140);
or U11297 (N_11297,N_10422,N_10581);
or U11298 (N_11298,N_10803,N_11064);
nor U11299 (N_11299,N_10633,N_10474);
nand U11300 (N_11300,N_10969,N_10819);
nand U11301 (N_11301,N_10649,N_10817);
nor U11302 (N_11302,N_10821,N_10659);
nor U11303 (N_11303,N_10948,N_10962);
and U11304 (N_11304,N_10955,N_11171);
or U11305 (N_11305,N_11073,N_10857);
or U11306 (N_11306,N_10594,N_10939);
or U11307 (N_11307,N_10852,N_10734);
and U11308 (N_11308,N_10883,N_11053);
nand U11309 (N_11309,N_10932,N_10546);
nor U11310 (N_11310,N_10648,N_10635);
nand U11311 (N_11311,N_10986,N_10956);
xor U11312 (N_11312,N_10554,N_11047);
nor U11313 (N_11313,N_10539,N_10628);
nor U11314 (N_11314,N_11149,N_10579);
nor U11315 (N_11315,N_10968,N_10851);
or U11316 (N_11316,N_11134,N_11110);
or U11317 (N_11317,N_11102,N_10732);
nor U11318 (N_11318,N_11157,N_10611);
xnor U11319 (N_11319,N_11106,N_10455);
or U11320 (N_11320,N_10914,N_10466);
nor U11321 (N_11321,N_11069,N_10421);
and U11322 (N_11322,N_11118,N_10761);
nor U11323 (N_11323,N_11129,N_11040);
and U11324 (N_11324,N_10597,N_10820);
xor U11325 (N_11325,N_10543,N_10950);
nor U11326 (N_11326,N_10668,N_10527);
nor U11327 (N_11327,N_10488,N_10901);
nor U11328 (N_11328,N_11015,N_10989);
or U11329 (N_11329,N_10686,N_10560);
nor U11330 (N_11330,N_10988,N_10810);
and U11331 (N_11331,N_11032,N_10963);
xnor U11332 (N_11332,N_11146,N_10440);
nand U11333 (N_11333,N_10607,N_10473);
or U11334 (N_11334,N_10831,N_10842);
or U11335 (N_11335,N_11041,N_10835);
and U11336 (N_11336,N_10480,N_10822);
and U11337 (N_11337,N_10760,N_10639);
nand U11338 (N_11338,N_10544,N_10589);
xor U11339 (N_11339,N_10503,N_11160);
or U11340 (N_11340,N_10524,N_10784);
nor U11341 (N_11341,N_10862,N_10954);
nand U11342 (N_11342,N_11121,N_10805);
nand U11343 (N_11343,N_10808,N_11155);
and U11344 (N_11344,N_10689,N_10870);
nand U11345 (N_11345,N_10551,N_11009);
xor U11346 (N_11346,N_10957,N_10708);
nand U11347 (N_11347,N_10571,N_11199);
or U11348 (N_11348,N_10869,N_10516);
nor U11349 (N_11349,N_10511,N_10787);
and U11350 (N_11350,N_11112,N_10814);
nand U11351 (N_11351,N_10773,N_10655);
nand U11352 (N_11352,N_11025,N_10839);
and U11353 (N_11353,N_10693,N_11187);
or U11354 (N_11354,N_10724,N_10723);
xnor U11355 (N_11355,N_10652,N_11198);
nand U11356 (N_11356,N_10971,N_10478);
and U11357 (N_11357,N_10519,N_10864);
nand U11358 (N_11358,N_11060,N_10645);
or U11359 (N_11359,N_11033,N_10902);
xor U11360 (N_11360,N_10677,N_11036);
xor U11361 (N_11361,N_11054,N_10929);
or U11362 (N_11362,N_10646,N_10493);
nand U11363 (N_11363,N_11159,N_11197);
nand U11364 (N_11364,N_10606,N_10577);
nand U11365 (N_11365,N_10829,N_10641);
xnor U11366 (N_11366,N_10624,N_10604);
or U11367 (N_11367,N_10502,N_10920);
or U11368 (N_11368,N_10906,N_10510);
and U11369 (N_11369,N_11099,N_11095);
nor U11370 (N_11370,N_10631,N_10926);
nand U11371 (N_11371,N_10783,N_11039);
or U11372 (N_11372,N_11006,N_10978);
and U11373 (N_11373,N_10779,N_10973);
nand U11374 (N_11374,N_10856,N_11013);
or U11375 (N_11375,N_11116,N_10743);
or U11376 (N_11376,N_11018,N_10497);
nand U11377 (N_11377,N_11137,N_11124);
or U11378 (N_11378,N_10746,N_10797);
xnor U11379 (N_11379,N_11089,N_10827);
or U11380 (N_11380,N_10726,N_10632);
or U11381 (N_11381,N_10443,N_11190);
nor U11382 (N_11382,N_11007,N_11061);
and U11383 (N_11383,N_11154,N_10413);
nand U11384 (N_11384,N_11144,N_10531);
nand U11385 (N_11385,N_10580,N_10952);
nand U11386 (N_11386,N_10462,N_11126);
nor U11387 (N_11387,N_10872,N_11091);
nor U11388 (N_11388,N_10995,N_11151);
xnor U11389 (N_11389,N_11076,N_11023);
nor U11390 (N_11390,N_10467,N_10584);
nand U11391 (N_11391,N_10690,N_10555);
and U11392 (N_11392,N_10845,N_10559);
nand U11393 (N_11393,N_11176,N_10927);
or U11394 (N_11394,N_10564,N_10702);
nor U11395 (N_11395,N_11030,N_10897);
xnor U11396 (N_11396,N_10737,N_10966);
and U11397 (N_11397,N_10896,N_11093);
nor U11398 (N_11398,N_10465,N_10816);
and U11399 (N_11399,N_10476,N_10776);
and U11400 (N_11400,N_11191,N_10840);
and U11401 (N_11401,N_11002,N_10941);
nor U11402 (N_11402,N_10998,N_11165);
nor U11403 (N_11403,N_10710,N_11020);
xnor U11404 (N_11404,N_10592,N_11108);
xnor U11405 (N_11405,N_10470,N_10664);
xnor U11406 (N_11406,N_10916,N_11044);
xnor U11407 (N_11407,N_10733,N_10640);
xnor U11408 (N_11408,N_10409,N_10904);
and U11409 (N_11409,N_11194,N_10898);
or U11410 (N_11410,N_11094,N_10918);
nor U11411 (N_11411,N_10938,N_11010);
nand U11412 (N_11412,N_10736,N_10917);
and U11413 (N_11413,N_10868,N_10700);
xor U11414 (N_11414,N_10781,N_10642);
xnor U11415 (N_11415,N_10999,N_10847);
nor U11416 (N_11416,N_10533,N_10841);
nor U11417 (N_11417,N_10537,N_10765);
nand U11418 (N_11418,N_10770,N_10930);
nor U11419 (N_11419,N_11085,N_10806);
xnor U11420 (N_11420,N_11065,N_11000);
nor U11421 (N_11421,N_11090,N_10411);
nor U11422 (N_11422,N_10501,N_10987);
nor U11423 (N_11423,N_10436,N_11092);
nor U11424 (N_11424,N_10698,N_10540);
nor U11425 (N_11425,N_10600,N_11114);
nand U11426 (N_11426,N_10570,N_10438);
or U11427 (N_11427,N_10515,N_10818);
or U11428 (N_11428,N_10729,N_10449);
or U11429 (N_11429,N_10975,N_10915);
xor U11430 (N_11430,N_10458,N_10699);
nor U11431 (N_11431,N_11051,N_10684);
and U11432 (N_11432,N_11172,N_11097);
xnor U11433 (N_11433,N_10454,N_11133);
xnor U11434 (N_11434,N_10406,N_10780);
nor U11435 (N_11435,N_10813,N_11167);
nor U11436 (N_11436,N_11048,N_10709);
or U11437 (N_11437,N_10880,N_10960);
nor U11438 (N_11438,N_11115,N_10587);
xnor U11439 (N_11439,N_10982,N_11096);
nor U11440 (N_11440,N_11175,N_10504);
or U11441 (N_11441,N_10573,N_10558);
nand U11442 (N_11442,N_10444,N_11082);
nor U11443 (N_11443,N_10450,N_10481);
xor U11444 (N_11444,N_11188,N_10498);
and U11445 (N_11445,N_10796,N_10582);
nand U11446 (N_11446,N_10716,N_10757);
nand U11447 (N_11447,N_10662,N_10935);
and U11448 (N_11448,N_11173,N_10855);
nand U11449 (N_11449,N_11179,N_11182);
xor U11450 (N_11450,N_11148,N_11086);
or U11451 (N_11451,N_11034,N_10886);
and U11452 (N_11452,N_10442,N_11168);
nor U11453 (N_11453,N_10913,N_10482);
xor U11454 (N_11454,N_10991,N_10672);
xor U11455 (N_11455,N_10725,N_10522);
nor U11456 (N_11456,N_10464,N_10644);
nand U11457 (N_11457,N_10643,N_10423);
and U11458 (N_11458,N_10425,N_11147);
nor U11459 (N_11459,N_10688,N_11120);
or U11460 (N_11460,N_10534,N_10919);
or U11461 (N_11461,N_10445,N_10807);
nor U11462 (N_11462,N_10890,N_10400);
or U11463 (N_11463,N_10961,N_10512);
nand U11464 (N_11464,N_10785,N_10542);
xor U11465 (N_11465,N_10484,N_10849);
nand U11466 (N_11466,N_10535,N_10728);
nor U11467 (N_11467,N_10778,N_10848);
nand U11468 (N_11468,N_11117,N_11049);
nand U11469 (N_11469,N_10414,N_10557);
nor U11470 (N_11470,N_10949,N_10457);
or U11471 (N_11471,N_10687,N_11136);
and U11472 (N_11472,N_10416,N_10426);
nor U11473 (N_11473,N_10500,N_10468);
nand U11474 (N_11474,N_11077,N_10647);
nor U11475 (N_11475,N_10891,N_11067);
or U11476 (N_11476,N_10925,N_10494);
nand U11477 (N_11477,N_10742,N_11008);
or U11478 (N_11478,N_10762,N_10745);
xor U11479 (N_11479,N_10658,N_10656);
nand U11480 (N_11480,N_10682,N_10981);
nor U11481 (N_11481,N_10630,N_11024);
or U11482 (N_11482,N_10614,N_10900);
or U11483 (N_11483,N_10885,N_10603);
and U11484 (N_11484,N_10574,N_11027);
xor U11485 (N_11485,N_11122,N_11101);
and U11486 (N_11486,N_10887,N_10435);
xor U11487 (N_11487,N_10674,N_10749);
xor U11488 (N_11488,N_10942,N_11128);
nand U11489 (N_11489,N_10590,N_10837);
nor U11490 (N_11490,N_11178,N_10408);
nor U11491 (N_11491,N_11145,N_10994);
and U11492 (N_11492,N_11169,N_11139);
nand U11493 (N_11493,N_11021,N_10853);
and U11494 (N_11494,N_10834,N_10824);
nand U11495 (N_11495,N_10882,N_10786);
or U11496 (N_11496,N_11011,N_10984);
or U11497 (N_11497,N_10767,N_11078);
xnor U11498 (N_11498,N_10405,N_10679);
or U11499 (N_11499,N_10789,N_10859);
nand U11500 (N_11500,N_10424,N_10730);
or U11501 (N_11501,N_10854,N_10448);
or U11502 (N_11502,N_10741,N_10871);
nand U11503 (N_11503,N_10657,N_10720);
xnor U11504 (N_11504,N_10951,N_10815);
xnor U11505 (N_11505,N_11150,N_10764);
or U11506 (N_11506,N_11130,N_10707);
nor U11507 (N_11507,N_10591,N_11125);
xor U11508 (N_11508,N_10922,N_10479);
nor U11509 (N_11509,N_11038,N_10626);
xnor U11510 (N_11510,N_10483,N_11003);
or U11511 (N_11511,N_10605,N_10608);
or U11512 (N_11512,N_10550,N_10972);
nand U11513 (N_11513,N_10958,N_10752);
xnor U11514 (N_11514,N_10496,N_10967);
or U11515 (N_11515,N_11163,N_10735);
or U11516 (N_11516,N_10826,N_11100);
nor U11517 (N_11517,N_10771,N_10615);
or U11518 (N_11518,N_10432,N_10623);
nand U11519 (N_11519,N_10809,N_10487);
and U11520 (N_11520,N_10905,N_11186);
nand U11521 (N_11521,N_10612,N_10650);
or U11522 (N_11522,N_10576,N_10506);
nand U11523 (N_11523,N_10541,N_11180);
and U11524 (N_11524,N_11059,N_10858);
and U11525 (N_11525,N_10980,N_10959);
or U11526 (N_11526,N_10782,N_10911);
xor U11527 (N_11527,N_10704,N_11192);
nor U11528 (N_11528,N_10675,N_11081);
or U11529 (N_11529,N_10431,N_10705);
and U11530 (N_11530,N_11004,N_10908);
xnor U11531 (N_11531,N_10489,N_10756);
and U11532 (N_11532,N_10703,N_10669);
nor U11533 (N_11533,N_10429,N_10596);
nor U11534 (N_11534,N_10439,N_10595);
or U11535 (N_11535,N_10812,N_10575);
xor U11536 (N_11536,N_10799,N_10486);
nor U11537 (N_11537,N_10924,N_10828);
and U11538 (N_11538,N_10879,N_10667);
nand U11539 (N_11539,N_10936,N_10884);
xnor U11540 (N_11540,N_10946,N_10976);
nand U11541 (N_11541,N_10873,N_10928);
nand U11542 (N_11542,N_11107,N_10530);
or U11543 (N_11543,N_10586,N_11070);
nor U11544 (N_11544,N_11193,N_10621);
nand U11545 (N_11545,N_10636,N_11174);
or U11546 (N_11546,N_11138,N_10562);
xor U11547 (N_11547,N_10620,N_10692);
nand U11548 (N_11548,N_10937,N_10520);
or U11549 (N_11549,N_10556,N_10718);
or U11550 (N_11550,N_10412,N_11017);
nor U11551 (N_11551,N_10654,N_10909);
nand U11552 (N_11552,N_10713,N_10683);
and U11553 (N_11553,N_10430,N_11181);
nor U11554 (N_11554,N_11195,N_10495);
and U11555 (N_11555,N_11152,N_10712);
and U11556 (N_11556,N_10452,N_10940);
or U11557 (N_11557,N_10715,N_10673);
and U11558 (N_11558,N_10404,N_11196);
xnor U11559 (N_11559,N_11135,N_10463);
nand U11560 (N_11560,N_11056,N_10525);
nand U11561 (N_11561,N_10788,N_10711);
xor U11562 (N_11562,N_10694,N_10447);
or U11563 (N_11563,N_10417,N_10610);
nand U11564 (N_11564,N_10651,N_11087);
or U11565 (N_11565,N_11050,N_10706);
xor U11566 (N_11566,N_10838,N_10619);
xnor U11567 (N_11567,N_10588,N_10420);
xnor U11568 (N_11568,N_10865,N_10602);
nand U11569 (N_11569,N_11035,N_10750);
or U11570 (N_11570,N_11075,N_10456);
nand U11571 (N_11571,N_10945,N_11111);
or U11572 (N_11572,N_10758,N_10567);
nand U11573 (N_11573,N_10791,N_10875);
nand U11574 (N_11574,N_10616,N_11031);
and U11575 (N_11575,N_10910,N_10696);
xnor U11576 (N_11576,N_10553,N_10634);
nor U11577 (N_11577,N_11045,N_10685);
nor U11578 (N_11578,N_11132,N_10747);
and U11579 (N_11579,N_11022,N_11066);
nor U11580 (N_11580,N_11104,N_10441);
and U11581 (N_11581,N_10599,N_10419);
nand U11582 (N_11582,N_10485,N_10681);
and U11583 (N_11583,N_11141,N_10844);
nor U11584 (N_11584,N_11055,N_10471);
or U11585 (N_11585,N_10895,N_10717);
and U11586 (N_11586,N_10823,N_11103);
nor U11587 (N_11587,N_10671,N_10751);
or U11588 (N_11588,N_10775,N_11026);
or U11589 (N_11589,N_10572,N_10437);
or U11590 (N_11590,N_10861,N_10997);
and U11591 (N_11591,N_10985,N_10830);
nor U11592 (N_11592,N_10451,N_10427);
and U11593 (N_11593,N_10428,N_11185);
nor U11594 (N_11594,N_10469,N_10714);
xor U11595 (N_11595,N_10697,N_10755);
nor U11596 (N_11596,N_10661,N_11088);
nand U11597 (N_11597,N_10490,N_10566);
nor U11598 (N_11598,N_10894,N_10893);
xor U11599 (N_11599,N_10561,N_11028);
xnor U11600 (N_11600,N_10620,N_10438);
xnor U11601 (N_11601,N_10714,N_10992);
and U11602 (N_11602,N_10538,N_11069);
nand U11603 (N_11603,N_10531,N_10994);
and U11604 (N_11604,N_11045,N_10743);
xor U11605 (N_11605,N_10953,N_10596);
xor U11606 (N_11606,N_10533,N_10493);
or U11607 (N_11607,N_10493,N_10924);
nor U11608 (N_11608,N_10712,N_10440);
or U11609 (N_11609,N_10551,N_10621);
nand U11610 (N_11610,N_10594,N_10992);
nand U11611 (N_11611,N_10595,N_10685);
nor U11612 (N_11612,N_10662,N_10812);
nor U11613 (N_11613,N_10587,N_10597);
nor U11614 (N_11614,N_10754,N_10707);
nand U11615 (N_11615,N_10491,N_10768);
xnor U11616 (N_11616,N_11046,N_10670);
and U11617 (N_11617,N_11108,N_10840);
and U11618 (N_11618,N_10732,N_10986);
or U11619 (N_11619,N_10539,N_11125);
nand U11620 (N_11620,N_10594,N_10697);
nand U11621 (N_11621,N_10717,N_10783);
or U11622 (N_11622,N_10691,N_11131);
and U11623 (N_11623,N_10845,N_10472);
xor U11624 (N_11624,N_11185,N_10877);
or U11625 (N_11625,N_10495,N_10991);
xnor U11626 (N_11626,N_10931,N_10660);
nand U11627 (N_11627,N_10568,N_11003);
or U11628 (N_11628,N_10844,N_10822);
xnor U11629 (N_11629,N_10962,N_10572);
or U11630 (N_11630,N_10595,N_10641);
nor U11631 (N_11631,N_10424,N_10978);
nand U11632 (N_11632,N_10817,N_10607);
nor U11633 (N_11633,N_10858,N_11150);
or U11634 (N_11634,N_10485,N_10566);
and U11635 (N_11635,N_10449,N_10437);
nand U11636 (N_11636,N_11172,N_11045);
xor U11637 (N_11637,N_10603,N_11090);
nor U11638 (N_11638,N_10937,N_11021);
and U11639 (N_11639,N_10416,N_10953);
xor U11640 (N_11640,N_10500,N_10746);
and U11641 (N_11641,N_10676,N_10881);
xnor U11642 (N_11642,N_10474,N_11046);
xnor U11643 (N_11643,N_10807,N_10697);
and U11644 (N_11644,N_11131,N_10575);
nand U11645 (N_11645,N_10746,N_10431);
nand U11646 (N_11646,N_10594,N_11051);
xor U11647 (N_11647,N_10931,N_11072);
nor U11648 (N_11648,N_10759,N_10703);
nor U11649 (N_11649,N_10962,N_11046);
nand U11650 (N_11650,N_10789,N_10696);
nor U11651 (N_11651,N_10568,N_11184);
nand U11652 (N_11652,N_11106,N_11046);
nand U11653 (N_11653,N_10941,N_10793);
xor U11654 (N_11654,N_10735,N_10928);
and U11655 (N_11655,N_10980,N_10935);
nor U11656 (N_11656,N_11118,N_10581);
and U11657 (N_11657,N_10548,N_11127);
and U11658 (N_11658,N_10704,N_10482);
xor U11659 (N_11659,N_10830,N_10696);
or U11660 (N_11660,N_10466,N_10475);
nand U11661 (N_11661,N_10809,N_11185);
or U11662 (N_11662,N_10622,N_10662);
xor U11663 (N_11663,N_10810,N_10857);
xor U11664 (N_11664,N_11054,N_10487);
and U11665 (N_11665,N_11047,N_10867);
xnor U11666 (N_11666,N_11169,N_10911);
and U11667 (N_11667,N_11192,N_10445);
xnor U11668 (N_11668,N_10486,N_10969);
nand U11669 (N_11669,N_11160,N_10980);
or U11670 (N_11670,N_10403,N_10991);
or U11671 (N_11671,N_10916,N_10407);
nor U11672 (N_11672,N_10418,N_10902);
nand U11673 (N_11673,N_11110,N_10566);
xnor U11674 (N_11674,N_11059,N_10473);
nor U11675 (N_11675,N_10638,N_10573);
nor U11676 (N_11676,N_10521,N_10662);
xor U11677 (N_11677,N_11010,N_11043);
nand U11678 (N_11678,N_10531,N_10787);
nand U11679 (N_11679,N_11013,N_11012);
nor U11680 (N_11680,N_10797,N_11117);
nor U11681 (N_11681,N_10658,N_11091);
nand U11682 (N_11682,N_10510,N_10448);
or U11683 (N_11683,N_10793,N_10576);
or U11684 (N_11684,N_10664,N_11061);
xor U11685 (N_11685,N_10583,N_11141);
xor U11686 (N_11686,N_11082,N_10608);
or U11687 (N_11687,N_10511,N_11015);
nand U11688 (N_11688,N_11118,N_10797);
xnor U11689 (N_11689,N_10723,N_10914);
and U11690 (N_11690,N_10577,N_10617);
and U11691 (N_11691,N_10828,N_11079);
and U11692 (N_11692,N_10430,N_10801);
xnor U11693 (N_11693,N_10976,N_11166);
nand U11694 (N_11694,N_10689,N_10942);
nor U11695 (N_11695,N_10603,N_10769);
or U11696 (N_11696,N_10622,N_11122);
and U11697 (N_11697,N_10572,N_10681);
nand U11698 (N_11698,N_10618,N_10549);
nand U11699 (N_11699,N_10894,N_10643);
or U11700 (N_11700,N_10654,N_10784);
or U11701 (N_11701,N_10939,N_10436);
nand U11702 (N_11702,N_10921,N_10725);
xor U11703 (N_11703,N_10698,N_10755);
or U11704 (N_11704,N_10638,N_11046);
or U11705 (N_11705,N_10916,N_10720);
or U11706 (N_11706,N_10987,N_10400);
xnor U11707 (N_11707,N_10482,N_10999);
and U11708 (N_11708,N_10755,N_10643);
or U11709 (N_11709,N_10478,N_11106);
nand U11710 (N_11710,N_11022,N_10522);
or U11711 (N_11711,N_11026,N_11163);
xnor U11712 (N_11712,N_10619,N_10967);
and U11713 (N_11713,N_10972,N_11179);
xor U11714 (N_11714,N_10992,N_10559);
nand U11715 (N_11715,N_10703,N_10871);
xor U11716 (N_11716,N_10704,N_10675);
xnor U11717 (N_11717,N_11085,N_10679);
xor U11718 (N_11718,N_10490,N_10929);
xor U11719 (N_11719,N_10655,N_10896);
and U11720 (N_11720,N_10596,N_10589);
or U11721 (N_11721,N_10819,N_10410);
and U11722 (N_11722,N_11143,N_10401);
and U11723 (N_11723,N_11025,N_10581);
or U11724 (N_11724,N_10884,N_11166);
nand U11725 (N_11725,N_11003,N_11189);
nor U11726 (N_11726,N_10556,N_10803);
or U11727 (N_11727,N_11030,N_11190);
nand U11728 (N_11728,N_10736,N_10578);
nor U11729 (N_11729,N_10999,N_10994);
and U11730 (N_11730,N_10986,N_10576);
and U11731 (N_11731,N_11188,N_10926);
xnor U11732 (N_11732,N_10754,N_10429);
and U11733 (N_11733,N_10612,N_11106);
xnor U11734 (N_11734,N_10433,N_10453);
xnor U11735 (N_11735,N_10929,N_10635);
and U11736 (N_11736,N_11039,N_10456);
and U11737 (N_11737,N_11090,N_10929);
or U11738 (N_11738,N_10927,N_10790);
xor U11739 (N_11739,N_11118,N_10689);
and U11740 (N_11740,N_10948,N_11012);
nand U11741 (N_11741,N_10562,N_10969);
xnor U11742 (N_11742,N_10514,N_11191);
nand U11743 (N_11743,N_10426,N_10677);
and U11744 (N_11744,N_10794,N_10680);
or U11745 (N_11745,N_10492,N_10729);
and U11746 (N_11746,N_11149,N_11055);
and U11747 (N_11747,N_10877,N_10695);
or U11748 (N_11748,N_10955,N_10917);
xnor U11749 (N_11749,N_10966,N_10902);
nand U11750 (N_11750,N_10406,N_10471);
xor U11751 (N_11751,N_11021,N_11162);
and U11752 (N_11752,N_10903,N_11172);
nor U11753 (N_11753,N_10842,N_10470);
or U11754 (N_11754,N_10415,N_10411);
xor U11755 (N_11755,N_10732,N_10748);
xor U11756 (N_11756,N_10881,N_10584);
nor U11757 (N_11757,N_10409,N_10953);
xor U11758 (N_11758,N_10614,N_10721);
nand U11759 (N_11759,N_10481,N_10500);
nor U11760 (N_11760,N_10931,N_11142);
nor U11761 (N_11761,N_10511,N_10683);
xor U11762 (N_11762,N_11074,N_10935);
nand U11763 (N_11763,N_10648,N_10746);
xnor U11764 (N_11764,N_10742,N_10754);
nand U11765 (N_11765,N_10483,N_11061);
nor U11766 (N_11766,N_11044,N_11110);
or U11767 (N_11767,N_10859,N_10800);
and U11768 (N_11768,N_10737,N_11132);
and U11769 (N_11769,N_10623,N_10681);
xor U11770 (N_11770,N_10783,N_10517);
nor U11771 (N_11771,N_10858,N_10773);
nor U11772 (N_11772,N_11084,N_11097);
xor U11773 (N_11773,N_10778,N_10966);
xor U11774 (N_11774,N_10750,N_10804);
and U11775 (N_11775,N_11124,N_10456);
and U11776 (N_11776,N_10792,N_11003);
nor U11777 (N_11777,N_10998,N_10537);
xnor U11778 (N_11778,N_10697,N_11031);
or U11779 (N_11779,N_11149,N_10551);
xnor U11780 (N_11780,N_11180,N_10748);
and U11781 (N_11781,N_11089,N_10447);
or U11782 (N_11782,N_10753,N_11001);
and U11783 (N_11783,N_11129,N_10640);
nor U11784 (N_11784,N_10574,N_10509);
nor U11785 (N_11785,N_10673,N_10887);
nand U11786 (N_11786,N_10743,N_10652);
or U11787 (N_11787,N_11048,N_11049);
nor U11788 (N_11788,N_10482,N_10895);
xor U11789 (N_11789,N_10943,N_10811);
nor U11790 (N_11790,N_10726,N_10860);
and U11791 (N_11791,N_10430,N_11129);
xnor U11792 (N_11792,N_11154,N_10723);
nand U11793 (N_11793,N_10406,N_10555);
nand U11794 (N_11794,N_11028,N_10455);
nor U11795 (N_11795,N_10432,N_10869);
or U11796 (N_11796,N_10576,N_10602);
xnor U11797 (N_11797,N_11019,N_11035);
nand U11798 (N_11798,N_11028,N_10731);
xnor U11799 (N_11799,N_11182,N_10798);
xor U11800 (N_11800,N_10643,N_11176);
or U11801 (N_11801,N_10725,N_10707);
nor U11802 (N_11802,N_10873,N_10708);
or U11803 (N_11803,N_10921,N_10481);
or U11804 (N_11804,N_11142,N_10429);
nand U11805 (N_11805,N_10422,N_10591);
nor U11806 (N_11806,N_11042,N_10445);
nor U11807 (N_11807,N_10803,N_10688);
and U11808 (N_11808,N_10772,N_10887);
or U11809 (N_11809,N_10447,N_11187);
or U11810 (N_11810,N_11102,N_11194);
nand U11811 (N_11811,N_11171,N_10884);
and U11812 (N_11812,N_11092,N_10759);
xor U11813 (N_11813,N_10407,N_11068);
and U11814 (N_11814,N_10651,N_10983);
or U11815 (N_11815,N_10678,N_10657);
or U11816 (N_11816,N_11143,N_10595);
or U11817 (N_11817,N_10498,N_11033);
and U11818 (N_11818,N_11186,N_11019);
or U11819 (N_11819,N_10546,N_10483);
nand U11820 (N_11820,N_11089,N_10915);
nand U11821 (N_11821,N_10790,N_11187);
or U11822 (N_11822,N_10509,N_11176);
or U11823 (N_11823,N_10498,N_10869);
or U11824 (N_11824,N_10880,N_10670);
xor U11825 (N_11825,N_10664,N_10592);
xnor U11826 (N_11826,N_10749,N_10476);
and U11827 (N_11827,N_10530,N_10991);
nand U11828 (N_11828,N_10729,N_11079);
and U11829 (N_11829,N_11043,N_10491);
or U11830 (N_11830,N_11056,N_10603);
or U11831 (N_11831,N_10633,N_11040);
and U11832 (N_11832,N_10467,N_10821);
nor U11833 (N_11833,N_10671,N_10774);
nor U11834 (N_11834,N_10827,N_11127);
nor U11835 (N_11835,N_11110,N_11020);
and U11836 (N_11836,N_10408,N_10679);
nor U11837 (N_11837,N_10404,N_10846);
and U11838 (N_11838,N_10431,N_11083);
xor U11839 (N_11839,N_10450,N_10767);
nor U11840 (N_11840,N_10915,N_10893);
or U11841 (N_11841,N_10753,N_10529);
xor U11842 (N_11842,N_11042,N_11001);
or U11843 (N_11843,N_10528,N_10552);
nand U11844 (N_11844,N_11171,N_10922);
nand U11845 (N_11845,N_11027,N_10470);
nor U11846 (N_11846,N_10423,N_10504);
nand U11847 (N_11847,N_10519,N_10580);
or U11848 (N_11848,N_11073,N_11118);
nand U11849 (N_11849,N_10677,N_11183);
xnor U11850 (N_11850,N_10449,N_10826);
nor U11851 (N_11851,N_10692,N_10573);
xor U11852 (N_11852,N_10820,N_10687);
nand U11853 (N_11853,N_11010,N_11108);
and U11854 (N_11854,N_10639,N_11085);
or U11855 (N_11855,N_11073,N_10823);
nand U11856 (N_11856,N_10918,N_11119);
nand U11857 (N_11857,N_10538,N_10868);
and U11858 (N_11858,N_10445,N_10460);
and U11859 (N_11859,N_11083,N_10608);
or U11860 (N_11860,N_11019,N_11138);
nor U11861 (N_11861,N_10428,N_10461);
nor U11862 (N_11862,N_10412,N_11198);
xnor U11863 (N_11863,N_11008,N_10472);
or U11864 (N_11864,N_10799,N_10631);
nor U11865 (N_11865,N_10571,N_10419);
and U11866 (N_11866,N_10600,N_10987);
nor U11867 (N_11867,N_10908,N_10677);
nand U11868 (N_11868,N_10681,N_10730);
nor U11869 (N_11869,N_10713,N_11115);
and U11870 (N_11870,N_11122,N_10516);
and U11871 (N_11871,N_10799,N_10573);
or U11872 (N_11872,N_10758,N_10680);
or U11873 (N_11873,N_10828,N_11103);
nand U11874 (N_11874,N_10866,N_10402);
xnor U11875 (N_11875,N_10921,N_10825);
and U11876 (N_11876,N_10608,N_10977);
xnor U11877 (N_11877,N_10441,N_10780);
xnor U11878 (N_11878,N_10735,N_10595);
and U11879 (N_11879,N_10848,N_10779);
nor U11880 (N_11880,N_10916,N_10892);
and U11881 (N_11881,N_11182,N_11160);
xor U11882 (N_11882,N_10754,N_10653);
or U11883 (N_11883,N_10598,N_11061);
nand U11884 (N_11884,N_11039,N_10564);
and U11885 (N_11885,N_10905,N_10887);
or U11886 (N_11886,N_10651,N_10687);
nor U11887 (N_11887,N_10621,N_10420);
and U11888 (N_11888,N_10434,N_11174);
and U11889 (N_11889,N_10736,N_11177);
or U11890 (N_11890,N_10517,N_10421);
xor U11891 (N_11891,N_10524,N_10611);
xnor U11892 (N_11892,N_11053,N_10555);
and U11893 (N_11893,N_10667,N_10488);
nor U11894 (N_11894,N_11060,N_10506);
or U11895 (N_11895,N_10715,N_10719);
xnor U11896 (N_11896,N_10830,N_10467);
and U11897 (N_11897,N_11179,N_10462);
or U11898 (N_11898,N_10667,N_10844);
nand U11899 (N_11899,N_10486,N_10490);
xnor U11900 (N_11900,N_10616,N_10845);
and U11901 (N_11901,N_10951,N_11096);
and U11902 (N_11902,N_10701,N_11059);
xnor U11903 (N_11903,N_10410,N_10714);
xor U11904 (N_11904,N_10832,N_11165);
xor U11905 (N_11905,N_10627,N_11119);
or U11906 (N_11906,N_10437,N_10687);
or U11907 (N_11907,N_11051,N_10475);
xor U11908 (N_11908,N_10741,N_10863);
nand U11909 (N_11909,N_11037,N_10863);
nor U11910 (N_11910,N_11045,N_10448);
xor U11911 (N_11911,N_11075,N_11146);
or U11912 (N_11912,N_11046,N_11055);
nor U11913 (N_11913,N_10578,N_11105);
or U11914 (N_11914,N_11003,N_11105);
xnor U11915 (N_11915,N_10633,N_10491);
and U11916 (N_11916,N_11195,N_10774);
nor U11917 (N_11917,N_10860,N_11182);
or U11918 (N_11918,N_10558,N_10616);
nand U11919 (N_11919,N_10720,N_10965);
nand U11920 (N_11920,N_11085,N_10912);
nor U11921 (N_11921,N_10448,N_10570);
or U11922 (N_11922,N_11190,N_11103);
nor U11923 (N_11923,N_11182,N_11161);
nor U11924 (N_11924,N_10741,N_10588);
xnor U11925 (N_11925,N_10979,N_10994);
xor U11926 (N_11926,N_10502,N_10516);
and U11927 (N_11927,N_10588,N_10851);
xnor U11928 (N_11928,N_11108,N_10555);
xnor U11929 (N_11929,N_10797,N_11114);
or U11930 (N_11930,N_10796,N_10579);
nor U11931 (N_11931,N_11143,N_11186);
nand U11932 (N_11932,N_10723,N_10554);
nand U11933 (N_11933,N_11022,N_11159);
and U11934 (N_11934,N_10541,N_10559);
xor U11935 (N_11935,N_10460,N_10789);
xor U11936 (N_11936,N_10455,N_10590);
or U11937 (N_11937,N_10551,N_10463);
nor U11938 (N_11938,N_10447,N_10429);
nand U11939 (N_11939,N_10669,N_10997);
and U11940 (N_11940,N_10875,N_10669);
or U11941 (N_11941,N_10758,N_10464);
xor U11942 (N_11942,N_10819,N_10994);
or U11943 (N_11943,N_10498,N_10820);
nor U11944 (N_11944,N_11060,N_11152);
or U11945 (N_11945,N_11147,N_11085);
nand U11946 (N_11946,N_10622,N_11063);
nand U11947 (N_11947,N_10425,N_10894);
xor U11948 (N_11948,N_10651,N_10989);
nor U11949 (N_11949,N_10662,N_10793);
xor U11950 (N_11950,N_10615,N_10791);
xnor U11951 (N_11951,N_11059,N_10453);
nand U11952 (N_11952,N_11070,N_11107);
xor U11953 (N_11953,N_11085,N_11072);
and U11954 (N_11954,N_10665,N_11113);
xnor U11955 (N_11955,N_10499,N_10493);
xnor U11956 (N_11956,N_10757,N_10820);
or U11957 (N_11957,N_11081,N_10497);
and U11958 (N_11958,N_10737,N_10529);
and U11959 (N_11959,N_10486,N_10921);
nand U11960 (N_11960,N_10686,N_10931);
nand U11961 (N_11961,N_10826,N_10954);
nand U11962 (N_11962,N_11075,N_11188);
nor U11963 (N_11963,N_11027,N_10925);
nand U11964 (N_11964,N_11039,N_10601);
or U11965 (N_11965,N_11183,N_10831);
and U11966 (N_11966,N_10496,N_10414);
nand U11967 (N_11967,N_10499,N_10960);
xnor U11968 (N_11968,N_10450,N_10435);
nand U11969 (N_11969,N_10425,N_11071);
nand U11970 (N_11970,N_10438,N_10820);
xnor U11971 (N_11971,N_10599,N_10593);
nand U11972 (N_11972,N_11003,N_11074);
nand U11973 (N_11973,N_11194,N_11197);
nor U11974 (N_11974,N_11052,N_11101);
and U11975 (N_11975,N_11018,N_10976);
xor U11976 (N_11976,N_10796,N_10994);
xnor U11977 (N_11977,N_10741,N_10421);
or U11978 (N_11978,N_10761,N_10846);
or U11979 (N_11979,N_11088,N_11163);
xnor U11980 (N_11980,N_10437,N_10965);
or U11981 (N_11981,N_10635,N_10781);
and U11982 (N_11982,N_10710,N_11149);
and U11983 (N_11983,N_11040,N_11087);
and U11984 (N_11984,N_10419,N_10569);
nor U11985 (N_11985,N_11004,N_10691);
or U11986 (N_11986,N_10920,N_10526);
or U11987 (N_11987,N_10822,N_11198);
and U11988 (N_11988,N_10406,N_10598);
nor U11989 (N_11989,N_10414,N_11198);
or U11990 (N_11990,N_11052,N_10530);
xor U11991 (N_11991,N_10737,N_10943);
or U11992 (N_11992,N_10798,N_10974);
or U11993 (N_11993,N_10458,N_10869);
xor U11994 (N_11994,N_11179,N_11164);
nor U11995 (N_11995,N_10682,N_10500);
and U11996 (N_11996,N_11063,N_10932);
and U11997 (N_11997,N_10480,N_11067);
or U11998 (N_11998,N_10523,N_10837);
nor U11999 (N_11999,N_10612,N_10915);
xor U12000 (N_12000,N_11525,N_11930);
or U12001 (N_12001,N_11751,N_11615);
nand U12002 (N_12002,N_11748,N_11923);
nand U12003 (N_12003,N_11733,N_11261);
nand U12004 (N_12004,N_11864,N_11595);
xor U12005 (N_12005,N_11391,N_11554);
or U12006 (N_12006,N_11549,N_11862);
or U12007 (N_12007,N_11987,N_11760);
nand U12008 (N_12008,N_11435,N_11646);
and U12009 (N_12009,N_11517,N_11800);
nand U12010 (N_12010,N_11260,N_11334);
or U12011 (N_12011,N_11815,N_11750);
nand U12012 (N_12012,N_11632,N_11227);
nand U12013 (N_12013,N_11870,N_11390);
or U12014 (N_12014,N_11233,N_11617);
and U12015 (N_12015,N_11639,N_11972);
nor U12016 (N_12016,N_11292,N_11231);
xnor U12017 (N_12017,N_11397,N_11339);
xnor U12018 (N_12018,N_11963,N_11844);
nor U12019 (N_12019,N_11867,N_11997);
and U12020 (N_12020,N_11542,N_11993);
and U12021 (N_12021,N_11341,N_11457);
nand U12022 (N_12022,N_11907,N_11775);
and U12023 (N_12023,N_11740,N_11774);
and U12024 (N_12024,N_11711,N_11316);
or U12025 (N_12025,N_11762,N_11620);
or U12026 (N_12026,N_11494,N_11265);
nand U12027 (N_12027,N_11582,N_11786);
or U12028 (N_12028,N_11256,N_11636);
and U12029 (N_12029,N_11217,N_11888);
xor U12030 (N_12030,N_11376,N_11369);
xnor U12031 (N_12031,N_11805,N_11484);
and U12032 (N_12032,N_11213,N_11251);
nand U12033 (N_12033,N_11979,N_11361);
nand U12034 (N_12034,N_11311,N_11258);
nor U12035 (N_12035,N_11429,N_11881);
and U12036 (N_12036,N_11282,N_11845);
nand U12037 (N_12037,N_11756,N_11934);
nand U12038 (N_12038,N_11736,N_11202);
and U12039 (N_12039,N_11710,N_11546);
nand U12040 (N_12040,N_11876,N_11555);
nand U12041 (N_12041,N_11797,N_11619);
nor U12042 (N_12042,N_11692,N_11204);
xor U12043 (N_12043,N_11970,N_11528);
and U12044 (N_12044,N_11268,N_11591);
and U12045 (N_12045,N_11698,N_11966);
or U12046 (N_12046,N_11912,N_11510);
xnor U12047 (N_12047,N_11214,N_11421);
and U12048 (N_12048,N_11332,N_11655);
or U12049 (N_12049,N_11223,N_11602);
nand U12050 (N_12050,N_11627,N_11380);
nor U12051 (N_12051,N_11454,N_11401);
or U12052 (N_12052,N_11821,N_11838);
and U12053 (N_12053,N_11833,N_11685);
nor U12054 (N_12054,N_11415,N_11588);
and U12055 (N_12055,N_11779,N_11348);
and U12056 (N_12056,N_11765,N_11737);
nand U12057 (N_12057,N_11696,N_11960);
and U12058 (N_12058,N_11402,N_11942);
nor U12059 (N_12059,N_11741,N_11221);
nand U12060 (N_12060,N_11622,N_11264);
nand U12061 (N_12061,N_11439,N_11477);
or U12062 (N_12062,N_11472,N_11530);
nand U12063 (N_12063,N_11850,N_11953);
or U12064 (N_12064,N_11495,N_11467);
nor U12065 (N_12065,N_11579,N_11531);
xnor U12066 (N_12066,N_11988,N_11427);
nand U12067 (N_12067,N_11940,N_11755);
or U12068 (N_12068,N_11676,N_11455);
or U12069 (N_12069,N_11854,N_11360);
xor U12070 (N_12070,N_11485,N_11875);
nand U12071 (N_12071,N_11941,N_11442);
xnor U12072 (N_12072,N_11347,N_11395);
and U12073 (N_12073,N_11813,N_11929);
nand U12074 (N_12074,N_11447,N_11414);
xor U12075 (N_12075,N_11802,N_11728);
or U12076 (N_12076,N_11583,N_11419);
nor U12077 (N_12077,N_11434,N_11708);
xnor U12078 (N_12078,N_11892,N_11468);
nor U12079 (N_12079,N_11416,N_11474);
nand U12080 (N_12080,N_11503,N_11314);
xnor U12081 (N_12081,N_11852,N_11443);
nor U12082 (N_12082,N_11350,N_11654);
nor U12083 (N_12083,N_11811,N_11705);
nand U12084 (N_12084,N_11629,N_11535);
or U12085 (N_12085,N_11568,N_11232);
or U12086 (N_12086,N_11521,N_11983);
or U12087 (N_12087,N_11663,N_11487);
nor U12088 (N_12088,N_11566,N_11518);
and U12089 (N_12089,N_11482,N_11859);
nand U12090 (N_12090,N_11349,N_11460);
xnor U12091 (N_12091,N_11355,N_11865);
and U12092 (N_12092,N_11352,N_11263);
nor U12093 (N_12093,N_11767,N_11976);
and U12094 (N_12094,N_11319,N_11229);
and U12095 (N_12095,N_11897,N_11304);
and U12096 (N_12096,N_11374,N_11280);
nand U12097 (N_12097,N_11593,N_11734);
or U12098 (N_12098,N_11808,N_11643);
and U12099 (N_12099,N_11954,N_11522);
nor U12100 (N_12100,N_11863,N_11597);
or U12101 (N_12101,N_11883,N_11921);
or U12102 (N_12102,N_11458,N_11365);
nand U12103 (N_12103,N_11650,N_11656);
or U12104 (N_12104,N_11475,N_11237);
nor U12105 (N_12105,N_11289,N_11450);
and U12106 (N_12106,N_11604,N_11999);
or U12107 (N_12107,N_11882,N_11356);
and U12108 (N_12108,N_11569,N_11224);
nor U12109 (N_12109,N_11307,N_11746);
xor U12110 (N_12110,N_11991,N_11978);
nand U12111 (N_12111,N_11625,N_11818);
or U12112 (N_12112,N_11473,N_11255);
or U12113 (N_12113,N_11877,N_11562);
or U12114 (N_12114,N_11284,N_11210);
xor U12115 (N_12115,N_11842,N_11955);
nand U12116 (N_12116,N_11861,N_11520);
and U12117 (N_12117,N_11533,N_11299);
nor U12118 (N_12118,N_11343,N_11290);
and U12119 (N_12119,N_11680,N_11441);
and U12120 (N_12120,N_11278,N_11652);
nand U12121 (N_12121,N_11285,N_11895);
nand U12122 (N_12122,N_11834,N_11302);
nor U12123 (N_12123,N_11889,N_11723);
or U12124 (N_12124,N_11313,N_11621);
nand U12125 (N_12125,N_11500,N_11668);
nor U12126 (N_12126,N_11684,N_11884);
nor U12127 (N_12127,N_11513,N_11325);
nand U12128 (N_12128,N_11644,N_11386);
or U12129 (N_12129,N_11287,N_11252);
xor U12130 (N_12130,N_11836,N_11981);
xnor U12131 (N_12131,N_11417,N_11234);
and U12132 (N_12132,N_11623,N_11523);
xnor U12133 (N_12133,N_11399,N_11968);
nor U12134 (N_12134,N_11911,N_11516);
nand U12135 (N_12135,N_11471,N_11727);
nand U12136 (N_12136,N_11248,N_11215);
xor U12137 (N_12137,N_11453,N_11274);
nand U12138 (N_12138,N_11939,N_11891);
nor U12139 (N_12139,N_11624,N_11661);
xnor U12140 (N_12140,N_11295,N_11470);
nand U12141 (N_12141,N_11456,N_11855);
nand U12142 (N_12142,N_11761,N_11943);
and U12143 (N_12143,N_11239,N_11605);
nor U12144 (N_12144,N_11216,N_11328);
and U12145 (N_12145,N_11373,N_11782);
nor U12146 (N_12146,N_11784,N_11406);
xor U12147 (N_12147,N_11823,N_11670);
or U12148 (N_12148,N_11409,N_11469);
nor U12149 (N_12149,N_11245,N_11275);
nor U12150 (N_12150,N_11411,N_11200);
nand U12151 (N_12151,N_11964,N_11683);
nor U12152 (N_12152,N_11686,N_11799);
and U12153 (N_12153,N_11587,N_11780);
xor U12154 (N_12154,N_11682,N_11671);
and U12155 (N_12155,N_11766,N_11336);
xor U12156 (N_12156,N_11543,N_11754);
and U12157 (N_12157,N_11388,N_11757);
nor U12158 (N_12158,N_11658,N_11504);
xnor U12159 (N_12159,N_11449,N_11281);
or U12160 (N_12160,N_11609,N_11707);
nor U12161 (N_12161,N_11956,N_11747);
and U12162 (N_12162,N_11207,N_11405);
nand U12163 (N_12163,N_11944,N_11916);
xnor U12164 (N_12164,N_11331,N_11666);
and U12165 (N_12165,N_11371,N_11791);
xor U12166 (N_12166,N_11556,N_11896);
xnor U12167 (N_12167,N_11222,N_11344);
xnor U12168 (N_12168,N_11236,N_11828);
xnor U12169 (N_12169,N_11545,N_11598);
nand U12170 (N_12170,N_11969,N_11947);
xor U12171 (N_12171,N_11228,N_11630);
xnor U12172 (N_12172,N_11716,N_11957);
xor U12173 (N_12173,N_11557,N_11835);
and U12174 (N_12174,N_11440,N_11327);
xor U12175 (N_12175,N_11631,N_11871);
and U12176 (N_12176,N_11948,N_11436);
nand U12177 (N_12177,N_11857,N_11493);
or U12178 (N_12178,N_11585,N_11269);
and U12179 (N_12179,N_11459,N_11403);
nor U12180 (N_12180,N_11846,N_11980);
nor U12181 (N_12181,N_11806,N_11490);
nor U12182 (N_12182,N_11667,N_11589);
or U12183 (N_12183,N_11770,N_11465);
xnor U12184 (N_12184,N_11301,N_11410);
nand U12185 (N_12185,N_11580,N_11553);
nand U12186 (N_12186,N_11206,N_11514);
or U12187 (N_12187,N_11426,N_11744);
and U12188 (N_12188,N_11719,N_11389);
nand U12189 (N_12189,N_11358,N_11959);
xor U12190 (N_12190,N_11574,N_11242);
and U12191 (N_12191,N_11437,N_11218);
xnor U12192 (N_12192,N_11985,N_11998);
and U12193 (N_12193,N_11481,N_11425);
xnor U12194 (N_12194,N_11669,N_11648);
or U12195 (N_12195,N_11396,N_11576);
and U12196 (N_12196,N_11428,N_11700);
xor U12197 (N_12197,N_11927,N_11407);
xor U12198 (N_12198,N_11653,N_11502);
nor U12199 (N_12199,N_11594,N_11938);
and U12200 (N_12200,N_11965,N_11253);
nand U12201 (N_12201,N_11759,N_11694);
nor U12202 (N_12202,N_11611,N_11730);
nor U12203 (N_12203,N_11789,N_11208);
or U12204 (N_12204,N_11312,N_11359);
nand U12205 (N_12205,N_11872,N_11946);
nor U12206 (N_12206,N_11873,N_11323);
xor U12207 (N_12207,N_11919,N_11558);
xnor U12208 (N_12208,N_11902,N_11527);
nor U12209 (N_12209,N_11431,N_11438);
or U12210 (N_12210,N_11788,N_11853);
nand U12211 (N_12211,N_11795,N_11259);
nor U12212 (N_12212,N_11749,N_11515);
nand U12213 (N_12213,N_11219,N_11420);
nor U12214 (N_12214,N_11778,N_11958);
nand U12215 (N_12215,N_11303,N_11660);
xor U12216 (N_12216,N_11793,N_11363);
and U12217 (N_12217,N_11404,N_11628);
nand U12218 (N_12218,N_11662,N_11909);
xnor U12219 (N_12219,N_11635,N_11771);
xnor U12220 (N_12220,N_11908,N_11507);
nand U12221 (N_12221,N_11308,N_11392);
nand U12222 (N_12222,N_11717,N_11509);
or U12223 (N_12223,N_11330,N_11952);
nand U12224 (N_12224,N_11989,N_11362);
or U12225 (N_12225,N_11364,N_11476);
xnor U12226 (N_12226,N_11764,N_11903);
nand U12227 (N_12227,N_11578,N_11320);
xnor U12228 (N_12228,N_11758,N_11715);
nor U12229 (N_12229,N_11353,N_11743);
or U12230 (N_12230,N_11878,N_11932);
nand U12231 (N_12231,N_11483,N_11918);
nand U12232 (N_12232,N_11905,N_11984);
and U12233 (N_12233,N_11840,N_11310);
and U12234 (N_12234,N_11928,N_11899);
xnor U12235 (N_12235,N_11935,N_11291);
or U12236 (N_12236,N_11581,N_11422);
and U12237 (N_12237,N_11492,N_11915);
and U12238 (N_12238,N_11967,N_11701);
nand U12239 (N_12239,N_11922,N_11277);
and U12240 (N_12240,N_11614,N_11512);
or U12241 (N_12241,N_11240,N_11423);
xor U12242 (N_12242,N_11276,N_11209);
xnor U12243 (N_12243,N_11709,N_11616);
nand U12244 (N_12244,N_11400,N_11641);
nand U12245 (N_12245,N_11296,N_11537);
nor U12246 (N_12246,N_11613,N_11849);
xnor U12247 (N_12247,N_11917,N_11739);
nand U12248 (N_12248,N_11488,N_11702);
and U12249 (N_12249,N_11445,N_11357);
xor U12250 (N_12250,N_11866,N_11982);
xor U12251 (N_12251,N_11212,N_11819);
and U12252 (N_12252,N_11830,N_11977);
or U12253 (N_12253,N_11571,N_11394);
nand U12254 (N_12254,N_11801,N_11642);
nor U12255 (N_12255,N_11412,N_11825);
nor U12256 (N_12256,N_11856,N_11713);
nand U12257 (N_12257,N_11637,N_11626);
xor U12258 (N_12258,N_11480,N_11270);
and U12259 (N_12259,N_11590,N_11781);
nor U12260 (N_12260,N_11726,N_11345);
nor U12261 (N_12261,N_11305,N_11651);
xor U12262 (N_12262,N_11393,N_11326);
nand U12263 (N_12263,N_11790,N_11783);
xor U12264 (N_12264,N_11550,N_11796);
and U12265 (N_12265,N_11563,N_11491);
nand U12266 (N_12266,N_11742,N_11203);
nor U12267 (N_12267,N_11890,N_11785);
nor U12268 (N_12268,N_11324,N_11674);
and U12269 (N_12269,N_11368,N_11634);
nand U12270 (N_12270,N_11600,N_11689);
nand U12271 (N_12271,N_11526,N_11945);
xor U12272 (N_12272,N_11949,N_11565);
nand U12273 (N_12273,N_11286,N_11794);
xor U12274 (N_12274,N_11432,N_11586);
nor U12275 (N_12275,N_11822,N_11894);
nor U12276 (N_12276,N_11317,N_11424);
xor U12277 (N_12277,N_11974,N_11552);
or U12278 (N_12278,N_11990,N_11267);
and U12279 (N_12279,N_11986,N_11868);
xnor U12280 (N_12280,N_11367,N_11886);
nor U12281 (N_12281,N_11448,N_11647);
nand U12282 (N_12282,N_11241,N_11596);
nor U12283 (N_12283,N_11321,N_11847);
or U12284 (N_12284,N_11486,N_11874);
or U12285 (N_12285,N_11592,N_11601);
or U12286 (N_12286,N_11675,N_11645);
or U12287 (N_12287,N_11254,N_11366);
xnor U12288 (N_12288,N_11372,N_11599);
xnor U12289 (N_12289,N_11539,N_11567);
nor U12290 (N_12290,N_11649,N_11379);
nor U12291 (N_12291,N_11848,N_11548);
or U12292 (N_12292,N_11288,N_11540);
nor U12293 (N_12293,N_11768,N_11377);
nor U12294 (N_12294,N_11387,N_11724);
nor U12295 (N_12295,N_11201,N_11817);
xor U12296 (N_12296,N_11272,N_11547);
nand U12297 (N_12297,N_11933,N_11704);
or U12298 (N_12298,N_11826,N_11688);
xnor U12299 (N_12299,N_11496,N_11773);
xor U12300 (N_12300,N_11519,N_11633);
nor U12301 (N_12301,N_11329,N_11497);
nand U12302 (N_12302,N_11887,N_11924);
nor U12303 (N_12303,N_11511,N_11839);
nand U12304 (N_12304,N_11293,N_11235);
xnor U12305 (N_12305,N_11505,N_11489);
nand U12306 (N_12306,N_11451,N_11745);
xnor U12307 (N_12307,N_11973,N_11936);
nand U12308 (N_12308,N_11225,N_11570);
nor U12309 (N_12309,N_11677,N_11430);
nor U12310 (N_12310,N_11478,N_11732);
xnor U12311 (N_12311,N_11678,N_11992);
xnor U12312 (N_12312,N_11573,N_11809);
or U12313 (N_12313,N_11792,N_11382);
and U12314 (N_12314,N_11753,N_11712);
and U12315 (N_12315,N_11257,N_11333);
nand U12316 (N_12316,N_11735,N_11342);
and U12317 (N_12317,N_11383,N_11309);
xor U12318 (N_12318,N_11338,N_11532);
or U12319 (N_12319,N_11381,N_11378);
and U12320 (N_12320,N_11971,N_11752);
and U12321 (N_12321,N_11879,N_11860);
nor U12322 (N_12322,N_11575,N_11577);
nand U12323 (N_12323,N_11603,N_11787);
xor U12324 (N_12324,N_11408,N_11725);
or U12325 (N_12325,N_11433,N_11205);
or U12326 (N_12326,N_11606,N_11807);
nor U12327 (N_12327,N_11300,N_11925);
xnor U12328 (N_12328,N_11306,N_11534);
xnor U12329 (N_12329,N_11699,N_11538);
nor U12330 (N_12330,N_11695,N_11370);
xor U12331 (N_12331,N_11832,N_11322);
nor U12332 (N_12332,N_11536,N_11803);
xor U12333 (N_12333,N_11893,N_11464);
nand U12334 (N_12334,N_11297,N_11901);
xor U12335 (N_12335,N_11837,N_11814);
nand U12336 (N_12336,N_11679,N_11729);
or U12337 (N_12337,N_11279,N_11950);
and U12338 (N_12338,N_11230,N_11452);
and U12339 (N_12339,N_11687,N_11243);
nand U12340 (N_12340,N_11226,N_11910);
or U12341 (N_12341,N_11346,N_11384);
and U12342 (N_12342,N_11858,N_11244);
or U12343 (N_12343,N_11385,N_11931);
and U12344 (N_12344,N_11463,N_11560);
or U12345 (N_12345,N_11610,N_11271);
xor U12346 (N_12346,N_11498,N_11898);
nor U12347 (N_12347,N_11996,N_11697);
nor U12348 (N_12348,N_11851,N_11354);
nor U12349 (N_12349,N_11584,N_11506);
and U12350 (N_12350,N_11718,N_11337);
nand U12351 (N_12351,N_11841,N_11827);
or U12352 (N_12352,N_11211,N_11398);
nor U12353 (N_12353,N_11246,N_11559);
nor U12354 (N_12354,N_11900,N_11444);
xnor U12355 (N_12355,N_11561,N_11816);
nor U12356 (N_12356,N_11479,N_11812);
xnor U12357 (N_12357,N_11722,N_11659);
or U12358 (N_12358,N_11564,N_11220);
nand U12359 (N_12359,N_11665,N_11769);
nand U12360 (N_12360,N_11951,N_11640);
or U12361 (N_12361,N_11681,N_11975);
or U12362 (N_12362,N_11529,N_11693);
nor U12363 (N_12363,N_11994,N_11466);
nor U12364 (N_12364,N_11618,N_11283);
and U12365 (N_12365,N_11720,N_11294);
nor U12366 (N_12366,N_11906,N_11721);
nand U12367 (N_12367,N_11691,N_11706);
nand U12368 (N_12368,N_11880,N_11829);
nor U12369 (N_12369,N_11413,N_11572);
nand U12370 (N_12370,N_11914,N_11501);
or U12371 (N_12371,N_11607,N_11315);
or U12372 (N_12372,N_11731,N_11962);
or U12373 (N_12373,N_11843,N_11926);
xor U12374 (N_12374,N_11738,N_11820);
nor U12375 (N_12375,N_11714,N_11508);
or U12376 (N_12376,N_11810,N_11351);
xor U12377 (N_12377,N_11541,N_11961);
xnor U12378 (N_12378,N_11247,N_11831);
xnor U12379 (N_12379,N_11551,N_11995);
and U12380 (N_12380,N_11340,N_11544);
and U12381 (N_12381,N_11776,N_11824);
and U12382 (N_12382,N_11920,N_11804);
and U12383 (N_12383,N_11446,N_11262);
and U12384 (N_12384,N_11904,N_11249);
and U12385 (N_12385,N_11612,N_11657);
nand U12386 (N_12386,N_11869,N_11703);
nor U12387 (N_12387,N_11250,N_11937);
xnor U12388 (N_12388,N_11638,N_11462);
xor U12389 (N_12389,N_11273,N_11266);
xor U12390 (N_12390,N_11690,N_11608);
and U12391 (N_12391,N_11763,N_11913);
or U12392 (N_12392,N_11499,N_11375);
and U12393 (N_12393,N_11461,N_11777);
nand U12394 (N_12394,N_11238,N_11418);
nor U12395 (N_12395,N_11772,N_11798);
and U12396 (N_12396,N_11524,N_11885);
xor U12397 (N_12397,N_11673,N_11672);
and U12398 (N_12398,N_11664,N_11335);
nor U12399 (N_12399,N_11298,N_11318);
nor U12400 (N_12400,N_11657,N_11925);
xor U12401 (N_12401,N_11439,N_11429);
nor U12402 (N_12402,N_11693,N_11883);
and U12403 (N_12403,N_11262,N_11835);
or U12404 (N_12404,N_11966,N_11596);
nand U12405 (N_12405,N_11597,N_11630);
or U12406 (N_12406,N_11980,N_11652);
nand U12407 (N_12407,N_11503,N_11270);
and U12408 (N_12408,N_11558,N_11357);
or U12409 (N_12409,N_11455,N_11721);
and U12410 (N_12410,N_11878,N_11463);
nor U12411 (N_12411,N_11220,N_11390);
and U12412 (N_12412,N_11455,N_11530);
nand U12413 (N_12413,N_11760,N_11279);
and U12414 (N_12414,N_11501,N_11207);
nand U12415 (N_12415,N_11954,N_11681);
or U12416 (N_12416,N_11657,N_11493);
xor U12417 (N_12417,N_11954,N_11281);
or U12418 (N_12418,N_11466,N_11744);
nor U12419 (N_12419,N_11704,N_11971);
nor U12420 (N_12420,N_11390,N_11788);
nand U12421 (N_12421,N_11756,N_11457);
nand U12422 (N_12422,N_11534,N_11840);
nor U12423 (N_12423,N_11652,N_11435);
nand U12424 (N_12424,N_11985,N_11297);
and U12425 (N_12425,N_11623,N_11719);
xor U12426 (N_12426,N_11631,N_11789);
nand U12427 (N_12427,N_11450,N_11759);
xor U12428 (N_12428,N_11206,N_11576);
or U12429 (N_12429,N_11666,N_11569);
nand U12430 (N_12430,N_11843,N_11906);
and U12431 (N_12431,N_11789,N_11861);
xor U12432 (N_12432,N_11236,N_11393);
and U12433 (N_12433,N_11277,N_11608);
or U12434 (N_12434,N_11679,N_11567);
and U12435 (N_12435,N_11372,N_11864);
nor U12436 (N_12436,N_11395,N_11704);
xor U12437 (N_12437,N_11974,N_11505);
xor U12438 (N_12438,N_11378,N_11809);
nor U12439 (N_12439,N_11671,N_11703);
nand U12440 (N_12440,N_11799,N_11612);
nand U12441 (N_12441,N_11798,N_11895);
xor U12442 (N_12442,N_11889,N_11608);
or U12443 (N_12443,N_11616,N_11225);
nor U12444 (N_12444,N_11648,N_11204);
nor U12445 (N_12445,N_11929,N_11669);
and U12446 (N_12446,N_11695,N_11907);
xnor U12447 (N_12447,N_11710,N_11847);
or U12448 (N_12448,N_11384,N_11800);
xnor U12449 (N_12449,N_11947,N_11925);
nand U12450 (N_12450,N_11946,N_11758);
nor U12451 (N_12451,N_11300,N_11674);
xnor U12452 (N_12452,N_11524,N_11619);
xor U12453 (N_12453,N_11703,N_11994);
nor U12454 (N_12454,N_11447,N_11928);
or U12455 (N_12455,N_11880,N_11247);
and U12456 (N_12456,N_11371,N_11206);
and U12457 (N_12457,N_11531,N_11353);
nand U12458 (N_12458,N_11461,N_11595);
nand U12459 (N_12459,N_11646,N_11492);
nor U12460 (N_12460,N_11630,N_11522);
nand U12461 (N_12461,N_11563,N_11667);
and U12462 (N_12462,N_11941,N_11994);
nand U12463 (N_12463,N_11970,N_11825);
nor U12464 (N_12464,N_11999,N_11948);
nand U12465 (N_12465,N_11882,N_11573);
or U12466 (N_12466,N_11605,N_11827);
xnor U12467 (N_12467,N_11466,N_11445);
nand U12468 (N_12468,N_11713,N_11547);
nand U12469 (N_12469,N_11359,N_11478);
xnor U12470 (N_12470,N_11660,N_11632);
and U12471 (N_12471,N_11358,N_11629);
nand U12472 (N_12472,N_11842,N_11683);
and U12473 (N_12473,N_11495,N_11958);
nor U12474 (N_12474,N_11380,N_11782);
and U12475 (N_12475,N_11886,N_11666);
and U12476 (N_12476,N_11694,N_11469);
nor U12477 (N_12477,N_11705,N_11953);
xor U12478 (N_12478,N_11888,N_11673);
nor U12479 (N_12479,N_11700,N_11682);
or U12480 (N_12480,N_11503,N_11887);
xor U12481 (N_12481,N_11531,N_11483);
and U12482 (N_12482,N_11482,N_11902);
xor U12483 (N_12483,N_11704,N_11826);
nand U12484 (N_12484,N_11683,N_11330);
xor U12485 (N_12485,N_11548,N_11379);
or U12486 (N_12486,N_11255,N_11380);
and U12487 (N_12487,N_11846,N_11735);
nor U12488 (N_12488,N_11209,N_11285);
nor U12489 (N_12489,N_11430,N_11322);
and U12490 (N_12490,N_11891,N_11547);
nor U12491 (N_12491,N_11210,N_11778);
or U12492 (N_12492,N_11448,N_11447);
nor U12493 (N_12493,N_11772,N_11318);
xnor U12494 (N_12494,N_11890,N_11983);
nand U12495 (N_12495,N_11448,N_11711);
nor U12496 (N_12496,N_11291,N_11410);
xor U12497 (N_12497,N_11480,N_11806);
or U12498 (N_12498,N_11641,N_11452);
nor U12499 (N_12499,N_11351,N_11224);
or U12500 (N_12500,N_11619,N_11842);
nor U12501 (N_12501,N_11533,N_11202);
nand U12502 (N_12502,N_11526,N_11795);
or U12503 (N_12503,N_11899,N_11208);
or U12504 (N_12504,N_11822,N_11348);
nand U12505 (N_12505,N_11628,N_11396);
or U12506 (N_12506,N_11698,N_11896);
and U12507 (N_12507,N_11859,N_11492);
nand U12508 (N_12508,N_11970,N_11729);
xor U12509 (N_12509,N_11258,N_11894);
nand U12510 (N_12510,N_11774,N_11891);
nand U12511 (N_12511,N_11409,N_11696);
or U12512 (N_12512,N_11437,N_11558);
nor U12513 (N_12513,N_11330,N_11720);
and U12514 (N_12514,N_11705,N_11463);
and U12515 (N_12515,N_11317,N_11598);
xor U12516 (N_12516,N_11345,N_11866);
nor U12517 (N_12517,N_11451,N_11237);
and U12518 (N_12518,N_11699,N_11774);
and U12519 (N_12519,N_11412,N_11213);
nor U12520 (N_12520,N_11811,N_11709);
or U12521 (N_12521,N_11770,N_11823);
nor U12522 (N_12522,N_11451,N_11309);
nand U12523 (N_12523,N_11596,N_11741);
nor U12524 (N_12524,N_11660,N_11595);
nor U12525 (N_12525,N_11638,N_11543);
nand U12526 (N_12526,N_11489,N_11930);
and U12527 (N_12527,N_11951,N_11645);
nand U12528 (N_12528,N_11717,N_11349);
and U12529 (N_12529,N_11623,N_11983);
nor U12530 (N_12530,N_11253,N_11202);
or U12531 (N_12531,N_11375,N_11240);
xor U12532 (N_12532,N_11862,N_11795);
xnor U12533 (N_12533,N_11381,N_11384);
and U12534 (N_12534,N_11540,N_11685);
nor U12535 (N_12535,N_11562,N_11869);
nand U12536 (N_12536,N_11629,N_11910);
nor U12537 (N_12537,N_11484,N_11449);
xnor U12538 (N_12538,N_11693,N_11918);
xnor U12539 (N_12539,N_11261,N_11561);
and U12540 (N_12540,N_11951,N_11564);
xor U12541 (N_12541,N_11440,N_11511);
xnor U12542 (N_12542,N_11578,N_11361);
and U12543 (N_12543,N_11851,N_11255);
or U12544 (N_12544,N_11760,N_11257);
and U12545 (N_12545,N_11785,N_11665);
xnor U12546 (N_12546,N_11880,N_11544);
nand U12547 (N_12547,N_11391,N_11614);
and U12548 (N_12548,N_11556,N_11541);
xnor U12549 (N_12549,N_11414,N_11743);
nand U12550 (N_12550,N_11812,N_11893);
xnor U12551 (N_12551,N_11998,N_11321);
nor U12552 (N_12552,N_11573,N_11353);
or U12553 (N_12553,N_11295,N_11469);
and U12554 (N_12554,N_11335,N_11712);
nor U12555 (N_12555,N_11539,N_11707);
nor U12556 (N_12556,N_11264,N_11279);
xnor U12557 (N_12557,N_11578,N_11257);
nor U12558 (N_12558,N_11295,N_11797);
and U12559 (N_12559,N_11262,N_11577);
and U12560 (N_12560,N_11635,N_11878);
or U12561 (N_12561,N_11287,N_11302);
and U12562 (N_12562,N_11572,N_11775);
xnor U12563 (N_12563,N_11302,N_11731);
or U12564 (N_12564,N_11665,N_11458);
nand U12565 (N_12565,N_11680,N_11848);
xnor U12566 (N_12566,N_11995,N_11473);
nor U12567 (N_12567,N_11905,N_11664);
and U12568 (N_12568,N_11928,N_11313);
or U12569 (N_12569,N_11967,N_11642);
or U12570 (N_12570,N_11475,N_11913);
and U12571 (N_12571,N_11539,N_11694);
xnor U12572 (N_12572,N_11823,N_11515);
nand U12573 (N_12573,N_11480,N_11344);
or U12574 (N_12574,N_11678,N_11857);
nand U12575 (N_12575,N_11700,N_11295);
and U12576 (N_12576,N_11247,N_11609);
nor U12577 (N_12577,N_11311,N_11757);
or U12578 (N_12578,N_11972,N_11277);
nand U12579 (N_12579,N_11372,N_11456);
nand U12580 (N_12580,N_11229,N_11939);
xnor U12581 (N_12581,N_11241,N_11641);
and U12582 (N_12582,N_11826,N_11230);
and U12583 (N_12583,N_11910,N_11874);
xnor U12584 (N_12584,N_11930,N_11377);
nor U12585 (N_12585,N_11258,N_11340);
nand U12586 (N_12586,N_11820,N_11846);
nand U12587 (N_12587,N_11558,N_11596);
xor U12588 (N_12588,N_11700,N_11602);
or U12589 (N_12589,N_11930,N_11295);
xor U12590 (N_12590,N_11777,N_11990);
or U12591 (N_12591,N_11489,N_11596);
xor U12592 (N_12592,N_11651,N_11792);
and U12593 (N_12593,N_11851,N_11425);
and U12594 (N_12594,N_11711,N_11737);
nor U12595 (N_12595,N_11284,N_11389);
nand U12596 (N_12596,N_11531,N_11303);
nor U12597 (N_12597,N_11936,N_11703);
xnor U12598 (N_12598,N_11584,N_11485);
nand U12599 (N_12599,N_11916,N_11397);
or U12600 (N_12600,N_11841,N_11759);
xor U12601 (N_12601,N_11522,N_11246);
xnor U12602 (N_12602,N_11604,N_11488);
xnor U12603 (N_12603,N_11940,N_11746);
and U12604 (N_12604,N_11652,N_11868);
nor U12605 (N_12605,N_11465,N_11208);
nor U12606 (N_12606,N_11764,N_11582);
and U12607 (N_12607,N_11384,N_11524);
xnor U12608 (N_12608,N_11356,N_11929);
nor U12609 (N_12609,N_11223,N_11724);
nor U12610 (N_12610,N_11314,N_11688);
nand U12611 (N_12611,N_11230,N_11674);
nand U12612 (N_12612,N_11894,N_11513);
and U12613 (N_12613,N_11227,N_11395);
nor U12614 (N_12614,N_11931,N_11532);
and U12615 (N_12615,N_11821,N_11293);
xor U12616 (N_12616,N_11998,N_11917);
and U12617 (N_12617,N_11576,N_11957);
nand U12618 (N_12618,N_11561,N_11372);
and U12619 (N_12619,N_11433,N_11430);
xnor U12620 (N_12620,N_11291,N_11791);
or U12621 (N_12621,N_11218,N_11390);
nor U12622 (N_12622,N_11520,N_11983);
xnor U12623 (N_12623,N_11800,N_11438);
nand U12624 (N_12624,N_11448,N_11436);
nand U12625 (N_12625,N_11592,N_11565);
or U12626 (N_12626,N_11548,N_11459);
nor U12627 (N_12627,N_11945,N_11886);
or U12628 (N_12628,N_11473,N_11354);
xor U12629 (N_12629,N_11385,N_11823);
nand U12630 (N_12630,N_11673,N_11948);
xnor U12631 (N_12631,N_11470,N_11675);
xor U12632 (N_12632,N_11348,N_11298);
nand U12633 (N_12633,N_11830,N_11337);
or U12634 (N_12634,N_11740,N_11823);
or U12635 (N_12635,N_11949,N_11795);
nor U12636 (N_12636,N_11670,N_11286);
and U12637 (N_12637,N_11361,N_11686);
xor U12638 (N_12638,N_11781,N_11389);
and U12639 (N_12639,N_11237,N_11626);
and U12640 (N_12640,N_11906,N_11218);
nor U12641 (N_12641,N_11301,N_11395);
nand U12642 (N_12642,N_11950,N_11484);
nand U12643 (N_12643,N_11968,N_11844);
and U12644 (N_12644,N_11925,N_11988);
and U12645 (N_12645,N_11853,N_11400);
nand U12646 (N_12646,N_11957,N_11502);
nor U12647 (N_12647,N_11697,N_11688);
or U12648 (N_12648,N_11659,N_11312);
or U12649 (N_12649,N_11759,N_11634);
or U12650 (N_12650,N_11384,N_11242);
and U12651 (N_12651,N_11825,N_11551);
xnor U12652 (N_12652,N_11635,N_11952);
xnor U12653 (N_12653,N_11554,N_11537);
or U12654 (N_12654,N_11934,N_11889);
xnor U12655 (N_12655,N_11213,N_11222);
nand U12656 (N_12656,N_11761,N_11717);
nand U12657 (N_12657,N_11477,N_11214);
nand U12658 (N_12658,N_11608,N_11804);
nand U12659 (N_12659,N_11885,N_11741);
and U12660 (N_12660,N_11880,N_11696);
or U12661 (N_12661,N_11301,N_11627);
or U12662 (N_12662,N_11219,N_11538);
xor U12663 (N_12663,N_11460,N_11820);
and U12664 (N_12664,N_11366,N_11320);
and U12665 (N_12665,N_11983,N_11845);
nor U12666 (N_12666,N_11576,N_11548);
and U12667 (N_12667,N_11792,N_11761);
nand U12668 (N_12668,N_11902,N_11298);
xor U12669 (N_12669,N_11763,N_11973);
or U12670 (N_12670,N_11421,N_11791);
xor U12671 (N_12671,N_11542,N_11517);
xor U12672 (N_12672,N_11929,N_11855);
and U12673 (N_12673,N_11486,N_11557);
nand U12674 (N_12674,N_11760,N_11974);
and U12675 (N_12675,N_11667,N_11397);
or U12676 (N_12676,N_11532,N_11747);
nand U12677 (N_12677,N_11713,N_11255);
xnor U12678 (N_12678,N_11895,N_11254);
nor U12679 (N_12679,N_11205,N_11574);
nand U12680 (N_12680,N_11670,N_11803);
or U12681 (N_12681,N_11286,N_11328);
nor U12682 (N_12682,N_11960,N_11272);
or U12683 (N_12683,N_11958,N_11353);
nor U12684 (N_12684,N_11795,N_11460);
nor U12685 (N_12685,N_11826,N_11763);
and U12686 (N_12686,N_11460,N_11410);
or U12687 (N_12687,N_11952,N_11725);
nand U12688 (N_12688,N_11517,N_11985);
nand U12689 (N_12689,N_11282,N_11527);
or U12690 (N_12690,N_11977,N_11276);
nor U12691 (N_12691,N_11383,N_11910);
or U12692 (N_12692,N_11280,N_11254);
nand U12693 (N_12693,N_11407,N_11449);
xnor U12694 (N_12694,N_11317,N_11531);
nor U12695 (N_12695,N_11496,N_11742);
xnor U12696 (N_12696,N_11317,N_11405);
nor U12697 (N_12697,N_11410,N_11933);
or U12698 (N_12698,N_11275,N_11260);
nand U12699 (N_12699,N_11303,N_11240);
nor U12700 (N_12700,N_11325,N_11752);
xnor U12701 (N_12701,N_11736,N_11726);
and U12702 (N_12702,N_11952,N_11236);
or U12703 (N_12703,N_11413,N_11524);
xor U12704 (N_12704,N_11860,N_11700);
and U12705 (N_12705,N_11304,N_11994);
nor U12706 (N_12706,N_11515,N_11396);
and U12707 (N_12707,N_11576,N_11861);
and U12708 (N_12708,N_11501,N_11489);
nand U12709 (N_12709,N_11714,N_11312);
nand U12710 (N_12710,N_11886,N_11833);
nand U12711 (N_12711,N_11743,N_11592);
nand U12712 (N_12712,N_11467,N_11723);
and U12713 (N_12713,N_11367,N_11323);
or U12714 (N_12714,N_11485,N_11264);
nor U12715 (N_12715,N_11246,N_11411);
and U12716 (N_12716,N_11236,N_11618);
xnor U12717 (N_12717,N_11875,N_11829);
or U12718 (N_12718,N_11553,N_11779);
and U12719 (N_12719,N_11872,N_11997);
xnor U12720 (N_12720,N_11801,N_11808);
and U12721 (N_12721,N_11590,N_11685);
nor U12722 (N_12722,N_11507,N_11994);
nor U12723 (N_12723,N_11844,N_11235);
nand U12724 (N_12724,N_11957,N_11821);
nand U12725 (N_12725,N_11925,N_11297);
xor U12726 (N_12726,N_11644,N_11855);
and U12727 (N_12727,N_11365,N_11338);
or U12728 (N_12728,N_11728,N_11933);
or U12729 (N_12729,N_11546,N_11467);
nor U12730 (N_12730,N_11761,N_11569);
and U12731 (N_12731,N_11380,N_11899);
or U12732 (N_12732,N_11964,N_11958);
or U12733 (N_12733,N_11620,N_11497);
xor U12734 (N_12734,N_11298,N_11243);
and U12735 (N_12735,N_11570,N_11858);
nor U12736 (N_12736,N_11297,N_11993);
nand U12737 (N_12737,N_11605,N_11832);
nor U12738 (N_12738,N_11852,N_11601);
nor U12739 (N_12739,N_11344,N_11378);
xnor U12740 (N_12740,N_11569,N_11360);
and U12741 (N_12741,N_11571,N_11748);
xnor U12742 (N_12742,N_11672,N_11421);
nand U12743 (N_12743,N_11822,N_11957);
xnor U12744 (N_12744,N_11769,N_11544);
and U12745 (N_12745,N_11233,N_11262);
nand U12746 (N_12746,N_11562,N_11542);
nor U12747 (N_12747,N_11902,N_11261);
or U12748 (N_12748,N_11517,N_11693);
nor U12749 (N_12749,N_11225,N_11889);
and U12750 (N_12750,N_11779,N_11962);
xnor U12751 (N_12751,N_11689,N_11375);
nor U12752 (N_12752,N_11849,N_11552);
xor U12753 (N_12753,N_11561,N_11736);
xor U12754 (N_12754,N_11926,N_11999);
or U12755 (N_12755,N_11543,N_11255);
and U12756 (N_12756,N_11854,N_11265);
and U12757 (N_12757,N_11246,N_11803);
xor U12758 (N_12758,N_11853,N_11898);
nand U12759 (N_12759,N_11449,N_11770);
xnor U12760 (N_12760,N_11536,N_11674);
or U12761 (N_12761,N_11280,N_11821);
and U12762 (N_12762,N_11946,N_11608);
or U12763 (N_12763,N_11605,N_11563);
nor U12764 (N_12764,N_11811,N_11903);
nor U12765 (N_12765,N_11928,N_11901);
xnor U12766 (N_12766,N_11455,N_11610);
nor U12767 (N_12767,N_11934,N_11826);
or U12768 (N_12768,N_11569,N_11517);
nand U12769 (N_12769,N_11838,N_11893);
or U12770 (N_12770,N_11477,N_11433);
and U12771 (N_12771,N_11296,N_11661);
xnor U12772 (N_12772,N_11873,N_11298);
nor U12773 (N_12773,N_11240,N_11931);
nand U12774 (N_12774,N_11478,N_11407);
nor U12775 (N_12775,N_11436,N_11571);
and U12776 (N_12776,N_11685,N_11876);
or U12777 (N_12777,N_11986,N_11508);
xnor U12778 (N_12778,N_11602,N_11494);
nand U12779 (N_12779,N_11528,N_11580);
nand U12780 (N_12780,N_11403,N_11425);
or U12781 (N_12781,N_11782,N_11570);
nor U12782 (N_12782,N_11363,N_11780);
xor U12783 (N_12783,N_11923,N_11903);
nand U12784 (N_12784,N_11688,N_11381);
and U12785 (N_12785,N_11227,N_11919);
xor U12786 (N_12786,N_11746,N_11664);
xnor U12787 (N_12787,N_11811,N_11953);
or U12788 (N_12788,N_11426,N_11898);
xor U12789 (N_12789,N_11908,N_11282);
xnor U12790 (N_12790,N_11782,N_11721);
or U12791 (N_12791,N_11954,N_11833);
nand U12792 (N_12792,N_11592,N_11253);
xnor U12793 (N_12793,N_11328,N_11403);
or U12794 (N_12794,N_11772,N_11536);
nor U12795 (N_12795,N_11639,N_11883);
nand U12796 (N_12796,N_11492,N_11433);
xor U12797 (N_12797,N_11993,N_11442);
and U12798 (N_12798,N_11204,N_11626);
nand U12799 (N_12799,N_11479,N_11881);
nand U12800 (N_12800,N_12388,N_12436);
xor U12801 (N_12801,N_12609,N_12769);
or U12802 (N_12802,N_12539,N_12641);
or U12803 (N_12803,N_12521,N_12125);
and U12804 (N_12804,N_12248,N_12040);
nand U12805 (N_12805,N_12008,N_12160);
xnor U12806 (N_12806,N_12785,N_12221);
nand U12807 (N_12807,N_12543,N_12045);
nand U12808 (N_12808,N_12283,N_12715);
nand U12809 (N_12809,N_12751,N_12084);
or U12810 (N_12810,N_12553,N_12727);
nand U12811 (N_12811,N_12281,N_12644);
nand U12812 (N_12812,N_12398,N_12441);
xnor U12813 (N_12813,N_12180,N_12113);
xor U12814 (N_12814,N_12597,N_12577);
and U12815 (N_12815,N_12695,N_12158);
nor U12816 (N_12816,N_12637,N_12691);
nand U12817 (N_12817,N_12055,N_12271);
or U12818 (N_12818,N_12462,N_12610);
nand U12819 (N_12819,N_12625,N_12519);
xnor U12820 (N_12820,N_12645,N_12209);
nand U12821 (N_12821,N_12781,N_12733);
or U12822 (N_12822,N_12147,N_12096);
nor U12823 (N_12823,N_12205,N_12512);
nor U12824 (N_12824,N_12674,N_12661);
nand U12825 (N_12825,N_12642,N_12511);
nand U12826 (N_12826,N_12282,N_12503);
or U12827 (N_12827,N_12707,N_12237);
xnor U12828 (N_12828,N_12138,N_12187);
and U12829 (N_12829,N_12446,N_12606);
or U12830 (N_12830,N_12599,N_12041);
nor U12831 (N_12831,N_12293,N_12002);
nor U12832 (N_12832,N_12465,N_12063);
xor U12833 (N_12833,N_12703,N_12582);
nor U12834 (N_12834,N_12693,N_12574);
or U12835 (N_12835,N_12506,N_12144);
and U12836 (N_12836,N_12662,N_12375);
xnor U12837 (N_12837,N_12302,N_12774);
or U12838 (N_12838,N_12342,N_12017);
or U12839 (N_12839,N_12027,N_12359);
and U12840 (N_12840,N_12530,N_12287);
and U12841 (N_12841,N_12292,N_12568);
xnor U12842 (N_12842,N_12548,N_12739);
and U12843 (N_12843,N_12748,N_12758);
nor U12844 (N_12844,N_12590,N_12267);
or U12845 (N_12845,N_12172,N_12333);
and U12846 (N_12846,N_12380,N_12690);
xor U12847 (N_12847,N_12663,N_12799);
and U12848 (N_12848,N_12572,N_12254);
nand U12849 (N_12849,N_12276,N_12341);
xnor U12850 (N_12850,N_12518,N_12304);
nand U12851 (N_12851,N_12497,N_12129);
or U12852 (N_12852,N_12598,N_12608);
nand U12853 (N_12853,N_12262,N_12155);
nand U12854 (N_12854,N_12128,N_12786);
and U12855 (N_12855,N_12257,N_12688);
xor U12856 (N_12856,N_12484,N_12225);
nor U12857 (N_12857,N_12194,N_12389);
xor U12858 (N_12858,N_12671,N_12569);
xnor U12859 (N_12859,N_12754,N_12629);
nor U12860 (N_12860,N_12760,N_12654);
and U12861 (N_12861,N_12470,N_12734);
nand U12862 (N_12862,N_12289,N_12090);
and U12863 (N_12863,N_12373,N_12356);
and U12864 (N_12864,N_12489,N_12330);
and U12865 (N_12865,N_12714,N_12717);
xor U12866 (N_12866,N_12583,N_12499);
or U12867 (N_12867,N_12097,N_12021);
and U12868 (N_12868,N_12584,N_12258);
nor U12869 (N_12869,N_12199,N_12475);
nand U12870 (N_12870,N_12686,N_12617);
nor U12871 (N_12871,N_12414,N_12186);
and U12872 (N_12872,N_12448,N_12025);
nor U12873 (N_12873,N_12526,N_12618);
nand U12874 (N_12874,N_12316,N_12740);
or U12875 (N_12875,N_12362,N_12153);
xnor U12876 (N_12876,N_12502,N_12451);
or U12877 (N_12877,N_12407,N_12188);
or U12878 (N_12878,N_12173,N_12633);
xor U12879 (N_12879,N_12500,N_12053);
and U12880 (N_12880,N_12058,N_12042);
nor U12881 (N_12881,N_12790,N_12131);
nand U12882 (N_12882,N_12393,N_12542);
nor U12883 (N_12883,N_12631,N_12249);
or U12884 (N_12884,N_12509,N_12770);
and U12885 (N_12885,N_12697,N_12615);
nand U12886 (N_12886,N_12551,N_12349);
and U12887 (N_12887,N_12562,N_12711);
and U12888 (N_12888,N_12396,N_12377);
xor U12889 (N_12889,N_12731,N_12732);
nor U12890 (N_12890,N_12034,N_12713);
and U12891 (N_12891,N_12259,N_12229);
or U12892 (N_12892,N_12746,N_12481);
nor U12893 (N_12893,N_12545,N_12296);
and U12894 (N_12894,N_12434,N_12080);
nor U12895 (N_12895,N_12060,N_12082);
nand U12896 (N_12896,N_12114,N_12167);
or U12897 (N_12897,N_12395,N_12412);
xor U12898 (N_12898,N_12202,N_12591);
nor U12899 (N_12899,N_12667,N_12496);
nor U12900 (N_12900,N_12555,N_12640);
nor U12901 (N_12901,N_12201,N_12438);
or U12902 (N_12902,N_12214,N_12603);
xnor U12903 (N_12903,N_12284,N_12386);
nor U12904 (N_12904,N_12531,N_12750);
and U12905 (N_12905,N_12309,N_12321);
nor U12906 (N_12906,N_12763,N_12081);
xnor U12907 (N_12907,N_12013,N_12263);
nor U12908 (N_12908,N_12533,N_12219);
xnor U12909 (N_12909,N_12437,N_12534);
nand U12910 (N_12910,N_12247,N_12652);
nor U12911 (N_12911,N_12657,N_12408);
nand U12912 (N_12912,N_12230,N_12520);
and U12913 (N_12913,N_12741,N_12235);
and U12914 (N_12914,N_12440,N_12651);
xor U12915 (N_12915,N_12239,N_12347);
and U12916 (N_12916,N_12211,N_12495);
or U12917 (N_12917,N_12007,N_12616);
xnor U12918 (N_12918,N_12505,N_12100);
nand U12919 (N_12919,N_12093,N_12557);
or U12920 (N_12920,N_12387,N_12277);
and U12921 (N_12921,N_12791,N_12384);
nand U12922 (N_12922,N_12265,N_12527);
xnor U12923 (N_12923,N_12112,N_12383);
and U12924 (N_12924,N_12464,N_12123);
or U12925 (N_12925,N_12579,N_12433);
and U12926 (N_12926,N_12317,N_12033);
nor U12927 (N_12927,N_12325,N_12655);
nor U12928 (N_12928,N_12665,N_12614);
nor U12929 (N_12929,N_12683,N_12793);
xor U12930 (N_12930,N_12626,N_12355);
xor U12931 (N_12931,N_12687,N_12723);
nand U12932 (N_12932,N_12454,N_12184);
nand U12933 (N_12933,N_12024,N_12189);
nor U12934 (N_12934,N_12547,N_12745);
nand U12935 (N_12935,N_12285,N_12392);
or U12936 (N_12936,N_12251,N_12623);
nor U12937 (N_12937,N_12587,N_12066);
nand U12938 (N_12938,N_12401,N_12728);
or U12939 (N_12939,N_12274,N_12327);
xnor U12940 (N_12940,N_12198,N_12191);
xor U12941 (N_12941,N_12213,N_12299);
nand U12942 (N_12942,N_12493,N_12491);
or U12943 (N_12943,N_12563,N_12098);
xor U12944 (N_12944,N_12541,N_12461);
or U12945 (N_12945,N_12567,N_12535);
or U12946 (N_12946,N_12789,N_12444);
nor U12947 (N_12947,N_12596,N_12212);
and U12948 (N_12948,N_12190,N_12658);
or U12949 (N_12949,N_12385,N_12056);
or U12950 (N_12950,N_12064,N_12312);
or U12951 (N_12951,N_12417,N_12656);
and U12952 (N_12952,N_12337,N_12668);
and U12953 (N_12953,N_12639,N_12515);
or U12954 (N_12954,N_12038,N_12694);
xnor U12955 (N_12955,N_12611,N_12650);
nor U12956 (N_12956,N_12540,N_12314);
nand U12957 (N_12957,N_12346,N_12692);
and U12958 (N_12958,N_12012,N_12738);
nor U12959 (N_12959,N_12099,N_12203);
xor U12960 (N_12960,N_12719,N_12702);
and U12961 (N_12961,N_12044,N_12605);
xnor U12962 (N_12962,N_12442,N_12195);
and U12963 (N_12963,N_12405,N_12394);
nor U12964 (N_12964,N_12571,N_12071);
nor U12965 (N_12965,N_12528,N_12415);
xnor U12966 (N_12966,N_12111,N_12701);
or U12967 (N_12967,N_12323,N_12266);
nor U12968 (N_12968,N_12788,N_12119);
or U12969 (N_12969,N_12704,N_12411);
nor U12970 (N_12970,N_12600,N_12218);
nand U12971 (N_12971,N_12028,N_12718);
and U12972 (N_12972,N_12091,N_12428);
nand U12973 (N_12973,N_12004,N_12369);
xor U12974 (N_12974,N_12196,N_12480);
and U12975 (N_12975,N_12592,N_12578);
or U12976 (N_12976,N_12143,N_12647);
xnor U12977 (N_12977,N_12653,N_12101);
nor U12978 (N_12978,N_12370,N_12242);
or U12979 (N_12979,N_12087,N_12179);
and U12980 (N_12980,N_12580,N_12636);
and U12981 (N_12981,N_12525,N_12675);
and U12982 (N_12982,N_12455,N_12275);
and U12983 (N_12983,N_12376,N_12332);
or U12984 (N_12984,N_12161,N_12065);
nand U12985 (N_12985,N_12443,N_12106);
nand U12986 (N_12986,N_12780,N_12260);
nand U12987 (N_12987,N_12456,N_12742);
or U12988 (N_12988,N_12104,N_12747);
and U12989 (N_12989,N_12241,N_12410);
nand U12990 (N_12990,N_12344,N_12059);
xor U12991 (N_12991,N_12326,N_12297);
nand U12992 (N_12992,N_12423,N_12372);
nor U12993 (N_12993,N_12245,N_12200);
nor U12994 (N_12994,N_12273,N_12418);
xor U12995 (N_12995,N_12607,N_12472);
nor U12996 (N_12996,N_12048,N_12593);
nand U12997 (N_12997,N_12320,N_12420);
and U12998 (N_12998,N_12779,N_12677);
xor U12999 (N_12999,N_12020,N_12014);
nor U13000 (N_13000,N_12560,N_12105);
nand U13001 (N_13001,N_12029,N_12336);
or U13002 (N_13002,N_12166,N_12117);
nor U13003 (N_13003,N_12351,N_12413);
or U13004 (N_13004,N_12223,N_12430);
xnor U13005 (N_13005,N_12238,N_12057);
nor U13006 (N_13006,N_12537,N_12146);
nand U13007 (N_13007,N_12797,N_12450);
xor U13008 (N_13008,N_12483,N_12368);
nor U13009 (N_13009,N_12796,N_12348);
and U13010 (N_13010,N_12030,N_12108);
nor U13011 (N_13011,N_12700,N_12737);
nand U13012 (N_13012,N_12233,N_12310);
nor U13013 (N_13013,N_12364,N_12795);
or U13014 (N_13014,N_12508,N_12306);
nor U13015 (N_13015,N_12141,N_12010);
nor U13016 (N_13016,N_12252,N_12552);
or U13017 (N_13017,N_12432,N_12234);
and U13018 (N_13018,N_12447,N_12749);
xor U13019 (N_13019,N_12102,N_12685);
nor U13020 (N_13020,N_12130,N_12178);
xor U13021 (N_13021,N_12126,N_12773);
or U13022 (N_13022,N_12517,N_12120);
xor U13023 (N_13023,N_12043,N_12089);
nand U13024 (N_13024,N_12268,N_12776);
and U13025 (N_13025,N_12513,N_12538);
and U13026 (N_13026,N_12291,N_12156);
and U13027 (N_13027,N_12335,N_12586);
nor U13028 (N_13028,N_12471,N_12744);
xnor U13029 (N_13029,N_12110,N_12624);
nand U13030 (N_13030,N_12649,N_12019);
and U13031 (N_13031,N_12094,N_12504);
or U13032 (N_13032,N_12382,N_12490);
xor U13033 (N_13033,N_12445,N_12487);
and U13034 (N_13034,N_12039,N_12075);
or U13035 (N_13035,N_12660,N_12666);
or U13036 (N_13036,N_12118,N_12595);
nand U13037 (N_13037,N_12003,N_12115);
nand U13038 (N_13038,N_12722,N_12708);
or U13039 (N_13039,N_12556,N_12208);
and U13040 (N_13040,N_12354,N_12255);
or U13041 (N_13041,N_12404,N_12689);
nor U13042 (N_13042,N_12232,N_12762);
and U13043 (N_13043,N_12575,N_12676);
nand U13044 (N_13044,N_12680,N_12185);
or U13045 (N_13045,N_12301,N_12710);
nand U13046 (N_13046,N_12062,N_12315);
nor U13047 (N_13047,N_12109,N_12127);
and U13048 (N_13048,N_12137,N_12116);
xor U13049 (N_13049,N_12678,N_12452);
nor U13050 (N_13050,N_12716,N_12240);
nand U13051 (N_13051,N_12357,N_12712);
and U13052 (N_13052,N_12148,N_12699);
and U13053 (N_13053,N_12630,N_12514);
nand U13054 (N_13054,N_12345,N_12107);
xor U13055 (N_13055,N_12510,N_12322);
nand U13056 (N_13056,N_12243,N_12253);
and U13057 (N_13057,N_12473,N_12778);
nand U13058 (N_13058,N_12554,N_12669);
and U13059 (N_13059,N_12244,N_12051);
xor U13060 (N_13060,N_12482,N_12278);
or U13061 (N_13061,N_12536,N_12588);
nand U13062 (N_13062,N_12050,N_12516);
xor U13063 (N_13063,N_12479,N_12022);
nor U13064 (N_13064,N_12005,N_12139);
and U13065 (N_13065,N_12132,N_12334);
or U13066 (N_13066,N_12419,N_12400);
and U13067 (N_13067,N_12145,N_12559);
xor U13068 (N_13068,N_12549,N_12054);
or U13069 (N_13069,N_12224,N_12206);
nand U13070 (N_13070,N_12544,N_12338);
and U13071 (N_13071,N_12318,N_12602);
nor U13072 (N_13072,N_12403,N_12366);
and U13073 (N_13073,N_12074,N_12648);
or U13074 (N_13074,N_12378,N_12416);
xor U13075 (N_13075,N_12288,N_12061);
nand U13076 (N_13076,N_12183,N_12726);
nand U13077 (N_13077,N_12049,N_12032);
xnor U13078 (N_13078,N_12492,N_12399);
or U13079 (N_13079,N_12072,N_12371);
or U13080 (N_13080,N_12016,N_12585);
xnor U13081 (N_13081,N_12724,N_12078);
and U13082 (N_13082,N_12467,N_12290);
nor U13083 (N_13083,N_12374,N_12365);
and U13084 (N_13084,N_12720,N_12092);
xnor U13085 (N_13085,N_12220,N_12397);
nor U13086 (N_13086,N_12681,N_12421);
and U13087 (N_13087,N_12231,N_12307);
or U13088 (N_13088,N_12460,N_12086);
xor U13089 (N_13089,N_12565,N_12000);
nor U13090 (N_13090,N_12226,N_12476);
nand U13091 (N_13091,N_12772,N_12498);
nor U13092 (N_13092,N_12705,N_12210);
xnor U13093 (N_13093,N_12133,N_12619);
xor U13094 (N_13094,N_12439,N_12798);
and U13095 (N_13095,N_12522,N_12477);
nand U13096 (N_13096,N_12328,N_12023);
xnor U13097 (N_13097,N_12573,N_12696);
or U13098 (N_13098,N_12402,N_12264);
and U13099 (N_13099,N_12069,N_12026);
xnor U13100 (N_13100,N_12735,N_12154);
nor U13101 (N_13101,N_12103,N_12164);
nor U13102 (N_13102,N_12435,N_12228);
and U13103 (N_13103,N_12766,N_12149);
nor U13104 (N_13104,N_12391,N_12706);
and U13105 (N_13105,N_12207,N_12634);
or U13106 (N_13106,N_12469,N_12163);
xor U13107 (N_13107,N_12725,N_12478);
or U13108 (N_13108,N_12169,N_12319);
nor U13109 (N_13109,N_12673,N_12601);
or U13110 (N_13110,N_12272,N_12083);
and U13111 (N_13111,N_12627,N_12331);
or U13112 (N_13112,N_12589,N_12635);
and U13113 (N_13113,N_12775,N_12759);
or U13114 (N_13114,N_12204,N_12682);
xor U13115 (N_13115,N_12488,N_12794);
xnor U13116 (N_13116,N_12494,N_12390);
or U13117 (N_13117,N_12379,N_12157);
xor U13118 (N_13118,N_12523,N_12581);
xnor U13119 (N_13119,N_12300,N_12426);
nand U13120 (N_13120,N_12621,N_12171);
or U13121 (N_13121,N_12270,N_12073);
nand U13122 (N_13122,N_12011,N_12070);
nand U13123 (N_13123,N_12136,N_12076);
or U13124 (N_13124,N_12679,N_12736);
nor U13125 (N_13125,N_12176,N_12729);
and U13126 (N_13126,N_12256,N_12095);
and U13127 (N_13127,N_12122,N_12767);
and U13128 (N_13128,N_12449,N_12558);
xnor U13129 (N_13129,N_12768,N_12215);
nor U13130 (N_13130,N_12771,N_12236);
or U13131 (N_13131,N_12646,N_12036);
xnor U13132 (N_13132,N_12339,N_12324);
xnor U13133 (N_13133,N_12546,N_12170);
or U13134 (N_13134,N_12177,N_12532);
and U13135 (N_13135,N_12564,N_12622);
and U13136 (N_13136,N_12353,N_12427);
xor U13137 (N_13137,N_12352,N_12612);
nor U13138 (N_13138,N_12018,N_12077);
or U13139 (N_13139,N_12250,N_12037);
xor U13140 (N_13140,N_12409,N_12782);
or U13141 (N_13141,N_12052,N_12761);
or U13142 (N_13142,N_12570,N_12361);
xor U13143 (N_13143,N_12604,N_12783);
and U13144 (N_13144,N_12670,N_12613);
and U13145 (N_13145,N_12643,N_12550);
nor U13146 (N_13146,N_12142,N_12261);
nor U13147 (N_13147,N_12381,N_12006);
xnor U13148 (N_13148,N_12684,N_12162);
nand U13149 (N_13149,N_12468,N_12295);
xor U13150 (N_13150,N_12458,N_12088);
nand U13151 (N_13151,N_12743,N_12672);
nand U13152 (N_13152,N_12193,N_12134);
nor U13153 (N_13153,N_12181,N_12507);
xor U13154 (N_13154,N_12709,N_12474);
nor U13155 (N_13155,N_12067,N_12311);
and U13156 (N_13156,N_12664,N_12730);
or U13157 (N_13157,N_12463,N_12457);
nand U13158 (N_13158,N_12001,N_12308);
nand U13159 (N_13159,N_12529,N_12217);
xor U13160 (N_13160,N_12182,N_12628);
nand U13161 (N_13161,N_12721,N_12561);
xor U13162 (N_13162,N_12298,N_12367);
nor U13163 (N_13163,N_12363,N_12046);
xor U13164 (N_13164,N_12175,N_12286);
nor U13165 (N_13165,N_12765,N_12485);
xor U13166 (N_13166,N_12752,N_12009);
or U13167 (N_13167,N_12360,N_12152);
xor U13168 (N_13168,N_12406,N_12159);
nand U13169 (N_13169,N_12632,N_12150);
or U13170 (N_13170,N_12168,N_12698);
or U13171 (N_13171,N_12305,N_12085);
nand U13172 (N_13172,N_12279,N_12429);
and U13173 (N_13173,N_12777,N_12784);
nand U13174 (N_13174,N_12047,N_12594);
nor U13175 (N_13175,N_12459,N_12486);
and U13176 (N_13176,N_12764,N_12329);
nor U13177 (N_13177,N_12174,N_12303);
or U13178 (N_13178,N_12197,N_12121);
nor U13179 (N_13179,N_12576,N_12424);
xor U13180 (N_13180,N_12358,N_12340);
xnor U13181 (N_13181,N_12135,N_12079);
nand U13182 (N_13182,N_12222,N_12753);
nand U13183 (N_13183,N_12638,N_12294);
or U13184 (N_13184,N_12453,N_12151);
nand U13185 (N_13185,N_12501,N_12269);
and U13186 (N_13186,N_12787,N_12165);
and U13187 (N_13187,N_12031,N_12140);
or U13188 (N_13188,N_12620,N_12466);
nor U13189 (N_13189,N_12192,N_12756);
and U13190 (N_13190,N_12422,N_12425);
and U13191 (N_13191,N_12068,N_12755);
nor U13192 (N_13192,N_12350,N_12313);
nor U13193 (N_13193,N_12659,N_12035);
or U13194 (N_13194,N_12227,N_12431);
or U13195 (N_13195,N_12015,N_12216);
nand U13196 (N_13196,N_12124,N_12566);
nand U13197 (N_13197,N_12524,N_12246);
or U13198 (N_13198,N_12757,N_12792);
and U13199 (N_13199,N_12280,N_12343);
nand U13200 (N_13200,N_12638,N_12022);
xnor U13201 (N_13201,N_12270,N_12263);
nor U13202 (N_13202,N_12146,N_12776);
nor U13203 (N_13203,N_12216,N_12043);
or U13204 (N_13204,N_12668,N_12203);
xnor U13205 (N_13205,N_12717,N_12162);
nand U13206 (N_13206,N_12248,N_12143);
nor U13207 (N_13207,N_12438,N_12266);
and U13208 (N_13208,N_12729,N_12498);
xor U13209 (N_13209,N_12384,N_12549);
and U13210 (N_13210,N_12096,N_12227);
xnor U13211 (N_13211,N_12265,N_12554);
xnor U13212 (N_13212,N_12639,N_12144);
xor U13213 (N_13213,N_12627,N_12794);
nor U13214 (N_13214,N_12205,N_12723);
or U13215 (N_13215,N_12779,N_12405);
or U13216 (N_13216,N_12123,N_12658);
nor U13217 (N_13217,N_12257,N_12284);
and U13218 (N_13218,N_12041,N_12791);
xnor U13219 (N_13219,N_12594,N_12678);
nor U13220 (N_13220,N_12044,N_12473);
and U13221 (N_13221,N_12498,N_12676);
and U13222 (N_13222,N_12273,N_12496);
or U13223 (N_13223,N_12741,N_12102);
or U13224 (N_13224,N_12377,N_12651);
and U13225 (N_13225,N_12410,N_12700);
or U13226 (N_13226,N_12074,N_12509);
nand U13227 (N_13227,N_12585,N_12326);
nand U13228 (N_13228,N_12116,N_12459);
nand U13229 (N_13229,N_12109,N_12344);
nand U13230 (N_13230,N_12145,N_12307);
nand U13231 (N_13231,N_12040,N_12096);
and U13232 (N_13232,N_12042,N_12073);
and U13233 (N_13233,N_12242,N_12404);
nand U13234 (N_13234,N_12492,N_12768);
and U13235 (N_13235,N_12174,N_12114);
xor U13236 (N_13236,N_12020,N_12190);
nor U13237 (N_13237,N_12205,N_12446);
xnor U13238 (N_13238,N_12447,N_12352);
xnor U13239 (N_13239,N_12140,N_12082);
or U13240 (N_13240,N_12784,N_12357);
and U13241 (N_13241,N_12136,N_12100);
nor U13242 (N_13242,N_12594,N_12299);
nor U13243 (N_13243,N_12326,N_12251);
nand U13244 (N_13244,N_12670,N_12535);
xnor U13245 (N_13245,N_12110,N_12658);
nor U13246 (N_13246,N_12605,N_12127);
xnor U13247 (N_13247,N_12183,N_12241);
or U13248 (N_13248,N_12145,N_12412);
xor U13249 (N_13249,N_12335,N_12394);
or U13250 (N_13250,N_12777,N_12618);
and U13251 (N_13251,N_12698,N_12341);
nand U13252 (N_13252,N_12659,N_12096);
nand U13253 (N_13253,N_12079,N_12364);
nand U13254 (N_13254,N_12293,N_12549);
nand U13255 (N_13255,N_12004,N_12482);
nand U13256 (N_13256,N_12261,N_12033);
nand U13257 (N_13257,N_12733,N_12491);
xor U13258 (N_13258,N_12596,N_12634);
or U13259 (N_13259,N_12466,N_12699);
xor U13260 (N_13260,N_12410,N_12020);
and U13261 (N_13261,N_12401,N_12332);
nor U13262 (N_13262,N_12075,N_12263);
and U13263 (N_13263,N_12346,N_12495);
nand U13264 (N_13264,N_12766,N_12610);
xnor U13265 (N_13265,N_12006,N_12251);
xor U13266 (N_13266,N_12107,N_12640);
or U13267 (N_13267,N_12217,N_12501);
or U13268 (N_13268,N_12003,N_12451);
nor U13269 (N_13269,N_12163,N_12785);
and U13270 (N_13270,N_12369,N_12041);
or U13271 (N_13271,N_12166,N_12729);
and U13272 (N_13272,N_12310,N_12757);
or U13273 (N_13273,N_12023,N_12029);
or U13274 (N_13274,N_12624,N_12056);
nand U13275 (N_13275,N_12676,N_12157);
or U13276 (N_13276,N_12047,N_12785);
and U13277 (N_13277,N_12747,N_12258);
xor U13278 (N_13278,N_12551,N_12644);
and U13279 (N_13279,N_12402,N_12475);
and U13280 (N_13280,N_12522,N_12591);
nor U13281 (N_13281,N_12218,N_12585);
and U13282 (N_13282,N_12215,N_12006);
xnor U13283 (N_13283,N_12452,N_12139);
nand U13284 (N_13284,N_12615,N_12571);
nand U13285 (N_13285,N_12037,N_12291);
and U13286 (N_13286,N_12170,N_12643);
and U13287 (N_13287,N_12414,N_12775);
xor U13288 (N_13288,N_12049,N_12793);
nand U13289 (N_13289,N_12681,N_12351);
and U13290 (N_13290,N_12467,N_12625);
and U13291 (N_13291,N_12561,N_12275);
nor U13292 (N_13292,N_12505,N_12223);
or U13293 (N_13293,N_12384,N_12632);
nand U13294 (N_13294,N_12535,N_12007);
nand U13295 (N_13295,N_12473,N_12236);
and U13296 (N_13296,N_12531,N_12020);
nor U13297 (N_13297,N_12007,N_12064);
or U13298 (N_13298,N_12184,N_12335);
nor U13299 (N_13299,N_12777,N_12019);
and U13300 (N_13300,N_12658,N_12170);
or U13301 (N_13301,N_12357,N_12559);
nor U13302 (N_13302,N_12520,N_12108);
nor U13303 (N_13303,N_12508,N_12401);
nor U13304 (N_13304,N_12643,N_12672);
nand U13305 (N_13305,N_12534,N_12525);
nand U13306 (N_13306,N_12769,N_12340);
or U13307 (N_13307,N_12369,N_12263);
or U13308 (N_13308,N_12487,N_12099);
nand U13309 (N_13309,N_12105,N_12532);
nand U13310 (N_13310,N_12212,N_12502);
nand U13311 (N_13311,N_12502,N_12723);
xor U13312 (N_13312,N_12616,N_12753);
or U13313 (N_13313,N_12156,N_12628);
nor U13314 (N_13314,N_12409,N_12681);
xnor U13315 (N_13315,N_12776,N_12294);
xor U13316 (N_13316,N_12345,N_12284);
or U13317 (N_13317,N_12109,N_12576);
nor U13318 (N_13318,N_12765,N_12368);
nand U13319 (N_13319,N_12465,N_12004);
nor U13320 (N_13320,N_12012,N_12167);
and U13321 (N_13321,N_12323,N_12686);
nand U13322 (N_13322,N_12407,N_12495);
xnor U13323 (N_13323,N_12311,N_12227);
or U13324 (N_13324,N_12142,N_12523);
and U13325 (N_13325,N_12163,N_12647);
nor U13326 (N_13326,N_12387,N_12549);
xor U13327 (N_13327,N_12227,N_12015);
xor U13328 (N_13328,N_12722,N_12576);
nand U13329 (N_13329,N_12442,N_12453);
and U13330 (N_13330,N_12557,N_12001);
or U13331 (N_13331,N_12647,N_12454);
nand U13332 (N_13332,N_12510,N_12559);
or U13333 (N_13333,N_12172,N_12266);
or U13334 (N_13334,N_12392,N_12749);
nor U13335 (N_13335,N_12586,N_12648);
nor U13336 (N_13336,N_12592,N_12034);
or U13337 (N_13337,N_12763,N_12748);
xor U13338 (N_13338,N_12232,N_12012);
nand U13339 (N_13339,N_12716,N_12095);
nand U13340 (N_13340,N_12106,N_12123);
xnor U13341 (N_13341,N_12635,N_12703);
nor U13342 (N_13342,N_12130,N_12332);
nand U13343 (N_13343,N_12698,N_12639);
or U13344 (N_13344,N_12173,N_12669);
and U13345 (N_13345,N_12198,N_12308);
and U13346 (N_13346,N_12183,N_12668);
and U13347 (N_13347,N_12232,N_12519);
nand U13348 (N_13348,N_12484,N_12753);
or U13349 (N_13349,N_12638,N_12178);
and U13350 (N_13350,N_12252,N_12422);
xnor U13351 (N_13351,N_12554,N_12282);
xor U13352 (N_13352,N_12249,N_12219);
nor U13353 (N_13353,N_12397,N_12459);
nor U13354 (N_13354,N_12679,N_12282);
or U13355 (N_13355,N_12131,N_12251);
or U13356 (N_13356,N_12545,N_12358);
xnor U13357 (N_13357,N_12590,N_12212);
nand U13358 (N_13358,N_12166,N_12238);
nor U13359 (N_13359,N_12023,N_12372);
and U13360 (N_13360,N_12505,N_12057);
nand U13361 (N_13361,N_12468,N_12486);
xor U13362 (N_13362,N_12648,N_12775);
and U13363 (N_13363,N_12599,N_12268);
or U13364 (N_13364,N_12185,N_12411);
xor U13365 (N_13365,N_12091,N_12110);
xnor U13366 (N_13366,N_12594,N_12435);
nand U13367 (N_13367,N_12350,N_12113);
or U13368 (N_13368,N_12714,N_12423);
nand U13369 (N_13369,N_12338,N_12068);
and U13370 (N_13370,N_12639,N_12286);
nand U13371 (N_13371,N_12087,N_12688);
nand U13372 (N_13372,N_12435,N_12691);
nand U13373 (N_13373,N_12150,N_12447);
nor U13374 (N_13374,N_12509,N_12722);
nand U13375 (N_13375,N_12395,N_12665);
xnor U13376 (N_13376,N_12397,N_12768);
or U13377 (N_13377,N_12766,N_12351);
nand U13378 (N_13378,N_12655,N_12351);
nor U13379 (N_13379,N_12368,N_12066);
xor U13380 (N_13380,N_12399,N_12398);
and U13381 (N_13381,N_12741,N_12451);
nand U13382 (N_13382,N_12583,N_12762);
or U13383 (N_13383,N_12198,N_12159);
and U13384 (N_13384,N_12762,N_12256);
nand U13385 (N_13385,N_12612,N_12037);
or U13386 (N_13386,N_12552,N_12669);
or U13387 (N_13387,N_12311,N_12438);
or U13388 (N_13388,N_12613,N_12341);
or U13389 (N_13389,N_12571,N_12562);
or U13390 (N_13390,N_12572,N_12213);
and U13391 (N_13391,N_12226,N_12777);
nand U13392 (N_13392,N_12234,N_12560);
or U13393 (N_13393,N_12601,N_12491);
and U13394 (N_13394,N_12553,N_12731);
nor U13395 (N_13395,N_12676,N_12051);
nor U13396 (N_13396,N_12798,N_12599);
nand U13397 (N_13397,N_12444,N_12470);
or U13398 (N_13398,N_12329,N_12780);
or U13399 (N_13399,N_12510,N_12281);
xnor U13400 (N_13400,N_12421,N_12158);
or U13401 (N_13401,N_12330,N_12205);
xnor U13402 (N_13402,N_12703,N_12730);
and U13403 (N_13403,N_12436,N_12091);
xnor U13404 (N_13404,N_12607,N_12301);
xor U13405 (N_13405,N_12681,N_12691);
nand U13406 (N_13406,N_12790,N_12009);
xnor U13407 (N_13407,N_12208,N_12363);
or U13408 (N_13408,N_12247,N_12451);
nand U13409 (N_13409,N_12410,N_12168);
and U13410 (N_13410,N_12730,N_12230);
and U13411 (N_13411,N_12163,N_12291);
nand U13412 (N_13412,N_12098,N_12188);
xor U13413 (N_13413,N_12735,N_12618);
xnor U13414 (N_13414,N_12736,N_12203);
and U13415 (N_13415,N_12764,N_12722);
and U13416 (N_13416,N_12668,N_12647);
or U13417 (N_13417,N_12182,N_12047);
nand U13418 (N_13418,N_12037,N_12046);
and U13419 (N_13419,N_12197,N_12333);
or U13420 (N_13420,N_12657,N_12074);
or U13421 (N_13421,N_12294,N_12527);
and U13422 (N_13422,N_12445,N_12677);
nor U13423 (N_13423,N_12172,N_12718);
or U13424 (N_13424,N_12448,N_12446);
or U13425 (N_13425,N_12065,N_12669);
xor U13426 (N_13426,N_12248,N_12623);
and U13427 (N_13427,N_12090,N_12554);
nor U13428 (N_13428,N_12495,N_12699);
or U13429 (N_13429,N_12639,N_12444);
xor U13430 (N_13430,N_12351,N_12794);
nor U13431 (N_13431,N_12180,N_12268);
nor U13432 (N_13432,N_12017,N_12285);
or U13433 (N_13433,N_12312,N_12164);
nor U13434 (N_13434,N_12631,N_12602);
and U13435 (N_13435,N_12140,N_12760);
or U13436 (N_13436,N_12713,N_12019);
nor U13437 (N_13437,N_12528,N_12542);
xnor U13438 (N_13438,N_12460,N_12189);
nor U13439 (N_13439,N_12746,N_12714);
nand U13440 (N_13440,N_12547,N_12082);
xnor U13441 (N_13441,N_12454,N_12378);
xnor U13442 (N_13442,N_12662,N_12668);
nand U13443 (N_13443,N_12252,N_12576);
nand U13444 (N_13444,N_12173,N_12557);
nand U13445 (N_13445,N_12017,N_12163);
and U13446 (N_13446,N_12713,N_12079);
xnor U13447 (N_13447,N_12688,N_12699);
and U13448 (N_13448,N_12227,N_12200);
xor U13449 (N_13449,N_12560,N_12723);
or U13450 (N_13450,N_12343,N_12673);
and U13451 (N_13451,N_12472,N_12481);
nand U13452 (N_13452,N_12613,N_12623);
or U13453 (N_13453,N_12468,N_12573);
nor U13454 (N_13454,N_12431,N_12219);
nor U13455 (N_13455,N_12352,N_12586);
or U13456 (N_13456,N_12183,N_12239);
nor U13457 (N_13457,N_12001,N_12014);
and U13458 (N_13458,N_12382,N_12668);
nor U13459 (N_13459,N_12729,N_12200);
nand U13460 (N_13460,N_12111,N_12283);
and U13461 (N_13461,N_12248,N_12036);
and U13462 (N_13462,N_12166,N_12506);
nor U13463 (N_13463,N_12673,N_12214);
and U13464 (N_13464,N_12296,N_12514);
nor U13465 (N_13465,N_12209,N_12678);
and U13466 (N_13466,N_12470,N_12562);
or U13467 (N_13467,N_12617,N_12108);
and U13468 (N_13468,N_12783,N_12742);
nor U13469 (N_13469,N_12276,N_12085);
nand U13470 (N_13470,N_12137,N_12006);
or U13471 (N_13471,N_12289,N_12228);
and U13472 (N_13472,N_12494,N_12675);
nor U13473 (N_13473,N_12269,N_12559);
nand U13474 (N_13474,N_12601,N_12187);
nand U13475 (N_13475,N_12674,N_12724);
or U13476 (N_13476,N_12345,N_12783);
or U13477 (N_13477,N_12373,N_12225);
xnor U13478 (N_13478,N_12323,N_12227);
nor U13479 (N_13479,N_12556,N_12359);
nand U13480 (N_13480,N_12518,N_12468);
and U13481 (N_13481,N_12367,N_12550);
or U13482 (N_13482,N_12362,N_12391);
nor U13483 (N_13483,N_12288,N_12290);
nor U13484 (N_13484,N_12753,N_12206);
nand U13485 (N_13485,N_12366,N_12326);
or U13486 (N_13486,N_12215,N_12244);
or U13487 (N_13487,N_12622,N_12596);
nor U13488 (N_13488,N_12016,N_12633);
nand U13489 (N_13489,N_12337,N_12523);
or U13490 (N_13490,N_12549,N_12351);
or U13491 (N_13491,N_12713,N_12707);
nand U13492 (N_13492,N_12406,N_12587);
and U13493 (N_13493,N_12701,N_12274);
and U13494 (N_13494,N_12329,N_12408);
nor U13495 (N_13495,N_12145,N_12551);
nor U13496 (N_13496,N_12128,N_12543);
nor U13497 (N_13497,N_12334,N_12583);
and U13498 (N_13498,N_12703,N_12489);
and U13499 (N_13499,N_12791,N_12067);
xnor U13500 (N_13500,N_12062,N_12635);
nand U13501 (N_13501,N_12538,N_12336);
nand U13502 (N_13502,N_12699,N_12687);
and U13503 (N_13503,N_12280,N_12341);
or U13504 (N_13504,N_12210,N_12103);
nand U13505 (N_13505,N_12676,N_12504);
or U13506 (N_13506,N_12176,N_12320);
or U13507 (N_13507,N_12124,N_12422);
or U13508 (N_13508,N_12500,N_12459);
nor U13509 (N_13509,N_12620,N_12125);
and U13510 (N_13510,N_12245,N_12793);
nor U13511 (N_13511,N_12772,N_12014);
nor U13512 (N_13512,N_12165,N_12522);
and U13513 (N_13513,N_12429,N_12672);
nor U13514 (N_13514,N_12259,N_12283);
nand U13515 (N_13515,N_12119,N_12706);
xor U13516 (N_13516,N_12617,N_12098);
and U13517 (N_13517,N_12427,N_12476);
or U13518 (N_13518,N_12034,N_12112);
nor U13519 (N_13519,N_12682,N_12008);
nand U13520 (N_13520,N_12146,N_12410);
nand U13521 (N_13521,N_12107,N_12350);
nor U13522 (N_13522,N_12402,N_12147);
nor U13523 (N_13523,N_12563,N_12602);
or U13524 (N_13524,N_12178,N_12022);
or U13525 (N_13525,N_12527,N_12684);
or U13526 (N_13526,N_12589,N_12571);
and U13527 (N_13527,N_12765,N_12089);
or U13528 (N_13528,N_12243,N_12462);
nand U13529 (N_13529,N_12142,N_12153);
nor U13530 (N_13530,N_12520,N_12356);
nor U13531 (N_13531,N_12047,N_12139);
or U13532 (N_13532,N_12117,N_12549);
nor U13533 (N_13533,N_12785,N_12533);
nor U13534 (N_13534,N_12693,N_12459);
or U13535 (N_13535,N_12583,N_12323);
or U13536 (N_13536,N_12142,N_12331);
and U13537 (N_13537,N_12625,N_12556);
or U13538 (N_13538,N_12631,N_12266);
and U13539 (N_13539,N_12348,N_12697);
nand U13540 (N_13540,N_12757,N_12431);
and U13541 (N_13541,N_12026,N_12790);
nand U13542 (N_13542,N_12774,N_12413);
nor U13543 (N_13543,N_12488,N_12174);
and U13544 (N_13544,N_12577,N_12485);
nor U13545 (N_13545,N_12222,N_12324);
nor U13546 (N_13546,N_12343,N_12547);
and U13547 (N_13547,N_12693,N_12053);
or U13548 (N_13548,N_12080,N_12653);
xnor U13549 (N_13549,N_12524,N_12673);
nand U13550 (N_13550,N_12692,N_12445);
or U13551 (N_13551,N_12692,N_12537);
and U13552 (N_13552,N_12216,N_12469);
or U13553 (N_13553,N_12379,N_12406);
or U13554 (N_13554,N_12416,N_12023);
nand U13555 (N_13555,N_12755,N_12692);
nor U13556 (N_13556,N_12365,N_12713);
xor U13557 (N_13557,N_12543,N_12004);
nor U13558 (N_13558,N_12138,N_12430);
and U13559 (N_13559,N_12237,N_12594);
nand U13560 (N_13560,N_12293,N_12744);
nand U13561 (N_13561,N_12211,N_12097);
and U13562 (N_13562,N_12416,N_12206);
and U13563 (N_13563,N_12196,N_12141);
nand U13564 (N_13564,N_12427,N_12551);
nor U13565 (N_13565,N_12661,N_12771);
nor U13566 (N_13566,N_12398,N_12177);
nand U13567 (N_13567,N_12231,N_12331);
or U13568 (N_13568,N_12545,N_12542);
nor U13569 (N_13569,N_12037,N_12123);
or U13570 (N_13570,N_12717,N_12724);
nor U13571 (N_13571,N_12655,N_12018);
xnor U13572 (N_13572,N_12556,N_12078);
and U13573 (N_13573,N_12560,N_12602);
and U13574 (N_13574,N_12505,N_12495);
or U13575 (N_13575,N_12576,N_12557);
or U13576 (N_13576,N_12079,N_12477);
or U13577 (N_13577,N_12136,N_12695);
nand U13578 (N_13578,N_12693,N_12669);
nor U13579 (N_13579,N_12705,N_12677);
and U13580 (N_13580,N_12114,N_12064);
xor U13581 (N_13581,N_12125,N_12536);
xor U13582 (N_13582,N_12600,N_12565);
nand U13583 (N_13583,N_12782,N_12066);
or U13584 (N_13584,N_12456,N_12349);
nand U13585 (N_13585,N_12048,N_12011);
and U13586 (N_13586,N_12444,N_12163);
or U13587 (N_13587,N_12059,N_12675);
xor U13588 (N_13588,N_12077,N_12166);
nor U13589 (N_13589,N_12515,N_12681);
nor U13590 (N_13590,N_12656,N_12653);
nor U13591 (N_13591,N_12245,N_12642);
xnor U13592 (N_13592,N_12207,N_12618);
and U13593 (N_13593,N_12326,N_12501);
or U13594 (N_13594,N_12412,N_12163);
and U13595 (N_13595,N_12733,N_12174);
xnor U13596 (N_13596,N_12044,N_12686);
and U13597 (N_13597,N_12513,N_12209);
xor U13598 (N_13598,N_12795,N_12578);
xnor U13599 (N_13599,N_12731,N_12723);
nand U13600 (N_13600,N_12915,N_13569);
nand U13601 (N_13601,N_12983,N_13336);
nand U13602 (N_13602,N_13510,N_13191);
nor U13603 (N_13603,N_12958,N_13523);
xor U13604 (N_13604,N_13036,N_13584);
and U13605 (N_13605,N_13274,N_13306);
nand U13606 (N_13606,N_13431,N_13023);
and U13607 (N_13607,N_13514,N_13102);
nand U13608 (N_13608,N_12828,N_12912);
xnor U13609 (N_13609,N_12898,N_13538);
nand U13610 (N_13610,N_13534,N_13333);
nand U13611 (N_13611,N_13511,N_12874);
xor U13612 (N_13612,N_13440,N_13019);
and U13613 (N_13613,N_12896,N_13087);
nor U13614 (N_13614,N_13299,N_12919);
and U13615 (N_13615,N_13117,N_13119);
nand U13616 (N_13616,N_13066,N_13383);
nand U13617 (N_13617,N_13152,N_13025);
or U13618 (N_13618,N_13298,N_13082);
or U13619 (N_13619,N_12990,N_13277);
xnor U13620 (N_13620,N_13002,N_13108);
xnor U13621 (N_13621,N_13240,N_13507);
and U13622 (N_13622,N_13582,N_13435);
or U13623 (N_13623,N_12895,N_13548);
nand U13624 (N_13624,N_13062,N_13357);
and U13625 (N_13625,N_13218,N_13140);
nor U13626 (N_13626,N_12893,N_13562);
xor U13627 (N_13627,N_13167,N_13091);
or U13628 (N_13628,N_13009,N_13234);
nor U13629 (N_13629,N_13047,N_13169);
nand U13630 (N_13630,N_13075,N_13519);
or U13631 (N_13631,N_13558,N_12993);
or U13632 (N_13632,N_13038,N_13463);
nand U13633 (N_13633,N_13184,N_13145);
nor U13634 (N_13634,N_13127,N_12873);
xor U13635 (N_13635,N_12859,N_12930);
and U13636 (N_13636,N_12812,N_13000);
nand U13637 (N_13637,N_12950,N_13100);
or U13638 (N_13638,N_13283,N_13202);
xor U13639 (N_13639,N_13549,N_13531);
and U13640 (N_13640,N_13280,N_12917);
nor U13641 (N_13641,N_13590,N_13288);
or U13642 (N_13642,N_12968,N_13592);
and U13643 (N_13643,N_13031,N_12823);
nand U13644 (N_13644,N_12988,N_13363);
xnor U13645 (N_13645,N_12967,N_12842);
nor U13646 (N_13646,N_13113,N_13198);
and U13647 (N_13647,N_13294,N_13057);
nand U13648 (N_13648,N_13226,N_12841);
or U13649 (N_13649,N_13556,N_13543);
xnor U13650 (N_13650,N_13493,N_13261);
and U13651 (N_13651,N_13587,N_13498);
xor U13652 (N_13652,N_12805,N_12889);
or U13653 (N_13653,N_13362,N_12867);
nor U13654 (N_13654,N_12811,N_13293);
nor U13655 (N_13655,N_12861,N_13407);
or U13656 (N_13656,N_12900,N_12853);
or U13657 (N_13657,N_13003,N_13395);
xor U13658 (N_13658,N_13273,N_13386);
and U13659 (N_13659,N_13500,N_12883);
and U13660 (N_13660,N_13034,N_13012);
nand U13661 (N_13661,N_13076,N_13227);
or U13662 (N_13662,N_12911,N_13301);
nor U13663 (N_13663,N_13143,N_13391);
nand U13664 (N_13664,N_13521,N_13422);
nor U13665 (N_13665,N_12979,N_13109);
nor U13666 (N_13666,N_13267,N_13216);
nor U13667 (N_13667,N_13461,N_13476);
and U13668 (N_13668,N_12852,N_13517);
nor U13669 (N_13669,N_13266,N_13134);
and U13670 (N_13670,N_13302,N_12864);
xnor U13671 (N_13671,N_13139,N_13397);
nand U13672 (N_13672,N_13300,N_13545);
and U13673 (N_13673,N_13453,N_13427);
or U13674 (N_13674,N_13532,N_13004);
or U13675 (N_13675,N_12872,N_13297);
or U13676 (N_13676,N_12845,N_13046);
or U13677 (N_13677,N_13369,N_13550);
and U13678 (N_13678,N_13092,N_13480);
and U13679 (N_13679,N_12963,N_13367);
and U13680 (N_13680,N_12858,N_13354);
or U13681 (N_13681,N_13473,N_12871);
nand U13682 (N_13682,N_13555,N_13284);
xnor U13683 (N_13683,N_13118,N_13450);
and U13684 (N_13684,N_13350,N_12816);
and U13685 (N_13685,N_13221,N_13196);
nand U13686 (N_13686,N_13518,N_12970);
nand U13687 (N_13687,N_13577,N_13501);
and U13688 (N_13688,N_13346,N_13137);
and U13689 (N_13689,N_13189,N_13268);
or U13690 (N_13690,N_13566,N_13232);
and U13691 (N_13691,N_13553,N_12847);
and U13692 (N_13692,N_12863,N_13123);
nor U13693 (N_13693,N_13467,N_13494);
nand U13694 (N_13694,N_13441,N_13250);
and U13695 (N_13695,N_13307,N_13116);
and U13696 (N_13696,N_13328,N_13131);
nor U13697 (N_13697,N_13182,N_13405);
nand U13698 (N_13698,N_12941,N_13579);
and U13699 (N_13699,N_13241,N_12857);
xor U13700 (N_13700,N_13394,N_13018);
and U13701 (N_13701,N_13275,N_12834);
nor U13702 (N_13702,N_12884,N_13387);
xor U13703 (N_13703,N_13502,N_12829);
xnor U13704 (N_13704,N_13291,N_13542);
nand U13705 (N_13705,N_13259,N_13599);
xnor U13706 (N_13706,N_13327,N_12945);
and U13707 (N_13707,N_12954,N_13376);
or U13708 (N_13708,N_13249,N_12817);
or U13709 (N_13709,N_13215,N_13110);
xnor U13710 (N_13710,N_12894,N_12955);
nor U13711 (N_13711,N_13505,N_12808);
nand U13712 (N_13712,N_12897,N_12980);
nor U13713 (N_13713,N_13225,N_13219);
nand U13714 (N_13714,N_13475,N_12860);
nor U13715 (N_13715,N_13311,N_13286);
xnor U13716 (N_13716,N_13035,N_13237);
xnor U13717 (N_13717,N_13213,N_13173);
or U13718 (N_13718,N_13375,N_13043);
xor U13719 (N_13719,N_13077,N_12998);
nand U13720 (N_13720,N_13398,N_13408);
nand U13721 (N_13721,N_13170,N_13314);
nor U13722 (N_13722,N_13437,N_12866);
and U13723 (N_13723,N_12856,N_12879);
xnor U13724 (N_13724,N_13103,N_13079);
and U13725 (N_13725,N_12985,N_13204);
and U13726 (N_13726,N_13222,N_13158);
nand U13727 (N_13727,N_12906,N_13029);
and U13728 (N_13728,N_13147,N_13088);
and U13729 (N_13729,N_13148,N_13159);
xor U13730 (N_13730,N_12903,N_13420);
and U13731 (N_13731,N_12885,N_13095);
and U13732 (N_13732,N_13146,N_13472);
nor U13733 (N_13733,N_13006,N_13200);
xor U13734 (N_13734,N_12913,N_12922);
and U13735 (N_13735,N_13474,N_13263);
and U13736 (N_13736,N_13128,N_12875);
nand U13737 (N_13737,N_13229,N_12962);
and U13738 (N_13738,N_13344,N_13197);
nand U13739 (N_13739,N_13180,N_13337);
or U13740 (N_13740,N_13488,N_13365);
xnor U13741 (N_13741,N_12914,N_12952);
or U13742 (N_13742,N_13008,N_13552);
nor U13743 (N_13743,N_13329,N_13413);
and U13744 (N_13744,N_13072,N_13432);
or U13745 (N_13745,N_13282,N_13099);
nor U13746 (N_13746,N_13345,N_12918);
or U13747 (N_13747,N_12830,N_12825);
and U13748 (N_13748,N_13506,N_13524);
nor U13749 (N_13749,N_13334,N_13192);
and U13750 (N_13750,N_13172,N_13425);
nor U13751 (N_13751,N_13591,N_13551);
nor U13752 (N_13752,N_13497,N_13439);
nand U13753 (N_13753,N_13338,N_13256);
xor U13754 (N_13754,N_13206,N_13522);
nand U13755 (N_13755,N_13205,N_13166);
nand U13756 (N_13756,N_13187,N_13086);
and U13757 (N_13757,N_13121,N_13112);
and U13758 (N_13758,N_13575,N_12840);
and U13759 (N_13759,N_12835,N_12965);
nand U13760 (N_13760,N_13588,N_13185);
xnor U13761 (N_13761,N_13352,N_13056);
xor U13762 (N_13762,N_13085,N_13157);
xnor U13763 (N_13763,N_13063,N_12844);
nand U13764 (N_13764,N_13257,N_13233);
and U13765 (N_13765,N_13404,N_13262);
or U13766 (N_13766,N_13203,N_13378);
nand U13767 (N_13767,N_13403,N_13212);
nand U13768 (N_13768,N_13144,N_13323);
nor U13769 (N_13769,N_13554,N_13305);
nor U13770 (N_13770,N_13392,N_13084);
nor U13771 (N_13771,N_13471,N_13245);
nand U13772 (N_13772,N_13456,N_12978);
and U13773 (N_13773,N_13013,N_13179);
xnor U13774 (N_13774,N_13050,N_13377);
nor U13775 (N_13775,N_13236,N_13595);
and U13776 (N_13776,N_13401,N_13341);
or U13777 (N_13777,N_13067,N_13135);
or U13778 (N_13778,N_13130,N_13083);
or U13779 (N_13779,N_13389,N_13570);
or U13780 (N_13780,N_13051,N_12821);
nor U13781 (N_13781,N_13574,N_13568);
nand U13782 (N_13782,N_13372,N_13269);
nor U13783 (N_13783,N_12907,N_13078);
nor U13784 (N_13784,N_13561,N_12868);
xor U13785 (N_13785,N_13010,N_12936);
and U13786 (N_13786,N_13381,N_13104);
and U13787 (N_13787,N_12891,N_13005);
or U13788 (N_13788,N_13483,N_13416);
and U13789 (N_13789,N_13559,N_13320);
and U13790 (N_13790,N_13155,N_13193);
nand U13791 (N_13791,N_12849,N_13512);
nand U13792 (N_13792,N_12887,N_13438);
xor U13793 (N_13793,N_13557,N_13513);
xnor U13794 (N_13794,N_13207,N_13281);
or U13795 (N_13795,N_12921,N_13356);
or U13796 (N_13796,N_13138,N_13547);
xnor U13797 (N_13797,N_13429,N_13271);
or U13798 (N_13798,N_12992,N_12905);
and U13799 (N_13799,N_13355,N_13028);
nor U13800 (N_13800,N_13445,N_13343);
or U13801 (N_13801,N_13322,N_13163);
nand U13802 (N_13802,N_13436,N_12947);
nor U13803 (N_13803,N_13089,N_13101);
xor U13804 (N_13804,N_13053,N_13452);
and U13805 (N_13805,N_13348,N_13258);
or U13806 (N_13806,N_12804,N_13370);
xnor U13807 (N_13807,N_13287,N_13011);
xor U13808 (N_13808,N_13541,N_13388);
or U13809 (N_13809,N_13421,N_13265);
xor U13810 (N_13810,N_13243,N_13544);
or U13811 (N_13811,N_12977,N_12809);
nand U13812 (N_13812,N_13492,N_12951);
nand U13813 (N_13813,N_13199,N_13396);
or U13814 (N_13814,N_13107,N_13161);
and U13815 (N_13815,N_12973,N_12882);
and U13816 (N_13816,N_13120,N_12961);
nor U13817 (N_13817,N_13424,N_13399);
nand U13818 (N_13818,N_13446,N_12981);
and U13819 (N_13819,N_13115,N_12939);
nand U13820 (N_13820,N_12803,N_13081);
nand U13821 (N_13821,N_13247,N_12953);
xor U13822 (N_13822,N_13385,N_13290);
and U13823 (N_13823,N_12940,N_13390);
nor U13824 (N_13824,N_13168,N_13252);
nand U13825 (N_13825,N_13528,N_13406);
and U13826 (N_13826,N_13358,N_12899);
and U13827 (N_13827,N_13419,N_13563);
nand U13828 (N_13828,N_12929,N_13393);
nor U13829 (N_13829,N_13540,N_13479);
nor U13830 (N_13830,N_12924,N_13276);
and U13831 (N_13831,N_13339,N_13330);
or U13832 (N_13832,N_12976,N_13593);
and U13833 (N_13833,N_13073,N_13535);
nor U13834 (N_13834,N_13228,N_13571);
xnor U13835 (N_13835,N_13585,N_12854);
nor U13836 (N_13836,N_13589,N_13596);
and U13837 (N_13837,N_13048,N_13317);
nor U13838 (N_13838,N_13162,N_12806);
and U13839 (N_13839,N_13141,N_12991);
nor U13840 (N_13840,N_13230,N_12886);
or U13841 (N_13841,N_13022,N_12920);
or U13842 (N_13842,N_13007,N_12937);
and U13843 (N_13843,N_13458,N_13171);
xor U13844 (N_13844,N_12902,N_12923);
nand U13845 (N_13845,N_13150,N_13014);
and U13846 (N_13846,N_13580,N_13310);
or U13847 (N_13847,N_13044,N_13321);
or U13848 (N_13848,N_13353,N_13254);
nor U13849 (N_13849,N_13183,N_12944);
and U13850 (N_13850,N_13032,N_13059);
xor U13851 (N_13851,N_13289,N_13264);
and U13852 (N_13852,N_13027,N_13485);
and U13853 (N_13853,N_12869,N_13454);
xor U13854 (N_13854,N_13361,N_13190);
or U13855 (N_13855,N_12862,N_13581);
or U13856 (N_13856,N_13484,N_13260);
nand U13857 (N_13857,N_13423,N_12901);
and U13858 (N_13858,N_12827,N_13495);
xnor U13859 (N_13859,N_12925,N_13373);
or U13860 (N_13860,N_13489,N_12904);
nor U13861 (N_13861,N_13251,N_13359);
xor U13862 (N_13862,N_13174,N_13176);
and U13863 (N_13863,N_13504,N_12974);
nand U13864 (N_13864,N_13149,N_13156);
nor U13865 (N_13865,N_13460,N_12987);
nor U13866 (N_13866,N_13016,N_13125);
and U13867 (N_13867,N_13520,N_13309);
nand U13868 (N_13868,N_13133,N_13160);
nand U13869 (N_13869,N_13126,N_13231);
and U13870 (N_13870,N_13217,N_13462);
nand U13871 (N_13871,N_13097,N_12819);
nand U13872 (N_13872,N_12999,N_13449);
and U13873 (N_13873,N_13576,N_13098);
nor U13874 (N_13874,N_12807,N_13055);
nand U13875 (N_13875,N_13090,N_13573);
and U13876 (N_13876,N_12935,N_12878);
nand U13877 (N_13877,N_13331,N_13459);
xor U13878 (N_13878,N_13209,N_12850);
nand U13879 (N_13879,N_13426,N_12948);
nor U13880 (N_13880,N_13069,N_13040);
nor U13881 (N_13881,N_12975,N_12932);
and U13882 (N_13882,N_13496,N_13351);
nor U13883 (N_13883,N_13129,N_13242);
or U13884 (N_13884,N_13379,N_13235);
or U13885 (N_13885,N_12831,N_13565);
nand U13886 (N_13886,N_13220,N_13175);
nor U13887 (N_13887,N_13560,N_13409);
nand U13888 (N_13888,N_12946,N_13384);
xnor U13889 (N_13889,N_13529,N_13165);
nor U13890 (N_13890,N_13537,N_13598);
xor U13891 (N_13891,N_13444,N_13536);
nor U13892 (N_13892,N_13238,N_12802);
nand U13893 (N_13893,N_13428,N_12964);
or U13894 (N_13894,N_13114,N_13349);
nor U13895 (N_13895,N_13325,N_13292);
and U13896 (N_13896,N_13296,N_13313);
or U13897 (N_13897,N_13021,N_12938);
or U13898 (N_13898,N_13061,N_13487);
xnor U13899 (N_13899,N_12851,N_13417);
xor U13900 (N_13900,N_12881,N_13415);
and U13901 (N_13901,N_13151,N_12995);
nor U13902 (N_13902,N_13042,N_13430);
nor U13903 (N_13903,N_13564,N_12956);
nor U13904 (N_13904,N_12926,N_13132);
xor U13905 (N_13905,N_13244,N_13410);
and U13906 (N_13906,N_12813,N_13223);
or U13907 (N_13907,N_13224,N_13527);
nand U13908 (N_13908,N_13360,N_13414);
nand U13909 (N_13909,N_13303,N_12865);
nand U13910 (N_13910,N_12890,N_13451);
and U13911 (N_13911,N_13382,N_12877);
nor U13912 (N_13912,N_13270,N_12888);
and U13913 (N_13913,N_13186,N_12908);
or U13914 (N_13914,N_13030,N_13332);
and U13915 (N_13915,N_12949,N_13026);
xnor U13916 (N_13916,N_12848,N_13368);
xor U13917 (N_13917,N_13515,N_13253);
nand U13918 (N_13918,N_13194,N_13464);
nor U13919 (N_13919,N_13448,N_13400);
or U13920 (N_13920,N_13074,N_13583);
and U13921 (N_13921,N_13094,N_12927);
or U13922 (N_13922,N_13326,N_12843);
xor U13923 (N_13923,N_13272,N_12994);
xor U13924 (N_13924,N_12928,N_13533);
xor U13925 (N_13925,N_13096,N_13466);
and U13926 (N_13926,N_13195,N_12839);
or U13927 (N_13927,N_13239,N_13246);
or U13928 (N_13928,N_13491,N_13153);
nor U13929 (N_13929,N_13068,N_13335);
nor U13930 (N_13930,N_13486,N_12876);
xor U13931 (N_13931,N_13106,N_12820);
or U13932 (N_13932,N_13526,N_13071);
or U13933 (N_13933,N_13080,N_13058);
or U13934 (N_13934,N_13015,N_13342);
and U13935 (N_13935,N_13065,N_13315);
and U13936 (N_13936,N_12880,N_13093);
nand U13937 (N_13937,N_13371,N_13364);
nand U13938 (N_13938,N_13465,N_12960);
nand U13939 (N_13939,N_12855,N_13470);
nor U13940 (N_13940,N_13312,N_13503);
nand U13941 (N_13941,N_12838,N_12933);
nor U13942 (N_13942,N_12910,N_13054);
and U13943 (N_13943,N_13039,N_13316);
or U13944 (N_13944,N_13340,N_13418);
nor U13945 (N_13945,N_12870,N_12931);
and U13946 (N_13946,N_13201,N_13530);
or U13947 (N_13947,N_13020,N_12942);
and U13948 (N_13948,N_13594,N_12801);
nand U13949 (N_13949,N_13278,N_12822);
or U13950 (N_13950,N_13154,N_13457);
xnor U13951 (N_13951,N_13001,N_13177);
or U13952 (N_13952,N_12846,N_13443);
xnor U13953 (N_13953,N_13041,N_13468);
xnor U13954 (N_13954,N_12800,N_13070);
or U13955 (N_13955,N_13164,N_13136);
and U13956 (N_13956,N_13586,N_12966);
or U13957 (N_13957,N_12943,N_13060);
xor U13958 (N_13958,N_13478,N_12836);
nand U13959 (N_13959,N_13049,N_12826);
xor U13960 (N_13960,N_12957,N_13210);
nor U13961 (N_13961,N_13380,N_12972);
nand U13962 (N_13962,N_13567,N_12837);
nor U13963 (N_13963,N_13304,N_12989);
and U13964 (N_13964,N_13017,N_13499);
xor U13965 (N_13965,N_13433,N_13308);
or U13966 (N_13966,N_13064,N_12818);
nor U13967 (N_13967,N_13295,N_13037);
and U13968 (N_13968,N_13578,N_13214);
or U13969 (N_13969,N_12824,N_13412);
and U13970 (N_13970,N_13447,N_13045);
nand U13971 (N_13971,N_13509,N_13469);
and U13972 (N_13972,N_12986,N_13181);
xor U13973 (N_13973,N_13366,N_13411);
nor U13974 (N_13974,N_13279,N_12892);
nand U13975 (N_13975,N_13516,N_12814);
or U13976 (N_13976,N_12815,N_12984);
nand U13977 (N_13977,N_13105,N_12997);
and U13978 (N_13978,N_13402,N_13255);
or U13979 (N_13979,N_13455,N_12833);
xor U13980 (N_13980,N_13539,N_12971);
and U13981 (N_13981,N_13347,N_13525);
nand U13982 (N_13982,N_12982,N_13374);
nor U13983 (N_13983,N_13052,N_13490);
and U13984 (N_13984,N_12934,N_13324);
xor U13985 (N_13985,N_13442,N_13285);
xnor U13986 (N_13986,N_13508,N_13482);
nor U13987 (N_13987,N_13248,N_13208);
or U13988 (N_13988,N_12916,N_12909);
xor U13989 (N_13989,N_12969,N_13033);
or U13990 (N_13990,N_13211,N_13319);
or U13991 (N_13991,N_13111,N_13572);
or U13992 (N_13992,N_13546,N_12810);
and U13993 (N_13993,N_13434,N_13178);
or U13994 (N_13994,N_12832,N_13597);
xor U13995 (N_13995,N_13122,N_13188);
or U13996 (N_13996,N_13481,N_12959);
nand U13997 (N_13997,N_13477,N_12996);
xor U13998 (N_13998,N_13318,N_13024);
nor U13999 (N_13999,N_13124,N_13142);
nor U14000 (N_14000,N_13009,N_13515);
xnor U14001 (N_14001,N_13123,N_13256);
nor U14002 (N_14002,N_12863,N_13031);
or U14003 (N_14003,N_13248,N_13445);
and U14004 (N_14004,N_13368,N_12976);
or U14005 (N_14005,N_12965,N_12802);
or U14006 (N_14006,N_13034,N_12857);
nor U14007 (N_14007,N_12891,N_13331);
and U14008 (N_14008,N_13148,N_12940);
and U14009 (N_14009,N_13373,N_13402);
nand U14010 (N_14010,N_13450,N_13108);
xor U14011 (N_14011,N_13373,N_13561);
xnor U14012 (N_14012,N_13538,N_12821);
nor U14013 (N_14013,N_13558,N_13085);
and U14014 (N_14014,N_13544,N_12872);
nor U14015 (N_14015,N_13370,N_13533);
nand U14016 (N_14016,N_12854,N_13489);
xnor U14017 (N_14017,N_13095,N_13105);
nor U14018 (N_14018,N_13285,N_13170);
xnor U14019 (N_14019,N_13208,N_13485);
nor U14020 (N_14020,N_13280,N_12882);
nand U14021 (N_14021,N_13182,N_13486);
nor U14022 (N_14022,N_13282,N_13062);
and U14023 (N_14023,N_13114,N_12918);
nor U14024 (N_14024,N_12957,N_12906);
xnor U14025 (N_14025,N_12902,N_13580);
nand U14026 (N_14026,N_13301,N_13120);
xnor U14027 (N_14027,N_13396,N_13540);
xor U14028 (N_14028,N_13321,N_13107);
and U14029 (N_14029,N_13083,N_12999);
xnor U14030 (N_14030,N_13252,N_13006);
nand U14031 (N_14031,N_12934,N_12825);
and U14032 (N_14032,N_13344,N_13451);
nor U14033 (N_14033,N_13320,N_13128);
or U14034 (N_14034,N_13031,N_13455);
and U14035 (N_14035,N_13262,N_12903);
and U14036 (N_14036,N_13434,N_13281);
nor U14037 (N_14037,N_13572,N_12801);
nor U14038 (N_14038,N_12947,N_13388);
or U14039 (N_14039,N_12872,N_13016);
nand U14040 (N_14040,N_13056,N_13344);
nor U14041 (N_14041,N_13145,N_13459);
nor U14042 (N_14042,N_13042,N_13089);
nand U14043 (N_14043,N_12832,N_12887);
or U14044 (N_14044,N_13003,N_13210);
nor U14045 (N_14045,N_12802,N_13388);
and U14046 (N_14046,N_13193,N_12876);
xnor U14047 (N_14047,N_13516,N_13480);
or U14048 (N_14048,N_12834,N_13339);
xor U14049 (N_14049,N_13049,N_12966);
and U14050 (N_14050,N_12816,N_13547);
nor U14051 (N_14051,N_12810,N_13399);
or U14052 (N_14052,N_13566,N_13441);
nor U14053 (N_14053,N_13096,N_13181);
nand U14054 (N_14054,N_13183,N_12834);
nor U14055 (N_14055,N_13490,N_13557);
nor U14056 (N_14056,N_13235,N_13117);
and U14057 (N_14057,N_13419,N_13048);
xor U14058 (N_14058,N_13054,N_13415);
or U14059 (N_14059,N_13089,N_13198);
and U14060 (N_14060,N_13549,N_13299);
xor U14061 (N_14061,N_12928,N_13055);
or U14062 (N_14062,N_13522,N_13170);
nand U14063 (N_14063,N_13458,N_13262);
or U14064 (N_14064,N_13581,N_13544);
nor U14065 (N_14065,N_13124,N_12882);
nand U14066 (N_14066,N_13190,N_13285);
xor U14067 (N_14067,N_13054,N_12934);
or U14068 (N_14068,N_13461,N_13415);
nand U14069 (N_14069,N_13025,N_13146);
and U14070 (N_14070,N_12892,N_12886);
nand U14071 (N_14071,N_12885,N_13262);
nor U14072 (N_14072,N_13234,N_12809);
nand U14073 (N_14073,N_13592,N_13465);
nand U14074 (N_14074,N_12847,N_13312);
nand U14075 (N_14075,N_13184,N_13047);
nand U14076 (N_14076,N_12885,N_13279);
xnor U14077 (N_14077,N_13286,N_12955);
nor U14078 (N_14078,N_13327,N_13537);
nand U14079 (N_14079,N_13332,N_13368);
and U14080 (N_14080,N_12888,N_13018);
or U14081 (N_14081,N_12909,N_12991);
nor U14082 (N_14082,N_13122,N_12897);
and U14083 (N_14083,N_12880,N_13192);
xor U14084 (N_14084,N_13068,N_13584);
xnor U14085 (N_14085,N_13109,N_13544);
nor U14086 (N_14086,N_13514,N_12859);
and U14087 (N_14087,N_13339,N_13424);
nand U14088 (N_14088,N_12975,N_13470);
or U14089 (N_14089,N_13489,N_13511);
xnor U14090 (N_14090,N_13337,N_13014);
or U14091 (N_14091,N_13049,N_13556);
xnor U14092 (N_14092,N_13165,N_12820);
xnor U14093 (N_14093,N_13021,N_13572);
xor U14094 (N_14094,N_13104,N_13069);
nor U14095 (N_14095,N_13035,N_13117);
nor U14096 (N_14096,N_13554,N_13021);
nand U14097 (N_14097,N_12926,N_12828);
or U14098 (N_14098,N_13274,N_13381);
nor U14099 (N_14099,N_13524,N_13337);
or U14100 (N_14100,N_12865,N_13263);
xnor U14101 (N_14101,N_13222,N_12941);
or U14102 (N_14102,N_12866,N_12991);
and U14103 (N_14103,N_12819,N_13010);
xor U14104 (N_14104,N_12808,N_13070);
or U14105 (N_14105,N_12982,N_13191);
xor U14106 (N_14106,N_13599,N_13033);
nand U14107 (N_14107,N_13301,N_13379);
or U14108 (N_14108,N_13107,N_13588);
nor U14109 (N_14109,N_13552,N_13304);
xnor U14110 (N_14110,N_12934,N_12811);
or U14111 (N_14111,N_13504,N_12847);
and U14112 (N_14112,N_13160,N_13283);
nor U14113 (N_14113,N_13456,N_12805);
or U14114 (N_14114,N_13547,N_13194);
xor U14115 (N_14115,N_13168,N_13045);
nand U14116 (N_14116,N_13070,N_12911);
nand U14117 (N_14117,N_13294,N_13396);
xor U14118 (N_14118,N_13004,N_13260);
nand U14119 (N_14119,N_13411,N_13400);
nand U14120 (N_14120,N_12930,N_13519);
and U14121 (N_14121,N_13113,N_12883);
xor U14122 (N_14122,N_13449,N_13322);
nor U14123 (N_14123,N_13019,N_13196);
nor U14124 (N_14124,N_13169,N_13413);
xnor U14125 (N_14125,N_12882,N_13335);
xor U14126 (N_14126,N_13087,N_12881);
and U14127 (N_14127,N_13274,N_13266);
nor U14128 (N_14128,N_13245,N_13178);
nor U14129 (N_14129,N_13011,N_13427);
nor U14130 (N_14130,N_12801,N_13506);
or U14131 (N_14131,N_13449,N_12976);
and U14132 (N_14132,N_13216,N_13260);
nor U14133 (N_14133,N_12983,N_13104);
nor U14134 (N_14134,N_13153,N_13587);
and U14135 (N_14135,N_13241,N_13403);
nor U14136 (N_14136,N_13329,N_12875);
and U14137 (N_14137,N_13075,N_13192);
nand U14138 (N_14138,N_13167,N_13598);
and U14139 (N_14139,N_13013,N_13437);
or U14140 (N_14140,N_12853,N_12848);
nand U14141 (N_14141,N_13053,N_13594);
or U14142 (N_14142,N_13585,N_13026);
nor U14143 (N_14143,N_12895,N_13420);
nand U14144 (N_14144,N_13108,N_12873);
xnor U14145 (N_14145,N_13275,N_13441);
nor U14146 (N_14146,N_13266,N_13093);
or U14147 (N_14147,N_13407,N_12961);
nand U14148 (N_14148,N_13528,N_13081);
xnor U14149 (N_14149,N_13328,N_13200);
xnor U14150 (N_14150,N_13459,N_13074);
nor U14151 (N_14151,N_12974,N_13488);
and U14152 (N_14152,N_13160,N_12910);
nor U14153 (N_14153,N_12978,N_13370);
and U14154 (N_14154,N_13097,N_13036);
and U14155 (N_14155,N_13278,N_13509);
nand U14156 (N_14156,N_12929,N_12878);
xor U14157 (N_14157,N_13569,N_12868);
and U14158 (N_14158,N_12808,N_13464);
nand U14159 (N_14159,N_13466,N_12948);
nor U14160 (N_14160,N_12978,N_12830);
xor U14161 (N_14161,N_13529,N_12918);
nor U14162 (N_14162,N_12884,N_13330);
nand U14163 (N_14163,N_13467,N_13043);
and U14164 (N_14164,N_13196,N_13246);
or U14165 (N_14165,N_13409,N_13438);
and U14166 (N_14166,N_12879,N_13363);
or U14167 (N_14167,N_12815,N_13459);
nor U14168 (N_14168,N_13147,N_13508);
and U14169 (N_14169,N_13192,N_13562);
xnor U14170 (N_14170,N_13250,N_13331);
or U14171 (N_14171,N_13481,N_13579);
or U14172 (N_14172,N_13549,N_13276);
nor U14173 (N_14173,N_13520,N_12800);
nor U14174 (N_14174,N_12827,N_12890);
or U14175 (N_14175,N_13350,N_12941);
xnor U14176 (N_14176,N_13248,N_13225);
nor U14177 (N_14177,N_13071,N_13086);
xor U14178 (N_14178,N_13413,N_13519);
nor U14179 (N_14179,N_13142,N_13115);
xor U14180 (N_14180,N_13144,N_13398);
or U14181 (N_14181,N_13253,N_13381);
nor U14182 (N_14182,N_13112,N_13026);
xor U14183 (N_14183,N_13472,N_13259);
nor U14184 (N_14184,N_13080,N_13033);
nand U14185 (N_14185,N_13097,N_12828);
nand U14186 (N_14186,N_13403,N_13444);
and U14187 (N_14187,N_13185,N_12947);
nor U14188 (N_14188,N_13517,N_12959);
nor U14189 (N_14189,N_12839,N_13015);
nor U14190 (N_14190,N_13417,N_13175);
nand U14191 (N_14191,N_13301,N_13217);
and U14192 (N_14192,N_13162,N_13317);
or U14193 (N_14193,N_13147,N_12828);
nand U14194 (N_14194,N_13052,N_12938);
xor U14195 (N_14195,N_12854,N_12891);
nand U14196 (N_14196,N_13595,N_12866);
or U14197 (N_14197,N_13096,N_12877);
or U14198 (N_14198,N_13335,N_13271);
nor U14199 (N_14199,N_13527,N_13306);
nand U14200 (N_14200,N_13090,N_13165);
nand U14201 (N_14201,N_13119,N_13081);
xnor U14202 (N_14202,N_13549,N_12861);
or U14203 (N_14203,N_13304,N_12855);
xor U14204 (N_14204,N_12890,N_13072);
xor U14205 (N_14205,N_12831,N_12921);
and U14206 (N_14206,N_12913,N_13337);
nand U14207 (N_14207,N_13285,N_13421);
xor U14208 (N_14208,N_12843,N_13131);
xnor U14209 (N_14209,N_13316,N_13161);
or U14210 (N_14210,N_13358,N_13364);
xnor U14211 (N_14211,N_12817,N_13535);
nor U14212 (N_14212,N_13587,N_13232);
and U14213 (N_14213,N_13128,N_13574);
or U14214 (N_14214,N_13146,N_13139);
and U14215 (N_14215,N_13268,N_13425);
nor U14216 (N_14216,N_12979,N_13457);
nand U14217 (N_14217,N_13565,N_13036);
nor U14218 (N_14218,N_12991,N_13384);
nor U14219 (N_14219,N_13597,N_12993);
nand U14220 (N_14220,N_13169,N_12980);
xor U14221 (N_14221,N_13496,N_13006);
or U14222 (N_14222,N_13352,N_13021);
nand U14223 (N_14223,N_12962,N_12848);
nand U14224 (N_14224,N_12900,N_12814);
or U14225 (N_14225,N_12917,N_12983);
or U14226 (N_14226,N_13272,N_13070);
nand U14227 (N_14227,N_13510,N_13092);
and U14228 (N_14228,N_13487,N_13464);
and U14229 (N_14229,N_13489,N_12877);
and U14230 (N_14230,N_13440,N_12939);
nor U14231 (N_14231,N_13254,N_13538);
nor U14232 (N_14232,N_13416,N_13384);
and U14233 (N_14233,N_12869,N_12939);
nor U14234 (N_14234,N_12959,N_13544);
nor U14235 (N_14235,N_12821,N_13211);
or U14236 (N_14236,N_13349,N_12865);
or U14237 (N_14237,N_13362,N_13414);
nand U14238 (N_14238,N_13242,N_13091);
or U14239 (N_14239,N_13061,N_13078);
or U14240 (N_14240,N_13163,N_12984);
nor U14241 (N_14241,N_13238,N_12826);
nand U14242 (N_14242,N_12906,N_13089);
xnor U14243 (N_14243,N_13481,N_13466);
xnor U14244 (N_14244,N_13308,N_13459);
nand U14245 (N_14245,N_13533,N_13079);
nor U14246 (N_14246,N_13330,N_13491);
or U14247 (N_14247,N_13117,N_13576);
and U14248 (N_14248,N_12931,N_13492);
nand U14249 (N_14249,N_12912,N_13038);
or U14250 (N_14250,N_13464,N_13088);
xor U14251 (N_14251,N_13559,N_12900);
xor U14252 (N_14252,N_12985,N_12995);
nor U14253 (N_14253,N_13483,N_13274);
xor U14254 (N_14254,N_12896,N_13451);
xnor U14255 (N_14255,N_13525,N_12978);
and U14256 (N_14256,N_13442,N_13059);
or U14257 (N_14257,N_13494,N_12817);
and U14258 (N_14258,N_13579,N_13391);
and U14259 (N_14259,N_13366,N_13341);
nand U14260 (N_14260,N_13103,N_13078);
or U14261 (N_14261,N_12908,N_12966);
nand U14262 (N_14262,N_13266,N_13547);
nand U14263 (N_14263,N_13448,N_12966);
and U14264 (N_14264,N_13366,N_13391);
nor U14265 (N_14265,N_13318,N_13008);
or U14266 (N_14266,N_12867,N_12978);
nor U14267 (N_14267,N_13267,N_13246);
nor U14268 (N_14268,N_12942,N_13345);
xnor U14269 (N_14269,N_13079,N_13580);
nor U14270 (N_14270,N_13048,N_13040);
nand U14271 (N_14271,N_13076,N_13244);
nor U14272 (N_14272,N_13490,N_13202);
or U14273 (N_14273,N_13052,N_13061);
and U14274 (N_14274,N_13178,N_13572);
and U14275 (N_14275,N_13261,N_12823);
nor U14276 (N_14276,N_13275,N_13438);
nand U14277 (N_14277,N_12936,N_13431);
xor U14278 (N_14278,N_12833,N_13210);
and U14279 (N_14279,N_13248,N_13036);
or U14280 (N_14280,N_13268,N_12896);
and U14281 (N_14281,N_13293,N_13281);
nand U14282 (N_14282,N_13505,N_13535);
and U14283 (N_14283,N_12942,N_12983);
and U14284 (N_14284,N_13078,N_13162);
nor U14285 (N_14285,N_12919,N_13252);
or U14286 (N_14286,N_13065,N_12854);
nand U14287 (N_14287,N_13182,N_12813);
nor U14288 (N_14288,N_13571,N_13562);
nand U14289 (N_14289,N_13250,N_13509);
nor U14290 (N_14290,N_13309,N_12852);
nor U14291 (N_14291,N_13338,N_13433);
nor U14292 (N_14292,N_12861,N_13097);
xor U14293 (N_14293,N_13091,N_13273);
nor U14294 (N_14294,N_13567,N_12844);
nand U14295 (N_14295,N_13230,N_13520);
or U14296 (N_14296,N_13037,N_13028);
nand U14297 (N_14297,N_13010,N_12927);
or U14298 (N_14298,N_12917,N_13196);
nand U14299 (N_14299,N_12934,N_13166);
nand U14300 (N_14300,N_13295,N_13474);
nor U14301 (N_14301,N_13368,N_12811);
nor U14302 (N_14302,N_13497,N_13173);
xor U14303 (N_14303,N_12908,N_13346);
and U14304 (N_14304,N_13427,N_13543);
or U14305 (N_14305,N_13597,N_13476);
nor U14306 (N_14306,N_13129,N_13509);
xor U14307 (N_14307,N_13598,N_12859);
and U14308 (N_14308,N_13230,N_13394);
nor U14309 (N_14309,N_12840,N_12974);
and U14310 (N_14310,N_12966,N_13237);
nand U14311 (N_14311,N_13100,N_13483);
nor U14312 (N_14312,N_12978,N_13282);
and U14313 (N_14313,N_12908,N_12946);
and U14314 (N_14314,N_13579,N_13441);
xor U14315 (N_14315,N_13004,N_13559);
or U14316 (N_14316,N_12801,N_13575);
nand U14317 (N_14317,N_12918,N_13062);
xnor U14318 (N_14318,N_12863,N_13014);
or U14319 (N_14319,N_13529,N_13191);
or U14320 (N_14320,N_13421,N_12961);
nand U14321 (N_14321,N_13593,N_13350);
xor U14322 (N_14322,N_13133,N_13422);
nand U14323 (N_14323,N_13163,N_13376);
nand U14324 (N_14324,N_13262,N_12806);
and U14325 (N_14325,N_13169,N_13232);
xor U14326 (N_14326,N_13342,N_13107);
and U14327 (N_14327,N_13071,N_13383);
or U14328 (N_14328,N_13241,N_12823);
xor U14329 (N_14329,N_13591,N_13371);
and U14330 (N_14330,N_13016,N_13104);
and U14331 (N_14331,N_13386,N_13283);
or U14332 (N_14332,N_13559,N_13068);
and U14333 (N_14333,N_13270,N_13401);
nand U14334 (N_14334,N_13311,N_13270);
and U14335 (N_14335,N_13599,N_13512);
xnor U14336 (N_14336,N_13363,N_12887);
nand U14337 (N_14337,N_13454,N_13354);
nand U14338 (N_14338,N_13010,N_12945);
xnor U14339 (N_14339,N_12878,N_13427);
nand U14340 (N_14340,N_12838,N_12944);
nor U14341 (N_14341,N_13428,N_13109);
nor U14342 (N_14342,N_13554,N_13242);
nand U14343 (N_14343,N_12946,N_13517);
xor U14344 (N_14344,N_13537,N_13265);
and U14345 (N_14345,N_13018,N_13149);
xor U14346 (N_14346,N_13446,N_12893);
and U14347 (N_14347,N_12928,N_13378);
xor U14348 (N_14348,N_13420,N_12805);
nand U14349 (N_14349,N_13176,N_12812);
and U14350 (N_14350,N_12927,N_12917);
or U14351 (N_14351,N_13237,N_13262);
or U14352 (N_14352,N_13177,N_12956);
or U14353 (N_14353,N_13424,N_13170);
and U14354 (N_14354,N_13588,N_12847);
or U14355 (N_14355,N_13166,N_13464);
nor U14356 (N_14356,N_13160,N_13074);
nor U14357 (N_14357,N_13165,N_12866);
xor U14358 (N_14358,N_12880,N_13370);
xor U14359 (N_14359,N_12849,N_13047);
nor U14360 (N_14360,N_13579,N_13583);
nor U14361 (N_14361,N_12871,N_12897);
nand U14362 (N_14362,N_13083,N_13066);
or U14363 (N_14363,N_13343,N_13263);
nor U14364 (N_14364,N_13407,N_13063);
and U14365 (N_14365,N_13455,N_13599);
nand U14366 (N_14366,N_12953,N_13200);
or U14367 (N_14367,N_13104,N_13447);
xor U14368 (N_14368,N_12974,N_13123);
nand U14369 (N_14369,N_13344,N_13007);
nor U14370 (N_14370,N_13590,N_13425);
nor U14371 (N_14371,N_13507,N_13489);
nand U14372 (N_14372,N_13412,N_13526);
nor U14373 (N_14373,N_13004,N_12853);
xnor U14374 (N_14374,N_13044,N_13067);
or U14375 (N_14375,N_13257,N_13544);
and U14376 (N_14376,N_13503,N_13598);
xor U14377 (N_14377,N_13529,N_13064);
and U14378 (N_14378,N_13001,N_13548);
nand U14379 (N_14379,N_13189,N_13243);
nand U14380 (N_14380,N_13015,N_13240);
xnor U14381 (N_14381,N_13499,N_12944);
and U14382 (N_14382,N_13068,N_12928);
xnor U14383 (N_14383,N_13169,N_12811);
nor U14384 (N_14384,N_13253,N_13096);
or U14385 (N_14385,N_12981,N_13143);
nand U14386 (N_14386,N_13424,N_12986);
or U14387 (N_14387,N_13117,N_13347);
and U14388 (N_14388,N_13038,N_13386);
and U14389 (N_14389,N_12951,N_13598);
xor U14390 (N_14390,N_12965,N_13240);
and U14391 (N_14391,N_13061,N_12808);
or U14392 (N_14392,N_13271,N_13364);
or U14393 (N_14393,N_13146,N_13457);
nor U14394 (N_14394,N_13098,N_13447);
and U14395 (N_14395,N_12856,N_13305);
xor U14396 (N_14396,N_13110,N_13242);
xnor U14397 (N_14397,N_13534,N_13596);
or U14398 (N_14398,N_12892,N_13143);
and U14399 (N_14399,N_13372,N_12968);
nor U14400 (N_14400,N_13998,N_13651);
nor U14401 (N_14401,N_13896,N_14304);
nor U14402 (N_14402,N_13795,N_14299);
nor U14403 (N_14403,N_13758,N_14210);
nand U14404 (N_14404,N_14390,N_13800);
or U14405 (N_14405,N_14115,N_13649);
or U14406 (N_14406,N_13618,N_14102);
and U14407 (N_14407,N_14131,N_14176);
xor U14408 (N_14408,N_13947,N_14193);
and U14409 (N_14409,N_13636,N_13619);
nand U14410 (N_14410,N_13993,N_14301);
xor U14411 (N_14411,N_13981,N_13767);
xnor U14412 (N_14412,N_13796,N_13970);
and U14413 (N_14413,N_14212,N_14114);
nor U14414 (N_14414,N_14024,N_13695);
and U14415 (N_14415,N_14388,N_13992);
xnor U14416 (N_14416,N_14311,N_13644);
or U14417 (N_14417,N_14044,N_14042);
nor U14418 (N_14418,N_13664,N_14209);
or U14419 (N_14419,N_13741,N_13804);
or U14420 (N_14420,N_13931,N_14262);
or U14421 (N_14421,N_14089,N_13916);
nand U14422 (N_14422,N_13726,N_13824);
or U14423 (N_14423,N_14256,N_13831);
or U14424 (N_14424,N_13703,N_14368);
xor U14425 (N_14425,N_14317,N_14218);
nand U14426 (N_14426,N_14387,N_14070);
or U14427 (N_14427,N_13958,N_14330);
or U14428 (N_14428,N_14118,N_14345);
nor U14429 (N_14429,N_13748,N_14075);
and U14430 (N_14430,N_14147,N_13754);
nor U14431 (N_14431,N_14276,N_13629);
nor U14432 (N_14432,N_14026,N_14049);
nand U14433 (N_14433,N_14116,N_14288);
and U14434 (N_14434,N_14383,N_14393);
nand U14435 (N_14435,N_13983,N_13708);
or U14436 (N_14436,N_14214,N_13766);
nor U14437 (N_14437,N_13728,N_13773);
and U14438 (N_14438,N_13731,N_13660);
xnor U14439 (N_14439,N_14028,N_13975);
and U14440 (N_14440,N_14015,N_14352);
or U14441 (N_14441,N_13980,N_14162);
and U14442 (N_14442,N_14012,N_13829);
and U14443 (N_14443,N_13878,N_13915);
or U14444 (N_14444,N_13871,N_14260);
nand U14445 (N_14445,N_14053,N_13968);
and U14446 (N_14446,N_14084,N_13909);
or U14447 (N_14447,N_13906,N_13682);
and U14448 (N_14448,N_13756,N_13976);
and U14449 (N_14449,N_13715,N_13768);
and U14450 (N_14450,N_13633,N_13605);
nand U14451 (N_14451,N_14341,N_13938);
nor U14452 (N_14452,N_14382,N_14291);
or U14453 (N_14453,N_14302,N_14211);
xor U14454 (N_14454,N_14106,N_13886);
or U14455 (N_14455,N_14050,N_13806);
nor U14456 (N_14456,N_13902,N_13784);
or U14457 (N_14457,N_14000,N_13630);
nand U14458 (N_14458,N_13600,N_14223);
xor U14459 (N_14459,N_14303,N_13639);
nand U14460 (N_14460,N_13617,N_13780);
or U14461 (N_14461,N_14006,N_14194);
and U14462 (N_14462,N_13716,N_14354);
nor U14463 (N_14463,N_13683,N_13720);
nor U14464 (N_14464,N_13872,N_13788);
xor U14465 (N_14465,N_13930,N_13765);
or U14466 (N_14466,N_13815,N_14229);
or U14467 (N_14467,N_14021,N_13620);
nor U14468 (N_14468,N_14230,N_13881);
and U14469 (N_14469,N_14280,N_14191);
nand U14470 (N_14470,N_14271,N_13727);
and U14471 (N_14471,N_14222,N_14142);
and U14472 (N_14472,N_13974,N_13949);
nand U14473 (N_14473,N_13862,N_14016);
nand U14474 (N_14474,N_13730,N_13899);
or U14475 (N_14475,N_14380,N_14134);
nand U14476 (N_14476,N_14047,N_14033);
and U14477 (N_14477,N_14083,N_14157);
or U14478 (N_14478,N_14346,N_14051);
xor U14479 (N_14479,N_13671,N_14321);
nor U14480 (N_14480,N_13696,N_14257);
xor U14481 (N_14481,N_14158,N_13688);
and U14482 (N_14482,N_14272,N_14248);
nor U14483 (N_14483,N_13616,N_14129);
nor U14484 (N_14484,N_13951,N_14367);
nand U14485 (N_14485,N_14150,N_14043);
or U14486 (N_14486,N_14245,N_13865);
nand U14487 (N_14487,N_14228,N_13857);
xor U14488 (N_14488,N_13954,N_13833);
or U14489 (N_14489,N_14067,N_13655);
or U14490 (N_14490,N_14079,N_14011);
nor U14491 (N_14491,N_14323,N_14001);
and U14492 (N_14492,N_14363,N_14225);
or U14493 (N_14493,N_14025,N_13609);
and U14494 (N_14494,N_13904,N_14105);
nand U14495 (N_14495,N_13681,N_14078);
and U14496 (N_14496,N_13685,N_14349);
nand U14497 (N_14497,N_13903,N_13747);
or U14498 (N_14498,N_14253,N_13739);
and U14499 (N_14499,N_13876,N_14278);
xor U14500 (N_14500,N_14018,N_13837);
or U14501 (N_14501,N_13613,N_14375);
or U14502 (N_14502,N_14156,N_13835);
and U14503 (N_14503,N_14076,N_14139);
and U14504 (N_14504,N_14263,N_13950);
and U14505 (N_14505,N_13694,N_13604);
nor U14506 (N_14506,N_14313,N_14013);
nor U14507 (N_14507,N_13999,N_13866);
nand U14508 (N_14508,N_13805,N_13812);
xor U14509 (N_14509,N_13803,N_13926);
or U14510 (N_14510,N_14316,N_13789);
nor U14511 (N_14511,N_13777,N_13661);
or U14512 (N_14512,N_13953,N_13973);
nor U14513 (N_14513,N_14241,N_14003);
or U14514 (N_14514,N_13791,N_13676);
nor U14515 (N_14515,N_14029,N_14334);
and U14516 (N_14516,N_13704,N_14054);
and U14517 (N_14517,N_14374,N_13891);
nor U14518 (N_14518,N_14154,N_13853);
nor U14519 (N_14519,N_13670,N_13971);
xnor U14520 (N_14520,N_13922,N_14133);
and U14521 (N_14521,N_13735,N_14231);
xnor U14522 (N_14522,N_14169,N_14037);
and U14523 (N_14523,N_13810,N_14357);
xnor U14524 (N_14524,N_14166,N_14252);
nand U14525 (N_14525,N_13924,N_14216);
nor U14526 (N_14526,N_13989,N_13624);
nand U14527 (N_14527,N_14200,N_14358);
xor U14528 (N_14528,N_14219,N_13729);
or U14529 (N_14529,N_13880,N_13920);
and U14530 (N_14530,N_14347,N_14127);
nor U14531 (N_14531,N_13850,N_13742);
nor U14532 (N_14532,N_13858,N_13937);
nand U14533 (N_14533,N_13634,N_14074);
or U14534 (N_14534,N_14058,N_13622);
xnor U14535 (N_14535,N_13801,N_14277);
nand U14536 (N_14536,N_13816,N_14395);
nand U14537 (N_14537,N_14073,N_14090);
nor U14538 (N_14538,N_14361,N_13840);
nor U14539 (N_14539,N_14233,N_14310);
xor U14540 (N_14540,N_13923,N_13625);
and U14541 (N_14541,N_14036,N_13652);
or U14542 (N_14542,N_14396,N_13867);
nand U14543 (N_14543,N_14199,N_13751);
nor U14544 (N_14544,N_13939,N_13809);
xor U14545 (N_14545,N_13641,N_14392);
or U14546 (N_14546,N_14389,N_14398);
and U14547 (N_14547,N_13952,N_13690);
and U14548 (N_14548,N_13884,N_14007);
and U14549 (N_14549,N_13781,N_14123);
nor U14550 (N_14550,N_14064,N_13897);
xor U14551 (N_14551,N_14226,N_14290);
xnor U14552 (N_14552,N_13755,N_13901);
or U14553 (N_14553,N_14017,N_14249);
nand U14554 (N_14554,N_14275,N_14195);
xor U14555 (N_14555,N_14239,N_14103);
nor U14556 (N_14556,N_13826,N_13945);
or U14557 (N_14557,N_13986,N_13602);
and U14558 (N_14558,N_13822,N_14250);
or U14559 (N_14559,N_13898,N_13817);
nor U14560 (N_14560,N_14258,N_14232);
and U14561 (N_14561,N_14152,N_13697);
and U14562 (N_14562,N_13699,N_14068);
and U14563 (N_14563,N_14356,N_14224);
nand U14564 (N_14564,N_14040,N_13763);
or U14565 (N_14565,N_13825,N_13959);
and U14566 (N_14566,N_13770,N_14034);
and U14567 (N_14567,N_13869,N_14052);
or U14568 (N_14568,N_13608,N_13813);
xnor U14569 (N_14569,N_13779,N_13911);
and U14570 (N_14570,N_13957,N_14082);
xor U14571 (N_14571,N_14085,N_13912);
or U14572 (N_14572,N_14137,N_13852);
nand U14573 (N_14573,N_13918,N_13787);
and U14574 (N_14574,N_14004,N_14181);
nor U14575 (N_14575,N_14071,N_14055);
and U14576 (N_14576,N_13928,N_13692);
xor U14577 (N_14577,N_14206,N_13994);
nor U14578 (N_14578,N_13723,N_13635);
nand U14579 (N_14579,N_13746,N_14038);
xor U14580 (N_14580,N_14178,N_13717);
nand U14581 (N_14581,N_13873,N_14238);
or U14582 (N_14582,N_14268,N_13962);
nor U14583 (N_14583,N_14148,N_14282);
and U14584 (N_14584,N_14295,N_13673);
xor U14585 (N_14585,N_14333,N_14377);
nand U14586 (N_14586,N_14014,N_14236);
xor U14587 (N_14587,N_14023,N_13819);
or U14588 (N_14588,N_13855,N_14286);
or U14589 (N_14589,N_13654,N_13894);
xnor U14590 (N_14590,N_14180,N_13653);
xnor U14591 (N_14591,N_13848,N_13790);
xnor U14592 (N_14592,N_13965,N_14237);
or U14593 (N_14593,N_14305,N_14246);
nor U14594 (N_14594,N_13701,N_13888);
and U14595 (N_14595,N_14332,N_13905);
or U14596 (N_14596,N_13693,N_14279);
and U14597 (N_14597,N_14360,N_13658);
nand U14598 (N_14598,N_13875,N_14160);
xnor U14599 (N_14599,N_13750,N_13808);
and U14600 (N_14600,N_14342,N_14110);
nand U14601 (N_14601,N_13623,N_13830);
nor U14602 (N_14602,N_14196,N_13882);
nand U14603 (N_14603,N_13709,N_13740);
xnor U14604 (N_14604,N_13745,N_14296);
nor U14605 (N_14605,N_14174,N_13979);
or U14606 (N_14606,N_14149,N_13820);
nor U14607 (N_14607,N_14065,N_13759);
nand U14608 (N_14608,N_14391,N_14124);
nand U14609 (N_14609,N_14372,N_13611);
nand U14610 (N_14610,N_13718,N_14066);
and U14611 (N_14611,N_14289,N_14130);
xnor U14612 (N_14612,N_13879,N_14045);
or U14613 (N_14613,N_14221,N_13985);
and U14614 (N_14614,N_14132,N_14264);
xnor U14615 (N_14615,N_14163,N_14183);
or U14616 (N_14616,N_13642,N_13782);
nand U14617 (N_14617,N_14088,N_14135);
xnor U14618 (N_14618,N_13821,N_13914);
xor U14619 (N_14619,N_13732,N_14030);
xnor U14620 (N_14620,N_13932,N_14096);
or U14621 (N_14621,N_14077,N_14197);
xnor U14622 (N_14622,N_14340,N_14143);
or U14623 (N_14623,N_13818,N_13849);
or U14624 (N_14624,N_14069,N_13612);
xnor U14625 (N_14625,N_13700,N_14121);
or U14626 (N_14626,N_13724,N_14370);
nand U14627 (N_14627,N_13771,N_13783);
and U14628 (N_14628,N_14318,N_14320);
and U14629 (N_14629,N_14161,N_13686);
nor U14630 (N_14630,N_13841,N_13778);
nand U14631 (N_14631,N_14274,N_13687);
or U14632 (N_14632,N_14351,N_13948);
nor U14633 (N_14633,N_13892,N_14273);
nand U14634 (N_14634,N_14104,N_13870);
and U14635 (N_14635,N_14022,N_14126);
nand U14636 (N_14636,N_14190,N_14101);
nand U14637 (N_14637,N_14270,N_13775);
or U14638 (N_14638,N_13793,N_13963);
nor U14639 (N_14639,N_13807,N_13843);
and U14640 (N_14640,N_13668,N_14172);
nor U14641 (N_14641,N_14329,N_14041);
xor U14642 (N_14642,N_13772,N_13764);
nand U14643 (N_14643,N_13721,N_13887);
and U14644 (N_14644,N_13614,N_14265);
and U14645 (N_14645,N_13969,N_13893);
and U14646 (N_14646,N_14005,N_13984);
and U14647 (N_14647,N_13917,N_14170);
and U14648 (N_14648,N_14056,N_13995);
nor U14649 (N_14649,N_14266,N_14240);
nand U14650 (N_14650,N_13761,N_14177);
or U14651 (N_14651,N_13854,N_13757);
nand U14652 (N_14652,N_13895,N_14086);
xnor U14653 (N_14653,N_14140,N_14173);
xor U14654 (N_14654,N_13705,N_13889);
xnor U14655 (N_14655,N_14300,N_14331);
xor U14656 (N_14656,N_14284,N_14365);
xor U14657 (N_14657,N_13603,N_14201);
nor U14658 (N_14658,N_13877,N_14247);
xor U14659 (N_14659,N_14027,N_14151);
or U14660 (N_14660,N_13734,N_13659);
nand U14661 (N_14661,N_14315,N_13799);
and U14662 (N_14662,N_14298,N_13846);
and U14663 (N_14663,N_14080,N_13900);
nand U14664 (N_14664,N_13972,N_14144);
nand U14665 (N_14665,N_13712,N_14307);
and U14666 (N_14666,N_13967,N_13607);
or U14667 (N_14667,N_14254,N_14324);
and U14668 (N_14668,N_14153,N_14048);
xnor U14669 (N_14669,N_13615,N_14159);
or U14670 (N_14670,N_13674,N_14009);
or U14671 (N_14671,N_14353,N_13811);
nor U14672 (N_14672,N_14063,N_13672);
nor U14673 (N_14673,N_13646,N_14060);
and U14674 (N_14674,N_14294,N_14072);
and U14675 (N_14675,N_13626,N_13794);
nor U14676 (N_14676,N_13698,N_13834);
and U14677 (N_14677,N_14386,N_13863);
nand U14678 (N_14678,N_14202,N_14235);
xor U14679 (N_14679,N_14204,N_14293);
nor U14680 (N_14680,N_13733,N_13785);
nand U14681 (N_14681,N_13844,N_14336);
nor U14682 (N_14682,N_14112,N_14283);
xor U14683 (N_14683,N_14227,N_13743);
nand U14684 (N_14684,N_13851,N_13944);
nor U14685 (N_14685,N_14255,N_14319);
nand U14686 (N_14686,N_14343,N_13946);
and U14687 (N_14687,N_13666,N_13606);
nand U14688 (N_14688,N_14095,N_13839);
and U14689 (N_14689,N_14186,N_14203);
and U14690 (N_14690,N_13722,N_14337);
xor U14691 (N_14691,N_14281,N_14269);
nor U14692 (N_14692,N_14355,N_14384);
nor U14693 (N_14693,N_13883,N_13689);
or U14694 (N_14694,N_13645,N_13838);
nor U14695 (N_14695,N_14192,N_14108);
nor U14696 (N_14696,N_13910,N_13956);
or U14697 (N_14697,N_14335,N_13991);
or U14698 (N_14698,N_13941,N_14189);
nand U14699 (N_14699,N_14394,N_13966);
and U14700 (N_14700,N_14184,N_13637);
and U14701 (N_14701,N_14168,N_13628);
or U14702 (N_14702,N_13977,N_14344);
xor U14703 (N_14703,N_13638,N_14031);
xnor U14704 (N_14704,N_13919,N_13913);
xor U14705 (N_14705,N_14285,N_14327);
xor U14706 (N_14706,N_14109,N_13921);
or U14707 (N_14707,N_14128,N_13665);
or U14708 (N_14708,N_14220,N_13943);
nor U14709 (N_14709,N_14259,N_14328);
or U14710 (N_14710,N_13885,N_13978);
and U14711 (N_14711,N_13601,N_14091);
or U14712 (N_14712,N_14008,N_14362);
xnor U14713 (N_14713,N_13610,N_13936);
nand U14714 (N_14714,N_14062,N_14338);
or U14715 (N_14715,N_13621,N_14187);
nor U14716 (N_14716,N_14155,N_14019);
nor U14717 (N_14717,N_13988,N_14039);
and U14718 (N_14718,N_13656,N_13760);
or U14719 (N_14719,N_13677,N_13842);
and U14720 (N_14720,N_13643,N_14359);
nand U14721 (N_14721,N_13996,N_13832);
nor U14722 (N_14722,N_13927,N_14164);
or U14723 (N_14723,N_13679,N_14242);
xnor U14724 (N_14724,N_14364,N_13762);
nand U14725 (N_14725,N_14297,N_13752);
nand U14726 (N_14726,N_14182,N_14100);
xnor U14727 (N_14727,N_14081,N_13738);
or U14728 (N_14728,N_14167,N_13702);
nand U14729 (N_14729,N_13907,N_14032);
and U14730 (N_14730,N_14120,N_13710);
nand U14731 (N_14731,N_14125,N_14308);
and U14732 (N_14732,N_14097,N_13859);
xnor U14733 (N_14733,N_13797,N_13814);
or U14734 (N_14734,N_14046,N_13935);
or U14735 (N_14735,N_13737,N_13908);
and U14736 (N_14736,N_14322,N_13802);
or U14737 (N_14737,N_14059,N_14035);
or U14738 (N_14738,N_13997,N_13684);
and U14739 (N_14739,N_14171,N_14205);
xor U14740 (N_14740,N_13990,N_14179);
nor U14741 (N_14741,N_13667,N_13934);
and U14742 (N_14742,N_13792,N_14371);
and U14743 (N_14743,N_13749,N_13964);
xnor U14744 (N_14744,N_14325,N_13678);
and U14745 (N_14745,N_14141,N_13982);
and U14746 (N_14746,N_14145,N_14348);
or U14747 (N_14747,N_13774,N_13933);
xor U14748 (N_14748,N_13657,N_14208);
xnor U14749 (N_14749,N_14350,N_13736);
nor U14750 (N_14750,N_14002,N_13868);
and U14751 (N_14751,N_14292,N_14381);
or U14752 (N_14752,N_14188,N_14113);
nor U14753 (N_14753,N_13675,N_14111);
xnor U14754 (N_14754,N_14314,N_14399);
xnor U14755 (N_14755,N_13827,N_14261);
nor U14756 (N_14756,N_14117,N_14185);
nand U14757 (N_14757,N_14138,N_14098);
or U14758 (N_14758,N_14020,N_13942);
xor U14759 (N_14759,N_13662,N_13856);
nand U14760 (N_14760,N_13961,N_14244);
and U14761 (N_14761,N_13627,N_13823);
nand U14762 (N_14762,N_14267,N_14366);
xnor U14763 (N_14763,N_14326,N_14339);
xnor U14764 (N_14764,N_14379,N_14369);
nand U14765 (N_14765,N_14234,N_13786);
and U14766 (N_14766,N_13860,N_14378);
nand U14767 (N_14767,N_14385,N_14213);
nor U14768 (N_14768,N_14122,N_14010);
nor U14769 (N_14769,N_14057,N_14099);
nand U14770 (N_14770,N_13874,N_14175);
and U14771 (N_14771,N_13776,N_13691);
nor U14772 (N_14772,N_13929,N_14092);
and U14773 (N_14773,N_14087,N_13719);
nor U14774 (N_14774,N_13650,N_13669);
nor U14775 (N_14775,N_13955,N_13714);
xor U14776 (N_14776,N_13890,N_13753);
or U14777 (N_14777,N_13632,N_13828);
xnor U14778 (N_14778,N_14312,N_14146);
nand U14779 (N_14779,N_13648,N_14094);
or U14780 (N_14780,N_14376,N_14198);
xor U14781 (N_14781,N_13847,N_13940);
and U14782 (N_14782,N_14309,N_13836);
xnor U14783 (N_14783,N_13663,N_13713);
or U14784 (N_14784,N_14207,N_14243);
nor U14785 (N_14785,N_13640,N_14251);
and U14786 (N_14786,N_13960,N_13744);
nand U14787 (N_14787,N_14397,N_14306);
nand U14788 (N_14788,N_13864,N_14061);
nand U14789 (N_14789,N_13861,N_14107);
xor U14790 (N_14790,N_14287,N_13707);
xnor U14791 (N_14791,N_13647,N_14119);
nand U14792 (N_14792,N_14165,N_14136);
or U14793 (N_14793,N_13680,N_13987);
xnor U14794 (N_14794,N_13725,N_13711);
or U14795 (N_14795,N_13706,N_14217);
and U14796 (N_14796,N_14373,N_14093);
nor U14797 (N_14797,N_14215,N_13631);
or U14798 (N_14798,N_13769,N_13925);
nor U14799 (N_14799,N_13845,N_13798);
and U14800 (N_14800,N_14374,N_14135);
xnor U14801 (N_14801,N_14345,N_13613);
nor U14802 (N_14802,N_13887,N_13655);
and U14803 (N_14803,N_13823,N_14317);
and U14804 (N_14804,N_14263,N_14366);
or U14805 (N_14805,N_14058,N_13919);
nor U14806 (N_14806,N_14247,N_13959);
xor U14807 (N_14807,N_13909,N_14088);
xor U14808 (N_14808,N_14228,N_13712);
xor U14809 (N_14809,N_13966,N_13839);
xor U14810 (N_14810,N_14065,N_13726);
xnor U14811 (N_14811,N_13755,N_13628);
xor U14812 (N_14812,N_13834,N_14049);
or U14813 (N_14813,N_14200,N_14221);
and U14814 (N_14814,N_14124,N_14269);
nand U14815 (N_14815,N_14234,N_14311);
xor U14816 (N_14816,N_13654,N_13975);
nor U14817 (N_14817,N_13666,N_14077);
or U14818 (N_14818,N_13673,N_14101);
and U14819 (N_14819,N_14062,N_14013);
nor U14820 (N_14820,N_14314,N_13872);
nand U14821 (N_14821,N_14205,N_14155);
nand U14822 (N_14822,N_13997,N_13770);
nand U14823 (N_14823,N_14341,N_13835);
or U14824 (N_14824,N_13708,N_14198);
or U14825 (N_14825,N_14173,N_14139);
and U14826 (N_14826,N_14025,N_13889);
or U14827 (N_14827,N_13668,N_13785);
or U14828 (N_14828,N_14163,N_13897);
nand U14829 (N_14829,N_13928,N_13849);
or U14830 (N_14830,N_14286,N_13609);
or U14831 (N_14831,N_14053,N_14026);
nor U14832 (N_14832,N_13948,N_14009);
nor U14833 (N_14833,N_13774,N_13824);
nand U14834 (N_14834,N_13773,N_13885);
or U14835 (N_14835,N_14184,N_13684);
nor U14836 (N_14836,N_13664,N_14357);
nand U14837 (N_14837,N_14283,N_14004);
xor U14838 (N_14838,N_13641,N_13870);
or U14839 (N_14839,N_14260,N_13625);
nor U14840 (N_14840,N_14074,N_13879);
and U14841 (N_14841,N_13980,N_13770);
and U14842 (N_14842,N_13760,N_13976);
nand U14843 (N_14843,N_14146,N_14205);
nand U14844 (N_14844,N_14296,N_13903);
nor U14845 (N_14845,N_13661,N_14115);
or U14846 (N_14846,N_14105,N_14219);
xor U14847 (N_14847,N_13685,N_13675);
and U14848 (N_14848,N_14257,N_14124);
nor U14849 (N_14849,N_13965,N_13949);
and U14850 (N_14850,N_13838,N_14280);
or U14851 (N_14851,N_13877,N_14249);
nor U14852 (N_14852,N_14325,N_13954);
nand U14853 (N_14853,N_13943,N_13854);
nor U14854 (N_14854,N_13976,N_13878);
xnor U14855 (N_14855,N_13803,N_14021);
or U14856 (N_14856,N_13924,N_14180);
nand U14857 (N_14857,N_14106,N_13882);
and U14858 (N_14858,N_13957,N_13817);
nor U14859 (N_14859,N_13843,N_13949);
nand U14860 (N_14860,N_13749,N_14047);
xnor U14861 (N_14861,N_13625,N_14212);
or U14862 (N_14862,N_13968,N_14280);
nor U14863 (N_14863,N_13730,N_13813);
nor U14864 (N_14864,N_13698,N_14314);
nor U14865 (N_14865,N_13623,N_13832);
and U14866 (N_14866,N_13831,N_13987);
or U14867 (N_14867,N_14241,N_14285);
and U14868 (N_14868,N_13691,N_13895);
nand U14869 (N_14869,N_13824,N_13901);
and U14870 (N_14870,N_13811,N_14074);
nand U14871 (N_14871,N_13706,N_14299);
and U14872 (N_14872,N_14117,N_14003);
nand U14873 (N_14873,N_13648,N_13921);
and U14874 (N_14874,N_13692,N_14148);
and U14875 (N_14875,N_13804,N_13870);
xor U14876 (N_14876,N_14283,N_13751);
nand U14877 (N_14877,N_13610,N_14119);
or U14878 (N_14878,N_13621,N_14262);
and U14879 (N_14879,N_14203,N_14369);
nand U14880 (N_14880,N_14324,N_14126);
xnor U14881 (N_14881,N_13709,N_14344);
xor U14882 (N_14882,N_13995,N_14220);
xnor U14883 (N_14883,N_13700,N_14250);
nand U14884 (N_14884,N_13672,N_13733);
xnor U14885 (N_14885,N_13891,N_13987);
xnor U14886 (N_14886,N_13956,N_14274);
nand U14887 (N_14887,N_14234,N_14302);
or U14888 (N_14888,N_14395,N_13661);
nand U14889 (N_14889,N_13873,N_13615);
xor U14890 (N_14890,N_14099,N_13727);
or U14891 (N_14891,N_13644,N_14249);
nand U14892 (N_14892,N_13997,N_13896);
and U14893 (N_14893,N_14301,N_13869);
xnor U14894 (N_14894,N_14351,N_14286);
xor U14895 (N_14895,N_13946,N_14007);
or U14896 (N_14896,N_14106,N_14118);
xor U14897 (N_14897,N_13950,N_13757);
nand U14898 (N_14898,N_13736,N_14136);
xnor U14899 (N_14899,N_13995,N_13788);
or U14900 (N_14900,N_14328,N_13846);
nand U14901 (N_14901,N_14269,N_14238);
nand U14902 (N_14902,N_13623,N_14149);
nand U14903 (N_14903,N_13901,N_13957);
or U14904 (N_14904,N_14143,N_14178);
xor U14905 (N_14905,N_13901,N_13635);
xor U14906 (N_14906,N_14234,N_13783);
xnor U14907 (N_14907,N_13809,N_14210);
or U14908 (N_14908,N_13607,N_13908);
xnor U14909 (N_14909,N_13862,N_14378);
and U14910 (N_14910,N_14215,N_13903);
and U14911 (N_14911,N_14323,N_13736);
xnor U14912 (N_14912,N_13741,N_14136);
nand U14913 (N_14913,N_14239,N_13777);
and U14914 (N_14914,N_14133,N_14186);
nand U14915 (N_14915,N_14061,N_13650);
nand U14916 (N_14916,N_13777,N_13709);
xor U14917 (N_14917,N_14070,N_13772);
nand U14918 (N_14918,N_14254,N_14164);
xnor U14919 (N_14919,N_13910,N_14324);
xnor U14920 (N_14920,N_13861,N_13993);
nand U14921 (N_14921,N_14398,N_13627);
nor U14922 (N_14922,N_14312,N_13994);
xor U14923 (N_14923,N_13711,N_14257);
or U14924 (N_14924,N_14062,N_14101);
nand U14925 (N_14925,N_13668,N_14055);
nor U14926 (N_14926,N_14321,N_13833);
and U14927 (N_14927,N_14004,N_13729);
xor U14928 (N_14928,N_13823,N_14028);
and U14929 (N_14929,N_14153,N_14141);
nand U14930 (N_14930,N_13630,N_13884);
and U14931 (N_14931,N_13895,N_14190);
nand U14932 (N_14932,N_13697,N_14171);
xnor U14933 (N_14933,N_14045,N_14358);
or U14934 (N_14934,N_14106,N_13759);
nor U14935 (N_14935,N_13609,N_13631);
and U14936 (N_14936,N_13612,N_14080);
nand U14937 (N_14937,N_13813,N_13827);
nand U14938 (N_14938,N_13799,N_14081);
nor U14939 (N_14939,N_13644,N_13791);
xnor U14940 (N_14940,N_13634,N_13771);
nand U14941 (N_14941,N_14198,N_14158);
nor U14942 (N_14942,N_13818,N_13948);
xor U14943 (N_14943,N_13907,N_13619);
nor U14944 (N_14944,N_13833,N_13610);
nand U14945 (N_14945,N_13904,N_13694);
nor U14946 (N_14946,N_14137,N_14260);
xnor U14947 (N_14947,N_13875,N_13911);
nand U14948 (N_14948,N_13790,N_14273);
or U14949 (N_14949,N_13721,N_14342);
and U14950 (N_14950,N_14360,N_13698);
and U14951 (N_14951,N_13728,N_14242);
and U14952 (N_14952,N_13879,N_13623);
xnor U14953 (N_14953,N_14012,N_14312);
xnor U14954 (N_14954,N_13883,N_14295);
nand U14955 (N_14955,N_14323,N_13993);
or U14956 (N_14956,N_13875,N_14042);
and U14957 (N_14957,N_14030,N_13993);
and U14958 (N_14958,N_13811,N_13996);
and U14959 (N_14959,N_14223,N_14069);
nor U14960 (N_14960,N_14328,N_14006);
xor U14961 (N_14961,N_14246,N_14141);
xnor U14962 (N_14962,N_13699,N_13779);
nor U14963 (N_14963,N_13857,N_14321);
nand U14964 (N_14964,N_14021,N_13720);
or U14965 (N_14965,N_13787,N_14085);
xnor U14966 (N_14966,N_13736,N_14111);
or U14967 (N_14967,N_13790,N_14334);
xor U14968 (N_14968,N_14171,N_14379);
nor U14969 (N_14969,N_13701,N_13742);
nand U14970 (N_14970,N_14131,N_14080);
nor U14971 (N_14971,N_14055,N_13649);
nor U14972 (N_14972,N_14267,N_13675);
xnor U14973 (N_14973,N_13979,N_13858);
nand U14974 (N_14974,N_14284,N_14171);
or U14975 (N_14975,N_14274,N_13952);
nor U14976 (N_14976,N_14359,N_13753);
and U14977 (N_14977,N_14303,N_13679);
or U14978 (N_14978,N_13845,N_14018);
or U14979 (N_14979,N_14299,N_13781);
and U14980 (N_14980,N_13605,N_13781);
or U14981 (N_14981,N_13846,N_13899);
nand U14982 (N_14982,N_13821,N_14318);
and U14983 (N_14983,N_14194,N_14229);
and U14984 (N_14984,N_13640,N_14092);
xnor U14985 (N_14985,N_13828,N_14319);
xnor U14986 (N_14986,N_14330,N_14257);
xnor U14987 (N_14987,N_14386,N_14314);
or U14988 (N_14988,N_13842,N_14188);
nand U14989 (N_14989,N_13941,N_14181);
and U14990 (N_14990,N_13855,N_14145);
xnor U14991 (N_14991,N_14159,N_13830);
nand U14992 (N_14992,N_14394,N_14224);
nor U14993 (N_14993,N_13972,N_13649);
nand U14994 (N_14994,N_13937,N_14049);
or U14995 (N_14995,N_14060,N_14248);
xnor U14996 (N_14996,N_13719,N_14244);
nand U14997 (N_14997,N_14227,N_14262);
and U14998 (N_14998,N_13954,N_13733);
nor U14999 (N_14999,N_14364,N_13920);
nor U15000 (N_15000,N_14192,N_13817);
or U15001 (N_15001,N_13659,N_13655);
nor U15002 (N_15002,N_13694,N_13985);
nand U15003 (N_15003,N_14050,N_14124);
or U15004 (N_15004,N_13780,N_14241);
nand U15005 (N_15005,N_14382,N_13819);
or U15006 (N_15006,N_14332,N_14031);
or U15007 (N_15007,N_14319,N_14317);
nand U15008 (N_15008,N_13724,N_13727);
and U15009 (N_15009,N_13956,N_14050);
nor U15010 (N_15010,N_13934,N_14364);
and U15011 (N_15011,N_13848,N_14232);
nor U15012 (N_15012,N_13847,N_13791);
and U15013 (N_15013,N_13607,N_14245);
nor U15014 (N_15014,N_13744,N_13623);
and U15015 (N_15015,N_14022,N_14337);
nand U15016 (N_15016,N_13808,N_14220);
and U15017 (N_15017,N_14101,N_13777);
nor U15018 (N_15018,N_13795,N_14290);
nand U15019 (N_15019,N_14234,N_14121);
nand U15020 (N_15020,N_14267,N_13965);
and U15021 (N_15021,N_13801,N_13947);
nor U15022 (N_15022,N_13649,N_13753);
and U15023 (N_15023,N_14049,N_13763);
or U15024 (N_15024,N_13759,N_14360);
nand U15025 (N_15025,N_13852,N_13656);
nor U15026 (N_15026,N_13846,N_14008);
or U15027 (N_15027,N_14280,N_13880);
nor U15028 (N_15028,N_13993,N_13945);
xor U15029 (N_15029,N_13693,N_14323);
xor U15030 (N_15030,N_14344,N_13846);
and U15031 (N_15031,N_14336,N_13849);
nor U15032 (N_15032,N_13756,N_14343);
and U15033 (N_15033,N_13853,N_14078);
and U15034 (N_15034,N_14071,N_13887);
and U15035 (N_15035,N_14243,N_13900);
and U15036 (N_15036,N_14157,N_14256);
xnor U15037 (N_15037,N_14230,N_13652);
xnor U15038 (N_15038,N_14296,N_14381);
and U15039 (N_15039,N_14295,N_14157);
nor U15040 (N_15040,N_13812,N_14073);
and U15041 (N_15041,N_13807,N_14249);
or U15042 (N_15042,N_13865,N_14122);
xor U15043 (N_15043,N_14076,N_13752);
xnor U15044 (N_15044,N_13628,N_13962);
nor U15045 (N_15045,N_14373,N_13894);
nor U15046 (N_15046,N_14289,N_14151);
xor U15047 (N_15047,N_13814,N_13691);
nand U15048 (N_15048,N_13749,N_14256);
or U15049 (N_15049,N_14255,N_14282);
xor U15050 (N_15050,N_14100,N_13835);
and U15051 (N_15051,N_13941,N_14155);
xnor U15052 (N_15052,N_14017,N_14132);
nor U15053 (N_15053,N_14356,N_14013);
nor U15054 (N_15054,N_14147,N_14062);
or U15055 (N_15055,N_14399,N_13858);
nor U15056 (N_15056,N_14248,N_14242);
and U15057 (N_15057,N_14152,N_14082);
nand U15058 (N_15058,N_14396,N_13993);
or U15059 (N_15059,N_13923,N_13816);
nand U15060 (N_15060,N_14310,N_13742);
and U15061 (N_15061,N_14319,N_14232);
or U15062 (N_15062,N_14129,N_14311);
or U15063 (N_15063,N_13981,N_13632);
xor U15064 (N_15064,N_14195,N_13760);
and U15065 (N_15065,N_14149,N_14060);
xnor U15066 (N_15066,N_14053,N_14300);
and U15067 (N_15067,N_14311,N_14008);
xor U15068 (N_15068,N_13931,N_14224);
nor U15069 (N_15069,N_13954,N_14209);
or U15070 (N_15070,N_14033,N_13952);
xor U15071 (N_15071,N_13897,N_14399);
xor U15072 (N_15072,N_14043,N_13764);
xnor U15073 (N_15073,N_13866,N_13703);
nor U15074 (N_15074,N_13608,N_14200);
xnor U15075 (N_15075,N_14319,N_14310);
nor U15076 (N_15076,N_14053,N_14155);
nand U15077 (N_15077,N_13817,N_13953);
and U15078 (N_15078,N_14374,N_13884);
xor U15079 (N_15079,N_13635,N_13684);
xor U15080 (N_15080,N_13919,N_14344);
nor U15081 (N_15081,N_13887,N_14052);
nand U15082 (N_15082,N_14229,N_13644);
nand U15083 (N_15083,N_13821,N_13626);
and U15084 (N_15084,N_14306,N_14344);
nand U15085 (N_15085,N_14251,N_14292);
xnor U15086 (N_15086,N_13972,N_13748);
nor U15087 (N_15087,N_14031,N_13641);
and U15088 (N_15088,N_14271,N_13933);
or U15089 (N_15089,N_13950,N_13789);
and U15090 (N_15090,N_13652,N_13675);
nor U15091 (N_15091,N_14302,N_14165);
nand U15092 (N_15092,N_14039,N_13721);
or U15093 (N_15093,N_14171,N_13965);
or U15094 (N_15094,N_14327,N_14188);
and U15095 (N_15095,N_13847,N_14196);
nand U15096 (N_15096,N_13774,N_14194);
xnor U15097 (N_15097,N_14367,N_13681);
xor U15098 (N_15098,N_14334,N_14077);
xnor U15099 (N_15099,N_13663,N_14201);
or U15100 (N_15100,N_14103,N_14366);
nand U15101 (N_15101,N_14343,N_13767);
xor U15102 (N_15102,N_13894,N_13792);
or U15103 (N_15103,N_14092,N_14151);
and U15104 (N_15104,N_14009,N_14262);
xor U15105 (N_15105,N_14042,N_13746);
nor U15106 (N_15106,N_14396,N_13615);
nor U15107 (N_15107,N_14343,N_13670);
nor U15108 (N_15108,N_13865,N_14272);
or U15109 (N_15109,N_13660,N_13766);
nor U15110 (N_15110,N_14060,N_13669);
nand U15111 (N_15111,N_13880,N_13678);
nor U15112 (N_15112,N_14139,N_14174);
or U15113 (N_15113,N_13799,N_13661);
nor U15114 (N_15114,N_14170,N_13921);
nor U15115 (N_15115,N_13714,N_13754);
and U15116 (N_15116,N_13789,N_13829);
xor U15117 (N_15117,N_13850,N_13764);
nand U15118 (N_15118,N_14159,N_14196);
nand U15119 (N_15119,N_13803,N_13746);
nand U15120 (N_15120,N_13690,N_13854);
and U15121 (N_15121,N_14130,N_14179);
or U15122 (N_15122,N_13900,N_14133);
and U15123 (N_15123,N_13843,N_13623);
xnor U15124 (N_15124,N_14274,N_13624);
nor U15125 (N_15125,N_13716,N_13647);
nand U15126 (N_15126,N_13997,N_13662);
or U15127 (N_15127,N_13774,N_13741);
xor U15128 (N_15128,N_13839,N_14009);
xnor U15129 (N_15129,N_14123,N_13746);
or U15130 (N_15130,N_14049,N_14234);
nand U15131 (N_15131,N_14012,N_13826);
or U15132 (N_15132,N_13977,N_14076);
or U15133 (N_15133,N_13960,N_14356);
nand U15134 (N_15134,N_14135,N_13608);
and U15135 (N_15135,N_14267,N_13831);
nor U15136 (N_15136,N_14347,N_14168);
nand U15137 (N_15137,N_14105,N_14240);
and U15138 (N_15138,N_13983,N_13852);
nand U15139 (N_15139,N_14359,N_14161);
xnor U15140 (N_15140,N_14325,N_14333);
xnor U15141 (N_15141,N_14232,N_14089);
or U15142 (N_15142,N_14344,N_14288);
nand U15143 (N_15143,N_14169,N_14206);
nor U15144 (N_15144,N_13736,N_13641);
or U15145 (N_15145,N_14241,N_14082);
xor U15146 (N_15146,N_13642,N_13665);
nor U15147 (N_15147,N_14257,N_14037);
or U15148 (N_15148,N_14030,N_14229);
and U15149 (N_15149,N_13916,N_13623);
nand U15150 (N_15150,N_14022,N_14330);
nand U15151 (N_15151,N_13780,N_13749);
nand U15152 (N_15152,N_13787,N_13695);
and U15153 (N_15153,N_13787,N_13711);
xnor U15154 (N_15154,N_14324,N_13813);
or U15155 (N_15155,N_13741,N_14019);
and U15156 (N_15156,N_13772,N_14360);
or U15157 (N_15157,N_14193,N_14048);
and U15158 (N_15158,N_14295,N_14239);
nor U15159 (N_15159,N_13796,N_14284);
nor U15160 (N_15160,N_14307,N_13819);
or U15161 (N_15161,N_13902,N_13816);
xnor U15162 (N_15162,N_14197,N_14151);
or U15163 (N_15163,N_13712,N_14331);
or U15164 (N_15164,N_13678,N_13974);
xnor U15165 (N_15165,N_13684,N_14192);
and U15166 (N_15166,N_13855,N_13601);
xnor U15167 (N_15167,N_13977,N_13851);
or U15168 (N_15168,N_14235,N_14350);
or U15169 (N_15169,N_13786,N_13783);
and U15170 (N_15170,N_13675,N_14341);
and U15171 (N_15171,N_13967,N_14296);
nor U15172 (N_15172,N_13621,N_13729);
nand U15173 (N_15173,N_13973,N_14219);
nor U15174 (N_15174,N_14274,N_14270);
and U15175 (N_15175,N_13891,N_14138);
nand U15176 (N_15176,N_14079,N_13665);
nor U15177 (N_15177,N_14399,N_13734);
nor U15178 (N_15178,N_13823,N_14319);
nor U15179 (N_15179,N_14107,N_13898);
nor U15180 (N_15180,N_13719,N_13873);
and U15181 (N_15181,N_13823,N_13642);
nand U15182 (N_15182,N_14274,N_13626);
nand U15183 (N_15183,N_14360,N_13996);
xnor U15184 (N_15184,N_13921,N_14054);
or U15185 (N_15185,N_13639,N_13649);
and U15186 (N_15186,N_14041,N_13811);
nor U15187 (N_15187,N_14056,N_13834);
xor U15188 (N_15188,N_13871,N_14377);
or U15189 (N_15189,N_14139,N_13761);
and U15190 (N_15190,N_14212,N_13772);
or U15191 (N_15191,N_14134,N_13888);
or U15192 (N_15192,N_13968,N_13803);
nand U15193 (N_15193,N_14325,N_13949);
xnor U15194 (N_15194,N_13848,N_14361);
nor U15195 (N_15195,N_14390,N_14312);
nor U15196 (N_15196,N_13959,N_13943);
and U15197 (N_15197,N_13790,N_13960);
nand U15198 (N_15198,N_13978,N_14095);
nand U15199 (N_15199,N_13984,N_14380);
and U15200 (N_15200,N_14876,N_14546);
nand U15201 (N_15201,N_15193,N_14492);
nand U15202 (N_15202,N_14771,N_15125);
xor U15203 (N_15203,N_14895,N_14669);
or U15204 (N_15204,N_14896,N_14735);
nor U15205 (N_15205,N_14841,N_14857);
nor U15206 (N_15206,N_14804,N_14974);
or U15207 (N_15207,N_14463,N_14464);
nand U15208 (N_15208,N_15181,N_14419);
and U15209 (N_15209,N_14973,N_15053);
or U15210 (N_15210,N_14545,N_14537);
nor U15211 (N_15211,N_15142,N_14527);
or U15212 (N_15212,N_14731,N_14903);
nor U15213 (N_15213,N_14885,N_14937);
xor U15214 (N_15214,N_14644,N_15051);
nor U15215 (N_15215,N_14913,N_14674);
or U15216 (N_15216,N_14760,N_15127);
or U15217 (N_15217,N_14708,N_15056);
nand U15218 (N_15218,N_14429,N_14749);
xnor U15219 (N_15219,N_14665,N_15138);
or U15220 (N_15220,N_14684,N_14963);
nand U15221 (N_15221,N_15197,N_14814);
nor U15222 (N_15222,N_14409,N_14411);
xnor U15223 (N_15223,N_15171,N_15044);
nor U15224 (N_15224,N_15072,N_14586);
nand U15225 (N_15225,N_14611,N_14483);
nor U15226 (N_15226,N_15050,N_15066);
xnor U15227 (N_15227,N_14740,N_14467);
xor U15228 (N_15228,N_14680,N_14757);
nand U15229 (N_15229,N_14931,N_15030);
xor U15230 (N_15230,N_15040,N_15163);
nand U15231 (N_15231,N_14968,N_15135);
or U15232 (N_15232,N_14512,N_14590);
and U15233 (N_15233,N_14621,N_14962);
nor U15234 (N_15234,N_14477,N_14957);
or U15235 (N_15235,N_14486,N_14981);
and U15236 (N_15236,N_14830,N_14979);
nor U15237 (N_15237,N_14671,N_14714);
and U15238 (N_15238,N_15005,N_14426);
nand U15239 (N_15239,N_15130,N_14566);
xor U15240 (N_15240,N_14883,N_14417);
nor U15241 (N_15241,N_14781,N_14449);
or U15242 (N_15242,N_15185,N_15158);
or U15243 (N_15243,N_14815,N_15132);
nand U15244 (N_15244,N_14940,N_15155);
nor U15245 (N_15245,N_15166,N_14461);
and U15246 (N_15246,N_14657,N_14718);
xnor U15247 (N_15247,N_14633,N_15182);
and U15248 (N_15248,N_14784,N_15134);
and U15249 (N_15249,N_14698,N_14787);
nand U15250 (N_15250,N_14648,N_14642);
nor U15251 (N_15251,N_15150,N_14686);
xnor U15252 (N_15252,N_14530,N_14614);
xor U15253 (N_15253,N_14475,N_15057);
nor U15254 (N_15254,N_14634,N_14859);
or U15255 (N_15255,N_14433,N_14776);
and U15256 (N_15256,N_14507,N_14427);
nor U15257 (N_15257,N_14676,N_15177);
nand U15258 (N_15258,N_14798,N_14988);
or U15259 (N_15259,N_15059,N_14478);
nor U15260 (N_15260,N_14679,N_15112);
nor U15261 (N_15261,N_15064,N_14910);
or U15262 (N_15262,N_14843,N_14966);
and U15263 (N_15263,N_15190,N_14908);
xor U15264 (N_15264,N_14923,N_15165);
nand U15265 (N_15265,N_14738,N_15115);
nand U15266 (N_15266,N_15060,N_14911);
and U15267 (N_15267,N_14816,N_14450);
or U15268 (N_15268,N_15162,N_15176);
xnor U15269 (N_15269,N_14422,N_14877);
or U15270 (N_15270,N_14799,N_15010);
xnor U15271 (N_15271,N_15023,N_14820);
nor U15272 (N_15272,N_15152,N_14889);
nand U15273 (N_15273,N_14746,N_15184);
xor U15274 (N_15274,N_14651,N_15080);
and U15275 (N_15275,N_14768,N_14649);
nand U15276 (N_15276,N_14709,N_14852);
nand U15277 (N_15277,N_14416,N_14995);
nor U15278 (N_15278,N_14608,N_14906);
nand U15279 (N_15279,N_14719,N_14456);
xnor U15280 (N_15280,N_14855,N_14965);
xor U15281 (N_15281,N_14888,N_14812);
nand U15282 (N_15282,N_14471,N_15042);
and U15283 (N_15283,N_15091,N_15031);
nor U15284 (N_15284,N_14505,N_14846);
or U15285 (N_15285,N_14543,N_15061);
or U15286 (N_15286,N_14402,N_14870);
and U15287 (N_15287,N_14504,N_14469);
xor U15288 (N_15288,N_14403,N_15062);
and U15289 (N_15289,N_14568,N_14440);
or U15290 (N_15290,N_14630,N_15033);
or U15291 (N_15291,N_14763,N_14598);
nand U15292 (N_15292,N_14861,N_14909);
xnor U15293 (N_15293,N_14547,N_14574);
nand U15294 (N_15294,N_14990,N_15029);
and U15295 (N_15295,N_14829,N_14999);
nand U15296 (N_15296,N_14622,N_14775);
nand U15297 (N_15297,N_14553,N_14444);
or U15298 (N_15298,N_14823,N_14796);
and U15299 (N_15299,N_14595,N_14828);
nand U15300 (N_15300,N_15109,N_15194);
xnor U15301 (N_15301,N_14953,N_14726);
nor U15302 (N_15302,N_14985,N_14993);
nand U15303 (N_15303,N_14460,N_14518);
xnor U15304 (N_15304,N_14654,N_15095);
and U15305 (N_15305,N_14720,N_15119);
and U15306 (N_15306,N_14701,N_14510);
or U15307 (N_15307,N_14922,N_14933);
nor U15308 (N_15308,N_15178,N_15167);
nand U15309 (N_15309,N_14792,N_14643);
and U15310 (N_15310,N_15035,N_14839);
xor U15311 (N_15311,N_14976,N_14620);
nand U15312 (N_15312,N_14805,N_14470);
xnor U15313 (N_15313,N_14756,N_15020);
xnor U15314 (N_15314,N_14869,N_15174);
or U15315 (N_15315,N_14951,N_14662);
xnor U15316 (N_15316,N_14754,N_14418);
and U15317 (N_15317,N_14540,N_14489);
nor U15318 (N_15318,N_14500,N_14693);
nand U15319 (N_15319,N_14646,N_15136);
nand U15320 (N_15320,N_15022,N_15169);
xor U15321 (N_15321,N_15039,N_14847);
xnor U15322 (N_15322,N_14958,N_14918);
nor U15323 (N_15323,N_14541,N_15086);
nor U15324 (N_15324,N_14700,N_14902);
nor U15325 (N_15325,N_14935,N_14459);
xor U15326 (N_15326,N_15137,N_15065);
or U15327 (N_15327,N_15045,N_14807);
nor U15328 (N_15328,N_15116,N_14840);
and U15329 (N_15329,N_14915,N_14410);
nand U15330 (N_15330,N_14890,N_14659);
or U15331 (N_15331,N_14837,N_14509);
and U15332 (N_15332,N_14549,N_14789);
nand U15333 (N_15333,N_14639,N_15107);
nor U15334 (N_15334,N_15101,N_14685);
nor U15335 (N_15335,N_14521,N_14865);
nand U15336 (N_15336,N_14623,N_15015);
xnor U15337 (N_15337,N_14508,N_14765);
and U15338 (N_15338,N_14743,N_14971);
xor U15339 (N_15339,N_15183,N_14635);
or U15340 (N_15340,N_14875,N_14564);
nor U15341 (N_15341,N_14597,N_14955);
xor U15342 (N_15342,N_14476,N_15102);
or U15343 (N_15343,N_15021,N_14548);
and U15344 (N_15344,N_15146,N_15006);
nand U15345 (N_15345,N_14739,N_14596);
nor U15346 (N_15346,N_14887,N_14975);
nand U15347 (N_15347,N_14443,N_14690);
nand U15348 (N_15348,N_14683,N_14939);
or U15349 (N_15349,N_14472,N_14882);
and U15350 (N_15350,N_15168,N_14400);
and U15351 (N_15351,N_14434,N_14678);
or U15352 (N_15352,N_15041,N_15007);
xnor U15353 (N_15353,N_14921,N_14579);
and U15354 (N_15354,N_14699,N_14414);
nor U15355 (N_15355,N_14984,N_14557);
or U15356 (N_15356,N_14406,N_14788);
and U15357 (N_15357,N_15099,N_14482);
nor U15358 (N_15358,N_14653,N_15110);
and U15359 (N_15359,N_14462,N_14632);
and U15360 (N_15360,N_14514,N_14961);
xor U15361 (N_15361,N_14986,N_15096);
nand U15362 (N_15362,N_14747,N_14725);
or U15363 (N_15363,N_14762,N_14930);
nor U15364 (N_15364,N_15188,N_14589);
and U15365 (N_15365,N_14948,N_15004);
nand U15366 (N_15366,N_14817,N_14905);
nor U15367 (N_15367,N_15052,N_14917);
nor U15368 (N_15368,N_15187,N_14465);
and U15369 (N_15369,N_14897,N_15055);
or U15370 (N_15370,N_14610,N_14919);
nand U15371 (N_15371,N_14980,N_14558);
and U15372 (N_15372,N_14484,N_14928);
nor U15373 (N_15373,N_14891,N_14866);
xnor U15374 (N_15374,N_14503,N_14535);
xnor U15375 (N_15375,N_14519,N_15104);
or U15376 (N_15376,N_14892,N_14501);
and U15377 (N_15377,N_14803,N_14451);
nor U15378 (N_15378,N_14592,N_14435);
xor U15379 (N_15379,N_14473,N_14533);
and U15380 (N_15380,N_14593,N_15047);
nor U15381 (N_15381,N_15172,N_14899);
nor U15382 (N_15382,N_14944,N_14569);
nand U15383 (N_15383,N_14878,N_14567);
nand U15384 (N_15384,N_14448,N_14607);
nor U15385 (N_15385,N_14702,N_14531);
and U15386 (N_15386,N_14577,N_15121);
nand U15387 (N_15387,N_14515,N_15084);
nand U15388 (N_15388,N_14544,N_14555);
and U15389 (N_15389,N_14538,N_14575);
and U15390 (N_15390,N_15100,N_14947);
and U15391 (N_15391,N_15122,N_15153);
or U15392 (N_15392,N_14942,N_15071);
nor U15393 (N_15393,N_14991,N_15049);
or U15394 (N_15394,N_15067,N_14802);
and U15395 (N_15395,N_14711,N_14526);
and U15396 (N_15396,N_14904,N_15199);
nand U15397 (N_15397,N_14570,N_14723);
xnor U15398 (N_15398,N_14864,N_14687);
nor U15399 (N_15399,N_14499,N_15151);
or U15400 (N_15400,N_14824,N_14627);
nor U15401 (N_15401,N_14927,N_15074);
xnor U15402 (N_15402,N_14806,N_15028);
and U15403 (N_15403,N_14525,N_15159);
and U15404 (N_15404,N_15088,N_14912);
nor U15405 (N_15405,N_14561,N_14728);
or U15406 (N_15406,N_14916,N_14932);
xor U15407 (N_15407,N_14582,N_14954);
xnor U15408 (N_15408,N_15038,N_14987);
nand U15409 (N_15409,N_14862,N_14934);
xnor U15410 (N_15410,N_14748,N_14445);
nand U15411 (N_15411,N_14481,N_14437);
xor U15412 (N_15412,N_14767,N_14801);
and U15413 (N_15413,N_14562,N_14438);
and U15414 (N_15414,N_14777,N_14613);
and U15415 (N_15415,N_14647,N_14485);
xnor U15416 (N_15416,N_14645,N_15008);
xnor U15417 (N_15417,N_14791,N_14832);
and U15418 (N_15418,N_14655,N_14523);
xor U15419 (N_15419,N_14867,N_14752);
xnor U15420 (N_15420,N_14428,N_14751);
or U15421 (N_15421,N_14759,N_14972);
or U15422 (N_15422,N_14554,N_14423);
nand U15423 (N_15423,N_15195,N_14640);
or U15424 (N_15424,N_14420,N_14556);
or U15425 (N_15425,N_14572,N_14736);
xnor U15426 (N_15426,N_14833,N_15189);
and U15427 (N_15427,N_15036,N_15173);
and U15428 (N_15428,N_14664,N_15012);
nand U15429 (N_15429,N_14636,N_14628);
and U15430 (N_15430,N_14407,N_15083);
or U15431 (N_15431,N_14844,N_14631);
and U15432 (N_15432,N_14415,N_14845);
xnor U15433 (N_15433,N_14641,N_15105);
xor U15434 (N_15434,N_14431,N_14658);
nand U15435 (N_15435,N_14490,N_14997);
xor U15436 (N_15436,N_15154,N_14929);
nand U15437 (N_15437,N_15017,N_15106);
or U15438 (N_15438,N_14964,N_14831);
nand U15439 (N_15439,N_15032,N_14532);
or U15440 (N_15440,N_14668,N_15140);
and U15441 (N_15441,N_15120,N_15126);
and U15442 (N_15442,N_14487,N_14848);
nand U15443 (N_15443,N_14809,N_14496);
xnor U15444 (N_15444,N_14790,N_14688);
and U15445 (N_15445,N_15037,N_14430);
xnor U15446 (N_15446,N_15186,N_14745);
or U15447 (N_15447,N_14498,N_14717);
xor U15448 (N_15448,N_15076,N_14774);
or U15449 (N_15449,N_15070,N_14949);
xnor U15450 (N_15450,N_14455,N_14779);
xor U15451 (N_15451,N_14907,N_14945);
nand U15452 (N_15452,N_14516,N_14727);
or U15453 (N_15453,N_14838,N_14825);
or U15454 (N_15454,N_15073,N_14425);
nand U15455 (N_15455,N_15075,N_14758);
xor U15456 (N_15456,N_15089,N_14778);
xnor U15457 (N_15457,N_14872,N_14681);
and U15458 (N_15458,N_15085,N_14401);
and U15459 (N_15459,N_14886,N_14615);
xor U15460 (N_15460,N_15175,N_14675);
xor U15461 (N_15461,N_14663,N_14969);
xor U15462 (N_15462,N_15016,N_14936);
and U15463 (N_15463,N_14692,N_14881);
and U15464 (N_15464,N_14697,N_14661);
and U15465 (N_15465,N_14488,N_14446);
or U15466 (N_15466,N_15124,N_14926);
xnor U15467 (N_15467,N_14694,N_14734);
nor U15468 (N_15468,N_14856,N_15113);
and U15469 (N_15469,N_14994,N_14696);
or U15470 (N_15470,N_15090,N_14529);
xnor U15471 (N_15471,N_14819,N_14713);
nor U15472 (N_15472,N_14453,N_14721);
and U15473 (N_15473,N_14591,N_14853);
nand U15474 (N_15474,N_14468,N_14712);
xnor U15475 (N_15475,N_14497,N_14925);
or U15476 (N_15476,N_14710,N_15148);
and U15477 (N_15477,N_14539,N_14629);
nand U15478 (N_15478,N_14528,N_14880);
and U15479 (N_15479,N_14894,N_14638);
nor U15480 (N_15480,N_14821,N_14625);
and U15481 (N_15481,N_14836,N_14893);
and U15482 (N_15482,N_15048,N_14952);
and U15483 (N_15483,N_14827,N_14573);
and U15484 (N_15484,N_14689,N_15043);
and U15485 (N_15485,N_14413,N_15003);
or U15486 (N_15486,N_14744,N_14956);
xnor U15487 (N_15487,N_14742,N_15196);
nor U15488 (N_15488,N_14599,N_14506);
nand U15489 (N_15489,N_14605,N_15068);
or U15490 (N_15490,N_14769,N_15114);
and U15491 (N_15491,N_15081,N_14732);
and U15492 (N_15492,N_14466,N_15018);
xor U15493 (N_15493,N_14666,N_14571);
or U15494 (N_15494,N_14452,N_15082);
or U15495 (N_15495,N_14616,N_14800);
nand U15496 (N_15496,N_15160,N_15094);
xnor U15497 (N_15497,N_14457,N_14860);
nand U15498 (N_15498,N_14436,N_14811);
or U15499 (N_15499,N_14578,N_14624);
nor U15500 (N_15500,N_14612,N_14729);
and U15501 (N_15501,N_14588,N_14458);
nand U15502 (N_15502,N_15079,N_15144);
and U15503 (N_15503,N_14849,N_14603);
xnor U15504 (N_15504,N_14782,N_14606);
nor U15505 (N_15505,N_14565,N_14677);
and U15506 (N_15506,N_15103,N_14924);
xor U15507 (N_15507,N_14874,N_14550);
nand U15508 (N_15508,N_15149,N_14996);
and U15509 (N_15509,N_15046,N_14741);
nor U15510 (N_15510,N_14863,N_14797);
nand U15511 (N_15511,N_14691,N_14619);
nand U15512 (N_15512,N_14673,N_14795);
and U15513 (N_15513,N_14650,N_14773);
nor U15514 (N_15514,N_14705,N_15054);
nand U15515 (N_15515,N_15097,N_14730);
and U15516 (N_15516,N_14842,N_15164);
nand U15517 (N_15517,N_15157,N_15161);
nand U15518 (N_15518,N_14835,N_14826);
xnor U15519 (N_15519,N_14536,N_15191);
or U15520 (N_15520,N_14682,N_15024);
or U15521 (N_15521,N_14959,N_14810);
or U15522 (N_15522,N_14667,N_14524);
nor U15523 (N_15523,N_15077,N_14601);
or U15524 (N_15524,N_14879,N_15139);
nor U15525 (N_15525,N_14502,N_14441);
and U15526 (N_15526,N_14670,N_14609);
nand U15527 (N_15527,N_14594,N_14583);
and U15528 (N_15528,N_14761,N_14943);
and U15529 (N_15529,N_15002,N_14672);
and U15530 (N_15530,N_14474,N_15128);
xor U15531 (N_15531,N_14766,N_14432);
nor U15532 (N_15532,N_14785,N_14580);
nor U15533 (N_15533,N_14424,N_15063);
nor U15534 (N_15534,N_14600,N_14920);
and U15535 (N_15535,N_15009,N_15179);
and U15536 (N_15536,N_14950,N_14439);
or U15537 (N_15537,N_15123,N_15143);
and U15538 (N_15538,N_14491,N_14818);
xor U15539 (N_15539,N_14584,N_15131);
xnor U15540 (N_15540,N_15034,N_15118);
nand U15541 (N_15541,N_14753,N_14660);
or U15542 (N_15542,N_14783,N_14914);
or U15543 (N_15543,N_14520,N_14868);
xor U15544 (N_15544,N_15000,N_14652);
xnor U15545 (N_15545,N_14970,N_14552);
or U15546 (N_15546,N_15019,N_14494);
and U15547 (N_15547,N_14941,N_14992);
xor U15548 (N_15548,N_14794,N_14834);
nor U15549 (N_15549,N_14576,N_14786);
and U15550 (N_15550,N_14618,N_14704);
and U15551 (N_15551,N_14513,N_14808);
and U15552 (N_15552,N_14998,N_14617);
nand U15553 (N_15553,N_14493,N_15133);
nand U15554 (N_15554,N_14637,N_14442);
or U15555 (N_15555,N_15011,N_14982);
nor U15556 (N_15556,N_15078,N_14511);
nor U15557 (N_15557,N_14850,N_15192);
xnor U15558 (N_15558,N_14989,N_14695);
and U15559 (N_15559,N_15027,N_14793);
xnor U15560 (N_15560,N_14522,N_14750);
nor U15561 (N_15561,N_15092,N_14733);
xnor U15562 (N_15562,N_14404,N_14534);
and U15563 (N_15563,N_14703,N_14560);
nand U15564 (N_15564,N_15147,N_15108);
and U15565 (N_15565,N_15001,N_14454);
or U15566 (N_15566,N_14764,N_14602);
xor U15567 (N_15567,N_14900,N_14551);
nor U15568 (N_15568,N_15087,N_15058);
nor U15569 (N_15569,N_15093,N_14977);
xor U15570 (N_15570,N_14898,N_14873);
xor U15571 (N_15571,N_14851,N_14854);
nand U15572 (N_15572,N_15141,N_14722);
nand U15573 (N_15573,N_14770,N_15014);
and U15574 (N_15574,N_14813,N_14858);
xor U15575 (N_15575,N_14960,N_14585);
and U15576 (N_15576,N_14967,N_14715);
xnor U15577 (N_15577,N_15117,N_14405);
nand U15578 (N_15578,N_14408,N_14581);
nand U15579 (N_15579,N_14755,N_15111);
or U15580 (N_15580,N_15098,N_14724);
nand U15581 (N_15581,N_14871,N_14447);
xor U15582 (N_15582,N_14707,N_14517);
and U15583 (N_15583,N_14587,N_14938);
xor U15584 (N_15584,N_14479,N_15198);
xor U15585 (N_15585,N_14884,N_14901);
or U15586 (N_15586,N_14780,N_14421);
or U15587 (N_15587,N_15026,N_14983);
nand U15588 (N_15588,N_15156,N_14495);
and U15589 (N_15589,N_15013,N_14656);
nor U15590 (N_15590,N_14772,N_14604);
nor U15591 (N_15591,N_14412,N_15170);
nand U15592 (N_15592,N_15025,N_14737);
xnor U15593 (N_15593,N_14978,N_14946);
nand U15594 (N_15594,N_14626,N_15145);
or U15595 (N_15595,N_14542,N_14706);
xnor U15596 (N_15596,N_14716,N_15069);
nor U15597 (N_15597,N_15180,N_14822);
nor U15598 (N_15598,N_14480,N_14559);
nand U15599 (N_15599,N_14563,N_15129);
xnor U15600 (N_15600,N_14537,N_15191);
xnor U15601 (N_15601,N_14980,N_14744);
xor U15602 (N_15602,N_14810,N_14575);
and U15603 (N_15603,N_14953,N_14989);
or U15604 (N_15604,N_15107,N_14738);
nand U15605 (N_15605,N_14483,N_14558);
nor U15606 (N_15606,N_14690,N_14952);
nand U15607 (N_15607,N_14438,N_15197);
nand U15608 (N_15608,N_14655,N_14499);
nand U15609 (N_15609,N_15060,N_14842);
nand U15610 (N_15610,N_15048,N_14611);
nand U15611 (N_15611,N_14811,N_15131);
xor U15612 (N_15612,N_14629,N_14784);
nor U15613 (N_15613,N_14824,N_14981);
and U15614 (N_15614,N_14666,N_14649);
nand U15615 (N_15615,N_14789,N_14527);
and U15616 (N_15616,N_15168,N_14818);
nand U15617 (N_15617,N_15087,N_14509);
nor U15618 (N_15618,N_15197,N_14542);
or U15619 (N_15619,N_14939,N_14988);
and U15620 (N_15620,N_14463,N_14600);
xor U15621 (N_15621,N_15030,N_14623);
nor U15622 (N_15622,N_15027,N_14613);
nand U15623 (N_15623,N_14917,N_14626);
or U15624 (N_15624,N_14779,N_14607);
nand U15625 (N_15625,N_14841,N_14715);
nor U15626 (N_15626,N_14862,N_14722);
nor U15627 (N_15627,N_14951,N_15009);
nand U15628 (N_15628,N_14919,N_14773);
or U15629 (N_15629,N_14712,N_14643);
or U15630 (N_15630,N_14576,N_14875);
and U15631 (N_15631,N_14723,N_14544);
xor U15632 (N_15632,N_14417,N_14493);
and U15633 (N_15633,N_15071,N_14695);
nor U15634 (N_15634,N_15027,N_14904);
nand U15635 (N_15635,N_14418,N_14977);
or U15636 (N_15636,N_15085,N_14560);
nor U15637 (N_15637,N_14899,N_14907);
nor U15638 (N_15638,N_15074,N_14432);
xor U15639 (N_15639,N_14637,N_14952);
nand U15640 (N_15640,N_14730,N_14726);
or U15641 (N_15641,N_14840,N_15102);
nand U15642 (N_15642,N_14626,N_14438);
and U15643 (N_15643,N_14986,N_14795);
or U15644 (N_15644,N_14685,N_15014);
and U15645 (N_15645,N_14429,N_14827);
and U15646 (N_15646,N_15110,N_14866);
xor U15647 (N_15647,N_14891,N_14715);
or U15648 (N_15648,N_15164,N_14925);
xor U15649 (N_15649,N_14668,N_14558);
or U15650 (N_15650,N_14732,N_15051);
and U15651 (N_15651,N_14577,N_14558);
nor U15652 (N_15652,N_14405,N_15197);
and U15653 (N_15653,N_14746,N_14638);
or U15654 (N_15654,N_15112,N_14526);
nand U15655 (N_15655,N_15020,N_14657);
nand U15656 (N_15656,N_14532,N_14640);
and U15657 (N_15657,N_15176,N_14785);
and U15658 (N_15658,N_15088,N_14784);
nor U15659 (N_15659,N_15199,N_14515);
nand U15660 (N_15660,N_14578,N_15010);
nand U15661 (N_15661,N_14746,N_14673);
nor U15662 (N_15662,N_14795,N_14752);
and U15663 (N_15663,N_14720,N_14658);
nand U15664 (N_15664,N_14410,N_14492);
or U15665 (N_15665,N_14933,N_14669);
or U15666 (N_15666,N_14992,N_14806);
xor U15667 (N_15667,N_14616,N_14406);
nand U15668 (N_15668,N_14882,N_14513);
nand U15669 (N_15669,N_14744,N_14528);
nand U15670 (N_15670,N_14610,N_14830);
nor U15671 (N_15671,N_14958,N_14431);
and U15672 (N_15672,N_14685,N_14907);
or U15673 (N_15673,N_14756,N_14648);
and U15674 (N_15674,N_14695,N_14713);
and U15675 (N_15675,N_14451,N_14594);
or U15676 (N_15676,N_14529,N_14675);
nand U15677 (N_15677,N_14670,N_15055);
nand U15678 (N_15678,N_15116,N_14648);
or U15679 (N_15679,N_14790,N_15199);
nand U15680 (N_15680,N_14763,N_14945);
or U15681 (N_15681,N_14916,N_15183);
and U15682 (N_15682,N_14740,N_14403);
nor U15683 (N_15683,N_14957,N_14655);
or U15684 (N_15684,N_14971,N_14468);
nand U15685 (N_15685,N_14796,N_15126);
or U15686 (N_15686,N_15060,N_14535);
xor U15687 (N_15687,N_14852,N_15182);
or U15688 (N_15688,N_14608,N_15097);
nand U15689 (N_15689,N_15176,N_14784);
and U15690 (N_15690,N_14944,N_15138);
or U15691 (N_15691,N_14453,N_14924);
and U15692 (N_15692,N_14447,N_14477);
nor U15693 (N_15693,N_15135,N_15081);
nand U15694 (N_15694,N_14943,N_14669);
or U15695 (N_15695,N_14783,N_14527);
or U15696 (N_15696,N_15049,N_14885);
and U15697 (N_15697,N_14832,N_15098);
xor U15698 (N_15698,N_14420,N_14670);
nand U15699 (N_15699,N_14796,N_14936);
or U15700 (N_15700,N_14909,N_15174);
nand U15701 (N_15701,N_14701,N_14534);
nor U15702 (N_15702,N_15156,N_14768);
nand U15703 (N_15703,N_14797,N_14670);
nand U15704 (N_15704,N_15134,N_14488);
or U15705 (N_15705,N_14615,N_14638);
xnor U15706 (N_15706,N_14542,N_14929);
nand U15707 (N_15707,N_14665,N_14474);
nor U15708 (N_15708,N_14860,N_14472);
nor U15709 (N_15709,N_14434,N_14999);
xnor U15710 (N_15710,N_14548,N_14720);
or U15711 (N_15711,N_14522,N_14757);
nor U15712 (N_15712,N_14776,N_15128);
nor U15713 (N_15713,N_15040,N_14795);
nor U15714 (N_15714,N_14569,N_14690);
nor U15715 (N_15715,N_15116,N_14461);
or U15716 (N_15716,N_14400,N_14617);
xor U15717 (N_15717,N_14743,N_14849);
xnor U15718 (N_15718,N_14677,N_14446);
or U15719 (N_15719,N_14514,N_14432);
xor U15720 (N_15720,N_14941,N_14587);
nand U15721 (N_15721,N_14421,N_14643);
or U15722 (N_15722,N_14623,N_14427);
or U15723 (N_15723,N_14570,N_14617);
and U15724 (N_15724,N_15015,N_15195);
nand U15725 (N_15725,N_14434,N_14967);
nand U15726 (N_15726,N_14990,N_15102);
and U15727 (N_15727,N_14880,N_15062);
and U15728 (N_15728,N_15066,N_14512);
or U15729 (N_15729,N_14957,N_14419);
xnor U15730 (N_15730,N_15071,N_14921);
or U15731 (N_15731,N_15067,N_14850);
nor U15732 (N_15732,N_15179,N_14543);
or U15733 (N_15733,N_14445,N_14414);
xor U15734 (N_15734,N_14744,N_15042);
nand U15735 (N_15735,N_15104,N_14469);
xor U15736 (N_15736,N_15192,N_15055);
nor U15737 (N_15737,N_14923,N_14418);
or U15738 (N_15738,N_14483,N_14586);
nand U15739 (N_15739,N_14471,N_15015);
or U15740 (N_15740,N_14551,N_15131);
nor U15741 (N_15741,N_14603,N_14923);
xor U15742 (N_15742,N_15187,N_15069);
nor U15743 (N_15743,N_14876,N_14899);
nand U15744 (N_15744,N_15143,N_14707);
nand U15745 (N_15745,N_14962,N_14864);
and U15746 (N_15746,N_14517,N_14899);
nor U15747 (N_15747,N_14807,N_14480);
xnor U15748 (N_15748,N_14542,N_14843);
and U15749 (N_15749,N_14606,N_15170);
nor U15750 (N_15750,N_14721,N_14812);
nor U15751 (N_15751,N_14790,N_14438);
or U15752 (N_15752,N_15197,N_14892);
and U15753 (N_15753,N_14858,N_15000);
and U15754 (N_15754,N_14467,N_14977);
xor U15755 (N_15755,N_14594,N_15187);
nand U15756 (N_15756,N_14751,N_14784);
or U15757 (N_15757,N_15039,N_14594);
xnor U15758 (N_15758,N_15033,N_15198);
nor U15759 (N_15759,N_14428,N_15116);
nor U15760 (N_15760,N_15162,N_14487);
nor U15761 (N_15761,N_15065,N_14853);
nor U15762 (N_15762,N_14884,N_14902);
and U15763 (N_15763,N_14654,N_15005);
nor U15764 (N_15764,N_14644,N_14492);
and U15765 (N_15765,N_14746,N_14892);
nor U15766 (N_15766,N_15040,N_14931);
nor U15767 (N_15767,N_14514,N_15177);
and U15768 (N_15768,N_15188,N_14919);
or U15769 (N_15769,N_15048,N_14618);
and U15770 (N_15770,N_14463,N_14729);
nor U15771 (N_15771,N_14799,N_14741);
and U15772 (N_15772,N_14818,N_14509);
nand U15773 (N_15773,N_14499,N_14469);
and U15774 (N_15774,N_14451,N_14631);
or U15775 (N_15775,N_15143,N_14476);
nor U15776 (N_15776,N_14870,N_14415);
nand U15777 (N_15777,N_14818,N_15042);
or U15778 (N_15778,N_14559,N_15016);
nor U15779 (N_15779,N_15195,N_15139);
or U15780 (N_15780,N_14894,N_15092);
and U15781 (N_15781,N_15020,N_14491);
nand U15782 (N_15782,N_14705,N_14951);
nand U15783 (N_15783,N_15146,N_14409);
or U15784 (N_15784,N_15199,N_14644);
xnor U15785 (N_15785,N_14937,N_14450);
nand U15786 (N_15786,N_14538,N_14946);
and U15787 (N_15787,N_14576,N_14436);
nor U15788 (N_15788,N_15099,N_14859);
nand U15789 (N_15789,N_14817,N_14917);
xnor U15790 (N_15790,N_14445,N_14866);
nand U15791 (N_15791,N_15193,N_14602);
or U15792 (N_15792,N_15102,N_14637);
and U15793 (N_15793,N_15152,N_14780);
and U15794 (N_15794,N_14574,N_15182);
nor U15795 (N_15795,N_14617,N_15107);
or U15796 (N_15796,N_14877,N_15056);
or U15797 (N_15797,N_14961,N_14864);
and U15798 (N_15798,N_14664,N_14414);
nand U15799 (N_15799,N_15167,N_15152);
or U15800 (N_15800,N_14948,N_14750);
nand U15801 (N_15801,N_14801,N_14510);
nand U15802 (N_15802,N_14506,N_14918);
or U15803 (N_15803,N_14555,N_14472);
nand U15804 (N_15804,N_15138,N_14781);
xnor U15805 (N_15805,N_15172,N_14837);
or U15806 (N_15806,N_14956,N_14413);
nor U15807 (N_15807,N_14820,N_14496);
nand U15808 (N_15808,N_14807,N_14552);
xnor U15809 (N_15809,N_14425,N_14463);
or U15810 (N_15810,N_14659,N_14882);
xnor U15811 (N_15811,N_14755,N_14970);
xor U15812 (N_15812,N_14670,N_15198);
xor U15813 (N_15813,N_14719,N_15058);
nand U15814 (N_15814,N_14489,N_14478);
nand U15815 (N_15815,N_14739,N_15094);
xor U15816 (N_15816,N_14728,N_14739);
xor U15817 (N_15817,N_14994,N_14805);
xor U15818 (N_15818,N_14589,N_15102);
xnor U15819 (N_15819,N_15179,N_15059);
and U15820 (N_15820,N_15132,N_14953);
and U15821 (N_15821,N_14517,N_14895);
xnor U15822 (N_15822,N_14637,N_14820);
or U15823 (N_15823,N_14688,N_15015);
or U15824 (N_15824,N_14708,N_14634);
or U15825 (N_15825,N_14966,N_14421);
xor U15826 (N_15826,N_15172,N_14913);
nor U15827 (N_15827,N_14941,N_14474);
and U15828 (N_15828,N_14883,N_14911);
nor U15829 (N_15829,N_14977,N_15023);
and U15830 (N_15830,N_14607,N_15179);
nand U15831 (N_15831,N_15089,N_15179);
nor U15832 (N_15832,N_14790,N_14726);
and U15833 (N_15833,N_14422,N_14472);
or U15834 (N_15834,N_14855,N_15008);
nand U15835 (N_15835,N_15194,N_14572);
xor U15836 (N_15836,N_14987,N_15094);
xor U15837 (N_15837,N_15072,N_14590);
nand U15838 (N_15838,N_14647,N_14857);
xor U15839 (N_15839,N_14682,N_14744);
or U15840 (N_15840,N_15133,N_14784);
nor U15841 (N_15841,N_15140,N_14744);
nand U15842 (N_15842,N_14812,N_15193);
xor U15843 (N_15843,N_14875,N_14798);
nor U15844 (N_15844,N_14874,N_14928);
xor U15845 (N_15845,N_14620,N_15014);
or U15846 (N_15846,N_14980,N_14455);
and U15847 (N_15847,N_14663,N_14832);
nand U15848 (N_15848,N_15060,N_15017);
nor U15849 (N_15849,N_14504,N_14982);
nor U15850 (N_15850,N_14632,N_15005);
nor U15851 (N_15851,N_14516,N_14661);
xnor U15852 (N_15852,N_14573,N_14426);
nand U15853 (N_15853,N_14815,N_14468);
nor U15854 (N_15854,N_14700,N_15156);
nor U15855 (N_15855,N_14565,N_14994);
or U15856 (N_15856,N_14741,N_14592);
xor U15857 (N_15857,N_14866,N_14629);
and U15858 (N_15858,N_15070,N_14950);
nor U15859 (N_15859,N_14503,N_14894);
and U15860 (N_15860,N_15135,N_14662);
or U15861 (N_15861,N_14780,N_14663);
xnor U15862 (N_15862,N_14448,N_14677);
and U15863 (N_15863,N_14533,N_15090);
nor U15864 (N_15864,N_14820,N_14805);
nor U15865 (N_15865,N_15127,N_14591);
xnor U15866 (N_15866,N_15049,N_14464);
and U15867 (N_15867,N_15027,N_14520);
nor U15868 (N_15868,N_15057,N_14982);
or U15869 (N_15869,N_14494,N_14927);
xnor U15870 (N_15870,N_14457,N_14772);
nand U15871 (N_15871,N_14516,N_14707);
and U15872 (N_15872,N_14938,N_15130);
and U15873 (N_15873,N_14962,N_14598);
xor U15874 (N_15874,N_15034,N_14694);
or U15875 (N_15875,N_15013,N_14785);
nand U15876 (N_15876,N_14472,N_14935);
nand U15877 (N_15877,N_14603,N_14856);
or U15878 (N_15878,N_15172,N_14758);
nor U15879 (N_15879,N_14506,N_15062);
and U15880 (N_15880,N_15179,N_14688);
and U15881 (N_15881,N_14641,N_15078);
or U15882 (N_15882,N_14405,N_14973);
nor U15883 (N_15883,N_14899,N_14434);
nor U15884 (N_15884,N_14636,N_15062);
nand U15885 (N_15885,N_14929,N_14868);
xor U15886 (N_15886,N_14618,N_14705);
or U15887 (N_15887,N_14783,N_14759);
nor U15888 (N_15888,N_15137,N_15093);
xor U15889 (N_15889,N_14881,N_14419);
nand U15890 (N_15890,N_14933,N_14582);
and U15891 (N_15891,N_15197,N_14877);
or U15892 (N_15892,N_15066,N_15115);
nor U15893 (N_15893,N_14648,N_14821);
and U15894 (N_15894,N_14930,N_14715);
nor U15895 (N_15895,N_15066,N_15147);
nor U15896 (N_15896,N_14538,N_14591);
or U15897 (N_15897,N_14508,N_14849);
and U15898 (N_15898,N_14427,N_14492);
and U15899 (N_15899,N_14931,N_14763);
and U15900 (N_15900,N_14706,N_15132);
xor U15901 (N_15901,N_14408,N_14637);
xor U15902 (N_15902,N_14634,N_15011);
or U15903 (N_15903,N_14536,N_15096);
or U15904 (N_15904,N_15176,N_14451);
nand U15905 (N_15905,N_14466,N_14475);
xnor U15906 (N_15906,N_14449,N_14590);
and U15907 (N_15907,N_14923,N_14649);
or U15908 (N_15908,N_14742,N_14936);
nor U15909 (N_15909,N_14430,N_14551);
xnor U15910 (N_15910,N_14585,N_15124);
or U15911 (N_15911,N_15017,N_14789);
nor U15912 (N_15912,N_14433,N_14741);
and U15913 (N_15913,N_14880,N_14810);
nand U15914 (N_15914,N_14584,N_14580);
xnor U15915 (N_15915,N_14743,N_14445);
nor U15916 (N_15916,N_14906,N_14820);
or U15917 (N_15917,N_15152,N_14925);
and U15918 (N_15918,N_15105,N_14945);
and U15919 (N_15919,N_14461,N_14765);
xor U15920 (N_15920,N_14964,N_14625);
or U15921 (N_15921,N_15113,N_15162);
or U15922 (N_15922,N_14477,N_14405);
or U15923 (N_15923,N_15087,N_14525);
nand U15924 (N_15924,N_14568,N_14513);
nor U15925 (N_15925,N_14882,N_14574);
nand U15926 (N_15926,N_14490,N_14574);
nor U15927 (N_15927,N_15109,N_14906);
nor U15928 (N_15928,N_14755,N_14674);
nor U15929 (N_15929,N_14786,N_14626);
nand U15930 (N_15930,N_14935,N_14913);
and U15931 (N_15931,N_14716,N_14735);
nor U15932 (N_15932,N_14636,N_14488);
xnor U15933 (N_15933,N_15020,N_14771);
and U15934 (N_15934,N_14457,N_14884);
or U15935 (N_15935,N_14583,N_14798);
nor U15936 (N_15936,N_14866,N_14627);
or U15937 (N_15937,N_14671,N_14510);
nand U15938 (N_15938,N_15051,N_14569);
xnor U15939 (N_15939,N_14885,N_14891);
nand U15940 (N_15940,N_14480,N_15045);
nand U15941 (N_15941,N_14874,N_14717);
or U15942 (N_15942,N_14905,N_14820);
nand U15943 (N_15943,N_15128,N_14700);
nor U15944 (N_15944,N_14928,N_15062);
or U15945 (N_15945,N_14439,N_14857);
nand U15946 (N_15946,N_15117,N_14507);
nor U15947 (N_15947,N_14791,N_14792);
and U15948 (N_15948,N_14534,N_15162);
nor U15949 (N_15949,N_14832,N_14904);
or U15950 (N_15950,N_14810,N_15015);
or U15951 (N_15951,N_14852,N_14994);
or U15952 (N_15952,N_14449,N_14927);
nand U15953 (N_15953,N_14720,N_15101);
or U15954 (N_15954,N_14693,N_14747);
and U15955 (N_15955,N_15151,N_14626);
nand U15956 (N_15956,N_14876,N_14880);
and U15957 (N_15957,N_14760,N_15012);
or U15958 (N_15958,N_14995,N_15169);
xnor U15959 (N_15959,N_14776,N_14508);
or U15960 (N_15960,N_14687,N_14681);
xor U15961 (N_15961,N_14963,N_14669);
nor U15962 (N_15962,N_15047,N_15057);
nand U15963 (N_15963,N_14874,N_14989);
xor U15964 (N_15964,N_15159,N_15190);
nor U15965 (N_15965,N_14979,N_14467);
nand U15966 (N_15966,N_14608,N_14548);
xor U15967 (N_15967,N_15142,N_15164);
xnor U15968 (N_15968,N_14614,N_14844);
nand U15969 (N_15969,N_15129,N_15084);
xnor U15970 (N_15970,N_15051,N_14862);
xnor U15971 (N_15971,N_14511,N_15095);
nor U15972 (N_15972,N_14608,N_14600);
nor U15973 (N_15973,N_14890,N_14424);
xnor U15974 (N_15974,N_14697,N_14794);
xor U15975 (N_15975,N_14928,N_14602);
nor U15976 (N_15976,N_14869,N_14723);
and U15977 (N_15977,N_14980,N_15153);
nand U15978 (N_15978,N_14722,N_15054);
nor U15979 (N_15979,N_15034,N_14685);
and U15980 (N_15980,N_14781,N_15151);
or U15981 (N_15981,N_15198,N_14929);
nand U15982 (N_15982,N_14511,N_15147);
nand U15983 (N_15983,N_14650,N_14735);
or U15984 (N_15984,N_14778,N_14688);
nand U15985 (N_15985,N_14808,N_15114);
nand U15986 (N_15986,N_14935,N_14626);
or U15987 (N_15987,N_14871,N_15109);
or U15988 (N_15988,N_15173,N_14917);
and U15989 (N_15989,N_14910,N_14595);
xor U15990 (N_15990,N_14772,N_14490);
nor U15991 (N_15991,N_14756,N_14950);
or U15992 (N_15992,N_14729,N_14608);
and U15993 (N_15993,N_14866,N_14521);
nand U15994 (N_15994,N_15043,N_15100);
nand U15995 (N_15995,N_14969,N_14983);
nand U15996 (N_15996,N_14401,N_14573);
nor U15997 (N_15997,N_14498,N_14537);
nand U15998 (N_15998,N_15186,N_15050);
nand U15999 (N_15999,N_14502,N_15057);
nand U16000 (N_16000,N_15503,N_15980);
nor U16001 (N_16001,N_15693,N_15886);
nor U16002 (N_16002,N_15700,N_15501);
nor U16003 (N_16003,N_15630,N_15297);
or U16004 (N_16004,N_15836,N_15466);
and U16005 (N_16005,N_15935,N_15916);
or U16006 (N_16006,N_15924,N_15462);
and U16007 (N_16007,N_15519,N_15629);
nor U16008 (N_16008,N_15239,N_15919);
nand U16009 (N_16009,N_15557,N_15270);
nand U16010 (N_16010,N_15614,N_15750);
nand U16011 (N_16011,N_15269,N_15400);
and U16012 (N_16012,N_15648,N_15995);
nor U16013 (N_16013,N_15350,N_15439);
xor U16014 (N_16014,N_15374,N_15522);
xnor U16015 (N_16015,N_15699,N_15384);
and U16016 (N_16016,N_15344,N_15786);
or U16017 (N_16017,N_15705,N_15277);
nand U16018 (N_16018,N_15500,N_15440);
xnor U16019 (N_16019,N_15704,N_15621);
nor U16020 (N_16020,N_15494,N_15562);
and U16021 (N_16021,N_15472,N_15229);
nor U16022 (N_16022,N_15335,N_15638);
nand U16023 (N_16023,N_15746,N_15302);
xor U16024 (N_16024,N_15727,N_15873);
xor U16025 (N_16025,N_15487,N_15837);
and U16026 (N_16026,N_15207,N_15352);
nand U16027 (N_16027,N_15737,N_15778);
xor U16028 (N_16028,N_15906,N_15917);
and U16029 (N_16029,N_15575,N_15251);
nor U16030 (N_16030,N_15521,N_15690);
and U16031 (N_16031,N_15976,N_15663);
nor U16032 (N_16032,N_15835,N_15734);
xnor U16033 (N_16033,N_15781,N_15530);
or U16034 (N_16034,N_15764,N_15831);
or U16035 (N_16035,N_15225,N_15801);
xor U16036 (N_16036,N_15461,N_15291);
nor U16037 (N_16037,N_15744,N_15210);
and U16038 (N_16038,N_15416,N_15850);
and U16039 (N_16039,N_15900,N_15565);
or U16040 (N_16040,N_15427,N_15459);
nand U16041 (N_16041,N_15814,N_15475);
xor U16042 (N_16042,N_15890,N_15369);
and U16043 (N_16043,N_15967,N_15798);
nand U16044 (N_16044,N_15852,N_15279);
nor U16045 (N_16045,N_15759,N_15767);
and U16046 (N_16046,N_15425,N_15482);
or U16047 (N_16047,N_15930,N_15914);
nand U16048 (N_16048,N_15548,N_15544);
nor U16049 (N_16049,N_15550,N_15212);
nand U16050 (N_16050,N_15288,N_15423);
nand U16051 (N_16051,N_15766,N_15318);
nand U16052 (N_16052,N_15576,N_15901);
and U16053 (N_16053,N_15345,N_15267);
xnor U16054 (N_16054,N_15419,N_15720);
and U16055 (N_16055,N_15712,N_15431);
xnor U16056 (N_16056,N_15992,N_15964);
xor U16057 (N_16057,N_15933,N_15396);
and U16058 (N_16058,N_15538,N_15249);
xor U16059 (N_16059,N_15853,N_15787);
xor U16060 (N_16060,N_15309,N_15960);
and U16061 (N_16061,N_15221,N_15594);
or U16062 (N_16062,N_15851,N_15246);
nor U16063 (N_16063,N_15686,N_15259);
and U16064 (N_16064,N_15479,N_15595);
xor U16065 (N_16065,N_15422,N_15637);
nor U16066 (N_16066,N_15862,N_15202);
xor U16067 (N_16067,N_15449,N_15512);
xor U16068 (N_16068,N_15551,N_15904);
or U16069 (N_16069,N_15633,N_15331);
or U16070 (N_16070,N_15962,N_15473);
xor U16071 (N_16071,N_15460,N_15793);
or U16072 (N_16072,N_15857,N_15819);
nor U16073 (N_16073,N_15628,N_15413);
nand U16074 (N_16074,N_15791,N_15278);
nor U16075 (N_16075,N_15478,N_15896);
or U16076 (N_16076,N_15321,N_15840);
and U16077 (N_16077,N_15861,N_15244);
xor U16078 (N_16078,N_15367,N_15817);
and U16079 (N_16079,N_15273,N_15553);
and U16080 (N_16080,N_15866,N_15903);
nor U16081 (N_16081,N_15932,N_15891);
or U16082 (N_16082,N_15841,N_15397);
nand U16083 (N_16083,N_15676,N_15540);
xor U16084 (N_16084,N_15560,N_15999);
or U16085 (N_16085,N_15796,N_15579);
and U16086 (N_16086,N_15597,N_15464);
and U16087 (N_16087,N_15457,N_15811);
or U16088 (N_16088,N_15523,N_15253);
xnor U16089 (N_16089,N_15966,N_15826);
nor U16090 (N_16090,N_15320,N_15592);
nor U16091 (N_16091,N_15739,N_15490);
nand U16092 (N_16092,N_15871,N_15788);
nor U16093 (N_16093,N_15784,N_15728);
and U16094 (N_16094,N_15343,N_15254);
xnor U16095 (N_16095,N_15405,N_15310);
xnor U16096 (N_16096,N_15542,N_15465);
or U16097 (N_16097,N_15589,N_15799);
nor U16098 (N_16098,N_15263,N_15359);
and U16099 (N_16099,N_15373,N_15392);
or U16100 (N_16100,N_15450,N_15453);
or U16101 (N_16101,N_15923,N_15566);
and U16102 (N_16102,N_15687,N_15527);
xnor U16103 (N_16103,N_15435,N_15447);
nand U16104 (N_16104,N_15902,N_15213);
nand U16105 (N_16105,N_15394,N_15701);
nor U16106 (N_16106,N_15326,N_15623);
nor U16107 (N_16107,N_15685,N_15681);
and U16108 (N_16108,N_15395,N_15651);
nor U16109 (N_16109,N_15642,N_15204);
and U16110 (N_16110,N_15771,N_15387);
and U16111 (N_16111,N_15883,N_15879);
nand U16112 (N_16112,N_15358,N_15554);
and U16113 (N_16113,N_15646,N_15806);
or U16114 (N_16114,N_15808,N_15418);
and U16115 (N_16115,N_15768,N_15751);
xor U16116 (N_16116,N_15371,N_15401);
nand U16117 (N_16117,N_15588,N_15430);
xor U16118 (N_16118,N_15558,N_15807);
and U16119 (N_16119,N_15242,N_15997);
and U16120 (N_16120,N_15481,N_15616);
and U16121 (N_16121,N_15934,N_15573);
nand U16122 (N_16122,N_15282,N_15828);
or U16123 (N_16123,N_15846,N_15293);
nor U16124 (N_16124,N_15234,N_15201);
and U16125 (N_16125,N_15668,N_15908);
or U16126 (N_16126,N_15514,N_15510);
xor U16127 (N_16127,N_15216,N_15314);
xnor U16128 (N_16128,N_15363,N_15518);
nand U16129 (N_16129,N_15477,N_15232);
xnor U16130 (N_16130,N_15657,N_15738);
nand U16131 (N_16131,N_15609,N_15617);
xor U16132 (N_16132,N_15532,N_15655);
nand U16133 (N_16133,N_15304,N_15390);
xor U16134 (N_16134,N_15910,N_15756);
or U16135 (N_16135,N_15794,N_15368);
xor U16136 (N_16136,N_15984,N_15695);
nor U16137 (N_16137,N_15236,N_15292);
nor U16138 (N_16138,N_15803,N_15349);
xnor U16139 (N_16139,N_15260,N_15590);
xor U16140 (N_16140,N_15446,N_15978);
or U16141 (N_16141,N_15949,N_15805);
or U16142 (N_16142,N_15892,N_15209);
or U16143 (N_16143,N_15876,N_15718);
or U16144 (N_16144,N_15287,N_15989);
and U16145 (N_16145,N_15333,N_15606);
or U16146 (N_16146,N_15240,N_15208);
nor U16147 (N_16147,N_15420,N_15280);
nand U16148 (N_16148,N_15535,N_15945);
xnor U16149 (N_16149,N_15337,N_15731);
nand U16150 (N_16150,N_15561,N_15568);
and U16151 (N_16151,N_15821,N_15290);
nor U16152 (N_16152,N_15328,N_15947);
nand U16153 (N_16153,N_15312,N_15436);
xnor U16154 (N_16154,N_15943,N_15858);
nand U16155 (N_16155,N_15958,N_15228);
xnor U16156 (N_16156,N_15211,N_15812);
nor U16157 (N_16157,N_15809,N_15383);
xnor U16158 (N_16158,N_15714,N_15563);
and U16159 (N_16159,N_15313,N_15596);
xnor U16160 (N_16160,N_15713,N_15719);
or U16161 (N_16161,N_15769,N_15643);
nand U16162 (N_16162,N_15878,N_15627);
xnor U16163 (N_16163,N_15275,N_15773);
and U16164 (N_16164,N_15777,N_15488);
nor U16165 (N_16165,N_15591,N_15533);
nand U16166 (N_16166,N_15804,N_15377);
nand U16167 (N_16167,N_15515,N_15990);
nand U16168 (N_16168,N_15889,N_15931);
and U16169 (N_16169,N_15770,N_15670);
nor U16170 (N_16170,N_15403,N_15336);
xor U16171 (N_16171,N_15775,N_15342);
and U16172 (N_16172,N_15379,N_15537);
nor U16173 (N_16173,N_15380,N_15939);
or U16174 (N_16174,N_15842,N_15559);
and U16175 (N_16175,N_15619,N_15707);
nand U16176 (N_16176,N_15755,N_15341);
nor U16177 (N_16177,N_15913,N_15255);
or U16178 (N_16178,N_15445,N_15956);
and U16179 (N_16179,N_15864,N_15790);
or U16180 (N_16180,N_15385,N_15742);
nor U16181 (N_16181,N_15970,N_15289);
nor U16182 (N_16182,N_15634,N_15417);
xor U16183 (N_16183,N_15856,N_15398);
xnor U16184 (N_16184,N_15581,N_15351);
nor U16185 (N_16185,N_15237,N_15758);
nand U16186 (N_16186,N_15894,N_15334);
nor U16187 (N_16187,N_15426,N_15206);
nand U16188 (N_16188,N_15415,N_15644);
and U16189 (N_16189,N_15584,N_15613);
and U16190 (N_16190,N_15959,N_15977);
nand U16191 (N_16191,N_15315,N_15492);
nor U16192 (N_16192,N_15441,N_15647);
or U16193 (N_16193,N_15907,N_15531);
nor U16194 (N_16194,N_15455,N_15872);
or U16195 (N_16195,N_15376,N_15496);
nor U16196 (N_16196,N_15528,N_15620);
nand U16197 (N_16197,N_15433,N_15607);
nor U16198 (N_16198,N_15982,N_15509);
nand U16199 (N_16199,N_15300,N_15414);
and U16200 (N_16200,N_15386,N_15583);
or U16201 (N_16201,N_15716,N_15372);
or U16202 (N_16202,N_15996,N_15513);
or U16203 (N_16203,N_15965,N_15498);
and U16204 (N_16204,N_15451,N_15823);
nand U16205 (N_16205,N_15732,N_15274);
or U16206 (N_16206,N_15493,N_15941);
nor U16207 (N_16207,N_15844,N_15863);
and U16208 (N_16208,N_15895,N_15677);
or U16209 (N_16209,N_15975,N_15929);
nand U16210 (N_16210,N_15258,N_15887);
xor U16211 (N_16211,N_15485,N_15968);
nand U16212 (N_16212,N_15832,N_15944);
xor U16213 (N_16213,N_15316,N_15480);
nor U16214 (N_16214,N_15231,N_15268);
or U16215 (N_16215,N_15653,N_15937);
nand U16216 (N_16216,N_15516,N_15950);
nand U16217 (N_16217,N_15323,N_15656);
and U16218 (N_16218,N_15438,N_15869);
nand U16219 (N_16219,N_15662,N_15536);
or U16220 (N_16220,N_15783,N_15985);
nor U16221 (N_16221,N_15322,N_15694);
nand U16222 (N_16222,N_15296,N_15816);
or U16223 (N_16223,N_15813,N_15649);
and U16224 (N_16224,N_15709,N_15424);
or U16225 (N_16225,N_15266,N_15303);
and U16226 (N_16226,N_15715,N_15262);
xnor U16227 (N_16227,N_15308,N_15672);
nand U16228 (N_16228,N_15993,N_15955);
and U16229 (N_16229,N_15332,N_15969);
nor U16230 (N_16230,N_15698,N_15586);
nand U16231 (N_16231,N_15833,N_15437);
nor U16232 (N_16232,N_15717,N_15612);
nor U16233 (N_16233,N_15257,N_15311);
or U16234 (N_16234,N_15870,N_15330);
or U16235 (N_16235,N_15603,N_15600);
nor U16236 (N_16236,N_15410,N_15608);
or U16237 (N_16237,N_15227,N_15381);
and U16238 (N_16238,N_15355,N_15725);
nand U16239 (N_16239,N_15624,N_15625);
and U16240 (N_16240,N_15505,N_15854);
and U16241 (N_16241,N_15782,N_15543);
nor U16242 (N_16242,N_15520,N_15529);
and U16243 (N_16243,N_15800,N_15248);
or U16244 (N_16244,N_15618,N_15382);
or U16245 (N_16245,N_15411,N_15598);
and U16246 (N_16246,N_15748,N_15795);
xor U16247 (N_16247,N_15261,N_15664);
nor U16248 (N_16248,N_15660,N_15703);
and U16249 (N_16249,N_15409,N_15294);
or U16250 (N_16250,N_15922,N_15679);
xor U16251 (N_16251,N_15972,N_15476);
nor U16252 (N_16252,N_15217,N_15688);
or U16253 (N_16253,N_15407,N_15868);
nor U16254 (N_16254,N_15245,N_15585);
and U16255 (N_16255,N_15843,N_15508);
xnor U16256 (N_16256,N_15752,N_15635);
or U16257 (N_16257,N_15406,N_15545);
nor U16258 (N_16258,N_15247,N_15789);
and U16259 (N_16259,N_15375,N_15348);
and U16260 (N_16260,N_15855,N_15525);
nand U16261 (N_16261,N_15730,N_15593);
and U16262 (N_16262,N_15658,N_15468);
nand U16263 (N_16263,N_15393,N_15983);
xnor U16264 (N_16264,N_15539,N_15489);
nand U16265 (N_16265,N_15745,N_15366);
nand U16266 (N_16266,N_15491,N_15675);
nand U16267 (N_16267,N_15541,N_15301);
or U16268 (N_16268,N_15546,N_15797);
nor U16269 (N_16269,N_15669,N_15741);
xnor U16270 (N_16270,N_15986,N_15306);
and U16271 (N_16271,N_15605,N_15953);
nand U16272 (N_16272,N_15325,N_15626);
and U16273 (N_16273,N_15684,N_15779);
xnor U16274 (N_16274,N_15827,N_15994);
nand U16275 (N_16275,N_15680,N_15495);
and U16276 (N_16276,N_15226,N_15243);
or U16277 (N_16277,N_15327,N_15942);
nand U16278 (N_16278,N_15517,N_15356);
and U16279 (N_16279,N_15250,N_15567);
nor U16280 (N_16280,N_15432,N_15428);
and U16281 (N_16281,N_15364,N_15859);
and U16282 (N_16282,N_15319,N_15346);
xor U16283 (N_16283,N_15448,N_15998);
and U16284 (N_16284,N_15483,N_15893);
nor U16285 (N_16285,N_15329,N_15927);
nand U16286 (N_16286,N_15574,N_15645);
nand U16287 (N_16287,N_15458,N_15404);
or U16288 (N_16288,N_15353,N_15421);
nor U16289 (N_16289,N_15682,N_15442);
nand U16290 (N_16290,N_15252,N_15979);
nand U16291 (N_16291,N_15761,N_15378);
or U16292 (N_16292,N_15285,N_15470);
and U16293 (N_16293,N_15912,N_15564);
nor U16294 (N_16294,N_15988,N_15921);
xnor U16295 (N_16295,N_15898,N_15722);
or U16296 (N_16296,N_15848,N_15763);
nor U16297 (N_16297,N_15641,N_15880);
and U16298 (N_16298,N_15578,N_15860);
and U16299 (N_16299,N_15954,N_15951);
nor U16300 (N_16300,N_15723,N_15471);
nor U16301 (N_16301,N_15678,N_15399);
nand U16302 (N_16302,N_15230,N_15760);
or U16303 (N_16303,N_15504,N_15610);
and U16304 (N_16304,N_15961,N_15365);
or U16305 (N_16305,N_15220,N_15203);
xnor U16306 (N_16306,N_15952,N_15830);
nand U16307 (N_16307,N_15264,N_15726);
nand U16308 (N_16308,N_15604,N_15486);
or U16309 (N_16309,N_15652,N_15469);
and U16310 (N_16310,N_15357,N_15911);
and U16311 (N_16311,N_15444,N_15456);
nor U16312 (N_16312,N_15205,N_15214);
or U16313 (N_16313,N_15391,N_15785);
or U16314 (N_16314,N_15671,N_15599);
xnor U16315 (N_16315,N_15283,N_15307);
and U16316 (N_16316,N_15733,N_15272);
xor U16317 (N_16317,N_15926,N_15877);
and U16318 (N_16318,N_15915,N_15340);
nand U16319 (N_16319,N_15347,N_15354);
xnor U16320 (N_16320,N_15666,N_15632);
nand U16321 (N_16321,N_15361,N_15936);
nand U16322 (N_16322,N_15697,N_15650);
nand U16323 (N_16323,N_15925,N_15569);
xor U16324 (N_16324,N_15888,N_15754);
nand U16325 (N_16325,N_15991,N_15434);
nand U16326 (N_16326,N_15780,N_15665);
xor U16327 (N_16327,N_15388,N_15654);
nand U16328 (N_16328,N_15463,N_15762);
or U16329 (N_16329,N_15281,N_15615);
nand U16330 (N_16330,N_15577,N_15484);
nand U16331 (N_16331,N_15729,N_15218);
xor U16332 (N_16332,N_15899,N_15526);
nand U16333 (N_16333,N_15305,N_15815);
xnor U16334 (N_16334,N_15611,N_15882);
and U16335 (N_16335,N_15757,N_15587);
nor U16336 (N_16336,N_15847,N_15667);
or U16337 (N_16337,N_15339,N_15572);
nor U16338 (N_16338,N_15838,N_15601);
and U16339 (N_16339,N_15219,N_15298);
and U16340 (N_16340,N_15412,N_15920);
xnor U16341 (N_16341,N_15256,N_15820);
or U16342 (N_16342,N_15834,N_15235);
or U16343 (N_16343,N_15511,N_15631);
nor U16344 (N_16344,N_15200,N_15223);
nor U16345 (N_16345,N_15948,N_15810);
and U16346 (N_16346,N_15580,N_15696);
and U16347 (N_16347,N_15659,N_15317);
and U16348 (N_16348,N_15776,N_15743);
or U16349 (N_16349,N_15940,N_15408);
or U16350 (N_16350,N_15556,N_15753);
nor U16351 (N_16351,N_15674,N_15822);
nand U16352 (N_16352,N_15443,N_15640);
and U16353 (N_16353,N_15324,N_15502);
nor U16354 (N_16354,N_15710,N_15711);
nor U16355 (N_16355,N_15222,N_15692);
nor U16356 (N_16356,N_15362,N_15338);
and U16357 (N_16357,N_15987,N_15845);
xnor U16358 (N_16358,N_15389,N_15499);
or U16359 (N_16359,N_15981,N_15849);
nand U16360 (N_16360,N_15973,N_15474);
nand U16361 (N_16361,N_15452,N_15467);
or U16362 (N_16362,N_15497,N_15691);
xor U16363 (N_16363,N_15885,N_15874);
nand U16364 (N_16364,N_15747,N_15772);
and U16365 (N_16365,N_15689,N_15881);
nand U16366 (N_16366,N_15286,N_15602);
nand U16367 (N_16367,N_15233,N_15524);
and U16368 (N_16368,N_15774,N_15549);
nor U16369 (N_16369,N_15839,N_15702);
nand U16370 (N_16370,N_15909,N_15946);
nor U16371 (N_16371,N_15271,N_15360);
xor U16372 (N_16372,N_15829,N_15276);
and U16373 (N_16373,N_15875,N_15765);
and U16374 (N_16374,N_15547,N_15215);
xor U16375 (N_16375,N_15534,N_15661);
nand U16376 (N_16376,N_15454,N_15636);
nor U16377 (N_16377,N_15818,N_15639);
or U16378 (N_16378,N_15867,N_15370);
or U16379 (N_16379,N_15708,N_15865);
and U16380 (N_16380,N_15429,N_15802);
xnor U16381 (N_16381,N_15971,N_15963);
nor U16382 (N_16382,N_15918,N_15792);
nand U16383 (N_16383,N_15724,N_15241);
xnor U16384 (N_16384,N_15905,N_15749);
nand U16385 (N_16385,N_15736,N_15552);
xor U16386 (N_16386,N_15571,N_15299);
or U16387 (N_16387,N_15884,N_15570);
or U16388 (N_16388,N_15582,N_15740);
xor U16389 (N_16389,N_15506,N_15402);
nor U16390 (N_16390,N_15555,N_15928);
or U16391 (N_16391,N_15295,N_15957);
or U16392 (N_16392,N_15224,N_15238);
xor U16393 (N_16393,N_15721,N_15897);
nor U16394 (N_16394,N_15284,N_15706);
xor U16395 (N_16395,N_15683,N_15825);
or U16396 (N_16396,N_15974,N_15824);
nand U16397 (N_16397,N_15673,N_15938);
nor U16398 (N_16398,N_15507,N_15265);
or U16399 (N_16399,N_15622,N_15735);
or U16400 (N_16400,N_15762,N_15697);
nor U16401 (N_16401,N_15923,N_15843);
nor U16402 (N_16402,N_15786,N_15793);
xor U16403 (N_16403,N_15731,N_15335);
nor U16404 (N_16404,N_15280,N_15249);
and U16405 (N_16405,N_15524,N_15924);
nand U16406 (N_16406,N_15344,N_15289);
nand U16407 (N_16407,N_15350,N_15390);
xnor U16408 (N_16408,N_15697,N_15785);
nor U16409 (N_16409,N_15467,N_15650);
and U16410 (N_16410,N_15749,N_15309);
nor U16411 (N_16411,N_15370,N_15488);
or U16412 (N_16412,N_15451,N_15400);
and U16413 (N_16413,N_15498,N_15603);
or U16414 (N_16414,N_15851,N_15206);
nor U16415 (N_16415,N_15818,N_15849);
and U16416 (N_16416,N_15387,N_15345);
and U16417 (N_16417,N_15927,N_15662);
nor U16418 (N_16418,N_15796,N_15751);
nand U16419 (N_16419,N_15760,N_15816);
xnor U16420 (N_16420,N_15504,N_15750);
and U16421 (N_16421,N_15954,N_15900);
nand U16422 (N_16422,N_15358,N_15794);
and U16423 (N_16423,N_15821,N_15651);
nand U16424 (N_16424,N_15955,N_15935);
nor U16425 (N_16425,N_15563,N_15831);
nor U16426 (N_16426,N_15955,N_15518);
nand U16427 (N_16427,N_15378,N_15467);
nor U16428 (N_16428,N_15929,N_15339);
and U16429 (N_16429,N_15840,N_15487);
or U16430 (N_16430,N_15233,N_15509);
nand U16431 (N_16431,N_15439,N_15438);
and U16432 (N_16432,N_15555,N_15993);
nor U16433 (N_16433,N_15771,N_15281);
and U16434 (N_16434,N_15408,N_15933);
nand U16435 (N_16435,N_15581,N_15705);
xor U16436 (N_16436,N_15537,N_15458);
xor U16437 (N_16437,N_15229,N_15298);
nand U16438 (N_16438,N_15971,N_15553);
and U16439 (N_16439,N_15773,N_15647);
or U16440 (N_16440,N_15300,N_15634);
nand U16441 (N_16441,N_15965,N_15271);
or U16442 (N_16442,N_15312,N_15250);
xnor U16443 (N_16443,N_15991,N_15239);
nor U16444 (N_16444,N_15410,N_15252);
nor U16445 (N_16445,N_15950,N_15208);
or U16446 (N_16446,N_15785,N_15214);
and U16447 (N_16447,N_15884,N_15241);
nand U16448 (N_16448,N_15845,N_15523);
or U16449 (N_16449,N_15313,N_15382);
xor U16450 (N_16450,N_15902,N_15973);
xor U16451 (N_16451,N_15564,N_15501);
xnor U16452 (N_16452,N_15699,N_15509);
nand U16453 (N_16453,N_15580,N_15564);
nand U16454 (N_16454,N_15407,N_15608);
xnor U16455 (N_16455,N_15544,N_15641);
nand U16456 (N_16456,N_15378,N_15465);
and U16457 (N_16457,N_15966,N_15675);
or U16458 (N_16458,N_15597,N_15773);
nor U16459 (N_16459,N_15399,N_15205);
nor U16460 (N_16460,N_15748,N_15540);
nor U16461 (N_16461,N_15405,N_15444);
nor U16462 (N_16462,N_15422,N_15513);
or U16463 (N_16463,N_15420,N_15522);
nand U16464 (N_16464,N_15872,N_15715);
xor U16465 (N_16465,N_15389,N_15916);
xnor U16466 (N_16466,N_15386,N_15375);
and U16467 (N_16467,N_15499,N_15393);
xor U16468 (N_16468,N_15970,N_15643);
nand U16469 (N_16469,N_15386,N_15707);
or U16470 (N_16470,N_15637,N_15222);
and U16471 (N_16471,N_15291,N_15863);
and U16472 (N_16472,N_15550,N_15413);
or U16473 (N_16473,N_15520,N_15543);
nor U16474 (N_16474,N_15695,N_15292);
and U16475 (N_16475,N_15505,N_15619);
and U16476 (N_16476,N_15688,N_15890);
and U16477 (N_16477,N_15982,N_15883);
nor U16478 (N_16478,N_15784,N_15478);
nand U16479 (N_16479,N_15431,N_15826);
nand U16480 (N_16480,N_15837,N_15444);
xor U16481 (N_16481,N_15996,N_15479);
nor U16482 (N_16482,N_15787,N_15941);
or U16483 (N_16483,N_15769,N_15433);
and U16484 (N_16484,N_15873,N_15297);
and U16485 (N_16485,N_15247,N_15607);
nor U16486 (N_16486,N_15449,N_15321);
nor U16487 (N_16487,N_15943,N_15364);
nand U16488 (N_16488,N_15337,N_15701);
xor U16489 (N_16489,N_15921,N_15266);
and U16490 (N_16490,N_15513,N_15216);
or U16491 (N_16491,N_15597,N_15406);
and U16492 (N_16492,N_15341,N_15800);
or U16493 (N_16493,N_15582,N_15661);
nand U16494 (N_16494,N_15936,N_15732);
xnor U16495 (N_16495,N_15600,N_15942);
nand U16496 (N_16496,N_15953,N_15392);
or U16497 (N_16497,N_15514,N_15393);
and U16498 (N_16498,N_15525,N_15688);
or U16499 (N_16499,N_15357,N_15642);
nor U16500 (N_16500,N_15974,N_15865);
xnor U16501 (N_16501,N_15499,N_15879);
and U16502 (N_16502,N_15482,N_15302);
nor U16503 (N_16503,N_15290,N_15221);
or U16504 (N_16504,N_15528,N_15882);
nor U16505 (N_16505,N_15593,N_15281);
xor U16506 (N_16506,N_15682,N_15291);
nand U16507 (N_16507,N_15666,N_15936);
nor U16508 (N_16508,N_15687,N_15723);
xor U16509 (N_16509,N_15684,N_15793);
xnor U16510 (N_16510,N_15479,N_15390);
nand U16511 (N_16511,N_15834,N_15696);
or U16512 (N_16512,N_15852,N_15654);
nor U16513 (N_16513,N_15252,N_15325);
nor U16514 (N_16514,N_15465,N_15898);
and U16515 (N_16515,N_15785,N_15711);
or U16516 (N_16516,N_15706,N_15787);
xor U16517 (N_16517,N_15255,N_15389);
or U16518 (N_16518,N_15452,N_15433);
nor U16519 (N_16519,N_15372,N_15819);
nor U16520 (N_16520,N_15222,N_15963);
nor U16521 (N_16521,N_15683,N_15831);
nor U16522 (N_16522,N_15942,N_15257);
nand U16523 (N_16523,N_15583,N_15965);
nand U16524 (N_16524,N_15612,N_15505);
nand U16525 (N_16525,N_15576,N_15877);
xor U16526 (N_16526,N_15357,N_15339);
nor U16527 (N_16527,N_15304,N_15326);
xor U16528 (N_16528,N_15287,N_15561);
nor U16529 (N_16529,N_15392,N_15879);
or U16530 (N_16530,N_15423,N_15765);
nor U16531 (N_16531,N_15531,N_15732);
and U16532 (N_16532,N_15589,N_15460);
or U16533 (N_16533,N_15330,N_15859);
xor U16534 (N_16534,N_15637,N_15257);
and U16535 (N_16535,N_15411,N_15340);
xnor U16536 (N_16536,N_15529,N_15456);
nand U16537 (N_16537,N_15569,N_15461);
and U16538 (N_16538,N_15342,N_15770);
and U16539 (N_16539,N_15763,N_15657);
or U16540 (N_16540,N_15696,N_15792);
nand U16541 (N_16541,N_15451,N_15968);
and U16542 (N_16542,N_15696,N_15924);
nand U16543 (N_16543,N_15205,N_15802);
nand U16544 (N_16544,N_15352,N_15745);
xnor U16545 (N_16545,N_15848,N_15434);
nand U16546 (N_16546,N_15630,N_15928);
and U16547 (N_16547,N_15306,N_15448);
nand U16548 (N_16548,N_15489,N_15950);
and U16549 (N_16549,N_15850,N_15705);
xor U16550 (N_16550,N_15780,N_15639);
xnor U16551 (N_16551,N_15561,N_15332);
nand U16552 (N_16552,N_15985,N_15427);
nand U16553 (N_16553,N_15474,N_15383);
or U16554 (N_16554,N_15783,N_15345);
or U16555 (N_16555,N_15542,N_15847);
or U16556 (N_16556,N_15561,N_15629);
and U16557 (N_16557,N_15490,N_15678);
nand U16558 (N_16558,N_15917,N_15327);
or U16559 (N_16559,N_15287,N_15867);
nor U16560 (N_16560,N_15537,N_15326);
nor U16561 (N_16561,N_15556,N_15405);
or U16562 (N_16562,N_15817,N_15316);
nor U16563 (N_16563,N_15654,N_15208);
or U16564 (N_16564,N_15530,N_15566);
nor U16565 (N_16565,N_15597,N_15811);
xnor U16566 (N_16566,N_15274,N_15366);
or U16567 (N_16567,N_15848,N_15222);
and U16568 (N_16568,N_15379,N_15787);
or U16569 (N_16569,N_15692,N_15953);
nor U16570 (N_16570,N_15916,N_15972);
and U16571 (N_16571,N_15991,N_15431);
nor U16572 (N_16572,N_15460,N_15279);
and U16573 (N_16573,N_15946,N_15520);
nand U16574 (N_16574,N_15369,N_15861);
nand U16575 (N_16575,N_15848,N_15803);
nand U16576 (N_16576,N_15982,N_15576);
nor U16577 (N_16577,N_15770,N_15703);
or U16578 (N_16578,N_15629,N_15489);
or U16579 (N_16579,N_15206,N_15357);
or U16580 (N_16580,N_15822,N_15725);
or U16581 (N_16581,N_15988,N_15342);
or U16582 (N_16582,N_15396,N_15853);
xnor U16583 (N_16583,N_15391,N_15343);
nand U16584 (N_16584,N_15358,N_15766);
and U16585 (N_16585,N_15334,N_15647);
nand U16586 (N_16586,N_15231,N_15739);
xor U16587 (N_16587,N_15417,N_15742);
nand U16588 (N_16588,N_15274,N_15929);
or U16589 (N_16589,N_15834,N_15688);
or U16590 (N_16590,N_15605,N_15822);
nor U16591 (N_16591,N_15770,N_15340);
xor U16592 (N_16592,N_15344,N_15247);
xnor U16593 (N_16593,N_15888,N_15473);
nor U16594 (N_16594,N_15998,N_15988);
xnor U16595 (N_16595,N_15354,N_15865);
or U16596 (N_16596,N_15344,N_15546);
nor U16597 (N_16597,N_15326,N_15824);
nor U16598 (N_16598,N_15781,N_15478);
or U16599 (N_16599,N_15447,N_15489);
and U16600 (N_16600,N_15358,N_15863);
nand U16601 (N_16601,N_15767,N_15927);
or U16602 (N_16602,N_15227,N_15994);
or U16603 (N_16603,N_15850,N_15528);
nand U16604 (N_16604,N_15486,N_15513);
or U16605 (N_16605,N_15407,N_15690);
nor U16606 (N_16606,N_15281,N_15673);
xor U16607 (N_16607,N_15822,N_15755);
nand U16608 (N_16608,N_15899,N_15211);
or U16609 (N_16609,N_15747,N_15514);
nand U16610 (N_16610,N_15864,N_15944);
nor U16611 (N_16611,N_15939,N_15546);
and U16612 (N_16612,N_15415,N_15476);
xnor U16613 (N_16613,N_15870,N_15517);
nor U16614 (N_16614,N_15434,N_15606);
xnor U16615 (N_16615,N_15303,N_15653);
nand U16616 (N_16616,N_15987,N_15890);
nor U16617 (N_16617,N_15958,N_15420);
and U16618 (N_16618,N_15541,N_15673);
and U16619 (N_16619,N_15757,N_15229);
nand U16620 (N_16620,N_15827,N_15211);
nor U16621 (N_16621,N_15226,N_15782);
and U16622 (N_16622,N_15313,N_15633);
and U16623 (N_16623,N_15870,N_15239);
xor U16624 (N_16624,N_15364,N_15825);
nand U16625 (N_16625,N_15799,N_15253);
xnor U16626 (N_16626,N_15705,N_15650);
xor U16627 (N_16627,N_15612,N_15854);
or U16628 (N_16628,N_15213,N_15601);
or U16629 (N_16629,N_15482,N_15698);
nor U16630 (N_16630,N_15546,N_15693);
nand U16631 (N_16631,N_15366,N_15873);
nor U16632 (N_16632,N_15447,N_15982);
and U16633 (N_16633,N_15895,N_15349);
nand U16634 (N_16634,N_15243,N_15954);
xor U16635 (N_16635,N_15816,N_15214);
nor U16636 (N_16636,N_15584,N_15357);
nand U16637 (N_16637,N_15302,N_15294);
or U16638 (N_16638,N_15850,N_15355);
nor U16639 (N_16639,N_15760,N_15363);
xor U16640 (N_16640,N_15443,N_15955);
or U16641 (N_16641,N_15979,N_15892);
nand U16642 (N_16642,N_15600,N_15926);
or U16643 (N_16643,N_15656,N_15809);
nor U16644 (N_16644,N_15574,N_15728);
or U16645 (N_16645,N_15296,N_15998);
nor U16646 (N_16646,N_15251,N_15239);
xor U16647 (N_16647,N_15591,N_15557);
or U16648 (N_16648,N_15661,N_15550);
xor U16649 (N_16649,N_15761,N_15548);
or U16650 (N_16650,N_15726,N_15205);
xor U16651 (N_16651,N_15894,N_15878);
nor U16652 (N_16652,N_15786,N_15726);
and U16653 (N_16653,N_15352,N_15313);
xnor U16654 (N_16654,N_15254,N_15689);
or U16655 (N_16655,N_15731,N_15616);
nor U16656 (N_16656,N_15863,N_15636);
nor U16657 (N_16657,N_15372,N_15961);
nand U16658 (N_16658,N_15238,N_15266);
and U16659 (N_16659,N_15725,N_15295);
or U16660 (N_16660,N_15573,N_15739);
or U16661 (N_16661,N_15834,N_15988);
nor U16662 (N_16662,N_15742,N_15998);
nor U16663 (N_16663,N_15466,N_15684);
and U16664 (N_16664,N_15604,N_15385);
nand U16665 (N_16665,N_15798,N_15814);
or U16666 (N_16666,N_15462,N_15852);
nor U16667 (N_16667,N_15237,N_15387);
nand U16668 (N_16668,N_15736,N_15814);
or U16669 (N_16669,N_15764,N_15439);
xnor U16670 (N_16670,N_15736,N_15267);
nor U16671 (N_16671,N_15759,N_15846);
and U16672 (N_16672,N_15316,N_15706);
and U16673 (N_16673,N_15406,N_15824);
nor U16674 (N_16674,N_15445,N_15601);
or U16675 (N_16675,N_15717,N_15973);
and U16676 (N_16676,N_15717,N_15592);
and U16677 (N_16677,N_15723,N_15632);
nor U16678 (N_16678,N_15959,N_15327);
or U16679 (N_16679,N_15502,N_15651);
xor U16680 (N_16680,N_15566,N_15279);
or U16681 (N_16681,N_15950,N_15892);
or U16682 (N_16682,N_15691,N_15612);
xor U16683 (N_16683,N_15813,N_15742);
nand U16684 (N_16684,N_15206,N_15374);
nand U16685 (N_16685,N_15451,N_15252);
nor U16686 (N_16686,N_15412,N_15547);
and U16687 (N_16687,N_15566,N_15652);
and U16688 (N_16688,N_15622,N_15632);
xor U16689 (N_16689,N_15467,N_15911);
xnor U16690 (N_16690,N_15980,N_15380);
or U16691 (N_16691,N_15731,N_15693);
or U16692 (N_16692,N_15613,N_15495);
and U16693 (N_16693,N_15588,N_15246);
and U16694 (N_16694,N_15891,N_15354);
nor U16695 (N_16695,N_15250,N_15750);
and U16696 (N_16696,N_15993,N_15945);
xnor U16697 (N_16697,N_15968,N_15692);
and U16698 (N_16698,N_15397,N_15891);
xor U16699 (N_16699,N_15856,N_15430);
xnor U16700 (N_16700,N_15989,N_15302);
or U16701 (N_16701,N_15525,N_15516);
and U16702 (N_16702,N_15738,N_15986);
and U16703 (N_16703,N_15459,N_15543);
or U16704 (N_16704,N_15913,N_15271);
or U16705 (N_16705,N_15979,N_15238);
nand U16706 (N_16706,N_15397,N_15303);
and U16707 (N_16707,N_15945,N_15955);
nor U16708 (N_16708,N_15320,N_15727);
nand U16709 (N_16709,N_15782,N_15538);
nand U16710 (N_16710,N_15361,N_15615);
or U16711 (N_16711,N_15540,N_15430);
xnor U16712 (N_16712,N_15556,N_15575);
or U16713 (N_16713,N_15463,N_15628);
nor U16714 (N_16714,N_15863,N_15217);
nand U16715 (N_16715,N_15896,N_15699);
nand U16716 (N_16716,N_15639,N_15837);
and U16717 (N_16717,N_15532,N_15836);
nor U16718 (N_16718,N_15339,N_15927);
or U16719 (N_16719,N_15267,N_15974);
nand U16720 (N_16720,N_15638,N_15512);
and U16721 (N_16721,N_15409,N_15218);
xor U16722 (N_16722,N_15569,N_15874);
and U16723 (N_16723,N_15291,N_15366);
nor U16724 (N_16724,N_15224,N_15678);
and U16725 (N_16725,N_15500,N_15741);
nor U16726 (N_16726,N_15205,N_15291);
or U16727 (N_16727,N_15898,N_15939);
or U16728 (N_16728,N_15220,N_15942);
nand U16729 (N_16729,N_15697,N_15834);
nand U16730 (N_16730,N_15837,N_15961);
nand U16731 (N_16731,N_15554,N_15703);
nor U16732 (N_16732,N_15272,N_15599);
xor U16733 (N_16733,N_15452,N_15896);
and U16734 (N_16734,N_15808,N_15329);
nor U16735 (N_16735,N_15961,N_15216);
nand U16736 (N_16736,N_15990,N_15513);
and U16737 (N_16737,N_15884,N_15960);
xnor U16738 (N_16738,N_15661,N_15861);
nand U16739 (N_16739,N_15694,N_15941);
nand U16740 (N_16740,N_15586,N_15982);
xor U16741 (N_16741,N_15531,N_15637);
nor U16742 (N_16742,N_15418,N_15815);
nor U16743 (N_16743,N_15333,N_15788);
nor U16744 (N_16744,N_15391,N_15449);
xor U16745 (N_16745,N_15503,N_15509);
or U16746 (N_16746,N_15724,N_15848);
xor U16747 (N_16747,N_15919,N_15677);
nand U16748 (N_16748,N_15535,N_15919);
and U16749 (N_16749,N_15609,N_15468);
xnor U16750 (N_16750,N_15877,N_15395);
nor U16751 (N_16751,N_15599,N_15838);
nor U16752 (N_16752,N_15469,N_15994);
nand U16753 (N_16753,N_15232,N_15252);
and U16754 (N_16754,N_15889,N_15243);
and U16755 (N_16755,N_15620,N_15539);
nand U16756 (N_16756,N_15569,N_15212);
or U16757 (N_16757,N_15359,N_15919);
and U16758 (N_16758,N_15789,N_15845);
xnor U16759 (N_16759,N_15926,N_15860);
nor U16760 (N_16760,N_15533,N_15515);
xnor U16761 (N_16761,N_15579,N_15986);
or U16762 (N_16762,N_15200,N_15468);
nor U16763 (N_16763,N_15703,N_15652);
nor U16764 (N_16764,N_15630,N_15442);
nand U16765 (N_16765,N_15822,N_15718);
nand U16766 (N_16766,N_15225,N_15721);
nand U16767 (N_16767,N_15618,N_15701);
nor U16768 (N_16768,N_15689,N_15877);
nand U16769 (N_16769,N_15860,N_15566);
or U16770 (N_16770,N_15801,N_15941);
nand U16771 (N_16771,N_15328,N_15214);
or U16772 (N_16772,N_15232,N_15875);
and U16773 (N_16773,N_15625,N_15508);
xnor U16774 (N_16774,N_15300,N_15970);
and U16775 (N_16775,N_15846,N_15991);
nand U16776 (N_16776,N_15656,N_15259);
xor U16777 (N_16777,N_15620,N_15597);
and U16778 (N_16778,N_15452,N_15836);
and U16779 (N_16779,N_15670,N_15538);
nand U16780 (N_16780,N_15224,N_15933);
or U16781 (N_16781,N_15380,N_15817);
nor U16782 (N_16782,N_15777,N_15609);
xor U16783 (N_16783,N_15967,N_15832);
xnor U16784 (N_16784,N_15931,N_15408);
nor U16785 (N_16785,N_15949,N_15417);
xnor U16786 (N_16786,N_15638,N_15771);
nor U16787 (N_16787,N_15725,N_15402);
xnor U16788 (N_16788,N_15671,N_15603);
nor U16789 (N_16789,N_15786,N_15798);
xor U16790 (N_16790,N_15337,N_15308);
xnor U16791 (N_16791,N_15972,N_15914);
xor U16792 (N_16792,N_15830,N_15852);
and U16793 (N_16793,N_15437,N_15954);
nand U16794 (N_16794,N_15302,N_15792);
nand U16795 (N_16795,N_15962,N_15904);
nand U16796 (N_16796,N_15278,N_15495);
and U16797 (N_16797,N_15798,N_15436);
or U16798 (N_16798,N_15728,N_15302);
nand U16799 (N_16799,N_15252,N_15962);
or U16800 (N_16800,N_16538,N_16069);
and U16801 (N_16801,N_16558,N_16425);
nand U16802 (N_16802,N_16470,N_16087);
and U16803 (N_16803,N_16413,N_16042);
and U16804 (N_16804,N_16549,N_16027);
nor U16805 (N_16805,N_16725,N_16784);
xor U16806 (N_16806,N_16169,N_16336);
or U16807 (N_16807,N_16318,N_16093);
and U16808 (N_16808,N_16401,N_16744);
xnor U16809 (N_16809,N_16384,N_16180);
nor U16810 (N_16810,N_16463,N_16755);
nor U16811 (N_16811,N_16740,N_16065);
xor U16812 (N_16812,N_16310,N_16721);
xor U16813 (N_16813,N_16489,N_16788);
or U16814 (N_16814,N_16698,N_16659);
nand U16815 (N_16815,N_16591,N_16535);
or U16816 (N_16816,N_16286,N_16412);
xor U16817 (N_16817,N_16016,N_16247);
nor U16818 (N_16818,N_16520,N_16737);
xnor U16819 (N_16819,N_16000,N_16732);
and U16820 (N_16820,N_16164,N_16051);
xnor U16821 (N_16821,N_16578,N_16296);
or U16822 (N_16822,N_16052,N_16224);
nand U16823 (N_16823,N_16213,N_16263);
or U16824 (N_16824,N_16143,N_16259);
nand U16825 (N_16825,N_16640,N_16102);
nor U16826 (N_16826,N_16273,N_16605);
nand U16827 (N_16827,N_16636,N_16472);
nor U16828 (N_16828,N_16211,N_16284);
or U16829 (N_16829,N_16025,N_16282);
xor U16830 (N_16830,N_16613,N_16394);
nor U16831 (N_16831,N_16332,N_16566);
or U16832 (N_16832,N_16618,N_16530);
xnor U16833 (N_16833,N_16473,N_16389);
and U16834 (N_16834,N_16419,N_16005);
and U16835 (N_16835,N_16722,N_16677);
nor U16836 (N_16836,N_16145,N_16307);
nor U16837 (N_16837,N_16778,N_16094);
and U16838 (N_16838,N_16351,N_16717);
or U16839 (N_16839,N_16794,N_16527);
nand U16840 (N_16840,N_16081,N_16250);
and U16841 (N_16841,N_16407,N_16643);
and U16842 (N_16842,N_16674,N_16562);
nand U16843 (N_16843,N_16540,N_16482);
or U16844 (N_16844,N_16376,N_16255);
or U16845 (N_16845,N_16751,N_16279);
nor U16846 (N_16846,N_16583,N_16156);
nand U16847 (N_16847,N_16555,N_16560);
and U16848 (N_16848,N_16458,N_16593);
nand U16849 (N_16849,N_16268,N_16360);
xor U16850 (N_16850,N_16035,N_16350);
xnor U16851 (N_16851,N_16132,N_16219);
or U16852 (N_16852,N_16104,N_16377);
xnor U16853 (N_16853,N_16793,N_16092);
and U16854 (N_16854,N_16074,N_16096);
xnor U16855 (N_16855,N_16446,N_16697);
or U16856 (N_16856,N_16604,N_16392);
and U16857 (N_16857,N_16232,N_16113);
nand U16858 (N_16858,N_16078,N_16528);
nand U16859 (N_16859,N_16603,N_16371);
xor U16860 (N_16860,N_16506,N_16017);
and U16861 (N_16861,N_16445,N_16203);
nand U16862 (N_16862,N_16423,N_16524);
nand U16863 (N_16863,N_16064,N_16786);
nor U16864 (N_16864,N_16466,N_16529);
nor U16865 (N_16865,N_16222,N_16465);
xor U16866 (N_16866,N_16624,N_16460);
and U16867 (N_16867,N_16253,N_16137);
and U16868 (N_16868,N_16041,N_16193);
and U16869 (N_16869,N_16038,N_16040);
or U16870 (N_16870,N_16690,N_16191);
or U16871 (N_16871,N_16430,N_16136);
or U16872 (N_16872,N_16714,N_16215);
nand U16873 (N_16873,N_16621,N_16707);
and U16874 (N_16874,N_16395,N_16452);
and U16875 (N_16875,N_16308,N_16571);
and U16876 (N_16876,N_16641,N_16183);
or U16877 (N_16877,N_16344,N_16607);
and U16878 (N_16878,N_16186,N_16107);
nor U16879 (N_16879,N_16544,N_16321);
nand U16880 (N_16880,N_16170,N_16030);
nor U16881 (N_16881,N_16587,N_16218);
nand U16882 (N_16882,N_16182,N_16105);
xnor U16883 (N_16883,N_16671,N_16650);
nor U16884 (N_16884,N_16763,N_16692);
nand U16885 (N_16885,N_16611,N_16316);
nand U16886 (N_16886,N_16476,N_16658);
xnor U16887 (N_16887,N_16333,N_16383);
or U16888 (N_16888,N_16303,N_16559);
and U16889 (N_16889,N_16483,N_16635);
nor U16890 (N_16890,N_16628,N_16475);
xor U16891 (N_16891,N_16339,N_16599);
nand U16892 (N_16892,N_16135,N_16187);
nor U16893 (N_16893,N_16154,N_16716);
nand U16894 (N_16894,N_16748,N_16724);
nand U16895 (N_16895,N_16759,N_16317);
and U16896 (N_16896,N_16311,N_16204);
nand U16897 (N_16897,N_16127,N_16620);
xnor U16898 (N_16898,N_16765,N_16297);
xor U16899 (N_16899,N_16500,N_16718);
nand U16900 (N_16900,N_16746,N_16711);
nand U16901 (N_16901,N_16457,N_16067);
nand U16902 (N_16902,N_16058,N_16543);
or U16903 (N_16903,N_16503,N_16736);
nor U16904 (N_16904,N_16433,N_16431);
and U16905 (N_16905,N_16043,N_16518);
or U16906 (N_16906,N_16071,N_16362);
xnor U16907 (N_16907,N_16046,N_16086);
and U16908 (N_16908,N_16235,N_16745);
nor U16909 (N_16909,N_16053,N_16777);
nand U16910 (N_16910,N_16150,N_16168);
xnor U16911 (N_16911,N_16660,N_16437);
xor U16912 (N_16912,N_16236,N_16299);
nand U16913 (N_16913,N_16396,N_16008);
xor U16914 (N_16914,N_16184,N_16032);
and U16915 (N_16915,N_16361,N_16664);
xnor U16916 (N_16916,N_16584,N_16764);
or U16917 (N_16917,N_16241,N_16009);
nand U16918 (N_16918,N_16020,N_16497);
and U16919 (N_16919,N_16670,N_16258);
xor U16920 (N_16920,N_16338,N_16428);
xnor U16921 (N_16921,N_16743,N_16240);
or U16922 (N_16922,N_16221,N_16228);
nor U16923 (N_16923,N_16254,N_16561);
and U16924 (N_16924,N_16403,N_16491);
nand U16925 (N_16925,N_16757,N_16516);
and U16926 (N_16926,N_16455,N_16696);
nand U16927 (N_16927,N_16539,N_16582);
xor U16928 (N_16928,N_16229,N_16651);
xnor U16929 (N_16929,N_16509,N_16122);
and U16930 (N_16930,N_16758,N_16410);
and U16931 (N_16931,N_16701,N_16178);
nand U16932 (N_16932,N_16368,N_16440);
and U16933 (N_16933,N_16700,N_16715);
nor U16934 (N_16934,N_16420,N_16220);
or U16935 (N_16935,N_16045,N_16075);
or U16936 (N_16936,N_16678,N_16631);
nor U16937 (N_16937,N_16792,N_16277);
xor U16938 (N_16938,N_16451,N_16270);
or U16939 (N_16939,N_16271,N_16144);
nand U16940 (N_16940,N_16496,N_16061);
and U16941 (N_16941,N_16598,N_16205);
nand U16942 (N_16942,N_16140,N_16672);
nand U16943 (N_16943,N_16161,N_16352);
nand U16944 (N_16944,N_16121,N_16626);
xor U16945 (N_16945,N_16153,N_16315);
or U16946 (N_16946,N_16068,N_16073);
and U16947 (N_16947,N_16126,N_16486);
or U16948 (N_16948,N_16272,N_16705);
nor U16949 (N_16949,N_16397,N_16444);
or U16950 (N_16950,N_16799,N_16123);
nor U16951 (N_16951,N_16275,N_16266);
and U16952 (N_16952,N_16098,N_16039);
xor U16953 (N_16953,N_16329,N_16726);
and U16954 (N_16954,N_16015,N_16487);
nor U16955 (N_16955,N_16312,N_16798);
or U16956 (N_16956,N_16111,N_16505);
or U16957 (N_16957,N_16526,N_16246);
nand U16958 (N_16958,N_16177,N_16124);
or U16959 (N_16959,N_16190,N_16602);
xor U16960 (N_16960,N_16265,N_16285);
xor U16961 (N_16961,N_16165,N_16449);
or U16962 (N_16962,N_16534,N_16762);
nand U16963 (N_16963,N_16325,N_16790);
and U16964 (N_16964,N_16432,N_16084);
and U16965 (N_16965,N_16484,N_16090);
xnor U16966 (N_16966,N_16185,N_16706);
and U16967 (N_16967,N_16490,N_16703);
and U16968 (N_16968,N_16531,N_16031);
nor U16969 (N_16969,N_16334,N_16378);
nor U16970 (N_16970,N_16057,N_16573);
and U16971 (N_16971,N_16062,N_16117);
and U16972 (N_16972,N_16588,N_16242);
and U16973 (N_16973,N_16536,N_16676);
xnor U16974 (N_16974,N_16456,N_16063);
and U16975 (N_16975,N_16160,N_16011);
nand U16976 (N_16976,N_16264,N_16429);
nand U16977 (N_16977,N_16210,N_16776);
xnor U16978 (N_16978,N_16357,N_16638);
and U16979 (N_16979,N_16498,N_16112);
or U16980 (N_16980,N_16194,N_16447);
and U16981 (N_16981,N_16044,N_16525);
nand U16982 (N_16982,N_16049,N_16385);
nand U16983 (N_16983,N_16454,N_16080);
nand U16984 (N_16984,N_16502,N_16149);
and U16985 (N_16985,N_16055,N_16633);
and U16986 (N_16986,N_16648,N_16304);
xnor U16987 (N_16987,N_16761,N_16320);
nand U16988 (N_16988,N_16655,N_16402);
and U16989 (N_16989,N_16129,N_16630);
nand U16990 (N_16990,N_16131,N_16018);
and U16991 (N_16991,N_16741,N_16499);
and U16992 (N_16992,N_16517,N_16089);
nor U16993 (N_16993,N_16479,N_16379);
and U16994 (N_16994,N_16467,N_16085);
or U16995 (N_16995,N_16106,N_16637);
nand U16996 (N_16996,N_16668,N_16314);
and U16997 (N_16997,N_16237,N_16217);
and U16998 (N_16998,N_16101,N_16667);
or U16999 (N_16999,N_16393,N_16550);
or U17000 (N_17000,N_16251,N_16688);
xor U17001 (N_17001,N_16290,N_16354);
xnor U17002 (N_17002,N_16034,N_16152);
and U17003 (N_17003,N_16363,N_16504);
or U17004 (N_17004,N_16581,N_16047);
and U17005 (N_17005,N_16114,N_16330);
and U17006 (N_17006,N_16797,N_16547);
nor U17007 (N_17007,N_16708,N_16557);
and U17008 (N_17008,N_16551,N_16056);
xnor U17009 (N_17009,N_16782,N_16374);
nor U17010 (N_17010,N_16596,N_16024);
and U17011 (N_17011,N_16292,N_16480);
xnor U17012 (N_17012,N_16709,N_16175);
nor U17013 (N_17013,N_16141,N_16305);
nand U17014 (N_17014,N_16645,N_16702);
nand U17015 (N_17015,N_16654,N_16408);
nand U17016 (N_17016,N_16586,N_16795);
nand U17017 (N_17017,N_16077,N_16597);
and U17018 (N_17018,N_16138,N_16048);
or U17019 (N_17019,N_16750,N_16225);
nand U17020 (N_17020,N_16033,N_16441);
nand U17021 (N_17021,N_16686,N_16280);
and U17022 (N_17022,N_16171,N_16002);
xor U17023 (N_17023,N_16181,N_16614);
nand U17024 (N_17024,N_16772,N_16589);
nor U17025 (N_17025,N_16208,N_16391);
and U17026 (N_17026,N_16448,N_16416);
nand U17027 (N_17027,N_16230,N_16546);
and U17028 (N_17028,N_16753,N_16545);
or U17029 (N_17029,N_16627,N_16601);
and U17030 (N_17030,N_16227,N_16507);
and U17031 (N_17031,N_16328,N_16026);
nor U17032 (N_17032,N_16249,N_16747);
or U17033 (N_17033,N_16533,N_16684);
or U17034 (N_17034,N_16612,N_16427);
nand U17035 (N_17035,N_16639,N_16116);
xnor U17036 (N_17036,N_16007,N_16644);
and U17037 (N_17037,N_16629,N_16577);
nor U17038 (N_17038,N_16151,N_16542);
or U17039 (N_17039,N_16459,N_16223);
xnor U17040 (N_17040,N_16775,N_16261);
nor U17041 (N_17041,N_16382,N_16343);
xnor U17042 (N_17042,N_16327,N_16120);
nor U17043 (N_17043,N_16590,N_16340);
nand U17044 (N_17044,N_16226,N_16142);
nor U17045 (N_17045,N_16563,N_16216);
and U17046 (N_17046,N_16592,N_16370);
nand U17047 (N_17047,N_16019,N_16733);
xor U17048 (N_17048,N_16685,N_16791);
nor U17049 (N_17049,N_16243,N_16097);
or U17050 (N_17050,N_16386,N_16512);
nor U17051 (N_17051,N_16373,N_16787);
nand U17052 (N_17052,N_16687,N_16346);
nor U17053 (N_17053,N_16521,N_16426);
or U17054 (N_17054,N_16569,N_16615);
and U17055 (N_17055,N_16146,N_16580);
nor U17056 (N_17056,N_16734,N_16439);
nor U17057 (N_17057,N_16207,N_16341);
nor U17058 (N_17058,N_16399,N_16585);
nor U17059 (N_17059,N_16720,N_16634);
xor U17060 (N_17060,N_16118,N_16257);
nor U17061 (N_17061,N_16231,N_16796);
nor U17062 (N_17062,N_16404,N_16189);
and U17063 (N_17063,N_16657,N_16435);
nor U17064 (N_17064,N_16622,N_16679);
and U17065 (N_17065,N_16625,N_16481);
nand U17066 (N_17066,N_16301,N_16158);
xnor U17067 (N_17067,N_16347,N_16478);
or U17068 (N_17068,N_16288,N_16760);
or U17069 (N_17069,N_16768,N_16477);
xnor U17070 (N_17070,N_16001,N_16174);
nor U17071 (N_17071,N_16442,N_16195);
xnor U17072 (N_17072,N_16730,N_16406);
or U17073 (N_17073,N_16157,N_16289);
or U17074 (N_17074,N_16004,N_16037);
and U17075 (N_17075,N_16206,N_16148);
and U17076 (N_17076,N_16511,N_16570);
or U17077 (N_17077,N_16617,N_16022);
xor U17078 (N_17078,N_16050,N_16453);
or U17079 (N_17079,N_16028,N_16147);
and U17080 (N_17080,N_16345,N_16749);
and U17081 (N_17081,N_16532,N_16364);
xnor U17082 (N_17082,N_16461,N_16119);
or U17083 (N_17083,N_16647,N_16695);
nor U17084 (N_17084,N_16681,N_16079);
and U17085 (N_17085,N_16783,N_16450);
and U17086 (N_17086,N_16474,N_16267);
nor U17087 (N_17087,N_16693,N_16492);
xnor U17088 (N_17088,N_16494,N_16493);
nor U17089 (N_17089,N_16245,N_16369);
nor U17090 (N_17090,N_16179,N_16198);
or U17091 (N_17091,N_16673,N_16262);
nand U17092 (N_17092,N_16335,N_16300);
nand U17093 (N_17093,N_16731,N_16537);
nor U17094 (N_17094,N_16485,N_16212);
xnor U17095 (N_17095,N_16554,N_16159);
and U17096 (N_17096,N_16661,N_16059);
and U17097 (N_17097,N_16682,N_16713);
nor U17098 (N_17098,N_16365,N_16779);
or U17099 (N_17099,N_16309,N_16752);
nor U17100 (N_17100,N_16699,N_16276);
and U17101 (N_17101,N_16469,N_16269);
nand U17102 (N_17102,N_16436,N_16110);
nor U17103 (N_17103,N_16214,N_16070);
nor U17104 (N_17104,N_16771,N_16774);
and U17105 (N_17105,N_16390,N_16510);
or U17106 (N_17106,N_16013,N_16066);
and U17107 (N_17107,N_16723,N_16322);
xnor U17108 (N_17108,N_16523,N_16632);
nand U17109 (N_17109,N_16417,N_16176);
nor U17110 (N_17110,N_16130,N_16541);
or U17111 (N_17111,N_16095,N_16209);
and U17112 (N_17112,N_16415,N_16471);
nor U17113 (N_17113,N_16381,N_16319);
nor U17114 (N_17114,N_16568,N_16349);
nor U17115 (N_17115,N_16501,N_16600);
and U17116 (N_17116,N_16785,N_16576);
or U17117 (N_17117,N_16293,N_16514);
xor U17118 (N_17118,N_16358,N_16754);
xnor U17119 (N_17119,N_16766,N_16552);
nand U17120 (N_17120,N_16133,N_16342);
or U17121 (N_17121,N_16574,N_16036);
and U17122 (N_17122,N_16619,N_16298);
nor U17123 (N_17123,N_16088,N_16662);
nor U17124 (N_17124,N_16252,N_16712);
xnor U17125 (N_17125,N_16029,N_16199);
and U17126 (N_17126,N_16443,N_16421);
and U17127 (N_17127,N_16515,N_16099);
and U17128 (N_17128,N_16767,N_16572);
xnor U17129 (N_17129,N_16739,N_16014);
and U17130 (N_17130,N_16278,N_16283);
and U17131 (N_17131,N_16414,N_16665);
and U17132 (N_17132,N_16579,N_16076);
or U17133 (N_17133,N_16166,N_16353);
nor U17134 (N_17134,N_16595,N_16462);
and U17135 (N_17135,N_16302,N_16438);
xor U17136 (N_17136,N_16653,N_16519);
nand U17137 (N_17137,N_16163,N_16359);
and U17138 (N_17138,N_16082,N_16109);
nand U17139 (N_17139,N_16367,N_16756);
xor U17140 (N_17140,N_16125,N_16719);
or U17141 (N_17141,N_16610,N_16201);
and U17142 (N_17142,N_16669,N_16380);
nand U17143 (N_17143,N_16256,N_16728);
nand U17144 (N_17144,N_16773,N_16162);
or U17145 (N_17145,N_16326,N_16239);
xnor U17146 (N_17146,N_16006,N_16704);
and U17147 (N_17147,N_16012,N_16060);
nand U17148 (N_17148,N_16128,N_16200);
nand U17149 (N_17149,N_16233,N_16424);
or U17150 (N_17150,N_16291,N_16274);
nand U17151 (N_17151,N_16003,N_16770);
and U17152 (N_17152,N_16649,N_16616);
and U17153 (N_17153,N_16398,N_16642);
nor U17154 (N_17154,N_16594,N_16234);
nor U17155 (N_17155,N_16323,N_16400);
nor U17156 (N_17156,N_16083,N_16623);
nand U17157 (N_17157,N_16238,N_16115);
nor U17158 (N_17158,N_16295,N_16355);
nor U17159 (N_17159,N_16689,N_16683);
nand U17160 (N_17160,N_16564,N_16780);
xor U17161 (N_17161,N_16680,N_16556);
nand U17162 (N_17162,N_16663,N_16260);
nor U17163 (N_17163,N_16735,N_16495);
nand U17164 (N_17164,N_16248,N_16324);
and U17165 (N_17165,N_16666,N_16072);
nor U17166 (N_17166,N_16348,N_16513);
and U17167 (N_17167,N_16139,N_16388);
nand U17168 (N_17168,N_16054,N_16694);
xnor U17169 (N_17169,N_16656,N_16738);
nor U17170 (N_17170,N_16434,N_16108);
nor U17171 (N_17171,N_16608,N_16567);
and U17172 (N_17172,N_16646,N_16313);
xnor U17173 (N_17173,N_16375,N_16418);
or U17174 (N_17174,N_16091,N_16411);
or U17175 (N_17175,N_16100,N_16010);
xor U17176 (N_17176,N_16196,N_16675);
or U17177 (N_17177,N_16103,N_16021);
and U17178 (N_17178,N_16727,N_16488);
or U17179 (N_17179,N_16553,N_16366);
xor U17180 (N_17180,N_16197,N_16729);
or U17181 (N_17181,N_16387,N_16464);
xor U17182 (N_17182,N_16548,N_16287);
xnor U17183 (N_17183,N_16188,N_16769);
and U17184 (N_17184,N_16522,N_16468);
and U17185 (N_17185,N_16710,N_16172);
xnor U17186 (N_17186,N_16565,N_16155);
and U17187 (N_17187,N_16609,N_16023);
nor U17188 (N_17188,N_16167,N_16331);
nand U17189 (N_17189,N_16173,N_16508);
or U17190 (N_17190,N_16244,N_16372);
and U17191 (N_17191,N_16337,N_16281);
nor U17192 (N_17192,N_16192,N_16691);
or U17193 (N_17193,N_16606,N_16575);
or U17194 (N_17194,N_16789,N_16422);
and U17195 (N_17195,N_16356,N_16405);
nand U17196 (N_17196,N_16202,N_16652);
nand U17197 (N_17197,N_16294,N_16306);
nand U17198 (N_17198,N_16409,N_16134);
and U17199 (N_17199,N_16742,N_16781);
and U17200 (N_17200,N_16380,N_16224);
nand U17201 (N_17201,N_16617,N_16202);
xnor U17202 (N_17202,N_16358,N_16781);
or U17203 (N_17203,N_16343,N_16263);
nor U17204 (N_17204,N_16014,N_16047);
xnor U17205 (N_17205,N_16124,N_16762);
xor U17206 (N_17206,N_16346,N_16317);
xor U17207 (N_17207,N_16185,N_16760);
nand U17208 (N_17208,N_16367,N_16671);
nor U17209 (N_17209,N_16261,N_16759);
or U17210 (N_17210,N_16420,N_16141);
nand U17211 (N_17211,N_16794,N_16208);
and U17212 (N_17212,N_16452,N_16421);
nand U17213 (N_17213,N_16313,N_16592);
and U17214 (N_17214,N_16289,N_16445);
and U17215 (N_17215,N_16544,N_16058);
nand U17216 (N_17216,N_16354,N_16704);
nor U17217 (N_17217,N_16712,N_16340);
xor U17218 (N_17218,N_16328,N_16534);
and U17219 (N_17219,N_16076,N_16058);
or U17220 (N_17220,N_16452,N_16276);
and U17221 (N_17221,N_16732,N_16469);
nor U17222 (N_17222,N_16469,N_16473);
and U17223 (N_17223,N_16283,N_16277);
or U17224 (N_17224,N_16794,N_16674);
nor U17225 (N_17225,N_16723,N_16109);
nand U17226 (N_17226,N_16319,N_16762);
or U17227 (N_17227,N_16268,N_16585);
xor U17228 (N_17228,N_16042,N_16075);
nor U17229 (N_17229,N_16147,N_16788);
and U17230 (N_17230,N_16116,N_16484);
xnor U17231 (N_17231,N_16366,N_16536);
nand U17232 (N_17232,N_16421,N_16395);
and U17233 (N_17233,N_16149,N_16053);
nand U17234 (N_17234,N_16410,N_16128);
nand U17235 (N_17235,N_16263,N_16404);
or U17236 (N_17236,N_16178,N_16564);
nor U17237 (N_17237,N_16493,N_16687);
xor U17238 (N_17238,N_16131,N_16177);
nor U17239 (N_17239,N_16712,N_16517);
or U17240 (N_17240,N_16563,N_16084);
nor U17241 (N_17241,N_16209,N_16601);
nand U17242 (N_17242,N_16285,N_16647);
xnor U17243 (N_17243,N_16176,N_16231);
or U17244 (N_17244,N_16592,N_16033);
xnor U17245 (N_17245,N_16710,N_16793);
or U17246 (N_17246,N_16742,N_16266);
xor U17247 (N_17247,N_16705,N_16234);
nand U17248 (N_17248,N_16556,N_16179);
nand U17249 (N_17249,N_16703,N_16177);
nand U17250 (N_17250,N_16459,N_16136);
and U17251 (N_17251,N_16651,N_16406);
or U17252 (N_17252,N_16654,N_16726);
nor U17253 (N_17253,N_16055,N_16578);
and U17254 (N_17254,N_16497,N_16545);
and U17255 (N_17255,N_16453,N_16008);
or U17256 (N_17256,N_16520,N_16767);
nand U17257 (N_17257,N_16622,N_16061);
and U17258 (N_17258,N_16718,N_16221);
and U17259 (N_17259,N_16401,N_16011);
xnor U17260 (N_17260,N_16185,N_16402);
and U17261 (N_17261,N_16335,N_16725);
and U17262 (N_17262,N_16535,N_16220);
and U17263 (N_17263,N_16318,N_16582);
xor U17264 (N_17264,N_16370,N_16700);
or U17265 (N_17265,N_16488,N_16299);
and U17266 (N_17266,N_16639,N_16270);
nor U17267 (N_17267,N_16482,N_16078);
nor U17268 (N_17268,N_16255,N_16547);
nor U17269 (N_17269,N_16137,N_16256);
nor U17270 (N_17270,N_16265,N_16092);
xnor U17271 (N_17271,N_16221,N_16750);
xor U17272 (N_17272,N_16226,N_16139);
nand U17273 (N_17273,N_16774,N_16176);
or U17274 (N_17274,N_16711,N_16362);
xnor U17275 (N_17275,N_16733,N_16532);
nand U17276 (N_17276,N_16102,N_16383);
and U17277 (N_17277,N_16235,N_16345);
nor U17278 (N_17278,N_16656,N_16323);
nand U17279 (N_17279,N_16419,N_16509);
xor U17280 (N_17280,N_16097,N_16232);
xor U17281 (N_17281,N_16543,N_16297);
nand U17282 (N_17282,N_16797,N_16158);
and U17283 (N_17283,N_16313,N_16206);
or U17284 (N_17284,N_16024,N_16398);
and U17285 (N_17285,N_16466,N_16640);
xor U17286 (N_17286,N_16520,N_16269);
xnor U17287 (N_17287,N_16025,N_16261);
nor U17288 (N_17288,N_16791,N_16736);
or U17289 (N_17289,N_16754,N_16770);
nor U17290 (N_17290,N_16668,N_16187);
xnor U17291 (N_17291,N_16121,N_16726);
nand U17292 (N_17292,N_16390,N_16525);
or U17293 (N_17293,N_16143,N_16486);
nor U17294 (N_17294,N_16543,N_16308);
or U17295 (N_17295,N_16735,N_16129);
or U17296 (N_17296,N_16387,N_16587);
or U17297 (N_17297,N_16644,N_16175);
xor U17298 (N_17298,N_16674,N_16672);
nor U17299 (N_17299,N_16593,N_16645);
and U17300 (N_17300,N_16557,N_16786);
xor U17301 (N_17301,N_16367,N_16250);
and U17302 (N_17302,N_16301,N_16523);
nand U17303 (N_17303,N_16386,N_16509);
and U17304 (N_17304,N_16589,N_16155);
and U17305 (N_17305,N_16120,N_16226);
nor U17306 (N_17306,N_16339,N_16153);
nand U17307 (N_17307,N_16199,N_16556);
nor U17308 (N_17308,N_16114,N_16179);
nor U17309 (N_17309,N_16706,N_16633);
and U17310 (N_17310,N_16645,N_16626);
or U17311 (N_17311,N_16533,N_16025);
and U17312 (N_17312,N_16604,N_16365);
or U17313 (N_17313,N_16692,N_16601);
or U17314 (N_17314,N_16358,N_16027);
nand U17315 (N_17315,N_16075,N_16547);
and U17316 (N_17316,N_16515,N_16266);
xnor U17317 (N_17317,N_16792,N_16227);
nor U17318 (N_17318,N_16565,N_16626);
and U17319 (N_17319,N_16617,N_16413);
nor U17320 (N_17320,N_16476,N_16441);
nand U17321 (N_17321,N_16205,N_16717);
and U17322 (N_17322,N_16670,N_16607);
and U17323 (N_17323,N_16053,N_16671);
nor U17324 (N_17324,N_16335,N_16013);
nor U17325 (N_17325,N_16025,N_16418);
nand U17326 (N_17326,N_16750,N_16367);
and U17327 (N_17327,N_16326,N_16375);
or U17328 (N_17328,N_16378,N_16592);
and U17329 (N_17329,N_16181,N_16592);
nand U17330 (N_17330,N_16293,N_16212);
or U17331 (N_17331,N_16692,N_16122);
and U17332 (N_17332,N_16301,N_16495);
xor U17333 (N_17333,N_16792,N_16440);
nor U17334 (N_17334,N_16033,N_16205);
or U17335 (N_17335,N_16760,N_16581);
or U17336 (N_17336,N_16531,N_16193);
nand U17337 (N_17337,N_16333,N_16316);
xnor U17338 (N_17338,N_16297,N_16528);
nand U17339 (N_17339,N_16759,N_16792);
nor U17340 (N_17340,N_16612,N_16668);
xnor U17341 (N_17341,N_16552,N_16139);
nand U17342 (N_17342,N_16057,N_16713);
or U17343 (N_17343,N_16407,N_16546);
and U17344 (N_17344,N_16557,N_16038);
nand U17345 (N_17345,N_16206,N_16405);
nand U17346 (N_17346,N_16613,N_16431);
nor U17347 (N_17347,N_16041,N_16055);
nor U17348 (N_17348,N_16693,N_16636);
or U17349 (N_17349,N_16122,N_16232);
nand U17350 (N_17350,N_16569,N_16408);
and U17351 (N_17351,N_16185,N_16477);
xnor U17352 (N_17352,N_16462,N_16676);
nor U17353 (N_17353,N_16285,N_16161);
or U17354 (N_17354,N_16102,N_16284);
or U17355 (N_17355,N_16340,N_16143);
and U17356 (N_17356,N_16757,N_16032);
xnor U17357 (N_17357,N_16626,N_16579);
nor U17358 (N_17358,N_16745,N_16242);
nor U17359 (N_17359,N_16166,N_16289);
and U17360 (N_17360,N_16589,N_16094);
nand U17361 (N_17361,N_16791,N_16152);
nor U17362 (N_17362,N_16457,N_16632);
xor U17363 (N_17363,N_16003,N_16018);
nor U17364 (N_17364,N_16654,N_16397);
or U17365 (N_17365,N_16665,N_16029);
nand U17366 (N_17366,N_16726,N_16628);
xnor U17367 (N_17367,N_16716,N_16779);
xor U17368 (N_17368,N_16151,N_16039);
nor U17369 (N_17369,N_16611,N_16288);
or U17370 (N_17370,N_16246,N_16122);
and U17371 (N_17371,N_16157,N_16532);
nand U17372 (N_17372,N_16157,N_16783);
or U17373 (N_17373,N_16207,N_16108);
nor U17374 (N_17374,N_16196,N_16270);
xnor U17375 (N_17375,N_16137,N_16556);
xnor U17376 (N_17376,N_16445,N_16139);
nand U17377 (N_17377,N_16718,N_16038);
and U17378 (N_17378,N_16489,N_16284);
nand U17379 (N_17379,N_16509,N_16111);
or U17380 (N_17380,N_16381,N_16273);
or U17381 (N_17381,N_16487,N_16298);
xor U17382 (N_17382,N_16254,N_16083);
nand U17383 (N_17383,N_16575,N_16586);
or U17384 (N_17384,N_16412,N_16084);
xnor U17385 (N_17385,N_16727,N_16085);
nor U17386 (N_17386,N_16563,N_16502);
nand U17387 (N_17387,N_16203,N_16128);
or U17388 (N_17388,N_16074,N_16452);
and U17389 (N_17389,N_16706,N_16738);
and U17390 (N_17390,N_16377,N_16024);
nor U17391 (N_17391,N_16557,N_16361);
or U17392 (N_17392,N_16576,N_16727);
or U17393 (N_17393,N_16360,N_16042);
and U17394 (N_17394,N_16526,N_16329);
and U17395 (N_17395,N_16128,N_16687);
xnor U17396 (N_17396,N_16522,N_16319);
nand U17397 (N_17397,N_16009,N_16713);
xnor U17398 (N_17398,N_16537,N_16573);
nand U17399 (N_17399,N_16470,N_16638);
nor U17400 (N_17400,N_16077,N_16759);
xnor U17401 (N_17401,N_16176,N_16770);
nor U17402 (N_17402,N_16794,N_16681);
or U17403 (N_17403,N_16042,N_16235);
and U17404 (N_17404,N_16617,N_16668);
xor U17405 (N_17405,N_16076,N_16742);
xnor U17406 (N_17406,N_16236,N_16275);
nor U17407 (N_17407,N_16594,N_16583);
xnor U17408 (N_17408,N_16528,N_16017);
xor U17409 (N_17409,N_16441,N_16789);
and U17410 (N_17410,N_16310,N_16683);
nor U17411 (N_17411,N_16754,N_16670);
and U17412 (N_17412,N_16201,N_16280);
or U17413 (N_17413,N_16793,N_16274);
or U17414 (N_17414,N_16770,N_16127);
and U17415 (N_17415,N_16557,N_16736);
and U17416 (N_17416,N_16033,N_16541);
or U17417 (N_17417,N_16366,N_16674);
nor U17418 (N_17418,N_16323,N_16763);
or U17419 (N_17419,N_16464,N_16405);
nand U17420 (N_17420,N_16091,N_16798);
nand U17421 (N_17421,N_16436,N_16093);
and U17422 (N_17422,N_16327,N_16182);
or U17423 (N_17423,N_16789,N_16195);
nor U17424 (N_17424,N_16093,N_16358);
or U17425 (N_17425,N_16275,N_16230);
and U17426 (N_17426,N_16517,N_16732);
and U17427 (N_17427,N_16427,N_16473);
nand U17428 (N_17428,N_16785,N_16449);
or U17429 (N_17429,N_16027,N_16374);
nand U17430 (N_17430,N_16189,N_16776);
xnor U17431 (N_17431,N_16029,N_16789);
nor U17432 (N_17432,N_16258,N_16277);
and U17433 (N_17433,N_16175,N_16534);
or U17434 (N_17434,N_16150,N_16035);
nand U17435 (N_17435,N_16774,N_16700);
xnor U17436 (N_17436,N_16095,N_16196);
xnor U17437 (N_17437,N_16449,N_16152);
and U17438 (N_17438,N_16277,N_16605);
and U17439 (N_17439,N_16672,N_16468);
nor U17440 (N_17440,N_16338,N_16283);
and U17441 (N_17441,N_16110,N_16241);
xor U17442 (N_17442,N_16026,N_16566);
nand U17443 (N_17443,N_16418,N_16372);
or U17444 (N_17444,N_16538,N_16226);
or U17445 (N_17445,N_16436,N_16252);
nor U17446 (N_17446,N_16600,N_16773);
xor U17447 (N_17447,N_16662,N_16669);
and U17448 (N_17448,N_16030,N_16666);
xnor U17449 (N_17449,N_16227,N_16588);
nor U17450 (N_17450,N_16224,N_16344);
nor U17451 (N_17451,N_16412,N_16225);
xor U17452 (N_17452,N_16133,N_16157);
and U17453 (N_17453,N_16692,N_16250);
and U17454 (N_17454,N_16462,N_16733);
nand U17455 (N_17455,N_16417,N_16651);
nand U17456 (N_17456,N_16653,N_16686);
and U17457 (N_17457,N_16743,N_16706);
and U17458 (N_17458,N_16502,N_16481);
nor U17459 (N_17459,N_16340,N_16727);
nand U17460 (N_17460,N_16585,N_16466);
nand U17461 (N_17461,N_16681,N_16065);
or U17462 (N_17462,N_16322,N_16422);
nand U17463 (N_17463,N_16586,N_16385);
and U17464 (N_17464,N_16440,N_16376);
or U17465 (N_17465,N_16184,N_16170);
nand U17466 (N_17466,N_16071,N_16194);
nand U17467 (N_17467,N_16552,N_16779);
and U17468 (N_17468,N_16215,N_16738);
or U17469 (N_17469,N_16251,N_16569);
xor U17470 (N_17470,N_16520,N_16521);
nor U17471 (N_17471,N_16418,N_16379);
xor U17472 (N_17472,N_16013,N_16015);
or U17473 (N_17473,N_16151,N_16540);
xnor U17474 (N_17474,N_16145,N_16557);
xnor U17475 (N_17475,N_16339,N_16061);
nand U17476 (N_17476,N_16532,N_16557);
or U17477 (N_17477,N_16031,N_16554);
nor U17478 (N_17478,N_16238,N_16142);
or U17479 (N_17479,N_16496,N_16241);
xnor U17480 (N_17480,N_16456,N_16556);
xor U17481 (N_17481,N_16584,N_16388);
and U17482 (N_17482,N_16765,N_16534);
or U17483 (N_17483,N_16701,N_16060);
or U17484 (N_17484,N_16619,N_16272);
xnor U17485 (N_17485,N_16449,N_16566);
and U17486 (N_17486,N_16373,N_16464);
nand U17487 (N_17487,N_16169,N_16635);
nor U17488 (N_17488,N_16520,N_16492);
nand U17489 (N_17489,N_16562,N_16315);
xor U17490 (N_17490,N_16720,N_16486);
xor U17491 (N_17491,N_16397,N_16458);
xor U17492 (N_17492,N_16247,N_16339);
xor U17493 (N_17493,N_16320,N_16216);
nor U17494 (N_17494,N_16521,N_16067);
nand U17495 (N_17495,N_16375,N_16683);
nand U17496 (N_17496,N_16374,N_16780);
xnor U17497 (N_17497,N_16743,N_16545);
or U17498 (N_17498,N_16560,N_16203);
or U17499 (N_17499,N_16603,N_16654);
xnor U17500 (N_17500,N_16628,N_16338);
xor U17501 (N_17501,N_16434,N_16014);
or U17502 (N_17502,N_16729,N_16281);
and U17503 (N_17503,N_16022,N_16788);
nor U17504 (N_17504,N_16743,N_16435);
or U17505 (N_17505,N_16631,N_16312);
nand U17506 (N_17506,N_16097,N_16347);
or U17507 (N_17507,N_16608,N_16506);
or U17508 (N_17508,N_16101,N_16785);
or U17509 (N_17509,N_16081,N_16656);
or U17510 (N_17510,N_16243,N_16709);
xnor U17511 (N_17511,N_16011,N_16036);
or U17512 (N_17512,N_16670,N_16326);
xnor U17513 (N_17513,N_16238,N_16659);
nand U17514 (N_17514,N_16623,N_16460);
nor U17515 (N_17515,N_16428,N_16703);
nand U17516 (N_17516,N_16110,N_16467);
and U17517 (N_17517,N_16081,N_16521);
nor U17518 (N_17518,N_16405,N_16229);
nand U17519 (N_17519,N_16587,N_16683);
nand U17520 (N_17520,N_16514,N_16463);
xnor U17521 (N_17521,N_16668,N_16277);
and U17522 (N_17522,N_16414,N_16529);
nand U17523 (N_17523,N_16207,N_16534);
nor U17524 (N_17524,N_16776,N_16149);
nor U17525 (N_17525,N_16665,N_16568);
nand U17526 (N_17526,N_16032,N_16748);
nor U17527 (N_17527,N_16236,N_16296);
nor U17528 (N_17528,N_16292,N_16482);
nand U17529 (N_17529,N_16293,N_16425);
nor U17530 (N_17530,N_16471,N_16668);
or U17531 (N_17531,N_16499,N_16349);
nor U17532 (N_17532,N_16602,N_16178);
and U17533 (N_17533,N_16433,N_16423);
xor U17534 (N_17534,N_16257,N_16493);
or U17535 (N_17535,N_16438,N_16755);
nand U17536 (N_17536,N_16799,N_16178);
or U17537 (N_17537,N_16163,N_16788);
xnor U17538 (N_17538,N_16758,N_16081);
or U17539 (N_17539,N_16079,N_16659);
nor U17540 (N_17540,N_16054,N_16360);
nor U17541 (N_17541,N_16187,N_16337);
nor U17542 (N_17542,N_16213,N_16211);
or U17543 (N_17543,N_16529,N_16147);
nand U17544 (N_17544,N_16052,N_16211);
or U17545 (N_17545,N_16494,N_16018);
nor U17546 (N_17546,N_16444,N_16080);
or U17547 (N_17547,N_16409,N_16677);
and U17548 (N_17548,N_16167,N_16170);
and U17549 (N_17549,N_16443,N_16449);
xnor U17550 (N_17550,N_16698,N_16024);
nand U17551 (N_17551,N_16359,N_16184);
nand U17552 (N_17552,N_16321,N_16708);
or U17553 (N_17553,N_16004,N_16707);
nand U17554 (N_17554,N_16603,N_16491);
and U17555 (N_17555,N_16385,N_16551);
xor U17556 (N_17556,N_16563,N_16368);
and U17557 (N_17557,N_16238,N_16031);
nand U17558 (N_17558,N_16540,N_16302);
xnor U17559 (N_17559,N_16372,N_16661);
nand U17560 (N_17560,N_16289,N_16413);
xor U17561 (N_17561,N_16229,N_16489);
nand U17562 (N_17562,N_16301,N_16027);
and U17563 (N_17563,N_16713,N_16429);
nand U17564 (N_17564,N_16463,N_16043);
xor U17565 (N_17565,N_16284,N_16723);
and U17566 (N_17566,N_16498,N_16685);
and U17567 (N_17567,N_16165,N_16600);
nor U17568 (N_17568,N_16169,N_16604);
xnor U17569 (N_17569,N_16735,N_16337);
or U17570 (N_17570,N_16782,N_16597);
or U17571 (N_17571,N_16029,N_16587);
nand U17572 (N_17572,N_16139,N_16405);
nand U17573 (N_17573,N_16746,N_16342);
nor U17574 (N_17574,N_16725,N_16317);
and U17575 (N_17575,N_16230,N_16550);
xor U17576 (N_17576,N_16755,N_16580);
and U17577 (N_17577,N_16438,N_16521);
xor U17578 (N_17578,N_16507,N_16168);
or U17579 (N_17579,N_16568,N_16167);
xnor U17580 (N_17580,N_16430,N_16235);
nand U17581 (N_17581,N_16545,N_16356);
and U17582 (N_17582,N_16017,N_16478);
nor U17583 (N_17583,N_16214,N_16696);
nand U17584 (N_17584,N_16280,N_16122);
xor U17585 (N_17585,N_16545,N_16507);
nor U17586 (N_17586,N_16022,N_16015);
and U17587 (N_17587,N_16062,N_16181);
xor U17588 (N_17588,N_16211,N_16651);
nand U17589 (N_17589,N_16213,N_16719);
nand U17590 (N_17590,N_16760,N_16243);
xnor U17591 (N_17591,N_16623,N_16725);
or U17592 (N_17592,N_16719,N_16179);
nand U17593 (N_17593,N_16290,N_16758);
and U17594 (N_17594,N_16720,N_16570);
or U17595 (N_17595,N_16349,N_16126);
and U17596 (N_17596,N_16676,N_16365);
nand U17597 (N_17597,N_16125,N_16272);
nor U17598 (N_17598,N_16486,N_16101);
xnor U17599 (N_17599,N_16352,N_16613);
or U17600 (N_17600,N_17066,N_17142);
and U17601 (N_17601,N_16831,N_17522);
xor U17602 (N_17602,N_17490,N_17435);
or U17603 (N_17603,N_16819,N_17588);
xor U17604 (N_17604,N_17068,N_16912);
nand U17605 (N_17605,N_17308,N_17237);
nand U17606 (N_17606,N_17331,N_16957);
nand U17607 (N_17607,N_17310,N_17302);
nor U17608 (N_17608,N_17055,N_17159);
and U17609 (N_17609,N_16808,N_17177);
or U17610 (N_17610,N_17321,N_17035);
xor U17611 (N_17611,N_17200,N_16940);
or U17612 (N_17612,N_16852,N_17556);
and U17613 (N_17613,N_17185,N_17313);
xnor U17614 (N_17614,N_17092,N_17328);
or U17615 (N_17615,N_17564,N_17131);
xnor U17616 (N_17616,N_16938,N_17444);
or U17617 (N_17617,N_16899,N_17501);
nand U17618 (N_17618,N_17195,N_17404);
and U17619 (N_17619,N_17259,N_17382);
xor U17620 (N_17620,N_17376,N_16875);
or U17621 (N_17621,N_17340,N_17231);
xor U17622 (N_17622,N_17080,N_16960);
nor U17623 (N_17623,N_17447,N_17593);
nand U17624 (N_17624,N_17081,N_16821);
nand U17625 (N_17625,N_16893,N_17000);
or U17626 (N_17626,N_17108,N_17175);
nor U17627 (N_17627,N_17364,N_16844);
or U17628 (N_17628,N_17220,N_16973);
nand U17629 (N_17629,N_16870,N_17106);
nor U17630 (N_17630,N_17184,N_17477);
nand U17631 (N_17631,N_17533,N_17458);
nor U17632 (N_17632,N_16931,N_17141);
xnor U17633 (N_17633,N_17069,N_16918);
nand U17634 (N_17634,N_17114,N_17459);
and U17635 (N_17635,N_16980,N_17309);
and U17636 (N_17636,N_17467,N_17329);
nor U17637 (N_17637,N_17421,N_17586);
and U17638 (N_17638,N_17552,N_17565);
and U17639 (N_17639,N_17377,N_17418);
and U17640 (N_17640,N_17074,N_16914);
and U17641 (N_17641,N_17219,N_17207);
nor U17642 (N_17642,N_17492,N_17059);
xor U17643 (N_17643,N_17233,N_17457);
nor U17644 (N_17644,N_17493,N_17222);
nand U17645 (N_17645,N_17428,N_17130);
nand U17646 (N_17646,N_17006,N_17167);
or U17647 (N_17647,N_17286,N_17359);
or U17648 (N_17648,N_17216,N_17266);
xor U17649 (N_17649,N_17496,N_16888);
and U17650 (N_17650,N_16959,N_17296);
or U17651 (N_17651,N_17532,N_17518);
nor U17652 (N_17652,N_16983,N_17137);
nor U17653 (N_17653,N_16845,N_17335);
or U17654 (N_17654,N_17127,N_17441);
nand U17655 (N_17655,N_17139,N_17476);
xnor U17656 (N_17656,N_17365,N_17483);
xnor U17657 (N_17657,N_17007,N_17390);
or U17658 (N_17658,N_16853,N_17230);
or U17659 (N_17659,N_16862,N_17361);
nor U17660 (N_17660,N_17555,N_16977);
nand U17661 (N_17661,N_17228,N_17126);
nand U17662 (N_17662,N_17383,N_17103);
nand U17663 (N_17663,N_17598,N_16811);
xor U17664 (N_17664,N_17057,N_17306);
and U17665 (N_17665,N_16967,N_17138);
nor U17666 (N_17666,N_17478,N_17115);
xnor U17667 (N_17667,N_17553,N_17579);
and U17668 (N_17668,N_17295,N_17014);
nand U17669 (N_17669,N_17503,N_17149);
nand U17670 (N_17670,N_17344,N_17443);
xnor U17671 (N_17671,N_17395,N_17368);
nand U17672 (N_17672,N_17509,N_16873);
or U17673 (N_17673,N_17086,N_17070);
nor U17674 (N_17674,N_16898,N_17456);
and U17675 (N_17675,N_17243,N_17168);
and U17676 (N_17676,N_17349,N_17363);
nand U17677 (N_17677,N_17119,N_17160);
nand U17678 (N_17678,N_17495,N_17537);
nor U17679 (N_17679,N_17357,N_17387);
xor U17680 (N_17680,N_17027,N_17234);
and U17681 (N_17681,N_17431,N_17193);
nand U17682 (N_17682,N_17013,N_17544);
nand U17683 (N_17683,N_17454,N_17320);
nor U17684 (N_17684,N_17560,N_17585);
or U17685 (N_17685,N_17209,N_17499);
xor U17686 (N_17686,N_17410,N_16849);
nor U17687 (N_17687,N_17225,N_17301);
nor U17688 (N_17688,N_17272,N_16840);
xor U17689 (N_17689,N_16805,N_17434);
and U17690 (N_17690,N_17534,N_17411);
or U17691 (N_17691,N_17021,N_17463);
xnor U17692 (N_17692,N_17455,N_17194);
nor U17693 (N_17693,N_17551,N_16908);
xor U17694 (N_17694,N_16939,N_16949);
nor U17695 (N_17695,N_17164,N_16901);
nand U17696 (N_17696,N_17392,N_17267);
nor U17697 (N_17697,N_17226,N_16824);
and U17698 (N_17698,N_17326,N_16857);
and U17699 (N_17699,N_17210,N_17214);
nor U17700 (N_17700,N_17022,N_17319);
or U17701 (N_17701,N_17337,N_17204);
xor U17702 (N_17702,N_17251,N_17072);
nor U17703 (N_17703,N_17051,N_16987);
or U17704 (N_17704,N_17017,N_17576);
and U17705 (N_17705,N_16815,N_17293);
or U17706 (N_17706,N_17557,N_17236);
and U17707 (N_17707,N_16814,N_17186);
nand U17708 (N_17708,N_17091,N_17113);
nor U17709 (N_17709,N_17474,N_16827);
or U17710 (N_17710,N_17386,N_17339);
nand U17711 (N_17711,N_17519,N_16843);
or U17712 (N_17712,N_16913,N_17547);
nor U17713 (N_17713,N_17545,N_16861);
nor U17714 (N_17714,N_17374,N_17062);
or U17715 (N_17715,N_16891,N_16934);
nand U17716 (N_17716,N_17128,N_16932);
nor U17717 (N_17717,N_16859,N_17394);
xor U17718 (N_17718,N_16975,N_17437);
xnor U17719 (N_17719,N_17054,N_17384);
nand U17720 (N_17720,N_17156,N_16904);
or U17721 (N_17721,N_17095,N_16919);
nor U17722 (N_17722,N_17120,N_16922);
nor U17723 (N_17723,N_16855,N_17292);
or U17724 (N_17724,N_17279,N_16955);
and U17725 (N_17725,N_17582,N_17248);
nor U17726 (N_17726,N_17379,N_17269);
or U17727 (N_17727,N_17527,N_17166);
nor U17728 (N_17728,N_17255,N_16945);
or U17729 (N_17729,N_17373,N_17439);
and U17730 (N_17730,N_16863,N_17351);
xnor U17731 (N_17731,N_16838,N_17132);
and U17732 (N_17732,N_17469,N_17366);
nor U17733 (N_17733,N_17152,N_16833);
xnor U17734 (N_17734,N_16905,N_16883);
nor U17735 (N_17735,N_17121,N_17050);
and U17736 (N_17736,N_17550,N_16995);
or U17737 (N_17737,N_17355,N_17278);
or U17738 (N_17738,N_17472,N_17155);
or U17739 (N_17739,N_17378,N_16807);
nor U17740 (N_17740,N_17283,N_17536);
and U17741 (N_17741,N_16981,N_17118);
nor U17742 (N_17742,N_17085,N_17165);
xnor U17743 (N_17743,N_17333,N_16956);
and U17744 (N_17744,N_16801,N_16816);
and U17745 (N_17745,N_17178,N_17073);
nand U17746 (N_17746,N_17133,N_17161);
and U17747 (N_17747,N_16884,N_16989);
xor U17748 (N_17748,N_16868,N_16818);
nand U17749 (N_17749,N_16900,N_17104);
nand U17750 (N_17750,N_17599,N_17354);
or U17751 (N_17751,N_16806,N_17526);
xnor U17752 (N_17752,N_17403,N_16910);
and U17753 (N_17753,N_16889,N_17083);
nor U17754 (N_17754,N_17360,N_17488);
or U17755 (N_17755,N_16860,N_17135);
nor U17756 (N_17756,N_17198,N_17004);
or U17757 (N_17757,N_17487,N_17049);
nand U17758 (N_17758,N_17399,N_17169);
xnor U17759 (N_17759,N_16974,N_17498);
nand U17760 (N_17760,N_17485,N_17427);
nor U17761 (N_17761,N_17569,N_17426);
or U17762 (N_17762,N_17117,N_16847);
xor U17763 (N_17763,N_17205,N_16856);
nor U17764 (N_17764,N_17046,N_17442);
or U17765 (N_17765,N_16924,N_17514);
xor U17766 (N_17766,N_17290,N_17034);
nor U17767 (N_17767,N_17516,N_16982);
xor U17768 (N_17768,N_17396,N_17018);
nand U17769 (N_17769,N_17330,N_17291);
nand U17770 (N_17770,N_17566,N_17572);
nor U17771 (N_17771,N_17523,N_17071);
xor U17772 (N_17772,N_17257,N_17239);
nor U17773 (N_17773,N_16866,N_17563);
nand U17774 (N_17774,N_17247,N_16990);
or U17775 (N_17775,N_17245,N_17024);
nand U17776 (N_17776,N_17388,N_17543);
and U17777 (N_17777,N_17494,N_17145);
xnor U17778 (N_17778,N_17093,N_17192);
or U17779 (N_17779,N_17419,N_17353);
or U17780 (N_17780,N_17486,N_16943);
or U17781 (N_17781,N_17078,N_17491);
and U17782 (N_17782,N_17263,N_16878);
and U17783 (N_17783,N_17256,N_17574);
nor U17784 (N_17784,N_17505,N_17067);
and U17785 (N_17785,N_17489,N_17546);
xnor U17786 (N_17786,N_16962,N_17208);
and U17787 (N_17787,N_16991,N_17541);
and U17788 (N_17788,N_17596,N_16950);
or U17789 (N_17789,N_16988,N_17438);
nor U17790 (N_17790,N_16882,N_16817);
xnor U17791 (N_17791,N_17273,N_17107);
and U17792 (N_17792,N_17285,N_17176);
and U17793 (N_17793,N_16892,N_17077);
nor U17794 (N_17794,N_17146,N_17500);
nand U17795 (N_17795,N_17450,N_17412);
nor U17796 (N_17796,N_16822,N_17398);
or U17797 (N_17797,N_16830,N_17023);
or U17798 (N_17798,N_17154,N_16851);
xor U17799 (N_17799,N_17451,N_17481);
nand U17800 (N_17800,N_17362,N_16823);
and U17801 (N_17801,N_17030,N_16804);
xnor U17802 (N_17802,N_16825,N_17352);
xor U17803 (N_17803,N_17568,N_17153);
and U17804 (N_17804,N_17162,N_17221);
xnor U17805 (N_17805,N_17482,N_16865);
nor U17806 (N_17806,N_17417,N_17033);
xor U17807 (N_17807,N_17042,N_16829);
nor U17808 (N_17808,N_17275,N_17510);
nand U17809 (N_17809,N_17157,N_17468);
and U17810 (N_17810,N_17520,N_17174);
or U17811 (N_17811,N_17199,N_17549);
xnor U17812 (N_17812,N_17422,N_17578);
and U17813 (N_17813,N_17590,N_16848);
xnor U17814 (N_17814,N_17241,N_17056);
nor U17815 (N_17815,N_16877,N_17090);
xor U17816 (N_17816,N_17372,N_17298);
nand U17817 (N_17817,N_17143,N_17334);
nand U17818 (N_17818,N_17327,N_17343);
nor U17819 (N_17819,N_17316,N_17587);
xnor U17820 (N_17820,N_16841,N_17045);
xor U17821 (N_17821,N_16944,N_17479);
and U17822 (N_17822,N_17448,N_16885);
nand U17823 (N_17823,N_17484,N_17538);
nand U17824 (N_17824,N_17271,N_17032);
xor U17825 (N_17825,N_17462,N_16994);
nor U17826 (N_17826,N_17274,N_17525);
xnor U17827 (N_17827,N_17129,N_16976);
nor U17828 (N_17828,N_17440,N_17089);
nand U17829 (N_17829,N_17163,N_17276);
xor U17830 (N_17830,N_17466,N_17594);
and U17831 (N_17831,N_16920,N_17406);
nor U17832 (N_17832,N_17511,N_16978);
xnor U17833 (N_17833,N_17539,N_17172);
and U17834 (N_17834,N_17179,N_16970);
nand U17835 (N_17835,N_17036,N_17196);
or U17836 (N_17836,N_16890,N_16813);
xor U17837 (N_17837,N_17227,N_17268);
and U17838 (N_17838,N_17350,N_17413);
nand U17839 (N_17839,N_17112,N_17063);
xnor U17840 (N_17840,N_17480,N_17088);
nor U17841 (N_17841,N_16923,N_16915);
xor U17842 (N_17842,N_17342,N_17173);
nand U17843 (N_17843,N_16926,N_17009);
and U17844 (N_17844,N_17506,N_17052);
nor U17845 (N_17845,N_16879,N_16828);
nand U17846 (N_17846,N_17453,N_17348);
and U17847 (N_17847,N_17109,N_17096);
xnor U17848 (N_17848,N_17215,N_16869);
xor U17849 (N_17849,N_17076,N_17529);
xnor U17850 (N_17850,N_17099,N_17452);
or U17851 (N_17851,N_17002,N_16952);
xnor U17852 (N_17852,N_17244,N_16903);
or U17853 (N_17853,N_16936,N_17048);
xnor U17854 (N_17854,N_16846,N_17264);
or U17855 (N_17855,N_17211,N_16812);
nand U17856 (N_17856,N_17515,N_17380);
and U17857 (N_17857,N_17280,N_17005);
nand U17858 (N_17858,N_17464,N_16842);
xor U17859 (N_17859,N_17561,N_17341);
xnor U17860 (N_17860,N_17581,N_16997);
and U17861 (N_17861,N_16937,N_17540);
nor U17862 (N_17862,N_17391,N_16902);
xnor U17863 (N_17863,N_17562,N_17213);
xor U17864 (N_17864,N_17583,N_16858);
xor U17865 (N_17865,N_17218,N_17147);
nor U17866 (N_17866,N_16880,N_16895);
and U17867 (N_17867,N_17430,N_17043);
nor U17868 (N_17868,N_17212,N_17202);
and U17869 (N_17869,N_17305,N_17345);
xor U17870 (N_17870,N_17038,N_17001);
and U17871 (N_17871,N_16809,N_17188);
or U17872 (N_17872,N_16927,N_17521);
or U17873 (N_17873,N_17317,N_17528);
xnor U17874 (N_17874,N_16925,N_16941);
xor U17875 (N_17875,N_17136,N_17206);
nand U17876 (N_17876,N_16948,N_17397);
xor U17877 (N_17877,N_17558,N_16906);
nor U17878 (N_17878,N_16993,N_17170);
nand U17879 (N_17879,N_17189,N_17182);
xnor U17880 (N_17880,N_17252,N_16954);
and U17881 (N_17881,N_17242,N_17318);
nor U17882 (N_17882,N_17250,N_16921);
and U17883 (N_17883,N_17294,N_16836);
xnor U17884 (N_17884,N_16896,N_16930);
and U17885 (N_17885,N_16942,N_17323);
nor U17886 (N_17886,N_16871,N_17436);
nor U17887 (N_17887,N_17371,N_17116);
or U17888 (N_17888,N_17031,N_17240);
xnor U17889 (N_17889,N_16837,N_17420);
xnor U17890 (N_17890,N_16886,N_16872);
nand U17891 (N_17891,N_16953,N_17571);
nor U17892 (N_17892,N_16916,N_17282);
and U17893 (N_17893,N_17589,N_17470);
or U17894 (N_17894,N_16826,N_16911);
and U17895 (N_17895,N_16933,N_17111);
and U17896 (N_17896,N_17098,N_17281);
xnor U17897 (N_17897,N_17148,N_17465);
and U17898 (N_17898,N_17535,N_16800);
and U17899 (N_17899,N_17284,N_17065);
xnor U17900 (N_17900,N_17082,N_16958);
and U17901 (N_17901,N_17249,N_16998);
nand U17902 (N_17902,N_17424,N_16835);
or U17903 (N_17903,N_17325,N_17580);
or U17904 (N_17904,N_17288,N_17414);
or U17905 (N_17905,N_17393,N_16996);
xor U17906 (N_17906,N_17389,N_17123);
nor U17907 (N_17907,N_17531,N_17203);
or U17908 (N_17908,N_17471,N_16832);
nand U17909 (N_17909,N_16968,N_17358);
xnor U17910 (N_17910,N_16907,N_17044);
nand U17911 (N_17911,N_16946,N_17449);
xnor U17912 (N_17912,N_17102,N_17064);
nor U17913 (N_17913,N_17084,N_16951);
nor U17914 (N_17914,N_17445,N_17235);
nor U17915 (N_17915,N_17332,N_17238);
or U17916 (N_17916,N_17338,N_17375);
and U17917 (N_17917,N_16985,N_16964);
nor U17918 (N_17918,N_16969,N_17554);
nor U17919 (N_17919,N_17559,N_17262);
nand U17920 (N_17920,N_16971,N_17461);
and U17921 (N_17921,N_17592,N_17101);
nand U17922 (N_17922,N_17415,N_17429);
nand U17923 (N_17923,N_17223,N_17094);
or U17924 (N_17924,N_17041,N_17407);
nand U17925 (N_17925,N_16874,N_16929);
or U17926 (N_17926,N_17507,N_16876);
nor U17927 (N_17927,N_17187,N_17058);
nor U17928 (N_17928,N_17597,N_16917);
or U17929 (N_17929,N_17003,N_17151);
xor U17930 (N_17930,N_17100,N_17019);
xnor U17931 (N_17931,N_17144,N_17181);
xor U17932 (N_17932,N_17020,N_16965);
xor U17933 (N_17933,N_17012,N_17190);
xnor U17934 (N_17934,N_17246,N_17171);
or U17935 (N_17935,N_16820,N_17577);
nor U17936 (N_17936,N_17265,N_17297);
nand U17937 (N_17937,N_17432,N_17409);
and U17938 (N_17938,N_16979,N_17307);
or U17939 (N_17939,N_17011,N_16897);
nand U17940 (N_17940,N_17567,N_17039);
nand U17941 (N_17941,N_17040,N_17258);
xnor U17942 (N_17942,N_17122,N_17158);
nand U17943 (N_17943,N_16802,N_17591);
and U17944 (N_17944,N_17315,N_17025);
xnor U17945 (N_17945,N_16972,N_17289);
xor U17946 (N_17946,N_16963,N_17497);
or U17947 (N_17947,N_17475,N_17134);
nor U17948 (N_17948,N_17400,N_17304);
and U17949 (N_17949,N_17584,N_17460);
or U17950 (N_17950,N_17303,N_17026);
nor U17951 (N_17951,N_17287,N_17508);
and U17952 (N_17952,N_17061,N_16947);
nand U17953 (N_17953,N_17370,N_17595);
nor U17954 (N_17954,N_17097,N_17401);
and U17955 (N_17955,N_17336,N_16961);
nand U17956 (N_17956,N_17110,N_16999);
nor U17957 (N_17957,N_17408,N_17312);
and U17958 (N_17958,N_17322,N_17053);
nor U17959 (N_17959,N_16887,N_16850);
or U17960 (N_17960,N_17029,N_17433);
nor U17961 (N_17961,N_17232,N_17311);
nand U17962 (N_17962,N_17548,N_17105);
xnor U17963 (N_17963,N_17369,N_17224);
xnor U17964 (N_17964,N_17517,N_17502);
and U17965 (N_17965,N_17015,N_17253);
and U17966 (N_17966,N_17524,N_16935);
or U17967 (N_17967,N_17446,N_16810);
nand U17968 (N_17968,N_17183,N_16864);
nor U17969 (N_17969,N_17079,N_17010);
or U17970 (N_17970,N_17473,N_17150);
xnor U17971 (N_17971,N_17047,N_17254);
and U17972 (N_17972,N_17028,N_16894);
nor U17973 (N_17973,N_17542,N_16966);
and U17974 (N_17974,N_17347,N_17324);
or U17975 (N_17975,N_17381,N_17201);
and U17976 (N_17976,N_17425,N_17367);
nand U17977 (N_17977,N_16867,N_17008);
nand U17978 (N_17978,N_16854,N_17217);
nand U17979 (N_17979,N_16986,N_16984);
or U17980 (N_17980,N_17570,N_17075);
xor U17981 (N_17981,N_16803,N_17346);
nor U17982 (N_17982,N_17037,N_17402);
xor U17983 (N_17983,N_17229,N_16839);
nor U17984 (N_17984,N_17513,N_17180);
xor U17985 (N_17985,N_17423,N_17356);
and U17986 (N_17986,N_17530,N_17405);
and U17987 (N_17987,N_16992,N_17124);
or U17988 (N_17988,N_17197,N_17416);
or U17989 (N_17989,N_17512,N_17261);
nand U17990 (N_17990,N_17016,N_16881);
nand U17991 (N_17991,N_17300,N_17277);
or U17992 (N_17992,N_17125,N_16834);
xor U17993 (N_17993,N_17060,N_17087);
or U17994 (N_17994,N_17314,N_17575);
xor U17995 (N_17995,N_17140,N_17573);
nand U17996 (N_17996,N_17191,N_17260);
and U17997 (N_17997,N_17385,N_16909);
nand U17998 (N_17998,N_17299,N_17504);
nor U17999 (N_17999,N_17270,N_16928);
and U18000 (N_18000,N_17095,N_17532);
nor U18001 (N_18001,N_17285,N_17256);
or U18002 (N_18002,N_16966,N_17420);
xnor U18003 (N_18003,N_17363,N_17252);
or U18004 (N_18004,N_17466,N_17009);
nand U18005 (N_18005,N_17446,N_17490);
nand U18006 (N_18006,N_16892,N_17365);
and U18007 (N_18007,N_16981,N_16978);
or U18008 (N_18008,N_17225,N_17502);
xnor U18009 (N_18009,N_17187,N_17085);
xor U18010 (N_18010,N_17483,N_16839);
nor U18011 (N_18011,N_17435,N_17307);
nand U18012 (N_18012,N_17558,N_17012);
nor U18013 (N_18013,N_16889,N_17161);
xor U18014 (N_18014,N_16975,N_17407);
or U18015 (N_18015,N_16927,N_17298);
xnor U18016 (N_18016,N_16832,N_17422);
xor U18017 (N_18017,N_17062,N_17422);
nor U18018 (N_18018,N_17401,N_17219);
nand U18019 (N_18019,N_16900,N_17183);
nand U18020 (N_18020,N_16953,N_17524);
nor U18021 (N_18021,N_17478,N_17373);
nor U18022 (N_18022,N_17138,N_17135);
or U18023 (N_18023,N_17063,N_17542);
or U18024 (N_18024,N_16826,N_17223);
nand U18025 (N_18025,N_17168,N_17154);
and U18026 (N_18026,N_16867,N_17102);
or U18027 (N_18027,N_17182,N_17185);
or U18028 (N_18028,N_17209,N_17302);
xor U18029 (N_18029,N_17002,N_17008);
or U18030 (N_18030,N_17255,N_17542);
nor U18031 (N_18031,N_17528,N_17149);
nand U18032 (N_18032,N_17573,N_17592);
nor U18033 (N_18033,N_16970,N_17059);
nor U18034 (N_18034,N_16969,N_17491);
nand U18035 (N_18035,N_17504,N_17210);
xor U18036 (N_18036,N_17040,N_17143);
or U18037 (N_18037,N_17124,N_16966);
nor U18038 (N_18038,N_16912,N_17346);
or U18039 (N_18039,N_16990,N_17323);
nand U18040 (N_18040,N_16924,N_17141);
nor U18041 (N_18041,N_17398,N_17395);
nand U18042 (N_18042,N_16956,N_17563);
nor U18043 (N_18043,N_17357,N_17531);
and U18044 (N_18044,N_17150,N_17551);
xnor U18045 (N_18045,N_16835,N_17358);
xor U18046 (N_18046,N_16971,N_17166);
nor U18047 (N_18047,N_17513,N_16918);
nand U18048 (N_18048,N_16873,N_17200);
nor U18049 (N_18049,N_16990,N_17042);
and U18050 (N_18050,N_17164,N_17166);
xnor U18051 (N_18051,N_17462,N_17558);
and U18052 (N_18052,N_16918,N_17076);
and U18053 (N_18053,N_17519,N_17054);
nand U18054 (N_18054,N_17118,N_17215);
or U18055 (N_18055,N_17055,N_17563);
and U18056 (N_18056,N_16824,N_17345);
xnor U18057 (N_18057,N_17569,N_17345);
xnor U18058 (N_18058,N_17270,N_16816);
nand U18059 (N_18059,N_17039,N_17374);
nand U18060 (N_18060,N_17159,N_17508);
and U18061 (N_18061,N_16815,N_17053);
nor U18062 (N_18062,N_16806,N_17018);
or U18063 (N_18063,N_17046,N_17459);
and U18064 (N_18064,N_17417,N_16806);
nor U18065 (N_18065,N_17307,N_17562);
nor U18066 (N_18066,N_17529,N_17525);
nand U18067 (N_18067,N_16894,N_17367);
xnor U18068 (N_18068,N_17063,N_17326);
and U18069 (N_18069,N_17085,N_17389);
xor U18070 (N_18070,N_17085,N_16842);
or U18071 (N_18071,N_17007,N_17487);
xor U18072 (N_18072,N_16950,N_17231);
nand U18073 (N_18073,N_16915,N_17099);
nand U18074 (N_18074,N_16996,N_17243);
or U18075 (N_18075,N_17537,N_17388);
and U18076 (N_18076,N_17376,N_16802);
xnor U18077 (N_18077,N_17245,N_17329);
and U18078 (N_18078,N_17244,N_17021);
nor U18079 (N_18079,N_17152,N_16809);
xor U18080 (N_18080,N_16944,N_16957);
and U18081 (N_18081,N_17558,N_17149);
xnor U18082 (N_18082,N_17552,N_17297);
nor U18083 (N_18083,N_17165,N_17054);
or U18084 (N_18084,N_17443,N_16840);
xor U18085 (N_18085,N_17295,N_16967);
nor U18086 (N_18086,N_17017,N_17331);
and U18087 (N_18087,N_17233,N_17055);
xnor U18088 (N_18088,N_16870,N_17305);
nand U18089 (N_18089,N_17247,N_16828);
and U18090 (N_18090,N_17106,N_17351);
xnor U18091 (N_18091,N_17291,N_17001);
or U18092 (N_18092,N_17465,N_17111);
xor U18093 (N_18093,N_16996,N_17060);
and U18094 (N_18094,N_17278,N_16952);
nor U18095 (N_18095,N_16900,N_17059);
or U18096 (N_18096,N_16882,N_17283);
nand U18097 (N_18097,N_17189,N_17517);
nor U18098 (N_18098,N_17017,N_17545);
or U18099 (N_18099,N_17189,N_17117);
nand U18100 (N_18100,N_17455,N_17045);
nor U18101 (N_18101,N_17526,N_17425);
nor U18102 (N_18102,N_17464,N_17327);
and U18103 (N_18103,N_16997,N_16831);
xor U18104 (N_18104,N_17011,N_16928);
xnor U18105 (N_18105,N_16813,N_17148);
and U18106 (N_18106,N_16975,N_17547);
and U18107 (N_18107,N_16966,N_17413);
or U18108 (N_18108,N_16824,N_17559);
or U18109 (N_18109,N_17311,N_17366);
or U18110 (N_18110,N_16826,N_16877);
xor U18111 (N_18111,N_17215,N_17066);
nand U18112 (N_18112,N_17208,N_17387);
xor U18113 (N_18113,N_16883,N_16824);
nand U18114 (N_18114,N_17338,N_17306);
and U18115 (N_18115,N_17433,N_17544);
or U18116 (N_18116,N_16956,N_16928);
nand U18117 (N_18117,N_17496,N_17551);
nand U18118 (N_18118,N_17241,N_17049);
and U18119 (N_18119,N_17467,N_16898);
xnor U18120 (N_18120,N_17196,N_17439);
nand U18121 (N_18121,N_17444,N_17517);
nand U18122 (N_18122,N_17315,N_17013);
xor U18123 (N_18123,N_17328,N_17313);
nand U18124 (N_18124,N_16885,N_16958);
or U18125 (N_18125,N_16924,N_17014);
and U18126 (N_18126,N_16871,N_16948);
and U18127 (N_18127,N_16881,N_17078);
nand U18128 (N_18128,N_17187,N_17109);
nor U18129 (N_18129,N_17030,N_16963);
nand U18130 (N_18130,N_17114,N_17054);
and U18131 (N_18131,N_17006,N_17323);
nand U18132 (N_18132,N_17358,N_17262);
or U18133 (N_18133,N_17241,N_17528);
xnor U18134 (N_18134,N_17131,N_17097);
and U18135 (N_18135,N_16826,N_16884);
xor U18136 (N_18136,N_16935,N_17483);
nor U18137 (N_18137,N_17259,N_17289);
nor U18138 (N_18138,N_17541,N_16895);
and U18139 (N_18139,N_17011,N_17197);
and U18140 (N_18140,N_17448,N_17308);
xor U18141 (N_18141,N_16806,N_17097);
nand U18142 (N_18142,N_17066,N_17140);
or U18143 (N_18143,N_17149,N_17460);
nor U18144 (N_18144,N_17367,N_17158);
or U18145 (N_18145,N_17275,N_17547);
and U18146 (N_18146,N_16905,N_17432);
nand U18147 (N_18147,N_16849,N_16867);
xnor U18148 (N_18148,N_17562,N_17297);
or U18149 (N_18149,N_17277,N_17185);
nor U18150 (N_18150,N_17339,N_17185);
nand U18151 (N_18151,N_17110,N_17117);
nor U18152 (N_18152,N_16880,N_17287);
nor U18153 (N_18153,N_17473,N_17423);
nor U18154 (N_18154,N_17406,N_16875);
nor U18155 (N_18155,N_17315,N_16927);
or U18156 (N_18156,N_17019,N_16935);
xor U18157 (N_18157,N_17570,N_17589);
nand U18158 (N_18158,N_17330,N_16837);
nand U18159 (N_18159,N_16851,N_16914);
and U18160 (N_18160,N_17024,N_17406);
and U18161 (N_18161,N_17109,N_16835);
xor U18162 (N_18162,N_17292,N_16871);
nor U18163 (N_18163,N_17475,N_16866);
xor U18164 (N_18164,N_17510,N_17076);
nand U18165 (N_18165,N_17334,N_17443);
or U18166 (N_18166,N_17065,N_17359);
or U18167 (N_18167,N_16925,N_17111);
nor U18168 (N_18168,N_16859,N_16964);
nor U18169 (N_18169,N_17396,N_17174);
xor U18170 (N_18170,N_17265,N_17432);
and U18171 (N_18171,N_17220,N_17277);
or U18172 (N_18172,N_17208,N_17288);
nor U18173 (N_18173,N_16861,N_17591);
or U18174 (N_18174,N_17296,N_16833);
nor U18175 (N_18175,N_17295,N_17440);
nand U18176 (N_18176,N_17399,N_17378);
xor U18177 (N_18177,N_17348,N_16897);
nor U18178 (N_18178,N_17033,N_17183);
and U18179 (N_18179,N_17525,N_17459);
xor U18180 (N_18180,N_16808,N_17473);
xor U18181 (N_18181,N_17405,N_16974);
or U18182 (N_18182,N_17316,N_17065);
nor U18183 (N_18183,N_17320,N_17181);
or U18184 (N_18184,N_17292,N_17233);
xnor U18185 (N_18185,N_17014,N_17324);
nand U18186 (N_18186,N_17449,N_17534);
and U18187 (N_18187,N_17442,N_16970);
nor U18188 (N_18188,N_17308,N_17399);
and U18189 (N_18189,N_17390,N_16898);
nor U18190 (N_18190,N_17210,N_17430);
nor U18191 (N_18191,N_17410,N_17255);
nand U18192 (N_18192,N_17240,N_17506);
xnor U18193 (N_18193,N_17381,N_16859);
nand U18194 (N_18194,N_17072,N_17034);
xnor U18195 (N_18195,N_16846,N_17219);
xor U18196 (N_18196,N_17159,N_17234);
nor U18197 (N_18197,N_17308,N_17278);
xnor U18198 (N_18198,N_17375,N_17317);
or U18199 (N_18199,N_17429,N_17171);
nand U18200 (N_18200,N_16850,N_17264);
xor U18201 (N_18201,N_16970,N_16809);
xnor U18202 (N_18202,N_17051,N_17556);
or U18203 (N_18203,N_17180,N_16975);
xnor U18204 (N_18204,N_17211,N_17290);
or U18205 (N_18205,N_17190,N_16852);
nand U18206 (N_18206,N_17519,N_17443);
nand U18207 (N_18207,N_16877,N_17500);
and U18208 (N_18208,N_17418,N_17416);
nand U18209 (N_18209,N_17447,N_17153);
nor U18210 (N_18210,N_17037,N_17060);
or U18211 (N_18211,N_16859,N_17338);
nand U18212 (N_18212,N_16872,N_16878);
nor U18213 (N_18213,N_17191,N_17500);
xor U18214 (N_18214,N_17251,N_17163);
or U18215 (N_18215,N_16987,N_17067);
or U18216 (N_18216,N_17270,N_17061);
nor U18217 (N_18217,N_17155,N_17539);
nor U18218 (N_18218,N_17574,N_17428);
and U18219 (N_18219,N_16958,N_16869);
and U18220 (N_18220,N_17463,N_17572);
nor U18221 (N_18221,N_16861,N_17342);
nor U18222 (N_18222,N_16961,N_17348);
or U18223 (N_18223,N_17347,N_16966);
or U18224 (N_18224,N_17346,N_17427);
nor U18225 (N_18225,N_16810,N_17280);
and U18226 (N_18226,N_16875,N_16905);
nand U18227 (N_18227,N_17131,N_17285);
nand U18228 (N_18228,N_17566,N_17309);
and U18229 (N_18229,N_17401,N_17307);
xor U18230 (N_18230,N_17116,N_17572);
or U18231 (N_18231,N_17495,N_16924);
or U18232 (N_18232,N_17315,N_16970);
and U18233 (N_18233,N_17418,N_17216);
and U18234 (N_18234,N_17225,N_17313);
xor U18235 (N_18235,N_16884,N_17121);
or U18236 (N_18236,N_17142,N_16922);
and U18237 (N_18237,N_17387,N_17032);
or U18238 (N_18238,N_17571,N_17090);
or U18239 (N_18239,N_17307,N_16998);
xnor U18240 (N_18240,N_17025,N_17260);
nand U18241 (N_18241,N_17341,N_17458);
and U18242 (N_18242,N_17435,N_17542);
and U18243 (N_18243,N_16923,N_16920);
or U18244 (N_18244,N_17145,N_17389);
and U18245 (N_18245,N_17536,N_17362);
nor U18246 (N_18246,N_17106,N_17297);
nand U18247 (N_18247,N_16917,N_17578);
or U18248 (N_18248,N_17283,N_17265);
or U18249 (N_18249,N_17377,N_17147);
nand U18250 (N_18250,N_17001,N_17456);
nor U18251 (N_18251,N_17149,N_17329);
nor U18252 (N_18252,N_17127,N_16819);
or U18253 (N_18253,N_17349,N_17126);
and U18254 (N_18254,N_17201,N_17339);
nor U18255 (N_18255,N_17476,N_17399);
nand U18256 (N_18256,N_17270,N_17389);
and U18257 (N_18257,N_16938,N_17376);
nor U18258 (N_18258,N_17258,N_17122);
and U18259 (N_18259,N_16935,N_16900);
xnor U18260 (N_18260,N_17494,N_16879);
and U18261 (N_18261,N_17036,N_17541);
and U18262 (N_18262,N_17180,N_16839);
xnor U18263 (N_18263,N_17482,N_16958);
nand U18264 (N_18264,N_17057,N_17533);
and U18265 (N_18265,N_17543,N_17238);
and U18266 (N_18266,N_17172,N_17481);
nand U18267 (N_18267,N_17308,N_17129);
xor U18268 (N_18268,N_17530,N_17243);
and U18269 (N_18269,N_16912,N_17591);
or U18270 (N_18270,N_17140,N_16950);
or U18271 (N_18271,N_17138,N_17123);
or U18272 (N_18272,N_16900,N_16990);
nand U18273 (N_18273,N_16969,N_17020);
xnor U18274 (N_18274,N_17492,N_16896);
nor U18275 (N_18275,N_17323,N_17173);
xor U18276 (N_18276,N_17512,N_17074);
nand U18277 (N_18277,N_16928,N_17151);
and U18278 (N_18278,N_17033,N_16968);
nor U18279 (N_18279,N_16864,N_17430);
xnor U18280 (N_18280,N_17145,N_17056);
nor U18281 (N_18281,N_17185,N_17156);
or U18282 (N_18282,N_16894,N_17066);
nand U18283 (N_18283,N_17202,N_17257);
nor U18284 (N_18284,N_17387,N_16912);
nor U18285 (N_18285,N_17348,N_16884);
nand U18286 (N_18286,N_17081,N_17019);
or U18287 (N_18287,N_16993,N_17239);
xnor U18288 (N_18288,N_17172,N_17405);
or U18289 (N_18289,N_17366,N_17224);
xnor U18290 (N_18290,N_16959,N_17125);
xor U18291 (N_18291,N_17560,N_16897);
nor U18292 (N_18292,N_16952,N_17014);
or U18293 (N_18293,N_17300,N_16800);
nor U18294 (N_18294,N_17128,N_16840);
nor U18295 (N_18295,N_17269,N_17359);
xnor U18296 (N_18296,N_17129,N_16952);
nand U18297 (N_18297,N_16842,N_17307);
and U18298 (N_18298,N_17089,N_17024);
nand U18299 (N_18299,N_17231,N_17543);
xnor U18300 (N_18300,N_17188,N_17237);
and U18301 (N_18301,N_17016,N_17406);
nor U18302 (N_18302,N_17217,N_17457);
xor U18303 (N_18303,N_17008,N_16810);
xnor U18304 (N_18304,N_17195,N_16853);
or U18305 (N_18305,N_17268,N_17370);
and U18306 (N_18306,N_17547,N_17284);
nor U18307 (N_18307,N_16829,N_17101);
xor U18308 (N_18308,N_17028,N_17084);
or U18309 (N_18309,N_17593,N_17051);
nand U18310 (N_18310,N_17264,N_17468);
nand U18311 (N_18311,N_17468,N_17269);
nor U18312 (N_18312,N_17428,N_17044);
or U18313 (N_18313,N_17219,N_17529);
or U18314 (N_18314,N_17525,N_17559);
nand U18315 (N_18315,N_17540,N_17353);
nand U18316 (N_18316,N_17459,N_17563);
nand U18317 (N_18317,N_17131,N_17140);
nand U18318 (N_18318,N_17592,N_17473);
and U18319 (N_18319,N_17372,N_16861);
nor U18320 (N_18320,N_16954,N_17326);
or U18321 (N_18321,N_17127,N_17399);
nor U18322 (N_18322,N_17523,N_17118);
xor U18323 (N_18323,N_17157,N_17061);
or U18324 (N_18324,N_17574,N_17041);
xnor U18325 (N_18325,N_17314,N_17582);
nor U18326 (N_18326,N_16959,N_17108);
nor U18327 (N_18327,N_17427,N_16934);
nand U18328 (N_18328,N_17499,N_17216);
and U18329 (N_18329,N_17198,N_17502);
or U18330 (N_18330,N_17210,N_17005);
nor U18331 (N_18331,N_17145,N_17249);
nand U18332 (N_18332,N_17022,N_17514);
xnor U18333 (N_18333,N_17070,N_17062);
nor U18334 (N_18334,N_17246,N_17326);
nor U18335 (N_18335,N_16852,N_17587);
xnor U18336 (N_18336,N_17291,N_17452);
nand U18337 (N_18337,N_17293,N_16833);
or U18338 (N_18338,N_17047,N_17103);
and U18339 (N_18339,N_17527,N_17556);
nand U18340 (N_18340,N_16917,N_17226);
nand U18341 (N_18341,N_17261,N_16801);
or U18342 (N_18342,N_17003,N_17497);
or U18343 (N_18343,N_17024,N_17295);
nand U18344 (N_18344,N_17237,N_17596);
xnor U18345 (N_18345,N_17323,N_17326);
and U18346 (N_18346,N_17435,N_16837);
or U18347 (N_18347,N_16827,N_17280);
nand U18348 (N_18348,N_17303,N_16819);
nor U18349 (N_18349,N_16986,N_17246);
xnor U18350 (N_18350,N_16848,N_17436);
xnor U18351 (N_18351,N_16892,N_17572);
or U18352 (N_18352,N_17211,N_17450);
nor U18353 (N_18353,N_17300,N_17251);
nand U18354 (N_18354,N_17369,N_17059);
nor U18355 (N_18355,N_17005,N_17206);
nor U18356 (N_18356,N_16988,N_17319);
xnor U18357 (N_18357,N_17404,N_17347);
or U18358 (N_18358,N_17206,N_17127);
or U18359 (N_18359,N_17003,N_17004);
xnor U18360 (N_18360,N_17298,N_16856);
nor U18361 (N_18361,N_16995,N_16817);
xor U18362 (N_18362,N_17196,N_17268);
and U18363 (N_18363,N_17168,N_17245);
xnor U18364 (N_18364,N_17414,N_17080);
and U18365 (N_18365,N_17347,N_17452);
or U18366 (N_18366,N_17438,N_17291);
xnor U18367 (N_18367,N_16995,N_17353);
and U18368 (N_18368,N_17094,N_17347);
xnor U18369 (N_18369,N_16974,N_17100);
nand U18370 (N_18370,N_17300,N_16904);
and U18371 (N_18371,N_17091,N_17544);
xnor U18372 (N_18372,N_17458,N_17079);
nand U18373 (N_18373,N_17260,N_17166);
or U18374 (N_18374,N_16868,N_16918);
nand U18375 (N_18375,N_16844,N_17105);
xnor U18376 (N_18376,N_17125,N_17134);
nand U18377 (N_18377,N_16898,N_17586);
and U18378 (N_18378,N_17565,N_16864);
or U18379 (N_18379,N_16849,N_17374);
or U18380 (N_18380,N_16993,N_16850);
nor U18381 (N_18381,N_17115,N_16991);
nand U18382 (N_18382,N_17045,N_16943);
and U18383 (N_18383,N_17431,N_17298);
and U18384 (N_18384,N_17521,N_16913);
or U18385 (N_18385,N_17100,N_17512);
or U18386 (N_18386,N_16863,N_16825);
nand U18387 (N_18387,N_17540,N_17396);
nor U18388 (N_18388,N_17211,N_17344);
or U18389 (N_18389,N_17099,N_17284);
and U18390 (N_18390,N_17179,N_16804);
or U18391 (N_18391,N_17525,N_17124);
nand U18392 (N_18392,N_17322,N_17530);
nand U18393 (N_18393,N_17171,N_16868);
or U18394 (N_18394,N_16840,N_16949);
xor U18395 (N_18395,N_16872,N_17302);
and U18396 (N_18396,N_16997,N_17508);
and U18397 (N_18397,N_17387,N_16972);
nor U18398 (N_18398,N_17398,N_17516);
or U18399 (N_18399,N_17265,N_17488);
nor U18400 (N_18400,N_18169,N_18216);
or U18401 (N_18401,N_17632,N_17733);
and U18402 (N_18402,N_18171,N_18243);
xor U18403 (N_18403,N_18362,N_18217);
and U18404 (N_18404,N_17824,N_18020);
nor U18405 (N_18405,N_17999,N_17896);
xor U18406 (N_18406,N_18140,N_17814);
xor U18407 (N_18407,N_18221,N_18040);
xnor U18408 (N_18408,N_18261,N_17683);
nand U18409 (N_18409,N_18110,N_17688);
xor U18410 (N_18410,N_18085,N_17846);
xnor U18411 (N_18411,N_17936,N_18181);
nand U18412 (N_18412,N_17926,N_18297);
nor U18413 (N_18413,N_18229,N_18190);
nand U18414 (N_18414,N_17704,N_18349);
and U18415 (N_18415,N_17728,N_18245);
xnor U18416 (N_18416,N_18026,N_17665);
and U18417 (N_18417,N_17785,N_17608);
or U18418 (N_18418,N_18271,N_18149);
xnor U18419 (N_18419,N_17695,N_17701);
nand U18420 (N_18420,N_18316,N_18058);
and U18421 (N_18421,N_18351,N_18253);
or U18422 (N_18422,N_17861,N_17744);
nor U18423 (N_18423,N_18055,N_18301);
xnor U18424 (N_18424,N_18017,N_18003);
or U18425 (N_18425,N_17952,N_18379);
and U18426 (N_18426,N_18376,N_18339);
and U18427 (N_18427,N_17789,N_18274);
or U18428 (N_18428,N_18014,N_18074);
nand U18429 (N_18429,N_18062,N_18302);
xnor U18430 (N_18430,N_17985,N_18358);
or U18431 (N_18431,N_18136,N_17800);
or U18432 (N_18432,N_17768,N_18178);
or U18433 (N_18433,N_18272,N_18319);
and U18434 (N_18434,N_17867,N_18044);
or U18435 (N_18435,N_18355,N_18115);
xor U18436 (N_18436,N_18341,N_18329);
or U18437 (N_18437,N_18255,N_18118);
and U18438 (N_18438,N_17812,N_18126);
xnor U18439 (N_18439,N_17663,N_18384);
nor U18440 (N_18440,N_18093,N_17705);
nor U18441 (N_18441,N_17901,N_18252);
or U18442 (N_18442,N_17965,N_17652);
nor U18443 (N_18443,N_18158,N_18005);
and U18444 (N_18444,N_17983,N_18064);
xor U18445 (N_18445,N_17915,N_18346);
and U18446 (N_18446,N_18097,N_17657);
or U18447 (N_18447,N_17868,N_18095);
nand U18448 (N_18448,N_18056,N_17754);
nand U18449 (N_18449,N_18264,N_18233);
xnor U18450 (N_18450,N_18087,N_17621);
nor U18451 (N_18451,N_18324,N_17964);
nor U18452 (N_18452,N_17892,N_17942);
or U18453 (N_18453,N_17816,N_17932);
xnor U18454 (N_18454,N_18286,N_17805);
and U18455 (N_18455,N_18353,N_17874);
xnor U18456 (N_18456,N_18021,N_17628);
or U18457 (N_18457,N_17742,N_18084);
nor U18458 (N_18458,N_17832,N_18198);
and U18459 (N_18459,N_17614,N_17623);
or U18460 (N_18460,N_18010,N_18065);
or U18461 (N_18461,N_17651,N_17792);
nor U18462 (N_18462,N_17869,N_17976);
or U18463 (N_18463,N_18340,N_18183);
nor U18464 (N_18464,N_17801,N_18269);
nor U18465 (N_18465,N_17904,N_18080);
xor U18466 (N_18466,N_17927,N_18082);
and U18467 (N_18467,N_18090,N_17756);
nand U18468 (N_18468,N_17712,N_18049);
nor U18469 (N_18469,N_18153,N_17931);
or U18470 (N_18470,N_17817,N_17618);
and U18471 (N_18471,N_17856,N_17886);
and U18472 (N_18472,N_17827,N_17626);
or U18473 (N_18473,N_17882,N_18394);
or U18474 (N_18474,N_17899,N_17716);
and U18475 (N_18475,N_18027,N_18280);
and U18476 (N_18476,N_18342,N_17720);
xor U18477 (N_18477,N_18235,N_17837);
or U18478 (N_18478,N_18392,N_17982);
xor U18479 (N_18479,N_18310,N_17786);
or U18480 (N_18480,N_18388,N_17831);
or U18481 (N_18481,N_18207,N_17708);
nand U18482 (N_18482,N_17828,N_18213);
xor U18483 (N_18483,N_17668,N_18244);
or U18484 (N_18484,N_17951,N_18038);
nor U18485 (N_18485,N_18396,N_18336);
nor U18486 (N_18486,N_17759,N_18367);
nand U18487 (N_18487,N_17803,N_18188);
or U18488 (N_18488,N_17878,N_18291);
and U18489 (N_18489,N_18222,N_18295);
xor U18490 (N_18490,N_17694,N_17909);
nor U18491 (N_18491,N_18385,N_17966);
and U18492 (N_18492,N_18315,N_17881);
nor U18493 (N_18493,N_18120,N_18366);
xnor U18494 (N_18494,N_18175,N_18139);
or U18495 (N_18495,N_17737,N_18210);
or U18496 (N_18496,N_18164,N_18125);
and U18497 (N_18497,N_17641,N_18386);
and U18498 (N_18498,N_17611,N_17911);
xnor U18499 (N_18499,N_17834,N_17849);
xnor U18500 (N_18500,N_17962,N_17703);
xor U18501 (N_18501,N_18240,N_18347);
xor U18502 (N_18502,N_17609,N_18278);
or U18503 (N_18503,N_18364,N_17760);
nand U18504 (N_18504,N_18144,N_18287);
and U18505 (N_18505,N_17889,N_18042);
nand U18506 (N_18506,N_17898,N_18022);
nand U18507 (N_18507,N_17808,N_18398);
and U18508 (N_18508,N_17725,N_17675);
or U18509 (N_18509,N_17635,N_18006);
nor U18510 (N_18510,N_17729,N_17910);
nand U18511 (N_18511,N_17689,N_17758);
nor U18512 (N_18512,N_18063,N_17813);
nor U18513 (N_18513,N_17988,N_17863);
or U18514 (N_18514,N_17778,N_18201);
nor U18515 (N_18515,N_17699,N_18350);
and U18516 (N_18516,N_17627,N_17859);
xor U18517 (N_18517,N_18079,N_18303);
nand U18518 (N_18518,N_17606,N_17843);
nor U18519 (N_18519,N_18224,N_17876);
or U18520 (N_18520,N_18104,N_18094);
xnor U18521 (N_18521,N_18275,N_17607);
nand U18522 (N_18522,N_18263,N_17745);
nand U18523 (N_18523,N_18039,N_18226);
and U18524 (N_18524,N_17809,N_17929);
and U18525 (N_18525,N_17616,N_17762);
and U18526 (N_18526,N_18293,N_17887);
and U18527 (N_18527,N_17734,N_17866);
or U18528 (N_18528,N_17921,N_17724);
and U18529 (N_18529,N_17862,N_17950);
nand U18530 (N_18530,N_18135,N_18331);
xnor U18531 (N_18531,N_17707,N_17885);
and U18532 (N_18532,N_18161,N_17902);
nand U18533 (N_18533,N_17897,N_17860);
and U18534 (N_18534,N_18051,N_18184);
nand U18535 (N_18535,N_17642,N_18177);
xor U18536 (N_18536,N_18028,N_18231);
nand U18537 (N_18537,N_18185,N_17600);
or U18538 (N_18538,N_18260,N_17907);
nor U18539 (N_18539,N_18061,N_17877);
nand U18540 (N_18540,N_17997,N_18209);
nor U18541 (N_18541,N_18053,N_17661);
nor U18542 (N_18542,N_18036,N_18294);
and U18543 (N_18543,N_18202,N_17957);
xor U18544 (N_18544,N_17680,N_18312);
or U18545 (N_18545,N_18156,N_18223);
or U18546 (N_18546,N_17920,N_17947);
or U18547 (N_18547,N_18111,N_17736);
nand U18548 (N_18548,N_17978,N_18119);
xor U18549 (N_18549,N_17631,N_17949);
or U18550 (N_18550,N_17672,N_18361);
and U18551 (N_18551,N_17650,N_17646);
and U18552 (N_18552,N_17740,N_17969);
nand U18553 (N_18553,N_18254,N_17836);
or U18554 (N_18554,N_18047,N_17908);
nand U18555 (N_18555,N_17996,N_17620);
nor U18556 (N_18556,N_18335,N_17658);
nand U18557 (N_18557,N_17764,N_18321);
and U18558 (N_18558,N_18377,N_18008);
xnor U18559 (N_18559,N_18208,N_18220);
nand U18560 (N_18560,N_17622,N_18289);
or U18561 (N_18561,N_18290,N_18155);
or U18562 (N_18562,N_17664,N_17682);
xor U18563 (N_18563,N_18241,N_18001);
xor U18564 (N_18564,N_18389,N_17829);
or U18565 (N_18565,N_18091,N_18180);
and U18566 (N_18566,N_18138,N_18197);
or U18567 (N_18567,N_18101,N_17763);
nand U18568 (N_18568,N_17780,N_17633);
and U18569 (N_18569,N_18107,N_18296);
xnor U18570 (N_18570,N_18334,N_17925);
and U18571 (N_18571,N_18071,N_17841);
and U18572 (N_18572,N_18285,N_18162);
nand U18573 (N_18573,N_17835,N_18133);
xnor U18574 (N_18574,N_18193,N_18311);
or U18575 (N_18575,N_17933,N_17944);
or U18576 (N_18576,N_17612,N_18251);
or U18577 (N_18577,N_18299,N_17706);
and U18578 (N_18578,N_17640,N_17795);
xor U18579 (N_18579,N_17986,N_18313);
and U18580 (N_18580,N_17830,N_18363);
and U18581 (N_18581,N_17719,N_17750);
or U18582 (N_18582,N_18189,N_18373);
nand U18583 (N_18583,N_18219,N_17919);
or U18584 (N_18584,N_17891,N_18106);
and U18585 (N_18585,N_17766,N_18077);
and U18586 (N_18586,N_18117,N_17603);
or U18587 (N_18587,N_17938,N_17960);
xnor U18588 (N_18588,N_18121,N_18371);
nor U18589 (N_18589,N_17848,N_17974);
xnor U18590 (N_18590,N_18069,N_17654);
or U18591 (N_18591,N_18168,N_17653);
xor U18592 (N_18592,N_18279,N_18143);
and U18593 (N_18593,N_17687,N_18011);
nor U18594 (N_18594,N_17784,N_18113);
xnor U18595 (N_18595,N_18199,N_17845);
and U18596 (N_18596,N_18035,N_18160);
or U18597 (N_18597,N_17840,N_18212);
nor U18598 (N_18598,N_18249,N_17604);
nand U18599 (N_18599,N_17782,N_17906);
nor U18600 (N_18600,N_18200,N_18018);
xnor U18601 (N_18601,N_17779,N_17787);
nand U18602 (N_18602,N_18309,N_18002);
or U18603 (N_18603,N_17850,N_17857);
or U18604 (N_18604,N_18086,N_18354);
nand U18605 (N_18605,N_17940,N_17970);
nand U18606 (N_18606,N_17751,N_18023);
xnor U18607 (N_18607,N_17659,N_18328);
or U18608 (N_18608,N_18259,N_18081);
xnor U18609 (N_18609,N_17799,N_17732);
nor U18610 (N_18610,N_17959,N_18151);
nor U18611 (N_18611,N_18172,N_17711);
nor U18612 (N_18612,N_18228,N_17776);
or U18613 (N_18613,N_18048,N_17772);
nand U18614 (N_18614,N_17775,N_18397);
nor U18615 (N_18615,N_17637,N_18214);
or U18616 (N_18616,N_17718,N_17880);
xor U18617 (N_18617,N_18225,N_17854);
xnor U18618 (N_18618,N_18330,N_17710);
or U18619 (N_18619,N_18173,N_17990);
nor U18620 (N_18620,N_17993,N_17773);
xnor U18621 (N_18621,N_18131,N_18196);
xor U18622 (N_18622,N_17922,N_17864);
nand U18623 (N_18623,N_17791,N_18165);
nand U18624 (N_18624,N_17987,N_17774);
nor U18625 (N_18625,N_18195,N_17771);
xnor U18626 (N_18626,N_18248,N_18194);
or U18627 (N_18627,N_17994,N_18325);
and U18628 (N_18628,N_18268,N_18075);
or U18629 (N_18629,N_18060,N_18134);
nor U18630 (N_18630,N_18032,N_17871);
and U18631 (N_18631,N_17660,N_17858);
or U18632 (N_18632,N_17681,N_18045);
xor U18633 (N_18633,N_18378,N_17671);
or U18634 (N_18634,N_18357,N_17722);
nor U18635 (N_18635,N_17638,N_18232);
and U18636 (N_18636,N_17666,N_17980);
nor U18637 (N_18637,N_18145,N_18154);
or U18638 (N_18638,N_18258,N_18150);
nor U18639 (N_18639,N_18344,N_17998);
or U18640 (N_18640,N_17713,N_17781);
xor U18641 (N_18641,N_17662,N_17839);
or U18642 (N_18642,N_17798,N_17746);
xnor U18643 (N_18643,N_18393,N_17818);
nand U18644 (N_18644,N_18015,N_17731);
xor U18645 (N_18645,N_18345,N_17967);
nor U18646 (N_18646,N_18163,N_18083);
xnor U18647 (N_18647,N_17679,N_17639);
xnor U18648 (N_18648,N_17793,N_17648);
and U18649 (N_18649,N_18218,N_18267);
nand U18650 (N_18650,N_17916,N_17804);
nor U18651 (N_18651,N_18326,N_18012);
or U18652 (N_18652,N_17924,N_17930);
xnor U18653 (N_18653,N_17678,N_17879);
and U18654 (N_18654,N_17625,N_17697);
or U18655 (N_18655,N_18307,N_17749);
and U18656 (N_18656,N_18333,N_17643);
nand U18657 (N_18657,N_18382,N_18170);
xor U18658 (N_18658,N_18332,N_18265);
nor U18659 (N_18659,N_17790,N_17700);
nand U18660 (N_18660,N_17847,N_17890);
xor U18661 (N_18661,N_18375,N_17823);
or U18662 (N_18662,N_17945,N_17844);
nor U18663 (N_18663,N_17755,N_17698);
nand U18664 (N_18664,N_18009,N_17702);
and U18665 (N_18665,N_18356,N_18322);
xor U18666 (N_18666,N_18211,N_17709);
or U18667 (N_18667,N_17838,N_17610);
nand U18668 (N_18668,N_18318,N_18387);
and U18669 (N_18669,N_17788,N_17870);
nor U18670 (N_18670,N_17872,N_18352);
or U18671 (N_18671,N_18266,N_17972);
xor U18672 (N_18672,N_18054,N_17636);
and U18673 (N_18673,N_18227,N_18238);
nand U18674 (N_18674,N_17981,N_18108);
nor U18675 (N_18675,N_18277,N_17963);
nor U18676 (N_18676,N_18298,N_18147);
and U18677 (N_18677,N_18176,N_17802);
and U18678 (N_18678,N_18076,N_17842);
or U18679 (N_18679,N_17696,N_18338);
and U18680 (N_18680,N_18380,N_18152);
xor U18681 (N_18681,N_18100,N_17973);
nor U18682 (N_18682,N_18166,N_18007);
xor U18683 (N_18683,N_18281,N_18369);
nor U18684 (N_18684,N_17723,N_18236);
nor U18685 (N_18685,N_18098,N_17943);
and U18686 (N_18686,N_17748,N_17649);
xnor U18687 (N_18687,N_17958,N_18034);
nand U18688 (N_18688,N_17677,N_18174);
or U18689 (N_18689,N_17691,N_17743);
nor U18690 (N_18690,N_17810,N_17955);
nor U18691 (N_18691,N_18073,N_18057);
and U18692 (N_18692,N_18317,N_18146);
nor U18693 (N_18693,N_18046,N_17634);
xnor U18694 (N_18694,N_17995,N_17865);
nor U18695 (N_18695,N_18025,N_18206);
nand U18696 (N_18696,N_17815,N_18204);
xor U18697 (N_18697,N_18368,N_18099);
or U18698 (N_18698,N_18041,N_17777);
nor U18699 (N_18699,N_18270,N_18273);
or U18700 (N_18700,N_17806,N_17769);
and U18701 (N_18701,N_17893,N_18129);
nand U18702 (N_18702,N_17797,N_17819);
or U18703 (N_18703,N_18300,N_18381);
xor U18704 (N_18704,N_17615,N_18159);
nand U18705 (N_18705,N_17912,N_18128);
xor U18706 (N_18706,N_17820,N_18096);
and U18707 (N_18707,N_18246,N_18066);
or U18708 (N_18708,N_17613,N_18102);
and U18709 (N_18709,N_18360,N_17968);
nand U18710 (N_18710,N_17647,N_18130);
nor U18711 (N_18711,N_18019,N_17913);
and U18712 (N_18712,N_17601,N_17852);
nand U18713 (N_18713,N_17727,N_17655);
xnor U18714 (N_18714,N_17726,N_18395);
xnor U18715 (N_18715,N_17914,N_17602);
xor U18716 (N_18716,N_17753,N_17741);
nand U18717 (N_18717,N_17630,N_18304);
nand U18718 (N_18718,N_18004,N_18239);
or U18719 (N_18719,N_18372,N_17923);
nor U18720 (N_18720,N_17989,N_18112);
and U18721 (N_18721,N_18203,N_18276);
nor U18722 (N_18722,N_17939,N_18391);
and U18723 (N_18723,N_18124,N_18186);
nor U18724 (N_18724,N_18359,N_18070);
or U18725 (N_18725,N_18013,N_17822);
xnor U18726 (N_18726,N_17605,N_18037);
nand U18727 (N_18727,N_18029,N_17783);
and U18728 (N_18728,N_18247,N_17961);
or U18729 (N_18729,N_18050,N_18192);
and U18730 (N_18730,N_18284,N_18103);
nor U18731 (N_18731,N_17676,N_17757);
and U18732 (N_18732,N_18283,N_18399);
nor U18733 (N_18733,N_17629,N_18142);
xnor U18734 (N_18734,N_18365,N_18191);
xor U18735 (N_18735,N_18157,N_17888);
xnor U18736 (N_18736,N_17935,N_17948);
nor U18737 (N_18737,N_18242,N_18257);
nor U18738 (N_18738,N_17794,N_17807);
nor U18739 (N_18739,N_17934,N_17883);
xnor U18740 (N_18740,N_18337,N_18105);
xnor U18741 (N_18741,N_17903,N_17894);
and U18742 (N_18742,N_17667,N_18030);
nor U18743 (N_18743,N_17656,N_17624);
or U18744 (N_18744,N_18067,N_17941);
and U18745 (N_18745,N_18072,N_18282);
or U18746 (N_18746,N_17670,N_18320);
xnor U18747 (N_18747,N_18000,N_18343);
or U18748 (N_18748,N_17984,N_17685);
and U18749 (N_18749,N_18078,N_18089);
nand U18750 (N_18750,N_17692,N_17875);
xor U18751 (N_18751,N_18390,N_18137);
or U18752 (N_18752,N_17918,N_17991);
or U18753 (N_18753,N_18292,N_18323);
and U18754 (N_18754,N_17730,N_18088);
nor U18755 (N_18755,N_17953,N_18370);
nor U18756 (N_18756,N_18116,N_17992);
xor U18757 (N_18757,N_18031,N_17855);
nor U18758 (N_18758,N_18205,N_17767);
and U18759 (N_18759,N_17825,N_17645);
and U18760 (N_18760,N_18182,N_17674);
and U18761 (N_18761,N_17747,N_17715);
xor U18762 (N_18762,N_17796,N_17644);
nor U18763 (N_18763,N_18288,N_18237);
or U18764 (N_18764,N_18179,N_17619);
or U18765 (N_18765,N_17971,N_17905);
and U18766 (N_18766,N_18092,N_17954);
or U18767 (N_18767,N_17895,N_18230);
nor U18768 (N_18768,N_17693,N_18127);
xnor U18769 (N_18769,N_18109,N_17937);
xnor U18770 (N_18770,N_18141,N_17821);
or U18771 (N_18771,N_17690,N_17811);
nand U18772 (N_18772,N_18306,N_17617);
and U18773 (N_18773,N_17975,N_18016);
and U18774 (N_18774,N_18033,N_18024);
nor U18775 (N_18775,N_18167,N_18234);
and U18776 (N_18776,N_18250,N_17739);
and U18777 (N_18777,N_17686,N_18114);
nand U18778 (N_18778,N_17977,N_18052);
xor U18779 (N_18779,N_17917,N_17735);
and U18780 (N_18780,N_17714,N_17900);
nor U18781 (N_18781,N_18374,N_18327);
nand U18782 (N_18782,N_18059,N_18123);
or U18783 (N_18783,N_17928,N_17884);
nand U18784 (N_18784,N_17752,N_17956);
nand U18785 (N_18785,N_18314,N_17684);
and U18786 (N_18786,N_18256,N_18132);
xor U18787 (N_18787,N_17738,N_17853);
and U18788 (N_18788,N_18122,N_18187);
or U18789 (N_18789,N_17765,N_18148);
xnor U18790 (N_18790,N_17851,N_18348);
nand U18791 (N_18791,N_17833,N_17826);
and U18792 (N_18792,N_18308,N_18043);
and U18793 (N_18793,N_17669,N_18262);
nor U18794 (N_18794,N_17761,N_18068);
xor U18795 (N_18795,N_17979,N_17721);
xor U18796 (N_18796,N_17673,N_18383);
nor U18797 (N_18797,N_17717,N_17946);
nand U18798 (N_18798,N_17770,N_17873);
nor U18799 (N_18799,N_18215,N_18305);
nand U18800 (N_18800,N_17927,N_18122);
xor U18801 (N_18801,N_17691,N_17821);
nand U18802 (N_18802,N_18208,N_17636);
and U18803 (N_18803,N_18230,N_18019);
nor U18804 (N_18804,N_17787,N_17689);
or U18805 (N_18805,N_17966,N_18242);
nor U18806 (N_18806,N_17781,N_17665);
xor U18807 (N_18807,N_18208,N_18177);
and U18808 (N_18808,N_17983,N_18107);
and U18809 (N_18809,N_17824,N_17600);
xor U18810 (N_18810,N_18083,N_17662);
xnor U18811 (N_18811,N_18041,N_18249);
nand U18812 (N_18812,N_17907,N_17748);
and U18813 (N_18813,N_17992,N_18375);
xor U18814 (N_18814,N_18172,N_17984);
xor U18815 (N_18815,N_17707,N_18255);
nand U18816 (N_18816,N_18153,N_17942);
nor U18817 (N_18817,N_18277,N_17912);
and U18818 (N_18818,N_17864,N_18022);
and U18819 (N_18819,N_17614,N_18316);
or U18820 (N_18820,N_18121,N_17634);
and U18821 (N_18821,N_18095,N_18188);
and U18822 (N_18822,N_18297,N_17734);
and U18823 (N_18823,N_17631,N_17886);
and U18824 (N_18824,N_18239,N_17891);
xnor U18825 (N_18825,N_18023,N_18342);
and U18826 (N_18826,N_18213,N_17674);
nand U18827 (N_18827,N_17625,N_17947);
nor U18828 (N_18828,N_18378,N_18240);
nand U18829 (N_18829,N_18233,N_17738);
and U18830 (N_18830,N_17831,N_18070);
xnor U18831 (N_18831,N_17900,N_18337);
nor U18832 (N_18832,N_17712,N_17640);
xnor U18833 (N_18833,N_17612,N_17897);
nand U18834 (N_18834,N_17871,N_17911);
nand U18835 (N_18835,N_18367,N_18117);
xor U18836 (N_18836,N_18295,N_18011);
xor U18837 (N_18837,N_17657,N_17683);
or U18838 (N_18838,N_18377,N_18342);
or U18839 (N_18839,N_17962,N_17835);
and U18840 (N_18840,N_17697,N_18317);
nand U18841 (N_18841,N_18237,N_18172);
and U18842 (N_18842,N_18066,N_18337);
xor U18843 (N_18843,N_17804,N_17955);
and U18844 (N_18844,N_17916,N_17846);
and U18845 (N_18845,N_18207,N_17924);
or U18846 (N_18846,N_18054,N_18186);
or U18847 (N_18847,N_18275,N_17611);
or U18848 (N_18848,N_17783,N_18051);
nor U18849 (N_18849,N_17617,N_18365);
nand U18850 (N_18850,N_18226,N_18022);
or U18851 (N_18851,N_18384,N_18368);
nor U18852 (N_18852,N_17647,N_18075);
xnor U18853 (N_18853,N_17748,N_17918);
and U18854 (N_18854,N_17701,N_18359);
xor U18855 (N_18855,N_17630,N_18011);
nor U18856 (N_18856,N_17877,N_17882);
xor U18857 (N_18857,N_18050,N_17975);
nand U18858 (N_18858,N_18168,N_17884);
nand U18859 (N_18859,N_18365,N_18248);
xor U18860 (N_18860,N_17946,N_17654);
nand U18861 (N_18861,N_18060,N_18319);
xor U18862 (N_18862,N_18201,N_18084);
or U18863 (N_18863,N_18321,N_17901);
and U18864 (N_18864,N_18348,N_18269);
nor U18865 (N_18865,N_18233,N_18102);
or U18866 (N_18866,N_18384,N_17774);
nand U18867 (N_18867,N_18015,N_17640);
or U18868 (N_18868,N_17632,N_18293);
nand U18869 (N_18869,N_17635,N_17975);
and U18870 (N_18870,N_17910,N_17605);
nor U18871 (N_18871,N_18109,N_18135);
nand U18872 (N_18872,N_18174,N_17721);
nand U18873 (N_18873,N_17995,N_17849);
xnor U18874 (N_18874,N_18203,N_17642);
nand U18875 (N_18875,N_17655,N_17929);
or U18876 (N_18876,N_18331,N_18254);
and U18877 (N_18877,N_18200,N_17921);
and U18878 (N_18878,N_17605,N_17968);
or U18879 (N_18879,N_17731,N_17814);
or U18880 (N_18880,N_17999,N_18201);
nand U18881 (N_18881,N_17760,N_17623);
or U18882 (N_18882,N_17767,N_18004);
and U18883 (N_18883,N_18105,N_18395);
xor U18884 (N_18884,N_17617,N_18386);
or U18885 (N_18885,N_17744,N_17672);
nor U18886 (N_18886,N_17747,N_17616);
or U18887 (N_18887,N_18260,N_17970);
or U18888 (N_18888,N_17890,N_18336);
and U18889 (N_18889,N_18017,N_18101);
nor U18890 (N_18890,N_17773,N_18204);
or U18891 (N_18891,N_18179,N_18166);
and U18892 (N_18892,N_18153,N_18337);
or U18893 (N_18893,N_18148,N_18307);
or U18894 (N_18894,N_17824,N_17983);
or U18895 (N_18895,N_17987,N_18228);
and U18896 (N_18896,N_17708,N_17957);
nand U18897 (N_18897,N_18183,N_18399);
nor U18898 (N_18898,N_18284,N_18094);
or U18899 (N_18899,N_18154,N_18360);
nand U18900 (N_18900,N_18173,N_18115);
or U18901 (N_18901,N_18096,N_18293);
and U18902 (N_18902,N_18142,N_17734);
nor U18903 (N_18903,N_17993,N_17829);
nand U18904 (N_18904,N_17755,N_18202);
nand U18905 (N_18905,N_17617,N_18136);
nand U18906 (N_18906,N_17654,N_17950);
nor U18907 (N_18907,N_18195,N_17864);
and U18908 (N_18908,N_17935,N_17825);
xnor U18909 (N_18909,N_18293,N_17987);
nand U18910 (N_18910,N_18129,N_18076);
nand U18911 (N_18911,N_18326,N_18163);
or U18912 (N_18912,N_18103,N_18264);
xor U18913 (N_18913,N_17727,N_18024);
or U18914 (N_18914,N_18121,N_18342);
and U18915 (N_18915,N_18004,N_17744);
nor U18916 (N_18916,N_17935,N_17889);
nand U18917 (N_18917,N_17907,N_18042);
nand U18918 (N_18918,N_17891,N_17972);
and U18919 (N_18919,N_18226,N_18172);
xnor U18920 (N_18920,N_17775,N_18077);
nand U18921 (N_18921,N_17976,N_18009);
and U18922 (N_18922,N_18312,N_17961);
xor U18923 (N_18923,N_18177,N_17969);
nor U18924 (N_18924,N_18346,N_17951);
xnor U18925 (N_18925,N_17830,N_18158);
nand U18926 (N_18926,N_18346,N_18230);
or U18927 (N_18927,N_18352,N_17867);
xnor U18928 (N_18928,N_18300,N_18029);
nor U18929 (N_18929,N_17878,N_17703);
nor U18930 (N_18930,N_17936,N_18012);
nand U18931 (N_18931,N_17878,N_17852);
and U18932 (N_18932,N_17735,N_18013);
or U18933 (N_18933,N_18352,N_17821);
or U18934 (N_18934,N_17930,N_18009);
or U18935 (N_18935,N_17971,N_18322);
xnor U18936 (N_18936,N_17891,N_17729);
and U18937 (N_18937,N_17617,N_18359);
or U18938 (N_18938,N_18171,N_18248);
xnor U18939 (N_18939,N_18246,N_18271);
nor U18940 (N_18940,N_18269,N_18369);
nor U18941 (N_18941,N_17852,N_18031);
and U18942 (N_18942,N_18175,N_17635);
or U18943 (N_18943,N_17983,N_17720);
or U18944 (N_18944,N_18276,N_18360);
or U18945 (N_18945,N_18055,N_17997);
xnor U18946 (N_18946,N_17639,N_18327);
or U18947 (N_18947,N_17773,N_17965);
and U18948 (N_18948,N_17643,N_18151);
nor U18949 (N_18949,N_18080,N_17942);
nor U18950 (N_18950,N_17931,N_17613);
or U18951 (N_18951,N_17816,N_18187);
nand U18952 (N_18952,N_17993,N_17782);
nor U18953 (N_18953,N_17921,N_18184);
and U18954 (N_18954,N_18151,N_17677);
and U18955 (N_18955,N_18289,N_18182);
or U18956 (N_18956,N_17724,N_18316);
nand U18957 (N_18957,N_17615,N_17774);
nand U18958 (N_18958,N_18027,N_18242);
or U18959 (N_18959,N_17792,N_17950);
or U18960 (N_18960,N_18276,N_17882);
or U18961 (N_18961,N_17779,N_17925);
nand U18962 (N_18962,N_17911,N_17677);
and U18963 (N_18963,N_18038,N_17803);
xnor U18964 (N_18964,N_18328,N_18366);
and U18965 (N_18965,N_18117,N_18339);
nor U18966 (N_18966,N_18282,N_17938);
and U18967 (N_18967,N_18274,N_18073);
or U18968 (N_18968,N_18329,N_18318);
nor U18969 (N_18969,N_18335,N_17794);
nand U18970 (N_18970,N_17897,N_18387);
nor U18971 (N_18971,N_17929,N_17960);
nor U18972 (N_18972,N_17608,N_17839);
xnor U18973 (N_18973,N_18089,N_18377);
and U18974 (N_18974,N_17751,N_17952);
and U18975 (N_18975,N_17970,N_17724);
and U18976 (N_18976,N_17871,N_17778);
and U18977 (N_18977,N_18059,N_18205);
and U18978 (N_18978,N_17720,N_18369);
and U18979 (N_18979,N_18179,N_18268);
or U18980 (N_18980,N_18120,N_17698);
or U18981 (N_18981,N_18119,N_17754);
xor U18982 (N_18982,N_18216,N_17969);
nand U18983 (N_18983,N_18278,N_18073);
and U18984 (N_18984,N_17703,N_17964);
nand U18985 (N_18985,N_17914,N_17644);
xor U18986 (N_18986,N_18199,N_18173);
or U18987 (N_18987,N_18053,N_17782);
and U18988 (N_18988,N_18156,N_17789);
xor U18989 (N_18989,N_18109,N_17695);
and U18990 (N_18990,N_18124,N_17946);
or U18991 (N_18991,N_18270,N_18238);
nor U18992 (N_18992,N_18318,N_17700);
xnor U18993 (N_18993,N_17639,N_17689);
and U18994 (N_18994,N_17601,N_18205);
xor U18995 (N_18995,N_18232,N_18239);
and U18996 (N_18996,N_18164,N_18005);
or U18997 (N_18997,N_18229,N_18341);
or U18998 (N_18998,N_17632,N_17657);
or U18999 (N_18999,N_18298,N_18001);
or U19000 (N_19000,N_17976,N_18140);
xor U19001 (N_19001,N_18157,N_18139);
nand U19002 (N_19002,N_18277,N_17792);
nand U19003 (N_19003,N_18063,N_18061);
or U19004 (N_19004,N_18387,N_18106);
xnor U19005 (N_19005,N_17734,N_18319);
nor U19006 (N_19006,N_18104,N_17907);
xor U19007 (N_19007,N_18074,N_17824);
nand U19008 (N_19008,N_18160,N_18240);
xnor U19009 (N_19009,N_18317,N_18262);
xnor U19010 (N_19010,N_17924,N_17680);
nand U19011 (N_19011,N_17966,N_17832);
or U19012 (N_19012,N_18079,N_18399);
or U19013 (N_19013,N_17922,N_18036);
nor U19014 (N_19014,N_17752,N_17797);
and U19015 (N_19015,N_17841,N_17736);
nand U19016 (N_19016,N_18026,N_17617);
nor U19017 (N_19017,N_17753,N_17923);
nand U19018 (N_19018,N_18230,N_17743);
nand U19019 (N_19019,N_17796,N_17899);
or U19020 (N_19020,N_17867,N_18394);
nor U19021 (N_19021,N_18047,N_18061);
or U19022 (N_19022,N_17770,N_18344);
or U19023 (N_19023,N_18168,N_17898);
xor U19024 (N_19024,N_17856,N_17678);
and U19025 (N_19025,N_17637,N_18197);
and U19026 (N_19026,N_18357,N_18094);
nand U19027 (N_19027,N_17951,N_18347);
xor U19028 (N_19028,N_17780,N_18311);
nor U19029 (N_19029,N_17721,N_18206);
or U19030 (N_19030,N_17608,N_17813);
nand U19031 (N_19031,N_17682,N_18159);
nand U19032 (N_19032,N_18253,N_18069);
or U19033 (N_19033,N_17820,N_17617);
and U19034 (N_19034,N_18126,N_18218);
nand U19035 (N_19035,N_18224,N_17689);
and U19036 (N_19036,N_18078,N_17760);
xor U19037 (N_19037,N_18145,N_17740);
nor U19038 (N_19038,N_17942,N_17682);
and U19039 (N_19039,N_17986,N_17881);
and U19040 (N_19040,N_18109,N_18266);
nor U19041 (N_19041,N_18348,N_18174);
and U19042 (N_19042,N_17886,N_18138);
nand U19043 (N_19043,N_18034,N_17804);
nand U19044 (N_19044,N_18165,N_17992);
nor U19045 (N_19045,N_17675,N_18356);
xor U19046 (N_19046,N_18152,N_17688);
nand U19047 (N_19047,N_18392,N_17722);
nand U19048 (N_19048,N_18234,N_17790);
and U19049 (N_19049,N_18011,N_18100);
xor U19050 (N_19050,N_18060,N_18038);
or U19051 (N_19051,N_17834,N_17692);
nand U19052 (N_19052,N_18184,N_18012);
and U19053 (N_19053,N_18013,N_17692);
xor U19054 (N_19054,N_18353,N_17644);
nand U19055 (N_19055,N_18022,N_18326);
nand U19056 (N_19056,N_17719,N_18035);
xnor U19057 (N_19057,N_18338,N_17896);
xor U19058 (N_19058,N_17826,N_18270);
nand U19059 (N_19059,N_18068,N_17928);
nor U19060 (N_19060,N_17710,N_17926);
or U19061 (N_19061,N_17709,N_18163);
nor U19062 (N_19062,N_18307,N_18127);
nand U19063 (N_19063,N_17728,N_18279);
and U19064 (N_19064,N_18258,N_17622);
nand U19065 (N_19065,N_17940,N_18083);
xor U19066 (N_19066,N_17995,N_18282);
nand U19067 (N_19067,N_18333,N_18055);
nand U19068 (N_19068,N_18043,N_18230);
nor U19069 (N_19069,N_17938,N_18215);
nor U19070 (N_19070,N_18228,N_18224);
and U19071 (N_19071,N_17702,N_18384);
nand U19072 (N_19072,N_18263,N_17622);
and U19073 (N_19073,N_18199,N_17759);
nand U19074 (N_19074,N_18141,N_18137);
and U19075 (N_19075,N_17847,N_17866);
and U19076 (N_19076,N_18036,N_17749);
and U19077 (N_19077,N_17816,N_18323);
and U19078 (N_19078,N_17787,N_17730);
and U19079 (N_19079,N_17717,N_18298);
nor U19080 (N_19080,N_17990,N_18180);
xnor U19081 (N_19081,N_17799,N_17935);
and U19082 (N_19082,N_17711,N_17904);
xor U19083 (N_19083,N_17803,N_18243);
xnor U19084 (N_19084,N_17801,N_18035);
and U19085 (N_19085,N_18068,N_17667);
nor U19086 (N_19086,N_17703,N_18345);
nand U19087 (N_19087,N_17973,N_18147);
nor U19088 (N_19088,N_18362,N_18388);
or U19089 (N_19089,N_17880,N_18206);
nor U19090 (N_19090,N_18395,N_18283);
or U19091 (N_19091,N_17718,N_17910);
xor U19092 (N_19092,N_17767,N_17742);
and U19093 (N_19093,N_18056,N_18074);
nor U19094 (N_19094,N_17742,N_18077);
xor U19095 (N_19095,N_17817,N_17859);
nand U19096 (N_19096,N_17858,N_18197);
and U19097 (N_19097,N_18082,N_17999);
and U19098 (N_19098,N_18151,N_18383);
nand U19099 (N_19099,N_18251,N_17682);
nor U19100 (N_19100,N_18092,N_17729);
nand U19101 (N_19101,N_17986,N_17966);
and U19102 (N_19102,N_17792,N_17794);
nand U19103 (N_19103,N_18366,N_17934);
nand U19104 (N_19104,N_18334,N_17897);
or U19105 (N_19105,N_17612,N_18203);
or U19106 (N_19106,N_18030,N_18396);
nor U19107 (N_19107,N_17836,N_17912);
nand U19108 (N_19108,N_18207,N_18213);
xnor U19109 (N_19109,N_18340,N_17968);
nor U19110 (N_19110,N_17974,N_17810);
xnor U19111 (N_19111,N_18296,N_17855);
nor U19112 (N_19112,N_18341,N_17993);
or U19113 (N_19113,N_18088,N_18230);
and U19114 (N_19114,N_18206,N_17751);
nand U19115 (N_19115,N_17629,N_18235);
xor U19116 (N_19116,N_18092,N_17704);
or U19117 (N_19117,N_17909,N_18232);
or U19118 (N_19118,N_18333,N_17912);
xor U19119 (N_19119,N_17816,N_17742);
or U19120 (N_19120,N_18087,N_17775);
xnor U19121 (N_19121,N_18280,N_18318);
and U19122 (N_19122,N_17815,N_18038);
nor U19123 (N_19123,N_18388,N_17625);
and U19124 (N_19124,N_18242,N_17669);
or U19125 (N_19125,N_17616,N_17953);
xor U19126 (N_19126,N_17874,N_17656);
and U19127 (N_19127,N_18269,N_18144);
nor U19128 (N_19128,N_17714,N_18066);
or U19129 (N_19129,N_18173,N_17744);
nand U19130 (N_19130,N_17770,N_17988);
nand U19131 (N_19131,N_17948,N_17722);
and U19132 (N_19132,N_17950,N_18043);
nand U19133 (N_19133,N_17660,N_18032);
and U19134 (N_19134,N_17631,N_18245);
and U19135 (N_19135,N_18066,N_18234);
and U19136 (N_19136,N_17896,N_17826);
xnor U19137 (N_19137,N_17875,N_17668);
xor U19138 (N_19138,N_17750,N_18107);
nand U19139 (N_19139,N_18112,N_18093);
xor U19140 (N_19140,N_17761,N_17629);
xnor U19141 (N_19141,N_18051,N_18152);
or U19142 (N_19142,N_18396,N_17664);
or U19143 (N_19143,N_18362,N_18212);
xor U19144 (N_19144,N_17881,N_18164);
or U19145 (N_19145,N_18234,N_17822);
nor U19146 (N_19146,N_17682,N_18368);
nor U19147 (N_19147,N_17901,N_18187);
nand U19148 (N_19148,N_18067,N_18355);
xor U19149 (N_19149,N_18157,N_17769);
or U19150 (N_19150,N_17738,N_18138);
or U19151 (N_19151,N_17801,N_17872);
or U19152 (N_19152,N_17612,N_18191);
and U19153 (N_19153,N_18310,N_17872);
or U19154 (N_19154,N_18195,N_17807);
nor U19155 (N_19155,N_17652,N_18370);
nand U19156 (N_19156,N_18092,N_18073);
or U19157 (N_19157,N_18059,N_18054);
nor U19158 (N_19158,N_17758,N_18096);
nand U19159 (N_19159,N_17659,N_18086);
xor U19160 (N_19160,N_17627,N_17684);
or U19161 (N_19161,N_17973,N_18372);
or U19162 (N_19162,N_18150,N_17775);
and U19163 (N_19163,N_18154,N_18052);
nor U19164 (N_19164,N_17972,N_17744);
nor U19165 (N_19165,N_18078,N_17973);
or U19166 (N_19166,N_17759,N_18173);
and U19167 (N_19167,N_18347,N_17652);
xor U19168 (N_19168,N_17884,N_18011);
and U19169 (N_19169,N_17646,N_18012);
and U19170 (N_19170,N_18073,N_17888);
and U19171 (N_19171,N_17895,N_18174);
and U19172 (N_19172,N_18219,N_18039);
nor U19173 (N_19173,N_17697,N_18166);
and U19174 (N_19174,N_18199,N_18317);
xor U19175 (N_19175,N_18164,N_18112);
or U19176 (N_19176,N_17905,N_17816);
nand U19177 (N_19177,N_17637,N_17627);
nand U19178 (N_19178,N_17983,N_18353);
xnor U19179 (N_19179,N_18116,N_17921);
and U19180 (N_19180,N_17939,N_17788);
and U19181 (N_19181,N_18047,N_18354);
nor U19182 (N_19182,N_18000,N_17763);
or U19183 (N_19183,N_18120,N_17768);
xnor U19184 (N_19184,N_18353,N_18187);
nand U19185 (N_19185,N_18112,N_18204);
nand U19186 (N_19186,N_18021,N_18264);
xor U19187 (N_19187,N_18270,N_17991);
nor U19188 (N_19188,N_17660,N_17713);
nand U19189 (N_19189,N_18210,N_18083);
nor U19190 (N_19190,N_18036,N_18141);
nor U19191 (N_19191,N_18029,N_18397);
and U19192 (N_19192,N_18341,N_17860);
and U19193 (N_19193,N_17667,N_18037);
xor U19194 (N_19194,N_17862,N_18095);
nand U19195 (N_19195,N_17987,N_18126);
nor U19196 (N_19196,N_18341,N_18228);
or U19197 (N_19197,N_18064,N_18285);
nand U19198 (N_19198,N_18197,N_18173);
or U19199 (N_19199,N_17810,N_18346);
and U19200 (N_19200,N_18636,N_18640);
nor U19201 (N_19201,N_18547,N_18579);
and U19202 (N_19202,N_19027,N_18578);
xnor U19203 (N_19203,N_18444,N_18482);
nand U19204 (N_19204,N_18416,N_18516);
nor U19205 (N_19205,N_18937,N_18822);
xor U19206 (N_19206,N_18779,N_18867);
or U19207 (N_19207,N_18964,N_19158);
or U19208 (N_19208,N_18989,N_18652);
xnor U19209 (N_19209,N_18703,N_18448);
nor U19210 (N_19210,N_18472,N_18474);
or U19211 (N_19211,N_18591,N_19160);
nand U19212 (N_19212,N_18506,N_18705);
or U19213 (N_19213,N_18771,N_18501);
or U19214 (N_19214,N_18632,N_18905);
nor U19215 (N_19215,N_18401,N_19035);
and U19216 (N_19216,N_18651,N_18864);
xor U19217 (N_19217,N_18819,N_18816);
nand U19218 (N_19218,N_18793,N_19077);
nand U19219 (N_19219,N_18828,N_18428);
nand U19220 (N_19220,N_18536,N_18443);
nand U19221 (N_19221,N_19179,N_19088);
nand U19222 (N_19222,N_18598,N_18689);
nand U19223 (N_19223,N_19149,N_18806);
nand U19224 (N_19224,N_18568,N_18934);
or U19225 (N_19225,N_18800,N_18635);
xnor U19226 (N_19226,N_18706,N_19128);
and U19227 (N_19227,N_18826,N_19113);
and U19228 (N_19228,N_18955,N_18456);
xnor U19229 (N_19229,N_18814,N_19022);
nand U19230 (N_19230,N_18559,N_19099);
nand U19231 (N_19231,N_19138,N_18714);
nand U19232 (N_19232,N_18941,N_18789);
xor U19233 (N_19233,N_18637,N_18875);
nand U19234 (N_19234,N_19172,N_18449);
nand U19235 (N_19235,N_18721,N_19168);
xor U19236 (N_19236,N_18719,N_19146);
or U19237 (N_19237,N_18969,N_18975);
and U19238 (N_19238,N_18597,N_18677);
nand U19239 (N_19239,N_18702,N_18557);
nor U19240 (N_19240,N_18611,N_18549);
nand U19241 (N_19241,N_19137,N_19165);
nand U19242 (N_19242,N_18972,N_19135);
nor U19243 (N_19243,N_19055,N_18490);
nand U19244 (N_19244,N_18788,N_18644);
and U19245 (N_19245,N_18987,N_18925);
and U19246 (N_19246,N_19100,N_18811);
and U19247 (N_19247,N_18731,N_18945);
nand U19248 (N_19248,N_19001,N_18833);
and U19249 (N_19249,N_19192,N_18497);
nor U19250 (N_19250,N_18571,N_19049);
nand U19251 (N_19251,N_19102,N_18863);
or U19252 (N_19252,N_18555,N_18510);
nand U19253 (N_19253,N_18754,N_18744);
nor U19254 (N_19254,N_18604,N_18954);
nand U19255 (N_19255,N_18874,N_19114);
nand U19256 (N_19256,N_18696,N_19072);
nor U19257 (N_19257,N_18647,N_19034);
or U19258 (N_19258,N_18468,N_19051);
or U19259 (N_19259,N_19081,N_18459);
xor U19260 (N_19260,N_19016,N_19039);
nor U19261 (N_19261,N_18500,N_18465);
nand U19262 (N_19262,N_18745,N_19038);
nor U19263 (N_19263,N_18939,N_18411);
and U19264 (N_19264,N_18629,N_18946);
and U19265 (N_19265,N_18515,N_18410);
xor U19266 (N_19266,N_19191,N_18626);
and U19267 (N_19267,N_18709,N_18633);
xnor U19268 (N_19268,N_18888,N_18612);
and U19269 (N_19269,N_18704,N_18792);
xnor U19270 (N_19270,N_19004,N_18861);
and U19271 (N_19271,N_18866,N_19107);
or U19272 (N_19272,N_18625,N_18913);
xor U19273 (N_19273,N_18736,N_18526);
nand U19274 (N_19274,N_18818,N_18440);
nor U19275 (N_19275,N_19150,N_19050);
or U19276 (N_19276,N_18406,N_18756);
and U19277 (N_19277,N_18796,N_18595);
xnor U19278 (N_19278,N_19196,N_18585);
nor U19279 (N_19279,N_18825,N_18802);
nor U19280 (N_19280,N_19032,N_18670);
xnor U19281 (N_19281,N_18948,N_18673);
nand U19282 (N_19282,N_18967,N_18622);
xnor U19283 (N_19283,N_18914,N_19154);
xnor U19284 (N_19284,N_18424,N_18880);
nand U19285 (N_19285,N_18458,N_18928);
nor U19286 (N_19286,N_18979,N_19166);
nor U19287 (N_19287,N_18577,N_19066);
or U19288 (N_19288,N_18537,N_19133);
nor U19289 (N_19289,N_18949,N_19025);
nor U19290 (N_19290,N_19047,N_18767);
xnor U19291 (N_19291,N_18518,N_18478);
xnor U19292 (N_19292,N_19093,N_18528);
nor U19293 (N_19293,N_18431,N_18879);
and U19294 (N_19294,N_18540,N_18694);
xor U19295 (N_19295,N_18881,N_18916);
xor U19296 (N_19296,N_18728,N_18760);
xor U19297 (N_19297,N_19112,N_18402);
or U19298 (N_19298,N_18603,N_18859);
xnor U19299 (N_19299,N_19056,N_18684);
nand U19300 (N_19300,N_18414,N_18730);
xor U19301 (N_19301,N_18587,N_18658);
xnor U19302 (N_19302,N_18533,N_19152);
xnor U19303 (N_19303,N_19111,N_18430);
and U19304 (N_19304,N_18952,N_18532);
xor U19305 (N_19305,N_19131,N_18734);
and U19306 (N_19306,N_19178,N_18556);
or U19307 (N_19307,N_18798,N_18463);
nor U19308 (N_19308,N_18817,N_18624);
nand U19309 (N_19309,N_18664,N_18682);
and U19310 (N_19310,N_19169,N_18727);
and U19311 (N_19311,N_18446,N_19141);
nand U19312 (N_19312,N_18769,N_18535);
or U19313 (N_19313,N_18906,N_18720);
or U19314 (N_19314,N_18433,N_18545);
and U19315 (N_19315,N_18742,N_18797);
and U19316 (N_19316,N_18417,N_18688);
or U19317 (N_19317,N_18643,N_18686);
xnor U19318 (N_19318,N_19030,N_18523);
xnor U19319 (N_19319,N_19068,N_18836);
or U19320 (N_19320,N_18824,N_18617);
nand U19321 (N_19321,N_18594,N_19078);
nand U19322 (N_19322,N_18755,N_18908);
xor U19323 (N_19323,N_18891,N_18495);
nor U19324 (N_19324,N_19082,N_19184);
or U19325 (N_19325,N_19124,N_18511);
and U19326 (N_19326,N_18509,N_19086);
nor U19327 (N_19327,N_18572,N_18639);
nand U19328 (N_19328,N_18872,N_19009);
or U19329 (N_19329,N_19143,N_18548);
and U19330 (N_19330,N_18968,N_18680);
and U19331 (N_19331,N_18685,N_19083);
and U19332 (N_19332,N_18672,N_19053);
xor U19333 (N_19333,N_18935,N_18641);
and U19334 (N_19334,N_18783,N_18567);
and U19335 (N_19335,N_18447,N_18821);
xor U19336 (N_19336,N_18854,N_18508);
or U19337 (N_19337,N_18971,N_18976);
nor U19338 (N_19338,N_18883,N_19110);
or U19339 (N_19339,N_18809,N_18623);
nor U19340 (N_19340,N_19084,N_18712);
and U19341 (N_19341,N_18912,N_18655);
nand U19342 (N_19342,N_18539,N_19017);
and U19343 (N_19343,N_18407,N_18884);
nor U19344 (N_19344,N_19041,N_18665);
xor U19345 (N_19345,N_18681,N_19136);
xnor U19346 (N_19346,N_18432,N_19060);
and U19347 (N_19347,N_18774,N_18451);
nor U19348 (N_19348,N_18580,N_18564);
nor U19349 (N_19349,N_19062,N_18661);
or U19350 (N_19350,N_18998,N_18846);
nor U19351 (N_19351,N_18606,N_18513);
and U19352 (N_19352,N_18710,N_18929);
nor U19353 (N_19353,N_18610,N_18885);
nand U19354 (N_19354,N_18507,N_18873);
xnor U19355 (N_19355,N_18958,N_18848);
or U19356 (N_19356,N_19183,N_18761);
xnor U19357 (N_19357,N_19155,N_18984);
and U19358 (N_19358,N_18415,N_18514);
xor U19359 (N_19359,N_18794,N_18882);
or U19360 (N_19360,N_18575,N_18426);
xnor U19361 (N_19361,N_18911,N_19079);
nand U19362 (N_19362,N_18951,N_18600);
nor U19363 (N_19363,N_19180,N_18910);
nand U19364 (N_19364,N_18413,N_18840);
nor U19365 (N_19365,N_18820,N_18412);
nand U19366 (N_19366,N_19046,N_18842);
and U19367 (N_19367,N_18887,N_18970);
nor U19368 (N_19368,N_19089,N_18534);
or U19369 (N_19369,N_19074,N_18570);
nand U19370 (N_19370,N_18835,N_18699);
nand U19371 (N_19371,N_18892,N_18542);
or U19372 (N_19372,N_19054,N_18743);
and U19373 (N_19373,N_19148,N_18483);
and U19374 (N_19374,N_19142,N_19123);
xnor U19375 (N_19375,N_18479,N_18749);
xnor U19376 (N_19376,N_18765,N_18654);
and U19377 (N_19377,N_18823,N_18886);
and U19378 (N_19378,N_18986,N_19194);
xor U19379 (N_19379,N_19023,N_18642);
or U19380 (N_19380,N_18697,N_18437);
or U19381 (N_19381,N_18865,N_18502);
nor U19382 (N_19382,N_18933,N_18438);
or U19383 (N_19383,N_19036,N_18663);
nand U19384 (N_19384,N_18810,N_18662);
xnor U19385 (N_19385,N_19162,N_19090);
nand U19386 (N_19386,N_18592,N_18420);
or U19387 (N_19387,N_18999,N_18997);
or U19388 (N_19388,N_18845,N_18834);
nand U19389 (N_19389,N_18405,N_18890);
nand U19390 (N_19390,N_18990,N_18676);
or U19391 (N_19391,N_18936,N_18860);
or U19392 (N_19392,N_18586,N_18876);
or U19393 (N_19393,N_18708,N_18544);
nor U19394 (N_19394,N_18425,N_18653);
or U19395 (N_19395,N_18832,N_19019);
xnor U19396 (N_19396,N_19134,N_18445);
or U19397 (N_19397,N_18576,N_18993);
and U19398 (N_19398,N_18870,N_18434);
xnor U19399 (N_19399,N_18487,N_18943);
and U19400 (N_19400,N_18505,N_18439);
and U19401 (N_19401,N_18926,N_19061);
and U19402 (N_19402,N_18877,N_18503);
nand U19403 (N_19403,N_18646,N_18609);
nand U19404 (N_19404,N_18748,N_18766);
xnor U19405 (N_19405,N_19188,N_18841);
and U19406 (N_19406,N_18992,N_19186);
or U19407 (N_19407,N_19024,N_18781);
xor U19408 (N_19408,N_18784,N_18768);
xnor U19409 (N_19409,N_18455,N_18650);
or U19410 (N_19410,N_19064,N_18581);
nor U19411 (N_19411,N_18675,N_18693);
or U19412 (N_19412,N_19052,N_18920);
nor U19413 (N_19413,N_18504,N_18961);
xnor U19414 (N_19414,N_18450,N_19000);
and U19415 (N_19415,N_18741,N_18775);
and U19416 (N_19416,N_18491,N_18752);
nor U19417 (N_19417,N_18400,N_18546);
and U19418 (N_19418,N_18452,N_18938);
nor U19419 (N_19419,N_18966,N_19119);
and U19420 (N_19420,N_18678,N_19042);
nand U19421 (N_19421,N_19120,N_18746);
or U19422 (N_19422,N_18616,N_18584);
nand U19423 (N_19423,N_18807,N_18895);
nand U19424 (N_19424,N_18956,N_18804);
nor U19425 (N_19425,N_18851,N_18957);
nand U19426 (N_19426,N_19031,N_18808);
or U19427 (N_19427,N_18486,N_19125);
nand U19428 (N_19428,N_19189,N_18715);
xor U19429 (N_19429,N_18960,N_19190);
and U19430 (N_19430,N_19085,N_18857);
or U19431 (N_19431,N_18674,N_19071);
xor U19432 (N_19432,N_18550,N_19067);
nand U19433 (N_19433,N_18470,N_18419);
or U19434 (N_19434,N_19014,N_18561);
xnor U19435 (N_19435,N_18493,N_19197);
or U19436 (N_19436,N_18525,N_18613);
and U19437 (N_19437,N_18837,N_18457);
nor U19438 (N_19438,N_19015,N_18750);
or U19439 (N_19439,N_18915,N_18722);
and U19440 (N_19440,N_19109,N_18805);
nand U19441 (N_19441,N_18460,N_18408);
and U19442 (N_19442,N_18441,N_18517);
nor U19443 (N_19443,N_18787,N_19117);
nor U19444 (N_19444,N_18475,N_18605);
or U19445 (N_19445,N_19013,N_18529);
nor U19446 (N_19446,N_18488,N_19005);
nand U19447 (N_19447,N_18563,N_18919);
or U19448 (N_19448,N_19126,N_18978);
nor U19449 (N_19449,N_18527,N_19103);
or U19450 (N_19450,N_18619,N_19040);
xor U19451 (N_19451,N_18893,N_18593);
and U19452 (N_19452,N_18778,N_18725);
nand U19453 (N_19453,N_18770,N_18422);
or U19454 (N_19454,N_19104,N_19106);
nand U19455 (N_19455,N_19116,N_18473);
and U19456 (N_19456,N_18812,N_19198);
or U19457 (N_19457,N_18522,N_18657);
nor U19458 (N_19458,N_18621,N_19156);
nor U19459 (N_19459,N_18738,N_18786);
nor U19460 (N_19460,N_18666,N_18649);
or U19461 (N_19461,N_18983,N_18973);
xor U19462 (N_19462,N_19069,N_18583);
nand U19463 (N_19463,N_19144,N_18790);
nand U19464 (N_19464,N_18852,N_18691);
and U19465 (N_19465,N_19012,N_18551);
xor U19466 (N_19466,N_19127,N_18695);
nor U19467 (N_19467,N_18485,N_18599);
and U19468 (N_19468,N_18780,N_19043);
and U19469 (N_19469,N_19118,N_19193);
nand U19470 (N_19470,N_18565,N_18889);
or U19471 (N_19471,N_18940,N_19045);
xor U19472 (N_19472,N_18862,N_19076);
or U19473 (N_19473,N_19181,N_18829);
and U19474 (N_19474,N_19026,N_18759);
nor U19475 (N_19475,N_18608,N_18902);
xor U19476 (N_19476,N_18762,N_18869);
nor U19477 (N_19477,N_18850,N_19182);
nand U19478 (N_19478,N_18453,N_18931);
or U19479 (N_19479,N_18977,N_19122);
xor U19480 (N_19480,N_18602,N_18573);
xor U19481 (N_19481,N_18645,N_18904);
xor U19482 (N_19482,N_18454,N_18962);
xnor U19483 (N_19483,N_18520,N_18659);
or U19484 (N_19484,N_18723,N_18950);
or U19485 (N_19485,N_18907,N_18531);
nor U19486 (N_19486,N_18648,N_18724);
nand U19487 (N_19487,N_18764,N_19185);
and U19488 (N_19488,N_19151,N_19170);
or U19489 (N_19489,N_18763,N_18436);
nor U19490 (N_19490,N_18732,N_18981);
or U19491 (N_19491,N_18707,N_18932);
nor U19492 (N_19492,N_18656,N_19174);
or U19493 (N_19493,N_18729,N_18494);
or U19494 (N_19494,N_18991,N_18669);
and U19495 (N_19495,N_19157,N_18521);
nor U19496 (N_19496,N_18512,N_18988);
or U19497 (N_19497,N_19011,N_18903);
and U19498 (N_19498,N_18442,N_18423);
xnor U19499 (N_19499,N_18898,N_18499);
or U19500 (N_19500,N_19167,N_18596);
xor U19501 (N_19501,N_18830,N_18582);
nor U19502 (N_19502,N_18484,N_19096);
nand U19503 (N_19503,N_18427,N_18660);
xnor U19504 (N_19504,N_18839,N_19097);
or U19505 (N_19505,N_18477,N_18801);
and U19506 (N_19506,N_19177,N_19115);
or U19507 (N_19507,N_18541,N_18985);
nand U19508 (N_19508,N_19048,N_19108);
nor U19509 (N_19509,N_18757,N_18530);
nor U19510 (N_19510,N_19075,N_18901);
and U19511 (N_19511,N_19140,N_18980);
nand U19512 (N_19512,N_19091,N_18461);
and U19513 (N_19513,N_18963,N_18858);
xor U19514 (N_19514,N_18553,N_18601);
nand U19515 (N_19515,N_19147,N_18687);
xor U19516 (N_19516,N_18588,N_18421);
nand U19517 (N_19517,N_18480,N_18927);
and U19518 (N_19518,N_18953,N_18607);
and U19519 (N_19519,N_19173,N_18923);
nor U19520 (N_19520,N_18492,N_18683);
xor U19521 (N_19521,N_18855,N_18713);
nor U19522 (N_19522,N_18469,N_18737);
nand U19523 (N_19523,N_19164,N_18429);
xnor U19524 (N_19524,N_18899,N_18844);
nor U19525 (N_19525,N_19058,N_18735);
xnor U19526 (N_19526,N_19098,N_18574);
nand U19527 (N_19527,N_18618,N_18853);
xor U19528 (N_19528,N_19010,N_18944);
nor U19529 (N_19529,N_18638,N_19006);
nand U19530 (N_19530,N_18942,N_18917);
or U19531 (N_19531,N_18897,N_18562);
nor U19532 (N_19532,N_18717,N_18776);
nand U19533 (N_19533,N_18996,N_18476);
nand U19534 (N_19534,N_18995,N_19176);
xnor U19535 (N_19535,N_19070,N_19159);
or U19536 (N_19536,N_18856,N_18569);
or U19537 (N_19537,N_19059,N_18849);
nand U19538 (N_19538,N_18753,N_18909);
or U19539 (N_19539,N_18813,N_19139);
nand U19540 (N_19540,N_19129,N_18519);
xnor U19541 (N_19541,N_18552,N_18740);
and U19542 (N_19542,N_18930,N_18466);
nand U19543 (N_19543,N_19063,N_18614);
xor U19544 (N_19544,N_19175,N_18671);
xnor U19545 (N_19545,N_19105,N_18894);
xnor U19546 (N_19546,N_19008,N_18922);
or U19547 (N_19547,N_18924,N_18489);
and U19548 (N_19548,N_18692,N_18524);
nor U19549 (N_19549,N_19044,N_18831);
xnor U19550 (N_19550,N_18772,N_18718);
nor U19551 (N_19551,N_19087,N_18711);
xor U19552 (N_19552,N_18959,N_18733);
nor U19553 (N_19553,N_18726,N_19020);
and U19554 (N_19554,N_18965,N_18690);
nor U19555 (N_19555,N_19130,N_18630);
or U19556 (N_19556,N_19101,N_18481);
nand U19557 (N_19557,N_18404,N_18974);
nor U19558 (N_19558,N_18698,N_19187);
nand U19559 (N_19559,N_18667,N_18815);
or U19560 (N_19560,N_18700,N_18634);
nand U19561 (N_19561,N_18878,N_18751);
nor U19562 (N_19562,N_18838,N_19073);
nand U19563 (N_19563,N_19065,N_18791);
or U19564 (N_19564,N_18496,N_18827);
nand U19565 (N_19565,N_18777,N_18795);
and U19566 (N_19566,N_19161,N_18994);
xnor U19567 (N_19567,N_18409,N_19121);
xor U19568 (N_19568,N_18871,N_18679);
or U19569 (N_19569,N_19094,N_18701);
or U19570 (N_19570,N_19003,N_18628);
nor U19571 (N_19571,N_18785,N_19007);
or U19572 (N_19572,N_18782,N_18418);
xnor U19573 (N_19573,N_19080,N_18747);
nand U19574 (N_19574,N_18538,N_19092);
xnor U19575 (N_19575,N_18847,N_18471);
nor U19576 (N_19576,N_19021,N_18896);
and U19577 (N_19577,N_18668,N_19195);
and U19578 (N_19578,N_19018,N_18554);
nor U19579 (N_19579,N_18558,N_18803);
nand U19580 (N_19580,N_18589,N_19028);
xor U19581 (N_19581,N_18918,N_19199);
nor U19582 (N_19582,N_19163,N_18464);
and U19583 (N_19583,N_18716,N_19153);
or U19584 (N_19584,N_19145,N_18435);
nor U19585 (N_19585,N_18947,N_19002);
or U19586 (N_19586,N_19037,N_18498);
and U19587 (N_19587,N_18620,N_19171);
xnor U19588 (N_19588,N_18627,N_18843);
xor U19589 (N_19589,N_19095,N_18467);
xnor U19590 (N_19590,N_18739,N_18462);
xor U19591 (N_19591,N_18615,N_18868);
xor U19592 (N_19592,N_18921,N_18773);
nand U19593 (N_19593,N_19132,N_18560);
or U19594 (N_19594,N_18631,N_18566);
and U19595 (N_19595,N_18543,N_18799);
and U19596 (N_19596,N_19057,N_18982);
nand U19597 (N_19597,N_18900,N_18590);
nor U19598 (N_19598,N_19033,N_18758);
nor U19599 (N_19599,N_19029,N_18403);
nand U19600 (N_19600,N_18400,N_18479);
xor U19601 (N_19601,N_18824,N_18662);
or U19602 (N_19602,N_18755,N_18895);
nand U19603 (N_19603,N_18676,N_18440);
xor U19604 (N_19604,N_18904,N_19048);
xor U19605 (N_19605,N_19188,N_18759);
and U19606 (N_19606,N_19019,N_18519);
xnor U19607 (N_19607,N_18766,N_18640);
xor U19608 (N_19608,N_18494,N_19198);
xnor U19609 (N_19609,N_18767,N_18823);
xor U19610 (N_19610,N_18960,N_19076);
or U19611 (N_19611,N_19033,N_18862);
xor U19612 (N_19612,N_18730,N_18931);
nand U19613 (N_19613,N_18794,N_19068);
and U19614 (N_19614,N_18613,N_19154);
nor U19615 (N_19615,N_18939,N_19079);
nand U19616 (N_19616,N_18519,N_18911);
nand U19617 (N_19617,N_18560,N_18705);
xnor U19618 (N_19618,N_18958,N_19103);
xor U19619 (N_19619,N_18430,N_18680);
nor U19620 (N_19620,N_19120,N_19079);
and U19621 (N_19621,N_18778,N_19057);
and U19622 (N_19622,N_18593,N_18606);
nand U19623 (N_19623,N_18985,N_18623);
and U19624 (N_19624,N_18431,N_18793);
or U19625 (N_19625,N_18583,N_18904);
and U19626 (N_19626,N_18993,N_18761);
nor U19627 (N_19627,N_18792,N_18645);
and U19628 (N_19628,N_18836,N_18785);
or U19629 (N_19629,N_18462,N_18811);
or U19630 (N_19630,N_18876,N_18533);
xnor U19631 (N_19631,N_18596,N_18765);
xor U19632 (N_19632,N_18434,N_18543);
xnor U19633 (N_19633,N_18632,N_19056);
or U19634 (N_19634,N_18813,N_18484);
nor U19635 (N_19635,N_18739,N_18914);
and U19636 (N_19636,N_18896,N_18836);
nand U19637 (N_19637,N_19019,N_18618);
and U19638 (N_19638,N_18615,N_18402);
or U19639 (N_19639,N_19081,N_18852);
nor U19640 (N_19640,N_19099,N_19044);
nand U19641 (N_19641,N_19074,N_19066);
and U19642 (N_19642,N_18430,N_18438);
nand U19643 (N_19643,N_18619,N_19187);
nor U19644 (N_19644,N_18950,N_19070);
nand U19645 (N_19645,N_18739,N_19188);
and U19646 (N_19646,N_18977,N_19173);
and U19647 (N_19647,N_19087,N_18757);
nand U19648 (N_19648,N_19125,N_19181);
xor U19649 (N_19649,N_18857,N_18643);
nand U19650 (N_19650,N_18496,N_18762);
and U19651 (N_19651,N_19003,N_19174);
and U19652 (N_19652,N_18973,N_18432);
and U19653 (N_19653,N_18980,N_18400);
or U19654 (N_19654,N_18942,N_18434);
xor U19655 (N_19655,N_18409,N_19084);
and U19656 (N_19656,N_19134,N_18602);
nor U19657 (N_19657,N_19133,N_18586);
and U19658 (N_19658,N_18707,N_19191);
nand U19659 (N_19659,N_19089,N_18805);
nor U19660 (N_19660,N_18784,N_18669);
and U19661 (N_19661,N_19181,N_18736);
or U19662 (N_19662,N_19016,N_18590);
xor U19663 (N_19663,N_18538,N_18964);
or U19664 (N_19664,N_19051,N_19075);
or U19665 (N_19665,N_19005,N_18682);
nor U19666 (N_19666,N_18466,N_19066);
nand U19667 (N_19667,N_18402,N_18747);
nand U19668 (N_19668,N_18832,N_18721);
xor U19669 (N_19669,N_18542,N_18571);
nor U19670 (N_19670,N_18871,N_18554);
or U19671 (N_19671,N_18551,N_18754);
and U19672 (N_19672,N_19182,N_18414);
nor U19673 (N_19673,N_18503,N_18702);
and U19674 (N_19674,N_18452,N_19120);
nor U19675 (N_19675,N_18979,N_18419);
nand U19676 (N_19676,N_19050,N_18898);
xnor U19677 (N_19677,N_18919,N_19066);
xnor U19678 (N_19678,N_19197,N_18878);
nor U19679 (N_19679,N_19131,N_18918);
xor U19680 (N_19680,N_18833,N_18510);
xor U19681 (N_19681,N_18436,N_18554);
xnor U19682 (N_19682,N_18569,N_19032);
and U19683 (N_19683,N_19065,N_19081);
nor U19684 (N_19684,N_18993,N_19176);
xor U19685 (N_19685,N_18769,N_18417);
nand U19686 (N_19686,N_18734,N_18724);
and U19687 (N_19687,N_18660,N_18935);
and U19688 (N_19688,N_18405,N_19184);
and U19689 (N_19689,N_19168,N_18617);
nor U19690 (N_19690,N_18615,N_18862);
and U19691 (N_19691,N_18400,N_18462);
or U19692 (N_19692,N_18704,N_18721);
xnor U19693 (N_19693,N_19180,N_18430);
xnor U19694 (N_19694,N_18584,N_18829);
and U19695 (N_19695,N_18974,N_18912);
and U19696 (N_19696,N_18801,N_18449);
and U19697 (N_19697,N_18989,N_18654);
or U19698 (N_19698,N_19024,N_19007);
nand U19699 (N_19699,N_18754,N_18615);
nand U19700 (N_19700,N_19029,N_18817);
xor U19701 (N_19701,N_18673,N_18835);
and U19702 (N_19702,N_18419,N_18926);
and U19703 (N_19703,N_18582,N_19119);
xnor U19704 (N_19704,N_18998,N_18635);
and U19705 (N_19705,N_18775,N_18979);
and U19706 (N_19706,N_18600,N_19169);
nand U19707 (N_19707,N_19142,N_18818);
xnor U19708 (N_19708,N_19124,N_19162);
xor U19709 (N_19709,N_18727,N_18551);
xor U19710 (N_19710,N_18406,N_18788);
and U19711 (N_19711,N_18643,N_18448);
nand U19712 (N_19712,N_18890,N_19013);
and U19713 (N_19713,N_18740,N_18685);
and U19714 (N_19714,N_18430,N_18694);
xor U19715 (N_19715,N_18920,N_19125);
xnor U19716 (N_19716,N_18735,N_18656);
xor U19717 (N_19717,N_19129,N_18499);
and U19718 (N_19718,N_18759,N_18682);
xor U19719 (N_19719,N_18619,N_18900);
xor U19720 (N_19720,N_18769,N_19193);
nor U19721 (N_19721,N_18574,N_18562);
nor U19722 (N_19722,N_19179,N_18827);
or U19723 (N_19723,N_18429,N_18712);
or U19724 (N_19724,N_18409,N_19174);
xor U19725 (N_19725,N_18407,N_19156);
and U19726 (N_19726,N_18741,N_18752);
xnor U19727 (N_19727,N_18429,N_19040);
nor U19728 (N_19728,N_18714,N_19016);
nor U19729 (N_19729,N_18898,N_18487);
xnor U19730 (N_19730,N_18940,N_18506);
or U19731 (N_19731,N_19156,N_19198);
or U19732 (N_19732,N_19072,N_18521);
nand U19733 (N_19733,N_18734,N_18595);
or U19734 (N_19734,N_19124,N_19076);
xor U19735 (N_19735,N_18532,N_18872);
xor U19736 (N_19736,N_18429,N_19064);
and U19737 (N_19737,N_18676,N_18506);
and U19738 (N_19738,N_18668,N_18492);
or U19739 (N_19739,N_18925,N_18691);
nand U19740 (N_19740,N_19033,N_18593);
xnor U19741 (N_19741,N_19106,N_18813);
xnor U19742 (N_19742,N_18417,N_18698);
nor U19743 (N_19743,N_19198,N_18955);
nand U19744 (N_19744,N_18435,N_18575);
nand U19745 (N_19745,N_18509,N_18525);
nor U19746 (N_19746,N_18690,N_18649);
and U19747 (N_19747,N_18788,N_18902);
nand U19748 (N_19748,N_18562,N_18619);
and U19749 (N_19749,N_19169,N_19124);
or U19750 (N_19750,N_19174,N_19084);
nand U19751 (N_19751,N_18964,N_18431);
xnor U19752 (N_19752,N_18730,N_18964);
xor U19753 (N_19753,N_18825,N_18929);
nand U19754 (N_19754,N_19177,N_19073);
and U19755 (N_19755,N_18939,N_18804);
or U19756 (N_19756,N_18931,N_18824);
xor U19757 (N_19757,N_18981,N_19040);
nor U19758 (N_19758,N_18511,N_18551);
xor U19759 (N_19759,N_18900,N_18782);
nand U19760 (N_19760,N_18432,N_18506);
or U19761 (N_19761,N_18430,N_18504);
xor U19762 (N_19762,N_19039,N_18645);
or U19763 (N_19763,N_18738,N_19042);
nor U19764 (N_19764,N_18825,N_18733);
nor U19765 (N_19765,N_19053,N_18714);
or U19766 (N_19766,N_18716,N_18843);
and U19767 (N_19767,N_18609,N_18411);
nor U19768 (N_19768,N_18535,N_18798);
nand U19769 (N_19769,N_18764,N_18563);
xor U19770 (N_19770,N_19132,N_19143);
nor U19771 (N_19771,N_18498,N_18993);
nor U19772 (N_19772,N_18846,N_18541);
nor U19773 (N_19773,N_18777,N_18638);
nand U19774 (N_19774,N_18942,N_18741);
nand U19775 (N_19775,N_18981,N_19116);
or U19776 (N_19776,N_18500,N_18453);
xnor U19777 (N_19777,N_18858,N_19068);
nor U19778 (N_19778,N_18604,N_18487);
or U19779 (N_19779,N_19065,N_18901);
nand U19780 (N_19780,N_19058,N_18912);
nor U19781 (N_19781,N_19059,N_18752);
nand U19782 (N_19782,N_18476,N_18433);
xnor U19783 (N_19783,N_18990,N_18614);
and U19784 (N_19784,N_18569,N_19132);
nand U19785 (N_19785,N_18676,N_18832);
or U19786 (N_19786,N_19022,N_19175);
or U19787 (N_19787,N_18519,N_18920);
or U19788 (N_19788,N_18830,N_18759);
nor U19789 (N_19789,N_19066,N_18888);
or U19790 (N_19790,N_18788,N_19043);
nand U19791 (N_19791,N_18487,N_18719);
nor U19792 (N_19792,N_19061,N_19070);
nand U19793 (N_19793,N_18429,N_18471);
or U19794 (N_19794,N_18462,N_19008);
and U19795 (N_19795,N_18510,N_18535);
or U19796 (N_19796,N_18674,N_18671);
or U19797 (N_19797,N_19088,N_18918);
nor U19798 (N_19798,N_18859,N_18438);
nand U19799 (N_19799,N_18945,N_18634);
nand U19800 (N_19800,N_18448,N_18725);
and U19801 (N_19801,N_18874,N_18465);
nand U19802 (N_19802,N_19179,N_18750);
xor U19803 (N_19803,N_18410,N_19158);
nand U19804 (N_19804,N_19063,N_18441);
or U19805 (N_19805,N_19056,N_18576);
nand U19806 (N_19806,N_19152,N_19080);
nor U19807 (N_19807,N_19155,N_18613);
nand U19808 (N_19808,N_19047,N_19068);
xor U19809 (N_19809,N_18486,N_18801);
or U19810 (N_19810,N_18743,N_18430);
nand U19811 (N_19811,N_19180,N_18873);
nor U19812 (N_19812,N_18809,N_18425);
and U19813 (N_19813,N_19011,N_18800);
nand U19814 (N_19814,N_18945,N_18479);
and U19815 (N_19815,N_18881,N_18610);
nand U19816 (N_19816,N_18688,N_18972);
nor U19817 (N_19817,N_18539,N_19125);
nor U19818 (N_19818,N_18683,N_18473);
xnor U19819 (N_19819,N_19091,N_18480);
and U19820 (N_19820,N_18686,N_18590);
or U19821 (N_19821,N_18796,N_18863);
or U19822 (N_19822,N_19109,N_19027);
or U19823 (N_19823,N_18847,N_19037);
nor U19824 (N_19824,N_18658,N_19192);
nand U19825 (N_19825,N_18884,N_18982);
and U19826 (N_19826,N_18991,N_18654);
xnor U19827 (N_19827,N_18753,N_19187);
or U19828 (N_19828,N_18423,N_19025);
nand U19829 (N_19829,N_18723,N_18567);
nor U19830 (N_19830,N_18624,N_18450);
nor U19831 (N_19831,N_18717,N_18870);
or U19832 (N_19832,N_18655,N_18567);
xnor U19833 (N_19833,N_18436,N_18703);
and U19834 (N_19834,N_18938,N_18720);
nand U19835 (N_19835,N_18933,N_18700);
nand U19836 (N_19836,N_18579,N_18723);
or U19837 (N_19837,N_18627,N_18400);
or U19838 (N_19838,N_18833,N_18508);
nor U19839 (N_19839,N_18746,N_18603);
nor U19840 (N_19840,N_18475,N_18828);
and U19841 (N_19841,N_19172,N_18506);
nor U19842 (N_19842,N_18458,N_18929);
nand U19843 (N_19843,N_18908,N_19007);
nor U19844 (N_19844,N_18801,N_18956);
xnor U19845 (N_19845,N_18743,N_19050);
nand U19846 (N_19846,N_18752,N_18942);
and U19847 (N_19847,N_19135,N_18550);
nor U19848 (N_19848,N_18457,N_18693);
or U19849 (N_19849,N_18450,N_18493);
xor U19850 (N_19850,N_18862,N_19153);
nand U19851 (N_19851,N_18992,N_18805);
and U19852 (N_19852,N_19136,N_19066);
nor U19853 (N_19853,N_18626,N_18900);
nor U19854 (N_19854,N_18965,N_18813);
nor U19855 (N_19855,N_18981,N_18498);
nor U19856 (N_19856,N_18494,N_18974);
xnor U19857 (N_19857,N_19114,N_19021);
nand U19858 (N_19858,N_18893,N_18527);
nand U19859 (N_19859,N_19011,N_18972);
xnor U19860 (N_19860,N_18580,N_19070);
nor U19861 (N_19861,N_18967,N_18876);
nor U19862 (N_19862,N_19030,N_18882);
nor U19863 (N_19863,N_18989,N_18410);
or U19864 (N_19864,N_18461,N_18585);
nor U19865 (N_19865,N_18792,N_18634);
nand U19866 (N_19866,N_19151,N_19174);
and U19867 (N_19867,N_18671,N_18416);
or U19868 (N_19868,N_18669,N_19066);
or U19869 (N_19869,N_18786,N_18526);
and U19870 (N_19870,N_18646,N_19004);
or U19871 (N_19871,N_18735,N_18622);
nand U19872 (N_19872,N_18731,N_19026);
nor U19873 (N_19873,N_18622,N_19121);
and U19874 (N_19874,N_19162,N_18895);
nor U19875 (N_19875,N_18530,N_18966);
xor U19876 (N_19876,N_18824,N_18903);
and U19877 (N_19877,N_18991,N_18913);
and U19878 (N_19878,N_18831,N_18802);
nor U19879 (N_19879,N_18848,N_19101);
and U19880 (N_19880,N_18844,N_18534);
nor U19881 (N_19881,N_18698,N_18400);
nand U19882 (N_19882,N_18823,N_18867);
or U19883 (N_19883,N_19099,N_18996);
nand U19884 (N_19884,N_18603,N_18589);
nand U19885 (N_19885,N_18597,N_19164);
and U19886 (N_19886,N_18495,N_18516);
nor U19887 (N_19887,N_19007,N_19137);
nand U19888 (N_19888,N_18554,N_18671);
nand U19889 (N_19889,N_18820,N_18547);
and U19890 (N_19890,N_18458,N_19072);
or U19891 (N_19891,N_18569,N_19070);
xnor U19892 (N_19892,N_19121,N_19011);
and U19893 (N_19893,N_18400,N_19080);
nand U19894 (N_19894,N_18727,N_18509);
nor U19895 (N_19895,N_18583,N_18513);
nand U19896 (N_19896,N_18472,N_18419);
nand U19897 (N_19897,N_18684,N_18769);
or U19898 (N_19898,N_18508,N_19001);
xor U19899 (N_19899,N_19014,N_18825);
nor U19900 (N_19900,N_19115,N_19051);
nand U19901 (N_19901,N_19075,N_18680);
and U19902 (N_19902,N_18579,N_18644);
xnor U19903 (N_19903,N_18620,N_18668);
nand U19904 (N_19904,N_18639,N_18522);
and U19905 (N_19905,N_19105,N_18736);
and U19906 (N_19906,N_18840,N_18937);
and U19907 (N_19907,N_18752,N_19078);
nand U19908 (N_19908,N_18818,N_19156);
nand U19909 (N_19909,N_19126,N_18864);
or U19910 (N_19910,N_18618,N_19092);
xnor U19911 (N_19911,N_19062,N_18487);
or U19912 (N_19912,N_19006,N_18469);
or U19913 (N_19913,N_18489,N_19106);
xnor U19914 (N_19914,N_18533,N_18848);
nor U19915 (N_19915,N_19014,N_19003);
nand U19916 (N_19916,N_18514,N_18717);
and U19917 (N_19917,N_18830,N_18913);
nor U19918 (N_19918,N_18609,N_18771);
nor U19919 (N_19919,N_18952,N_19049);
or U19920 (N_19920,N_18506,N_19104);
nand U19921 (N_19921,N_18520,N_18996);
or U19922 (N_19922,N_18810,N_18411);
nor U19923 (N_19923,N_18592,N_18832);
xor U19924 (N_19924,N_19068,N_19101);
or U19925 (N_19925,N_18822,N_18707);
and U19926 (N_19926,N_18602,N_18895);
and U19927 (N_19927,N_19103,N_19135);
or U19928 (N_19928,N_19190,N_19144);
nand U19929 (N_19929,N_18637,N_18876);
nor U19930 (N_19930,N_18929,N_18573);
or U19931 (N_19931,N_19121,N_19072);
xnor U19932 (N_19932,N_18769,N_18546);
nor U19933 (N_19933,N_19027,N_18968);
nor U19934 (N_19934,N_18748,N_18896);
nor U19935 (N_19935,N_18607,N_18518);
or U19936 (N_19936,N_19189,N_18666);
nor U19937 (N_19937,N_19163,N_18937);
nor U19938 (N_19938,N_18420,N_19014);
or U19939 (N_19939,N_19038,N_18781);
xor U19940 (N_19940,N_18481,N_18433);
nor U19941 (N_19941,N_19154,N_18673);
or U19942 (N_19942,N_18686,N_19132);
or U19943 (N_19943,N_19146,N_18992);
xor U19944 (N_19944,N_18640,N_18597);
and U19945 (N_19945,N_18748,N_18922);
nand U19946 (N_19946,N_18717,N_18716);
nor U19947 (N_19947,N_18606,N_18698);
or U19948 (N_19948,N_19194,N_18868);
xor U19949 (N_19949,N_18868,N_19115);
nor U19950 (N_19950,N_19023,N_18631);
and U19951 (N_19951,N_18935,N_18436);
and U19952 (N_19952,N_18742,N_18926);
xor U19953 (N_19953,N_18958,N_18585);
xor U19954 (N_19954,N_18992,N_18873);
nor U19955 (N_19955,N_19019,N_18438);
nand U19956 (N_19956,N_18455,N_19185);
or U19957 (N_19957,N_19059,N_18572);
nor U19958 (N_19958,N_19071,N_18806);
nor U19959 (N_19959,N_18797,N_18911);
nand U19960 (N_19960,N_18716,N_18837);
nand U19961 (N_19961,N_18847,N_18511);
and U19962 (N_19962,N_18774,N_18635);
nand U19963 (N_19963,N_18761,N_18515);
nand U19964 (N_19964,N_18529,N_19007);
nor U19965 (N_19965,N_19114,N_18714);
nand U19966 (N_19966,N_18702,N_19104);
nand U19967 (N_19967,N_19015,N_19027);
xor U19968 (N_19968,N_18884,N_18635);
or U19969 (N_19969,N_19003,N_18764);
nor U19970 (N_19970,N_18433,N_18503);
or U19971 (N_19971,N_19008,N_19029);
and U19972 (N_19972,N_18876,N_18433);
nor U19973 (N_19973,N_18946,N_18443);
and U19974 (N_19974,N_19143,N_19055);
nand U19975 (N_19975,N_18404,N_18586);
or U19976 (N_19976,N_18528,N_18566);
or U19977 (N_19977,N_19060,N_19149);
and U19978 (N_19978,N_18822,N_19176);
nand U19979 (N_19979,N_18450,N_18671);
or U19980 (N_19980,N_18854,N_19179);
xor U19981 (N_19981,N_19172,N_18624);
nor U19982 (N_19982,N_18862,N_18917);
nor U19983 (N_19983,N_18806,N_18691);
or U19984 (N_19984,N_18462,N_18672);
nor U19985 (N_19985,N_18415,N_18696);
nor U19986 (N_19986,N_18719,N_19092);
and U19987 (N_19987,N_18490,N_18935);
or U19988 (N_19988,N_18579,N_18524);
xnor U19989 (N_19989,N_19125,N_18808);
and U19990 (N_19990,N_18410,N_19026);
xor U19991 (N_19991,N_18923,N_19109);
nor U19992 (N_19992,N_18585,N_18777);
xnor U19993 (N_19993,N_18511,N_18618);
and U19994 (N_19994,N_19042,N_18875);
xnor U19995 (N_19995,N_18963,N_18723);
xor U19996 (N_19996,N_18593,N_18447);
and U19997 (N_19997,N_18839,N_18424);
nand U19998 (N_19998,N_18618,N_18922);
xnor U19999 (N_19999,N_18938,N_18897);
nand UO_0 (O_0,N_19856,N_19463);
and UO_1 (O_1,N_19716,N_19666);
and UO_2 (O_2,N_19350,N_19571);
or UO_3 (O_3,N_19524,N_19864);
nor UO_4 (O_4,N_19830,N_19767);
xor UO_5 (O_5,N_19436,N_19410);
and UO_6 (O_6,N_19668,N_19734);
xor UO_7 (O_7,N_19260,N_19663);
xor UO_8 (O_8,N_19619,N_19355);
nand UO_9 (O_9,N_19318,N_19375);
xor UO_10 (O_10,N_19758,N_19428);
or UO_11 (O_11,N_19839,N_19865);
xor UO_12 (O_12,N_19433,N_19304);
or UO_13 (O_13,N_19937,N_19849);
xnor UO_14 (O_14,N_19422,N_19944);
nand UO_15 (O_15,N_19217,N_19890);
and UO_16 (O_16,N_19623,N_19307);
nor UO_17 (O_17,N_19413,N_19998);
xor UO_18 (O_18,N_19662,N_19387);
nand UO_19 (O_19,N_19746,N_19905);
nand UO_20 (O_20,N_19957,N_19687);
nor UO_21 (O_21,N_19540,N_19869);
and UO_22 (O_22,N_19693,N_19395);
nor UO_23 (O_23,N_19978,N_19925);
or UO_24 (O_24,N_19807,N_19381);
and UO_25 (O_25,N_19562,N_19382);
or UO_26 (O_26,N_19589,N_19425);
and UO_27 (O_27,N_19363,N_19234);
nor UO_28 (O_28,N_19765,N_19251);
nor UO_29 (O_29,N_19986,N_19518);
nor UO_30 (O_30,N_19711,N_19760);
or UO_31 (O_31,N_19919,N_19982);
nand UO_32 (O_32,N_19831,N_19641);
and UO_33 (O_33,N_19420,N_19288);
or UO_34 (O_34,N_19759,N_19983);
or UO_35 (O_35,N_19652,N_19582);
or UO_36 (O_36,N_19888,N_19501);
nor UO_37 (O_37,N_19333,N_19223);
nand UO_38 (O_38,N_19719,N_19536);
nand UO_39 (O_39,N_19591,N_19301);
xnor UO_40 (O_40,N_19908,N_19928);
nand UO_41 (O_41,N_19277,N_19399);
nand UO_42 (O_42,N_19930,N_19400);
xor UO_43 (O_43,N_19336,N_19263);
nor UO_44 (O_44,N_19927,N_19955);
xor UO_45 (O_45,N_19423,N_19601);
nor UO_46 (O_46,N_19238,N_19655);
nand UO_47 (O_47,N_19945,N_19384);
nand UO_48 (O_48,N_19300,N_19320);
nor UO_49 (O_49,N_19622,N_19292);
and UO_50 (O_50,N_19611,N_19871);
and UO_51 (O_51,N_19431,N_19337);
nor UO_52 (O_52,N_19850,N_19366);
or UO_53 (O_53,N_19672,N_19441);
nand UO_54 (O_54,N_19684,N_19513);
nand UO_55 (O_55,N_19946,N_19820);
xnor UO_56 (O_56,N_19340,N_19812);
and UO_57 (O_57,N_19502,N_19570);
or UO_58 (O_58,N_19305,N_19416);
or UO_59 (O_59,N_19694,N_19806);
nand UO_60 (O_60,N_19299,N_19326);
nand UO_61 (O_61,N_19907,N_19948);
and UO_62 (O_62,N_19763,N_19893);
or UO_63 (O_63,N_19804,N_19607);
xnor UO_64 (O_64,N_19226,N_19979);
and UO_65 (O_65,N_19915,N_19862);
nor UO_66 (O_66,N_19426,N_19965);
and UO_67 (O_67,N_19389,N_19418);
and UO_68 (O_68,N_19278,N_19397);
and UO_69 (O_69,N_19303,N_19692);
nand UO_70 (O_70,N_19459,N_19421);
nand UO_71 (O_71,N_19933,N_19963);
or UO_72 (O_72,N_19916,N_19887);
or UO_73 (O_73,N_19229,N_19755);
nor UO_74 (O_74,N_19493,N_19659);
and UO_75 (O_75,N_19374,N_19510);
xor UO_76 (O_76,N_19360,N_19764);
nor UO_77 (O_77,N_19247,N_19624);
or UO_78 (O_78,N_19857,N_19654);
xnor UO_79 (O_79,N_19786,N_19492);
and UO_80 (O_80,N_19789,N_19784);
nand UO_81 (O_81,N_19590,N_19265);
or UO_82 (O_82,N_19310,N_19816);
xor UO_83 (O_83,N_19579,N_19991);
or UO_84 (O_84,N_19519,N_19832);
xnor UO_85 (O_85,N_19696,N_19473);
xor UO_86 (O_86,N_19942,N_19914);
xnor UO_87 (O_87,N_19995,N_19508);
nand UO_88 (O_88,N_19828,N_19396);
nor UO_89 (O_89,N_19721,N_19772);
and UO_90 (O_90,N_19625,N_19718);
or UO_91 (O_91,N_19600,N_19621);
or UO_92 (O_92,N_19818,N_19636);
or UO_93 (O_93,N_19253,N_19594);
nor UO_94 (O_94,N_19456,N_19559);
nand UO_95 (O_95,N_19637,N_19385);
and UO_96 (O_96,N_19270,N_19489);
or UO_97 (O_97,N_19439,N_19380);
or UO_98 (O_98,N_19639,N_19327);
or UO_99 (O_99,N_19909,N_19227);
xor UO_100 (O_100,N_19671,N_19936);
nand UO_101 (O_101,N_19911,N_19731);
xnor UO_102 (O_102,N_19324,N_19701);
and UO_103 (O_103,N_19574,N_19403);
xnor UO_104 (O_104,N_19939,N_19285);
and UO_105 (O_105,N_19612,N_19412);
or UO_106 (O_106,N_19297,N_19640);
and UO_107 (O_107,N_19975,N_19537);
nor UO_108 (O_108,N_19530,N_19709);
xnor UO_109 (O_109,N_19593,N_19823);
or UO_110 (O_110,N_19988,N_19279);
or UO_111 (O_111,N_19921,N_19917);
xnor UO_112 (O_112,N_19923,N_19321);
nand UO_113 (O_113,N_19809,N_19458);
nor UO_114 (O_114,N_19268,N_19861);
xnor UO_115 (O_115,N_19878,N_19203);
and UO_116 (O_116,N_19884,N_19616);
nor UO_117 (O_117,N_19686,N_19770);
or UO_118 (O_118,N_19368,N_19854);
or UO_119 (O_119,N_19649,N_19653);
and UO_120 (O_120,N_19523,N_19323);
xor UO_121 (O_121,N_19977,N_19450);
and UO_122 (O_122,N_19408,N_19967);
xor UO_123 (O_123,N_19596,N_19932);
xor UO_124 (O_124,N_19386,N_19660);
or UO_125 (O_125,N_19214,N_19880);
xor UO_126 (O_126,N_19240,N_19796);
and UO_127 (O_127,N_19533,N_19442);
nor UO_128 (O_128,N_19252,N_19401);
nor UO_129 (O_129,N_19514,N_19475);
nor UO_130 (O_130,N_19896,N_19209);
nor UO_131 (O_131,N_19218,N_19264);
or UO_132 (O_132,N_19414,N_19296);
or UO_133 (O_133,N_19542,N_19656);
nor UO_134 (O_134,N_19605,N_19364);
or UO_135 (O_135,N_19840,N_19406);
or UO_136 (O_136,N_19996,N_19308);
nor UO_137 (O_137,N_19695,N_19526);
nand UO_138 (O_138,N_19319,N_19648);
nor UO_139 (O_139,N_19561,N_19273);
nor UO_140 (O_140,N_19785,N_19434);
nor UO_141 (O_141,N_19328,N_19868);
and UO_142 (O_142,N_19555,N_19630);
nand UO_143 (O_143,N_19883,N_19311);
nor UO_144 (O_144,N_19244,N_19259);
and UO_145 (O_145,N_19951,N_19383);
and UO_146 (O_146,N_19280,N_19200);
nor UO_147 (O_147,N_19245,N_19920);
xnor UO_148 (O_148,N_19969,N_19494);
nand UO_149 (O_149,N_19315,N_19257);
nor UO_150 (O_150,N_19306,N_19312);
or UO_151 (O_151,N_19903,N_19215);
nand UO_152 (O_152,N_19521,N_19943);
nand UO_153 (O_153,N_19713,N_19778);
or UO_154 (O_154,N_19810,N_19237);
and UO_155 (O_155,N_19528,N_19973);
or UO_156 (O_156,N_19626,N_19405);
or UO_157 (O_157,N_19814,N_19954);
xnor UO_158 (O_158,N_19730,N_19503);
or UO_159 (O_159,N_19912,N_19833);
or UO_160 (O_160,N_19469,N_19614);
and UO_161 (O_161,N_19790,N_19344);
or UO_162 (O_162,N_19747,N_19958);
xor UO_163 (O_163,N_19870,N_19782);
nor UO_164 (O_164,N_19815,N_19783);
xor UO_165 (O_165,N_19525,N_19348);
nand UO_166 (O_166,N_19733,N_19262);
nand UO_167 (O_167,N_19242,N_19918);
and UO_168 (O_168,N_19225,N_19873);
or UO_169 (O_169,N_19438,N_19404);
nand UO_170 (O_170,N_19287,N_19803);
nor UO_171 (O_171,N_19678,N_19239);
xor UO_172 (O_172,N_19726,N_19276);
and UO_173 (O_173,N_19291,N_19867);
or UO_174 (O_174,N_19346,N_19752);
nor UO_175 (O_175,N_19699,N_19343);
xnor UO_176 (O_176,N_19429,N_19222);
or UO_177 (O_177,N_19361,N_19827);
xor UO_178 (O_178,N_19956,N_19522);
nor UO_179 (O_179,N_19775,N_19787);
and UO_180 (O_180,N_19517,N_19959);
nand UO_181 (O_181,N_19462,N_19283);
nor UO_182 (O_182,N_19609,N_19367);
nor UO_183 (O_183,N_19424,N_19681);
and UO_184 (O_184,N_19881,N_19651);
nand UO_185 (O_185,N_19506,N_19885);
xnor UO_186 (O_186,N_19970,N_19643);
xnor UO_187 (O_187,N_19577,N_19520);
nand UO_188 (O_188,N_19388,N_19208);
nand UO_189 (O_189,N_19398,N_19795);
nand UO_190 (O_190,N_19698,N_19750);
nand UO_191 (O_191,N_19606,N_19531);
nor UO_192 (O_192,N_19595,N_19682);
and UO_193 (O_193,N_19586,N_19427);
nand UO_194 (O_194,N_19771,N_19766);
xor UO_195 (O_195,N_19232,N_19359);
nand UO_196 (O_196,N_19373,N_19339);
nand UO_197 (O_197,N_19558,N_19900);
or UO_198 (O_198,N_19634,N_19675);
xor UO_199 (O_199,N_19723,N_19309);
nor UO_200 (O_200,N_19910,N_19560);
nand UO_201 (O_201,N_19712,N_19415);
or UO_202 (O_202,N_19892,N_19485);
and UO_203 (O_203,N_19466,N_19365);
or UO_204 (O_204,N_19357,N_19739);
nor UO_205 (O_205,N_19842,N_19569);
and UO_206 (O_206,N_19875,N_19894);
xor UO_207 (O_207,N_19735,N_19322);
nand UO_208 (O_208,N_19255,N_19479);
or UO_209 (O_209,N_19216,N_19592);
and UO_210 (O_210,N_19940,N_19836);
and UO_211 (O_211,N_19897,N_19211);
xnor UO_212 (O_212,N_19886,N_19379);
nand UO_213 (O_213,N_19566,N_19353);
or UO_214 (O_214,N_19825,N_19358);
nand UO_215 (O_215,N_19669,N_19302);
xor UO_216 (O_216,N_19876,N_19556);
nand UO_217 (O_217,N_19511,N_19706);
or UO_218 (O_218,N_19529,N_19547);
and UO_219 (O_219,N_19204,N_19821);
nand UO_220 (O_220,N_19749,N_19443);
nor UO_221 (O_221,N_19349,N_19805);
xnor UO_222 (O_222,N_19352,N_19314);
nand UO_223 (O_223,N_19550,N_19507);
xnor UO_224 (O_224,N_19604,N_19347);
or UO_225 (O_225,N_19779,N_19271);
and UO_226 (O_226,N_19847,N_19235);
nor UO_227 (O_227,N_19551,N_19464);
nand UO_228 (O_228,N_19497,N_19851);
or UO_229 (O_229,N_19976,N_19674);
or UO_230 (O_230,N_19793,N_19286);
or UO_231 (O_231,N_19947,N_19440);
nor UO_232 (O_232,N_19476,N_19356);
nor UO_233 (O_233,N_19393,N_19563);
nand UO_234 (O_234,N_19535,N_19802);
and UO_235 (O_235,N_19205,N_19435);
or UO_236 (O_236,N_19811,N_19748);
nand UO_237 (O_237,N_19295,N_19859);
and UO_238 (O_238,N_19598,N_19834);
and UO_239 (O_239,N_19791,N_19822);
xor UO_240 (O_240,N_19829,N_19498);
or UO_241 (O_241,N_19342,N_19902);
and UO_242 (O_242,N_19838,N_19906);
xnor UO_243 (O_243,N_19534,N_19743);
nand UO_244 (O_244,N_19950,N_19482);
and UO_245 (O_245,N_19557,N_19960);
and UO_246 (O_246,N_19581,N_19231);
nand UO_247 (O_247,N_19275,N_19646);
and UO_248 (O_248,N_19757,N_19904);
nand UO_249 (O_249,N_19505,N_19797);
nand UO_250 (O_250,N_19568,N_19372);
and UO_251 (O_251,N_19298,N_19632);
nand UO_252 (O_252,N_19889,N_19202);
and UO_253 (O_253,N_19572,N_19629);
xor UO_254 (O_254,N_19362,N_19994);
or UO_255 (O_255,N_19484,N_19329);
nor UO_256 (O_256,N_19817,N_19544);
nand UO_257 (O_257,N_19670,N_19207);
nand UO_258 (O_258,N_19931,N_19448);
or UO_259 (O_259,N_19487,N_19858);
and UO_260 (O_260,N_19685,N_19341);
or UO_261 (O_261,N_19844,N_19788);
nor UO_262 (O_262,N_19377,N_19941);
xnor UO_263 (O_263,N_19345,N_19631);
nor UO_264 (O_264,N_19691,N_19575);
nor UO_265 (O_265,N_19243,N_19700);
or UO_266 (O_266,N_19578,N_19898);
xnor UO_267 (O_267,N_19588,N_19576);
nor UO_268 (O_268,N_19628,N_19432);
and UO_269 (O_269,N_19446,N_19325);
nand UO_270 (O_270,N_19256,N_19756);
nor UO_271 (O_271,N_19742,N_19866);
nand UO_272 (O_272,N_19650,N_19813);
and UO_273 (O_273,N_19290,N_19638);
nor UO_274 (O_274,N_19603,N_19705);
nand UO_275 (O_275,N_19781,N_19564);
or UO_276 (O_276,N_19872,N_19673);
nor UO_277 (O_277,N_19732,N_19258);
nand UO_278 (O_278,N_19527,N_19679);
or UO_279 (O_279,N_19644,N_19437);
or UO_280 (O_280,N_19267,N_19798);
and UO_281 (O_281,N_19210,N_19860);
nand UO_282 (O_282,N_19667,N_19411);
or UO_283 (O_283,N_19233,N_19879);
nor UO_284 (O_284,N_19773,N_19661);
and UO_285 (O_285,N_19477,N_19332);
nor UO_286 (O_286,N_19799,N_19997);
nor UO_287 (O_287,N_19585,N_19455);
nand UO_288 (O_288,N_19676,N_19338);
nand UO_289 (O_289,N_19740,N_19539);
nor UO_290 (O_290,N_19468,N_19330);
or UO_291 (O_291,N_19647,N_19454);
or UO_292 (O_292,N_19272,N_19274);
xnor UO_293 (O_293,N_19753,N_19516);
nor UO_294 (O_294,N_19608,N_19457);
nor UO_295 (O_295,N_19481,N_19972);
nand UO_296 (O_296,N_19220,N_19714);
nor UO_297 (O_297,N_19702,N_19736);
or UO_298 (O_298,N_19488,N_19664);
nand UO_299 (O_299,N_19776,N_19370);
nand UO_300 (O_300,N_19938,N_19369);
nand UO_301 (O_301,N_19495,N_19419);
or UO_302 (O_302,N_19724,N_19250);
xnor UO_303 (O_303,N_19848,N_19835);
xor UO_304 (O_304,N_19819,N_19390);
xnor UO_305 (O_305,N_19248,N_19284);
nand UO_306 (O_306,N_19690,N_19587);
and UO_307 (O_307,N_19853,N_19549);
xor UO_308 (O_308,N_19877,N_19824);
nand UO_309 (O_309,N_19926,N_19780);
and UO_310 (O_310,N_19597,N_19874);
xor UO_311 (O_311,N_19212,N_19470);
or UO_312 (O_312,N_19567,N_19583);
or UO_313 (O_313,N_19990,N_19725);
and UO_314 (O_314,N_19720,N_19683);
and UO_315 (O_315,N_19491,N_19792);
nand UO_316 (O_316,N_19837,N_19472);
nor UO_317 (O_317,N_19460,N_19762);
and UO_318 (O_318,N_19613,N_19254);
and UO_319 (O_319,N_19855,N_19981);
nor UO_320 (O_320,N_19545,N_19985);
and UO_321 (O_321,N_19509,N_19610);
nor UO_322 (O_322,N_19444,N_19891);
xnor UO_323 (O_323,N_19962,N_19445);
or UO_324 (O_324,N_19228,N_19407);
or UO_325 (O_325,N_19335,N_19417);
or UO_326 (O_326,N_19769,N_19707);
and UO_327 (O_327,N_19741,N_19289);
or UO_328 (O_328,N_19313,N_19738);
or UO_329 (O_329,N_19452,N_19236);
xnor UO_330 (O_330,N_19354,N_19635);
and UO_331 (O_331,N_19515,N_19961);
nand UO_332 (O_332,N_19548,N_19573);
or UO_333 (O_333,N_19658,N_19845);
or UO_334 (O_334,N_19704,N_19899);
or UO_335 (O_335,N_19924,N_19378);
nor UO_336 (O_336,N_19371,N_19901);
nor UO_337 (O_337,N_19774,N_19934);
nand UO_338 (O_338,N_19453,N_19727);
nand UO_339 (O_339,N_19953,N_19677);
and UO_340 (O_340,N_19294,N_19984);
nor UO_341 (O_341,N_19580,N_19852);
or UO_342 (O_342,N_19543,N_19922);
nand UO_343 (O_343,N_19728,N_19841);
and UO_344 (O_344,N_19751,N_19949);
and UO_345 (O_345,N_19863,N_19717);
nor UO_346 (O_346,N_19602,N_19689);
nand UO_347 (O_347,N_19447,N_19615);
or UO_348 (O_348,N_19552,N_19241);
nor UO_349 (O_349,N_19708,N_19281);
nor UO_350 (O_350,N_19964,N_19627);
nor UO_351 (O_351,N_19565,N_19499);
nor UO_352 (O_352,N_19843,N_19409);
nand UO_353 (O_353,N_19657,N_19971);
nor UO_354 (O_354,N_19761,N_19989);
nor UO_355 (O_355,N_19993,N_19645);
or UO_356 (O_356,N_19293,N_19554);
and UO_357 (O_357,N_19715,N_19496);
and UO_358 (O_358,N_19584,N_19430);
nand UO_359 (O_359,N_19490,N_19754);
nor UO_360 (O_360,N_19992,N_19968);
xnor UO_361 (O_361,N_19317,N_19794);
xnor UO_362 (O_362,N_19697,N_19478);
and UO_363 (O_363,N_19282,N_19541);
xnor UO_364 (O_364,N_19201,N_19471);
and UO_365 (O_365,N_19744,N_19800);
and UO_366 (O_366,N_19246,N_19249);
and UO_367 (O_367,N_19480,N_19665);
nor UO_368 (O_368,N_19376,N_19688);
nor UO_369 (O_369,N_19546,N_19737);
xnor UO_370 (O_370,N_19966,N_19451);
and UO_371 (O_371,N_19777,N_19710);
or UO_372 (O_372,N_19895,N_19999);
nand UO_373 (O_373,N_19980,N_19261);
and UO_374 (O_374,N_19538,N_19483);
or UO_375 (O_375,N_19826,N_19392);
or UO_376 (O_376,N_19882,N_19213);
nand UO_377 (O_377,N_19620,N_19449);
and UO_378 (O_378,N_19846,N_19935);
xnor UO_379 (O_379,N_19266,N_19722);
nand UO_380 (O_380,N_19224,N_19219);
and UO_381 (O_381,N_19394,N_19331);
and UO_382 (O_382,N_19532,N_19929);
nor UO_383 (O_383,N_19269,N_19402);
nor UO_384 (O_384,N_19974,N_19913);
xnor UO_385 (O_385,N_19553,N_19486);
and UO_386 (O_386,N_19745,N_19461);
and UO_387 (O_387,N_19467,N_19987);
xor UO_388 (O_388,N_19801,N_19474);
nor UO_389 (O_389,N_19500,N_19391);
nand UO_390 (O_390,N_19768,N_19642);
and UO_391 (O_391,N_19618,N_19729);
or UO_392 (O_392,N_19680,N_19230);
nand UO_393 (O_393,N_19808,N_19351);
xnor UO_394 (O_394,N_19316,N_19633);
and UO_395 (O_395,N_19334,N_19465);
nand UO_396 (O_396,N_19703,N_19952);
nor UO_397 (O_397,N_19206,N_19599);
and UO_398 (O_398,N_19617,N_19512);
nor UO_399 (O_399,N_19221,N_19504);
xnor UO_400 (O_400,N_19454,N_19628);
xor UO_401 (O_401,N_19642,N_19997);
xnor UO_402 (O_402,N_19258,N_19806);
nand UO_403 (O_403,N_19926,N_19864);
nor UO_404 (O_404,N_19880,N_19746);
xor UO_405 (O_405,N_19260,N_19761);
or UO_406 (O_406,N_19286,N_19530);
and UO_407 (O_407,N_19658,N_19481);
or UO_408 (O_408,N_19300,N_19765);
or UO_409 (O_409,N_19259,N_19923);
nand UO_410 (O_410,N_19853,N_19783);
and UO_411 (O_411,N_19823,N_19308);
nand UO_412 (O_412,N_19442,N_19335);
or UO_413 (O_413,N_19401,N_19896);
or UO_414 (O_414,N_19988,N_19315);
or UO_415 (O_415,N_19282,N_19268);
nor UO_416 (O_416,N_19708,N_19565);
or UO_417 (O_417,N_19931,N_19218);
nand UO_418 (O_418,N_19998,N_19394);
xnor UO_419 (O_419,N_19258,N_19929);
nor UO_420 (O_420,N_19373,N_19900);
and UO_421 (O_421,N_19759,N_19752);
and UO_422 (O_422,N_19255,N_19376);
or UO_423 (O_423,N_19670,N_19310);
xor UO_424 (O_424,N_19325,N_19372);
xor UO_425 (O_425,N_19492,N_19380);
xnor UO_426 (O_426,N_19550,N_19580);
xnor UO_427 (O_427,N_19696,N_19499);
xor UO_428 (O_428,N_19787,N_19765);
nor UO_429 (O_429,N_19426,N_19894);
nor UO_430 (O_430,N_19382,N_19432);
xor UO_431 (O_431,N_19873,N_19677);
nand UO_432 (O_432,N_19667,N_19315);
or UO_433 (O_433,N_19753,N_19965);
and UO_434 (O_434,N_19555,N_19659);
or UO_435 (O_435,N_19410,N_19796);
nor UO_436 (O_436,N_19352,N_19906);
or UO_437 (O_437,N_19582,N_19869);
or UO_438 (O_438,N_19980,N_19902);
nor UO_439 (O_439,N_19215,N_19300);
xor UO_440 (O_440,N_19805,N_19315);
and UO_441 (O_441,N_19850,N_19796);
or UO_442 (O_442,N_19200,N_19376);
and UO_443 (O_443,N_19907,N_19414);
xor UO_444 (O_444,N_19343,N_19223);
or UO_445 (O_445,N_19284,N_19448);
xnor UO_446 (O_446,N_19514,N_19648);
and UO_447 (O_447,N_19827,N_19437);
nand UO_448 (O_448,N_19754,N_19918);
and UO_449 (O_449,N_19946,N_19736);
xor UO_450 (O_450,N_19313,N_19937);
xnor UO_451 (O_451,N_19961,N_19940);
nand UO_452 (O_452,N_19519,N_19308);
nor UO_453 (O_453,N_19276,N_19775);
xnor UO_454 (O_454,N_19754,N_19433);
nor UO_455 (O_455,N_19777,N_19630);
nor UO_456 (O_456,N_19249,N_19571);
nand UO_457 (O_457,N_19853,N_19648);
and UO_458 (O_458,N_19760,N_19777);
or UO_459 (O_459,N_19930,N_19833);
and UO_460 (O_460,N_19272,N_19475);
nor UO_461 (O_461,N_19403,N_19290);
and UO_462 (O_462,N_19556,N_19340);
xor UO_463 (O_463,N_19483,N_19933);
nor UO_464 (O_464,N_19280,N_19615);
nand UO_465 (O_465,N_19200,N_19595);
and UO_466 (O_466,N_19743,N_19429);
or UO_467 (O_467,N_19236,N_19605);
and UO_468 (O_468,N_19431,N_19444);
nor UO_469 (O_469,N_19891,N_19732);
and UO_470 (O_470,N_19900,N_19846);
or UO_471 (O_471,N_19678,N_19417);
or UO_472 (O_472,N_19912,N_19941);
xor UO_473 (O_473,N_19291,N_19966);
or UO_474 (O_474,N_19860,N_19548);
nor UO_475 (O_475,N_19482,N_19303);
and UO_476 (O_476,N_19225,N_19912);
nand UO_477 (O_477,N_19923,N_19993);
nor UO_478 (O_478,N_19289,N_19487);
nand UO_479 (O_479,N_19693,N_19357);
and UO_480 (O_480,N_19893,N_19977);
or UO_481 (O_481,N_19253,N_19728);
nand UO_482 (O_482,N_19487,N_19892);
or UO_483 (O_483,N_19231,N_19208);
xor UO_484 (O_484,N_19807,N_19274);
nand UO_485 (O_485,N_19205,N_19862);
nor UO_486 (O_486,N_19550,N_19764);
nand UO_487 (O_487,N_19787,N_19301);
or UO_488 (O_488,N_19453,N_19882);
or UO_489 (O_489,N_19542,N_19635);
nand UO_490 (O_490,N_19780,N_19984);
or UO_491 (O_491,N_19740,N_19252);
xnor UO_492 (O_492,N_19660,N_19869);
xnor UO_493 (O_493,N_19260,N_19379);
and UO_494 (O_494,N_19676,N_19320);
and UO_495 (O_495,N_19384,N_19222);
and UO_496 (O_496,N_19835,N_19487);
nand UO_497 (O_497,N_19829,N_19824);
or UO_498 (O_498,N_19317,N_19930);
nor UO_499 (O_499,N_19879,N_19960);
or UO_500 (O_500,N_19823,N_19674);
and UO_501 (O_501,N_19648,N_19457);
or UO_502 (O_502,N_19226,N_19852);
nand UO_503 (O_503,N_19290,N_19487);
xnor UO_504 (O_504,N_19583,N_19560);
nor UO_505 (O_505,N_19576,N_19590);
nand UO_506 (O_506,N_19736,N_19859);
or UO_507 (O_507,N_19790,N_19297);
xor UO_508 (O_508,N_19863,N_19450);
xor UO_509 (O_509,N_19593,N_19963);
xor UO_510 (O_510,N_19981,N_19433);
xor UO_511 (O_511,N_19421,N_19410);
xnor UO_512 (O_512,N_19670,N_19999);
xnor UO_513 (O_513,N_19725,N_19970);
nor UO_514 (O_514,N_19304,N_19880);
or UO_515 (O_515,N_19985,N_19660);
xor UO_516 (O_516,N_19688,N_19568);
nand UO_517 (O_517,N_19822,N_19260);
nand UO_518 (O_518,N_19636,N_19885);
and UO_519 (O_519,N_19850,N_19745);
nor UO_520 (O_520,N_19607,N_19407);
nor UO_521 (O_521,N_19331,N_19365);
nand UO_522 (O_522,N_19531,N_19216);
xnor UO_523 (O_523,N_19513,N_19748);
or UO_524 (O_524,N_19390,N_19583);
nor UO_525 (O_525,N_19407,N_19317);
nand UO_526 (O_526,N_19479,N_19793);
and UO_527 (O_527,N_19617,N_19838);
or UO_528 (O_528,N_19924,N_19224);
or UO_529 (O_529,N_19574,N_19445);
nor UO_530 (O_530,N_19373,N_19593);
nor UO_531 (O_531,N_19425,N_19493);
xnor UO_532 (O_532,N_19722,N_19438);
xnor UO_533 (O_533,N_19781,N_19829);
nand UO_534 (O_534,N_19792,N_19974);
xor UO_535 (O_535,N_19758,N_19532);
nand UO_536 (O_536,N_19605,N_19927);
nand UO_537 (O_537,N_19391,N_19886);
nand UO_538 (O_538,N_19975,N_19971);
xor UO_539 (O_539,N_19735,N_19878);
nand UO_540 (O_540,N_19720,N_19269);
xnor UO_541 (O_541,N_19742,N_19898);
nor UO_542 (O_542,N_19276,N_19325);
nand UO_543 (O_543,N_19325,N_19725);
xnor UO_544 (O_544,N_19302,N_19312);
nand UO_545 (O_545,N_19314,N_19766);
and UO_546 (O_546,N_19759,N_19373);
and UO_547 (O_547,N_19954,N_19607);
or UO_548 (O_548,N_19962,N_19559);
and UO_549 (O_549,N_19789,N_19451);
or UO_550 (O_550,N_19925,N_19331);
and UO_551 (O_551,N_19645,N_19523);
nor UO_552 (O_552,N_19428,N_19213);
nand UO_553 (O_553,N_19489,N_19496);
nand UO_554 (O_554,N_19594,N_19343);
and UO_555 (O_555,N_19699,N_19968);
xor UO_556 (O_556,N_19726,N_19633);
xor UO_557 (O_557,N_19677,N_19820);
nor UO_558 (O_558,N_19476,N_19912);
nor UO_559 (O_559,N_19216,N_19596);
xnor UO_560 (O_560,N_19459,N_19356);
xor UO_561 (O_561,N_19780,N_19718);
nand UO_562 (O_562,N_19306,N_19417);
or UO_563 (O_563,N_19228,N_19482);
and UO_564 (O_564,N_19550,N_19430);
or UO_565 (O_565,N_19615,N_19834);
xor UO_566 (O_566,N_19805,N_19661);
and UO_567 (O_567,N_19548,N_19769);
nand UO_568 (O_568,N_19789,N_19532);
nor UO_569 (O_569,N_19313,N_19484);
or UO_570 (O_570,N_19396,N_19975);
nand UO_571 (O_571,N_19906,N_19253);
or UO_572 (O_572,N_19784,N_19202);
nand UO_573 (O_573,N_19277,N_19762);
or UO_574 (O_574,N_19459,N_19825);
and UO_575 (O_575,N_19986,N_19660);
or UO_576 (O_576,N_19849,N_19695);
or UO_577 (O_577,N_19313,N_19762);
nand UO_578 (O_578,N_19290,N_19457);
xnor UO_579 (O_579,N_19845,N_19778);
xor UO_580 (O_580,N_19387,N_19353);
xnor UO_581 (O_581,N_19639,N_19254);
xor UO_582 (O_582,N_19539,N_19967);
and UO_583 (O_583,N_19877,N_19349);
nand UO_584 (O_584,N_19907,N_19371);
nor UO_585 (O_585,N_19541,N_19648);
and UO_586 (O_586,N_19694,N_19685);
xnor UO_587 (O_587,N_19915,N_19264);
nor UO_588 (O_588,N_19328,N_19309);
xor UO_589 (O_589,N_19819,N_19957);
nor UO_590 (O_590,N_19910,N_19388);
nor UO_591 (O_591,N_19651,N_19224);
nor UO_592 (O_592,N_19922,N_19875);
nor UO_593 (O_593,N_19659,N_19738);
nor UO_594 (O_594,N_19561,N_19993);
nand UO_595 (O_595,N_19844,N_19606);
xnor UO_596 (O_596,N_19774,N_19773);
xnor UO_597 (O_597,N_19761,N_19288);
nor UO_598 (O_598,N_19302,N_19203);
xor UO_599 (O_599,N_19289,N_19922);
or UO_600 (O_600,N_19487,N_19631);
and UO_601 (O_601,N_19977,N_19422);
or UO_602 (O_602,N_19590,N_19699);
xnor UO_603 (O_603,N_19978,N_19903);
xnor UO_604 (O_604,N_19534,N_19477);
nand UO_605 (O_605,N_19325,N_19415);
or UO_606 (O_606,N_19628,N_19771);
or UO_607 (O_607,N_19697,N_19552);
nand UO_608 (O_608,N_19207,N_19972);
or UO_609 (O_609,N_19305,N_19283);
or UO_610 (O_610,N_19262,N_19778);
nand UO_611 (O_611,N_19321,N_19747);
xor UO_612 (O_612,N_19223,N_19381);
nor UO_613 (O_613,N_19273,N_19292);
xnor UO_614 (O_614,N_19615,N_19537);
xnor UO_615 (O_615,N_19338,N_19373);
nand UO_616 (O_616,N_19508,N_19493);
nand UO_617 (O_617,N_19664,N_19895);
nor UO_618 (O_618,N_19634,N_19261);
nor UO_619 (O_619,N_19709,N_19466);
and UO_620 (O_620,N_19700,N_19240);
or UO_621 (O_621,N_19647,N_19919);
nor UO_622 (O_622,N_19914,N_19967);
or UO_623 (O_623,N_19720,N_19897);
and UO_624 (O_624,N_19626,N_19533);
xor UO_625 (O_625,N_19906,N_19931);
xnor UO_626 (O_626,N_19279,N_19830);
nand UO_627 (O_627,N_19941,N_19457);
xnor UO_628 (O_628,N_19360,N_19920);
nand UO_629 (O_629,N_19408,N_19833);
and UO_630 (O_630,N_19487,N_19484);
nor UO_631 (O_631,N_19706,N_19699);
nor UO_632 (O_632,N_19605,N_19756);
and UO_633 (O_633,N_19600,N_19620);
or UO_634 (O_634,N_19573,N_19671);
nor UO_635 (O_635,N_19996,N_19809);
and UO_636 (O_636,N_19753,N_19400);
nand UO_637 (O_637,N_19244,N_19715);
nor UO_638 (O_638,N_19360,N_19251);
nor UO_639 (O_639,N_19954,N_19713);
xor UO_640 (O_640,N_19443,N_19725);
nand UO_641 (O_641,N_19793,N_19330);
nor UO_642 (O_642,N_19245,N_19945);
and UO_643 (O_643,N_19474,N_19583);
nor UO_644 (O_644,N_19307,N_19276);
nand UO_645 (O_645,N_19951,N_19282);
nor UO_646 (O_646,N_19888,N_19528);
and UO_647 (O_647,N_19397,N_19415);
nor UO_648 (O_648,N_19598,N_19247);
or UO_649 (O_649,N_19861,N_19750);
or UO_650 (O_650,N_19604,N_19265);
nand UO_651 (O_651,N_19868,N_19743);
and UO_652 (O_652,N_19950,N_19580);
nor UO_653 (O_653,N_19960,N_19584);
or UO_654 (O_654,N_19961,N_19701);
and UO_655 (O_655,N_19676,N_19335);
nand UO_656 (O_656,N_19855,N_19202);
or UO_657 (O_657,N_19849,N_19844);
nand UO_658 (O_658,N_19836,N_19772);
xnor UO_659 (O_659,N_19682,N_19699);
or UO_660 (O_660,N_19269,N_19369);
nand UO_661 (O_661,N_19777,N_19977);
and UO_662 (O_662,N_19409,N_19864);
and UO_663 (O_663,N_19974,N_19873);
nor UO_664 (O_664,N_19432,N_19725);
or UO_665 (O_665,N_19303,N_19495);
xnor UO_666 (O_666,N_19641,N_19915);
nor UO_667 (O_667,N_19802,N_19894);
xor UO_668 (O_668,N_19875,N_19495);
nand UO_669 (O_669,N_19202,N_19631);
nand UO_670 (O_670,N_19930,N_19480);
nand UO_671 (O_671,N_19791,N_19437);
nor UO_672 (O_672,N_19872,N_19295);
xnor UO_673 (O_673,N_19277,N_19239);
xor UO_674 (O_674,N_19591,N_19640);
or UO_675 (O_675,N_19244,N_19939);
and UO_676 (O_676,N_19713,N_19901);
xor UO_677 (O_677,N_19373,N_19402);
or UO_678 (O_678,N_19436,N_19295);
or UO_679 (O_679,N_19922,N_19821);
nand UO_680 (O_680,N_19710,N_19891);
nand UO_681 (O_681,N_19287,N_19282);
or UO_682 (O_682,N_19949,N_19327);
or UO_683 (O_683,N_19539,N_19459);
and UO_684 (O_684,N_19216,N_19632);
nor UO_685 (O_685,N_19887,N_19953);
and UO_686 (O_686,N_19720,N_19446);
and UO_687 (O_687,N_19240,N_19948);
nand UO_688 (O_688,N_19872,N_19568);
or UO_689 (O_689,N_19670,N_19465);
or UO_690 (O_690,N_19659,N_19824);
xor UO_691 (O_691,N_19879,N_19985);
and UO_692 (O_692,N_19580,N_19910);
and UO_693 (O_693,N_19431,N_19521);
xor UO_694 (O_694,N_19317,N_19257);
and UO_695 (O_695,N_19260,N_19475);
or UO_696 (O_696,N_19737,N_19340);
xor UO_697 (O_697,N_19702,N_19232);
xnor UO_698 (O_698,N_19483,N_19404);
nand UO_699 (O_699,N_19546,N_19265);
xor UO_700 (O_700,N_19972,N_19290);
nand UO_701 (O_701,N_19253,N_19403);
nand UO_702 (O_702,N_19750,N_19486);
nand UO_703 (O_703,N_19777,N_19381);
and UO_704 (O_704,N_19525,N_19439);
or UO_705 (O_705,N_19826,N_19905);
and UO_706 (O_706,N_19555,N_19224);
nand UO_707 (O_707,N_19522,N_19918);
nand UO_708 (O_708,N_19371,N_19625);
or UO_709 (O_709,N_19433,N_19356);
nor UO_710 (O_710,N_19801,N_19384);
nor UO_711 (O_711,N_19693,N_19537);
or UO_712 (O_712,N_19284,N_19270);
or UO_713 (O_713,N_19332,N_19468);
or UO_714 (O_714,N_19253,N_19913);
and UO_715 (O_715,N_19663,N_19329);
nand UO_716 (O_716,N_19559,N_19800);
nand UO_717 (O_717,N_19458,N_19229);
or UO_718 (O_718,N_19224,N_19666);
nand UO_719 (O_719,N_19814,N_19629);
nor UO_720 (O_720,N_19545,N_19293);
or UO_721 (O_721,N_19752,N_19852);
or UO_722 (O_722,N_19257,N_19541);
and UO_723 (O_723,N_19382,N_19402);
or UO_724 (O_724,N_19265,N_19202);
nor UO_725 (O_725,N_19551,N_19843);
nor UO_726 (O_726,N_19266,N_19481);
nor UO_727 (O_727,N_19379,N_19610);
or UO_728 (O_728,N_19746,N_19517);
xor UO_729 (O_729,N_19909,N_19304);
and UO_730 (O_730,N_19239,N_19800);
nor UO_731 (O_731,N_19682,N_19322);
nand UO_732 (O_732,N_19816,N_19272);
and UO_733 (O_733,N_19332,N_19308);
xnor UO_734 (O_734,N_19235,N_19313);
or UO_735 (O_735,N_19493,N_19502);
or UO_736 (O_736,N_19665,N_19221);
and UO_737 (O_737,N_19447,N_19235);
nand UO_738 (O_738,N_19786,N_19366);
nor UO_739 (O_739,N_19776,N_19536);
xnor UO_740 (O_740,N_19549,N_19316);
nand UO_741 (O_741,N_19301,N_19342);
xnor UO_742 (O_742,N_19614,N_19404);
xnor UO_743 (O_743,N_19714,N_19701);
or UO_744 (O_744,N_19608,N_19407);
nand UO_745 (O_745,N_19471,N_19315);
nor UO_746 (O_746,N_19349,N_19205);
nor UO_747 (O_747,N_19594,N_19572);
or UO_748 (O_748,N_19660,N_19433);
nor UO_749 (O_749,N_19883,N_19972);
nand UO_750 (O_750,N_19689,N_19447);
or UO_751 (O_751,N_19223,N_19613);
nand UO_752 (O_752,N_19785,N_19605);
and UO_753 (O_753,N_19526,N_19955);
nor UO_754 (O_754,N_19252,N_19626);
and UO_755 (O_755,N_19621,N_19692);
and UO_756 (O_756,N_19342,N_19461);
xnor UO_757 (O_757,N_19334,N_19748);
xnor UO_758 (O_758,N_19551,N_19918);
xnor UO_759 (O_759,N_19421,N_19647);
or UO_760 (O_760,N_19683,N_19427);
nor UO_761 (O_761,N_19919,N_19783);
nand UO_762 (O_762,N_19609,N_19765);
xor UO_763 (O_763,N_19858,N_19788);
or UO_764 (O_764,N_19768,N_19359);
and UO_765 (O_765,N_19585,N_19746);
xor UO_766 (O_766,N_19830,N_19361);
nand UO_767 (O_767,N_19218,N_19948);
or UO_768 (O_768,N_19960,N_19633);
and UO_769 (O_769,N_19792,N_19947);
nand UO_770 (O_770,N_19922,N_19478);
and UO_771 (O_771,N_19273,N_19753);
nand UO_772 (O_772,N_19808,N_19219);
xnor UO_773 (O_773,N_19536,N_19417);
or UO_774 (O_774,N_19752,N_19445);
and UO_775 (O_775,N_19394,N_19629);
or UO_776 (O_776,N_19595,N_19980);
and UO_777 (O_777,N_19701,N_19408);
nand UO_778 (O_778,N_19449,N_19829);
or UO_779 (O_779,N_19434,N_19964);
or UO_780 (O_780,N_19365,N_19227);
or UO_781 (O_781,N_19463,N_19284);
or UO_782 (O_782,N_19372,N_19395);
and UO_783 (O_783,N_19870,N_19461);
or UO_784 (O_784,N_19481,N_19339);
nand UO_785 (O_785,N_19263,N_19602);
nand UO_786 (O_786,N_19960,N_19256);
or UO_787 (O_787,N_19214,N_19786);
and UO_788 (O_788,N_19909,N_19551);
and UO_789 (O_789,N_19229,N_19355);
nor UO_790 (O_790,N_19955,N_19727);
nand UO_791 (O_791,N_19987,N_19526);
nor UO_792 (O_792,N_19220,N_19739);
nand UO_793 (O_793,N_19987,N_19952);
or UO_794 (O_794,N_19881,N_19934);
xnor UO_795 (O_795,N_19865,N_19727);
nand UO_796 (O_796,N_19804,N_19582);
nand UO_797 (O_797,N_19776,N_19527);
xor UO_798 (O_798,N_19820,N_19461);
and UO_799 (O_799,N_19717,N_19256);
and UO_800 (O_800,N_19679,N_19545);
nor UO_801 (O_801,N_19431,N_19614);
nand UO_802 (O_802,N_19912,N_19404);
or UO_803 (O_803,N_19734,N_19454);
xnor UO_804 (O_804,N_19413,N_19923);
nand UO_805 (O_805,N_19461,N_19624);
nor UO_806 (O_806,N_19617,N_19995);
or UO_807 (O_807,N_19367,N_19445);
nor UO_808 (O_808,N_19329,N_19268);
xor UO_809 (O_809,N_19977,N_19670);
nand UO_810 (O_810,N_19571,N_19272);
and UO_811 (O_811,N_19445,N_19891);
nand UO_812 (O_812,N_19701,N_19563);
nand UO_813 (O_813,N_19295,N_19631);
or UO_814 (O_814,N_19809,N_19360);
or UO_815 (O_815,N_19866,N_19753);
nor UO_816 (O_816,N_19435,N_19831);
nand UO_817 (O_817,N_19867,N_19205);
xnor UO_818 (O_818,N_19736,N_19209);
nand UO_819 (O_819,N_19756,N_19203);
or UO_820 (O_820,N_19387,N_19451);
nor UO_821 (O_821,N_19892,N_19265);
or UO_822 (O_822,N_19319,N_19650);
or UO_823 (O_823,N_19583,N_19329);
nor UO_824 (O_824,N_19616,N_19326);
or UO_825 (O_825,N_19959,N_19327);
nand UO_826 (O_826,N_19621,N_19948);
xnor UO_827 (O_827,N_19509,N_19713);
nand UO_828 (O_828,N_19383,N_19241);
nand UO_829 (O_829,N_19932,N_19902);
nand UO_830 (O_830,N_19839,N_19981);
or UO_831 (O_831,N_19877,N_19508);
nand UO_832 (O_832,N_19368,N_19291);
and UO_833 (O_833,N_19455,N_19982);
nand UO_834 (O_834,N_19438,N_19380);
and UO_835 (O_835,N_19696,N_19780);
xor UO_836 (O_836,N_19637,N_19691);
xor UO_837 (O_837,N_19988,N_19340);
nor UO_838 (O_838,N_19804,N_19389);
nor UO_839 (O_839,N_19903,N_19513);
and UO_840 (O_840,N_19369,N_19854);
or UO_841 (O_841,N_19403,N_19987);
and UO_842 (O_842,N_19672,N_19859);
nand UO_843 (O_843,N_19295,N_19610);
xor UO_844 (O_844,N_19209,N_19812);
or UO_845 (O_845,N_19767,N_19871);
or UO_846 (O_846,N_19609,N_19280);
xnor UO_847 (O_847,N_19993,N_19822);
or UO_848 (O_848,N_19906,N_19959);
nor UO_849 (O_849,N_19433,N_19939);
and UO_850 (O_850,N_19456,N_19539);
or UO_851 (O_851,N_19785,N_19758);
or UO_852 (O_852,N_19966,N_19641);
and UO_853 (O_853,N_19214,N_19763);
and UO_854 (O_854,N_19662,N_19476);
xor UO_855 (O_855,N_19903,N_19645);
xor UO_856 (O_856,N_19410,N_19432);
nand UO_857 (O_857,N_19880,N_19707);
and UO_858 (O_858,N_19474,N_19448);
nand UO_859 (O_859,N_19466,N_19837);
xor UO_860 (O_860,N_19565,N_19420);
xor UO_861 (O_861,N_19526,N_19697);
xnor UO_862 (O_862,N_19615,N_19628);
and UO_863 (O_863,N_19713,N_19897);
and UO_864 (O_864,N_19682,N_19795);
nor UO_865 (O_865,N_19829,N_19535);
or UO_866 (O_866,N_19367,N_19264);
and UO_867 (O_867,N_19651,N_19371);
nor UO_868 (O_868,N_19428,N_19970);
nor UO_869 (O_869,N_19923,N_19253);
xnor UO_870 (O_870,N_19686,N_19893);
nor UO_871 (O_871,N_19613,N_19915);
nor UO_872 (O_872,N_19396,N_19247);
or UO_873 (O_873,N_19810,N_19699);
and UO_874 (O_874,N_19831,N_19680);
nand UO_875 (O_875,N_19232,N_19917);
nor UO_876 (O_876,N_19958,N_19549);
or UO_877 (O_877,N_19804,N_19896);
nor UO_878 (O_878,N_19389,N_19796);
xor UO_879 (O_879,N_19286,N_19503);
nand UO_880 (O_880,N_19529,N_19860);
or UO_881 (O_881,N_19689,N_19856);
xnor UO_882 (O_882,N_19930,N_19579);
and UO_883 (O_883,N_19559,N_19413);
nor UO_884 (O_884,N_19783,N_19657);
xnor UO_885 (O_885,N_19306,N_19628);
and UO_886 (O_886,N_19619,N_19591);
and UO_887 (O_887,N_19651,N_19940);
nor UO_888 (O_888,N_19798,N_19274);
or UO_889 (O_889,N_19960,N_19278);
or UO_890 (O_890,N_19457,N_19317);
or UO_891 (O_891,N_19454,N_19799);
nand UO_892 (O_892,N_19305,N_19378);
nand UO_893 (O_893,N_19631,N_19891);
nand UO_894 (O_894,N_19987,N_19477);
nand UO_895 (O_895,N_19342,N_19489);
nand UO_896 (O_896,N_19339,N_19270);
or UO_897 (O_897,N_19568,N_19802);
xnor UO_898 (O_898,N_19714,N_19781);
xor UO_899 (O_899,N_19706,N_19814);
and UO_900 (O_900,N_19614,N_19627);
nor UO_901 (O_901,N_19247,N_19480);
xor UO_902 (O_902,N_19668,N_19482);
nor UO_903 (O_903,N_19516,N_19304);
or UO_904 (O_904,N_19834,N_19216);
nand UO_905 (O_905,N_19818,N_19357);
nand UO_906 (O_906,N_19521,N_19567);
and UO_907 (O_907,N_19902,N_19839);
xnor UO_908 (O_908,N_19634,N_19862);
nor UO_909 (O_909,N_19614,N_19802);
or UO_910 (O_910,N_19251,N_19728);
xnor UO_911 (O_911,N_19336,N_19203);
nor UO_912 (O_912,N_19313,N_19460);
and UO_913 (O_913,N_19400,N_19409);
or UO_914 (O_914,N_19718,N_19600);
or UO_915 (O_915,N_19797,N_19858);
nor UO_916 (O_916,N_19741,N_19672);
xnor UO_917 (O_917,N_19200,N_19423);
or UO_918 (O_918,N_19226,N_19668);
xor UO_919 (O_919,N_19233,N_19460);
and UO_920 (O_920,N_19851,N_19419);
or UO_921 (O_921,N_19389,N_19857);
and UO_922 (O_922,N_19345,N_19589);
nor UO_923 (O_923,N_19683,N_19536);
nand UO_924 (O_924,N_19476,N_19837);
or UO_925 (O_925,N_19329,N_19660);
xnor UO_926 (O_926,N_19548,N_19431);
nand UO_927 (O_927,N_19831,N_19340);
nand UO_928 (O_928,N_19257,N_19547);
nor UO_929 (O_929,N_19876,N_19323);
xnor UO_930 (O_930,N_19244,N_19352);
nor UO_931 (O_931,N_19497,N_19647);
and UO_932 (O_932,N_19385,N_19527);
and UO_933 (O_933,N_19833,N_19330);
or UO_934 (O_934,N_19219,N_19839);
nand UO_935 (O_935,N_19794,N_19427);
or UO_936 (O_936,N_19292,N_19823);
and UO_937 (O_937,N_19840,N_19592);
nor UO_938 (O_938,N_19881,N_19532);
and UO_939 (O_939,N_19395,N_19359);
and UO_940 (O_940,N_19858,N_19220);
or UO_941 (O_941,N_19935,N_19498);
xor UO_942 (O_942,N_19701,N_19343);
or UO_943 (O_943,N_19300,N_19293);
or UO_944 (O_944,N_19386,N_19796);
or UO_945 (O_945,N_19262,N_19354);
xor UO_946 (O_946,N_19967,N_19907);
nand UO_947 (O_947,N_19519,N_19532);
nand UO_948 (O_948,N_19544,N_19664);
and UO_949 (O_949,N_19893,N_19497);
xnor UO_950 (O_950,N_19970,N_19818);
and UO_951 (O_951,N_19313,N_19362);
nand UO_952 (O_952,N_19298,N_19734);
nand UO_953 (O_953,N_19345,N_19358);
nor UO_954 (O_954,N_19603,N_19783);
nor UO_955 (O_955,N_19730,N_19800);
and UO_956 (O_956,N_19795,N_19352);
nand UO_957 (O_957,N_19833,N_19710);
or UO_958 (O_958,N_19852,N_19203);
nor UO_959 (O_959,N_19669,N_19639);
nand UO_960 (O_960,N_19794,N_19334);
and UO_961 (O_961,N_19598,N_19692);
xnor UO_962 (O_962,N_19220,N_19888);
or UO_963 (O_963,N_19431,N_19466);
and UO_964 (O_964,N_19882,N_19377);
and UO_965 (O_965,N_19225,N_19593);
nand UO_966 (O_966,N_19486,N_19490);
nor UO_967 (O_967,N_19211,N_19811);
nand UO_968 (O_968,N_19877,N_19718);
or UO_969 (O_969,N_19424,N_19798);
xnor UO_970 (O_970,N_19335,N_19541);
or UO_971 (O_971,N_19548,N_19355);
nor UO_972 (O_972,N_19697,N_19644);
or UO_973 (O_973,N_19474,N_19841);
nor UO_974 (O_974,N_19780,N_19860);
nand UO_975 (O_975,N_19351,N_19419);
nor UO_976 (O_976,N_19839,N_19540);
nor UO_977 (O_977,N_19249,N_19356);
nor UO_978 (O_978,N_19999,N_19367);
nor UO_979 (O_979,N_19422,N_19780);
nand UO_980 (O_980,N_19852,N_19787);
nand UO_981 (O_981,N_19886,N_19409);
nor UO_982 (O_982,N_19297,N_19863);
or UO_983 (O_983,N_19674,N_19626);
xor UO_984 (O_984,N_19543,N_19578);
nand UO_985 (O_985,N_19982,N_19225);
nor UO_986 (O_986,N_19603,N_19547);
nand UO_987 (O_987,N_19584,N_19226);
nor UO_988 (O_988,N_19678,N_19609);
xor UO_989 (O_989,N_19439,N_19748);
xor UO_990 (O_990,N_19371,N_19246);
and UO_991 (O_991,N_19473,N_19702);
nor UO_992 (O_992,N_19966,N_19375);
nand UO_993 (O_993,N_19968,N_19562);
and UO_994 (O_994,N_19437,N_19350);
nor UO_995 (O_995,N_19974,N_19640);
nor UO_996 (O_996,N_19834,N_19866);
or UO_997 (O_997,N_19881,N_19883);
nor UO_998 (O_998,N_19427,N_19502);
or UO_999 (O_999,N_19814,N_19480);
nand UO_1000 (O_1000,N_19421,N_19691);
nand UO_1001 (O_1001,N_19268,N_19633);
or UO_1002 (O_1002,N_19212,N_19414);
or UO_1003 (O_1003,N_19972,N_19202);
nor UO_1004 (O_1004,N_19866,N_19527);
nor UO_1005 (O_1005,N_19884,N_19312);
nor UO_1006 (O_1006,N_19760,N_19820);
xnor UO_1007 (O_1007,N_19575,N_19318);
and UO_1008 (O_1008,N_19353,N_19579);
nand UO_1009 (O_1009,N_19844,N_19824);
or UO_1010 (O_1010,N_19911,N_19767);
or UO_1011 (O_1011,N_19208,N_19792);
nor UO_1012 (O_1012,N_19400,N_19910);
nand UO_1013 (O_1013,N_19351,N_19857);
nand UO_1014 (O_1014,N_19859,N_19925);
nor UO_1015 (O_1015,N_19217,N_19655);
nor UO_1016 (O_1016,N_19931,N_19645);
nor UO_1017 (O_1017,N_19643,N_19575);
and UO_1018 (O_1018,N_19770,N_19874);
or UO_1019 (O_1019,N_19595,N_19524);
nand UO_1020 (O_1020,N_19573,N_19380);
and UO_1021 (O_1021,N_19825,N_19883);
nand UO_1022 (O_1022,N_19678,N_19891);
xnor UO_1023 (O_1023,N_19272,N_19948);
nand UO_1024 (O_1024,N_19605,N_19845);
nand UO_1025 (O_1025,N_19725,N_19536);
xnor UO_1026 (O_1026,N_19557,N_19297);
or UO_1027 (O_1027,N_19970,N_19863);
and UO_1028 (O_1028,N_19242,N_19833);
or UO_1029 (O_1029,N_19739,N_19287);
and UO_1030 (O_1030,N_19888,N_19757);
nand UO_1031 (O_1031,N_19720,N_19337);
or UO_1032 (O_1032,N_19851,N_19412);
xnor UO_1033 (O_1033,N_19677,N_19716);
nor UO_1034 (O_1034,N_19301,N_19862);
and UO_1035 (O_1035,N_19595,N_19885);
nor UO_1036 (O_1036,N_19642,N_19674);
or UO_1037 (O_1037,N_19762,N_19394);
nor UO_1038 (O_1038,N_19366,N_19319);
xor UO_1039 (O_1039,N_19245,N_19374);
nor UO_1040 (O_1040,N_19522,N_19570);
xnor UO_1041 (O_1041,N_19651,N_19699);
and UO_1042 (O_1042,N_19421,N_19572);
and UO_1043 (O_1043,N_19322,N_19407);
nor UO_1044 (O_1044,N_19443,N_19673);
or UO_1045 (O_1045,N_19503,N_19924);
or UO_1046 (O_1046,N_19844,N_19699);
nor UO_1047 (O_1047,N_19883,N_19364);
nor UO_1048 (O_1048,N_19399,N_19677);
or UO_1049 (O_1049,N_19990,N_19738);
nor UO_1050 (O_1050,N_19248,N_19218);
xor UO_1051 (O_1051,N_19267,N_19880);
nand UO_1052 (O_1052,N_19284,N_19304);
and UO_1053 (O_1053,N_19898,N_19758);
or UO_1054 (O_1054,N_19302,N_19625);
and UO_1055 (O_1055,N_19415,N_19315);
or UO_1056 (O_1056,N_19767,N_19430);
nand UO_1057 (O_1057,N_19367,N_19340);
nor UO_1058 (O_1058,N_19797,N_19906);
or UO_1059 (O_1059,N_19663,N_19368);
and UO_1060 (O_1060,N_19327,N_19973);
and UO_1061 (O_1061,N_19705,N_19926);
nand UO_1062 (O_1062,N_19389,N_19525);
or UO_1063 (O_1063,N_19808,N_19270);
nor UO_1064 (O_1064,N_19677,N_19649);
nor UO_1065 (O_1065,N_19670,N_19377);
nand UO_1066 (O_1066,N_19403,N_19516);
or UO_1067 (O_1067,N_19993,N_19880);
or UO_1068 (O_1068,N_19513,N_19812);
xor UO_1069 (O_1069,N_19887,N_19231);
nand UO_1070 (O_1070,N_19480,N_19589);
or UO_1071 (O_1071,N_19753,N_19459);
nor UO_1072 (O_1072,N_19519,N_19455);
nand UO_1073 (O_1073,N_19569,N_19876);
nor UO_1074 (O_1074,N_19989,N_19931);
and UO_1075 (O_1075,N_19464,N_19539);
nor UO_1076 (O_1076,N_19714,N_19821);
nand UO_1077 (O_1077,N_19468,N_19570);
nor UO_1078 (O_1078,N_19472,N_19313);
nand UO_1079 (O_1079,N_19552,N_19483);
xnor UO_1080 (O_1080,N_19676,N_19204);
nand UO_1081 (O_1081,N_19291,N_19448);
nand UO_1082 (O_1082,N_19989,N_19728);
nor UO_1083 (O_1083,N_19325,N_19859);
and UO_1084 (O_1084,N_19582,N_19224);
and UO_1085 (O_1085,N_19248,N_19604);
xnor UO_1086 (O_1086,N_19777,N_19913);
xnor UO_1087 (O_1087,N_19658,N_19478);
nand UO_1088 (O_1088,N_19656,N_19458);
xor UO_1089 (O_1089,N_19479,N_19359);
nor UO_1090 (O_1090,N_19798,N_19762);
nor UO_1091 (O_1091,N_19740,N_19511);
or UO_1092 (O_1092,N_19644,N_19290);
and UO_1093 (O_1093,N_19269,N_19528);
nand UO_1094 (O_1094,N_19959,N_19782);
or UO_1095 (O_1095,N_19460,N_19712);
xor UO_1096 (O_1096,N_19973,N_19453);
nand UO_1097 (O_1097,N_19689,N_19935);
xnor UO_1098 (O_1098,N_19879,N_19651);
nand UO_1099 (O_1099,N_19637,N_19405);
and UO_1100 (O_1100,N_19332,N_19427);
xnor UO_1101 (O_1101,N_19748,N_19905);
nor UO_1102 (O_1102,N_19831,N_19266);
and UO_1103 (O_1103,N_19675,N_19622);
xnor UO_1104 (O_1104,N_19530,N_19871);
nor UO_1105 (O_1105,N_19229,N_19617);
xnor UO_1106 (O_1106,N_19405,N_19814);
and UO_1107 (O_1107,N_19731,N_19568);
nand UO_1108 (O_1108,N_19895,N_19309);
nand UO_1109 (O_1109,N_19715,N_19942);
nor UO_1110 (O_1110,N_19549,N_19589);
nand UO_1111 (O_1111,N_19499,N_19804);
or UO_1112 (O_1112,N_19893,N_19470);
xor UO_1113 (O_1113,N_19242,N_19320);
xor UO_1114 (O_1114,N_19904,N_19694);
and UO_1115 (O_1115,N_19218,N_19265);
xor UO_1116 (O_1116,N_19374,N_19459);
xor UO_1117 (O_1117,N_19843,N_19426);
nor UO_1118 (O_1118,N_19834,N_19809);
nand UO_1119 (O_1119,N_19241,N_19231);
or UO_1120 (O_1120,N_19730,N_19770);
and UO_1121 (O_1121,N_19799,N_19977);
nor UO_1122 (O_1122,N_19769,N_19259);
xnor UO_1123 (O_1123,N_19530,N_19505);
xnor UO_1124 (O_1124,N_19457,N_19711);
nand UO_1125 (O_1125,N_19984,N_19378);
nand UO_1126 (O_1126,N_19866,N_19347);
and UO_1127 (O_1127,N_19740,N_19696);
xnor UO_1128 (O_1128,N_19267,N_19424);
nor UO_1129 (O_1129,N_19726,N_19349);
and UO_1130 (O_1130,N_19884,N_19762);
and UO_1131 (O_1131,N_19230,N_19479);
and UO_1132 (O_1132,N_19388,N_19675);
or UO_1133 (O_1133,N_19590,N_19839);
xnor UO_1134 (O_1134,N_19852,N_19267);
nor UO_1135 (O_1135,N_19417,N_19275);
nand UO_1136 (O_1136,N_19831,N_19700);
nor UO_1137 (O_1137,N_19640,N_19455);
or UO_1138 (O_1138,N_19620,N_19949);
or UO_1139 (O_1139,N_19824,N_19483);
nor UO_1140 (O_1140,N_19433,N_19956);
or UO_1141 (O_1141,N_19274,N_19634);
nor UO_1142 (O_1142,N_19815,N_19454);
xor UO_1143 (O_1143,N_19377,N_19569);
xnor UO_1144 (O_1144,N_19356,N_19464);
and UO_1145 (O_1145,N_19463,N_19632);
xnor UO_1146 (O_1146,N_19422,N_19504);
nand UO_1147 (O_1147,N_19700,N_19426);
or UO_1148 (O_1148,N_19978,N_19758);
nand UO_1149 (O_1149,N_19410,N_19512);
and UO_1150 (O_1150,N_19946,N_19715);
and UO_1151 (O_1151,N_19488,N_19621);
nor UO_1152 (O_1152,N_19944,N_19269);
nor UO_1153 (O_1153,N_19370,N_19242);
and UO_1154 (O_1154,N_19685,N_19435);
and UO_1155 (O_1155,N_19489,N_19464);
or UO_1156 (O_1156,N_19615,N_19295);
xor UO_1157 (O_1157,N_19783,N_19992);
or UO_1158 (O_1158,N_19749,N_19891);
nand UO_1159 (O_1159,N_19538,N_19692);
and UO_1160 (O_1160,N_19208,N_19851);
nand UO_1161 (O_1161,N_19469,N_19959);
and UO_1162 (O_1162,N_19238,N_19892);
xor UO_1163 (O_1163,N_19693,N_19377);
nand UO_1164 (O_1164,N_19360,N_19648);
nand UO_1165 (O_1165,N_19334,N_19506);
and UO_1166 (O_1166,N_19759,N_19553);
xor UO_1167 (O_1167,N_19361,N_19471);
and UO_1168 (O_1168,N_19616,N_19211);
xnor UO_1169 (O_1169,N_19894,N_19825);
or UO_1170 (O_1170,N_19945,N_19612);
nor UO_1171 (O_1171,N_19534,N_19576);
nand UO_1172 (O_1172,N_19739,N_19494);
nand UO_1173 (O_1173,N_19222,N_19398);
or UO_1174 (O_1174,N_19947,N_19651);
xnor UO_1175 (O_1175,N_19725,N_19695);
xnor UO_1176 (O_1176,N_19651,N_19435);
nand UO_1177 (O_1177,N_19535,N_19990);
nor UO_1178 (O_1178,N_19430,N_19736);
nand UO_1179 (O_1179,N_19779,N_19919);
nor UO_1180 (O_1180,N_19510,N_19263);
or UO_1181 (O_1181,N_19588,N_19469);
nand UO_1182 (O_1182,N_19471,N_19498);
xor UO_1183 (O_1183,N_19933,N_19309);
xnor UO_1184 (O_1184,N_19584,N_19706);
and UO_1185 (O_1185,N_19877,N_19282);
nor UO_1186 (O_1186,N_19990,N_19638);
nor UO_1187 (O_1187,N_19345,N_19864);
nand UO_1188 (O_1188,N_19587,N_19994);
nand UO_1189 (O_1189,N_19509,N_19546);
nand UO_1190 (O_1190,N_19747,N_19478);
nor UO_1191 (O_1191,N_19892,N_19779);
nor UO_1192 (O_1192,N_19830,N_19922);
xor UO_1193 (O_1193,N_19539,N_19607);
or UO_1194 (O_1194,N_19798,N_19995);
and UO_1195 (O_1195,N_19948,N_19912);
nand UO_1196 (O_1196,N_19751,N_19765);
nand UO_1197 (O_1197,N_19593,N_19227);
and UO_1198 (O_1198,N_19240,N_19600);
nor UO_1199 (O_1199,N_19644,N_19289);
and UO_1200 (O_1200,N_19993,N_19597);
nand UO_1201 (O_1201,N_19827,N_19819);
nor UO_1202 (O_1202,N_19962,N_19853);
nor UO_1203 (O_1203,N_19404,N_19263);
nand UO_1204 (O_1204,N_19349,N_19264);
or UO_1205 (O_1205,N_19346,N_19274);
and UO_1206 (O_1206,N_19775,N_19551);
or UO_1207 (O_1207,N_19202,N_19619);
xnor UO_1208 (O_1208,N_19805,N_19819);
or UO_1209 (O_1209,N_19702,N_19817);
or UO_1210 (O_1210,N_19481,N_19271);
and UO_1211 (O_1211,N_19687,N_19458);
and UO_1212 (O_1212,N_19701,N_19545);
nand UO_1213 (O_1213,N_19235,N_19393);
nand UO_1214 (O_1214,N_19343,N_19553);
nand UO_1215 (O_1215,N_19400,N_19859);
or UO_1216 (O_1216,N_19425,N_19267);
nand UO_1217 (O_1217,N_19252,N_19883);
or UO_1218 (O_1218,N_19702,N_19521);
nor UO_1219 (O_1219,N_19995,N_19738);
nand UO_1220 (O_1220,N_19219,N_19583);
nand UO_1221 (O_1221,N_19674,N_19580);
nor UO_1222 (O_1222,N_19770,N_19294);
xor UO_1223 (O_1223,N_19589,N_19279);
nand UO_1224 (O_1224,N_19940,N_19990);
xnor UO_1225 (O_1225,N_19936,N_19372);
xor UO_1226 (O_1226,N_19688,N_19269);
nor UO_1227 (O_1227,N_19253,N_19628);
nand UO_1228 (O_1228,N_19746,N_19455);
and UO_1229 (O_1229,N_19808,N_19222);
and UO_1230 (O_1230,N_19688,N_19897);
or UO_1231 (O_1231,N_19305,N_19718);
or UO_1232 (O_1232,N_19736,N_19626);
xor UO_1233 (O_1233,N_19370,N_19482);
and UO_1234 (O_1234,N_19512,N_19474);
and UO_1235 (O_1235,N_19968,N_19257);
or UO_1236 (O_1236,N_19673,N_19343);
or UO_1237 (O_1237,N_19543,N_19678);
nand UO_1238 (O_1238,N_19535,N_19988);
xnor UO_1239 (O_1239,N_19323,N_19864);
xnor UO_1240 (O_1240,N_19826,N_19232);
xor UO_1241 (O_1241,N_19264,N_19294);
nand UO_1242 (O_1242,N_19395,N_19648);
nor UO_1243 (O_1243,N_19751,N_19623);
nor UO_1244 (O_1244,N_19275,N_19988);
nor UO_1245 (O_1245,N_19757,N_19897);
nand UO_1246 (O_1246,N_19633,N_19214);
or UO_1247 (O_1247,N_19629,N_19794);
nor UO_1248 (O_1248,N_19299,N_19691);
nand UO_1249 (O_1249,N_19578,N_19922);
and UO_1250 (O_1250,N_19454,N_19810);
xor UO_1251 (O_1251,N_19904,N_19429);
nand UO_1252 (O_1252,N_19765,N_19465);
xnor UO_1253 (O_1253,N_19616,N_19234);
or UO_1254 (O_1254,N_19221,N_19429);
nor UO_1255 (O_1255,N_19885,N_19917);
and UO_1256 (O_1256,N_19615,N_19272);
and UO_1257 (O_1257,N_19608,N_19329);
and UO_1258 (O_1258,N_19590,N_19832);
and UO_1259 (O_1259,N_19261,N_19941);
nor UO_1260 (O_1260,N_19311,N_19967);
nor UO_1261 (O_1261,N_19831,N_19555);
nand UO_1262 (O_1262,N_19993,N_19574);
nand UO_1263 (O_1263,N_19451,N_19454);
or UO_1264 (O_1264,N_19349,N_19242);
and UO_1265 (O_1265,N_19869,N_19845);
nand UO_1266 (O_1266,N_19991,N_19974);
and UO_1267 (O_1267,N_19242,N_19684);
or UO_1268 (O_1268,N_19527,N_19792);
or UO_1269 (O_1269,N_19961,N_19401);
nand UO_1270 (O_1270,N_19311,N_19338);
nand UO_1271 (O_1271,N_19786,N_19408);
and UO_1272 (O_1272,N_19581,N_19911);
xnor UO_1273 (O_1273,N_19573,N_19269);
nand UO_1274 (O_1274,N_19625,N_19602);
nand UO_1275 (O_1275,N_19791,N_19674);
xor UO_1276 (O_1276,N_19272,N_19593);
or UO_1277 (O_1277,N_19236,N_19304);
nor UO_1278 (O_1278,N_19314,N_19356);
nand UO_1279 (O_1279,N_19778,N_19310);
nor UO_1280 (O_1280,N_19338,N_19719);
xnor UO_1281 (O_1281,N_19849,N_19810);
or UO_1282 (O_1282,N_19848,N_19867);
or UO_1283 (O_1283,N_19372,N_19526);
and UO_1284 (O_1284,N_19524,N_19417);
nor UO_1285 (O_1285,N_19301,N_19413);
xnor UO_1286 (O_1286,N_19827,N_19646);
or UO_1287 (O_1287,N_19821,N_19528);
xor UO_1288 (O_1288,N_19532,N_19701);
and UO_1289 (O_1289,N_19413,N_19801);
nor UO_1290 (O_1290,N_19739,N_19568);
nor UO_1291 (O_1291,N_19588,N_19649);
and UO_1292 (O_1292,N_19275,N_19389);
or UO_1293 (O_1293,N_19618,N_19853);
nor UO_1294 (O_1294,N_19346,N_19571);
xnor UO_1295 (O_1295,N_19726,N_19275);
nor UO_1296 (O_1296,N_19865,N_19960);
nand UO_1297 (O_1297,N_19942,N_19896);
nand UO_1298 (O_1298,N_19390,N_19509);
xor UO_1299 (O_1299,N_19889,N_19371);
xnor UO_1300 (O_1300,N_19387,N_19360);
xor UO_1301 (O_1301,N_19383,N_19697);
nand UO_1302 (O_1302,N_19598,N_19912);
and UO_1303 (O_1303,N_19796,N_19214);
and UO_1304 (O_1304,N_19394,N_19317);
xor UO_1305 (O_1305,N_19640,N_19941);
nor UO_1306 (O_1306,N_19365,N_19588);
nor UO_1307 (O_1307,N_19200,N_19665);
nand UO_1308 (O_1308,N_19930,N_19420);
nand UO_1309 (O_1309,N_19391,N_19205);
nor UO_1310 (O_1310,N_19643,N_19664);
nor UO_1311 (O_1311,N_19604,N_19808);
nand UO_1312 (O_1312,N_19865,N_19864);
nand UO_1313 (O_1313,N_19919,N_19903);
nand UO_1314 (O_1314,N_19397,N_19799);
xnor UO_1315 (O_1315,N_19627,N_19752);
nand UO_1316 (O_1316,N_19748,N_19465);
xnor UO_1317 (O_1317,N_19559,N_19621);
or UO_1318 (O_1318,N_19317,N_19444);
xnor UO_1319 (O_1319,N_19577,N_19663);
xor UO_1320 (O_1320,N_19451,N_19461);
or UO_1321 (O_1321,N_19722,N_19411);
nor UO_1322 (O_1322,N_19848,N_19892);
and UO_1323 (O_1323,N_19606,N_19829);
or UO_1324 (O_1324,N_19335,N_19688);
or UO_1325 (O_1325,N_19541,N_19755);
nor UO_1326 (O_1326,N_19342,N_19770);
nand UO_1327 (O_1327,N_19546,N_19426);
or UO_1328 (O_1328,N_19689,N_19432);
or UO_1329 (O_1329,N_19477,N_19759);
or UO_1330 (O_1330,N_19911,N_19826);
nand UO_1331 (O_1331,N_19294,N_19918);
nand UO_1332 (O_1332,N_19301,N_19430);
and UO_1333 (O_1333,N_19841,N_19621);
and UO_1334 (O_1334,N_19227,N_19214);
and UO_1335 (O_1335,N_19518,N_19308);
or UO_1336 (O_1336,N_19979,N_19723);
xor UO_1337 (O_1337,N_19310,N_19748);
or UO_1338 (O_1338,N_19250,N_19635);
and UO_1339 (O_1339,N_19957,N_19230);
or UO_1340 (O_1340,N_19450,N_19580);
or UO_1341 (O_1341,N_19576,N_19851);
xnor UO_1342 (O_1342,N_19594,N_19331);
or UO_1343 (O_1343,N_19933,N_19654);
xnor UO_1344 (O_1344,N_19577,N_19718);
xnor UO_1345 (O_1345,N_19371,N_19379);
nand UO_1346 (O_1346,N_19990,N_19982);
nand UO_1347 (O_1347,N_19495,N_19340);
and UO_1348 (O_1348,N_19952,N_19477);
or UO_1349 (O_1349,N_19928,N_19233);
or UO_1350 (O_1350,N_19443,N_19476);
or UO_1351 (O_1351,N_19981,N_19534);
or UO_1352 (O_1352,N_19650,N_19412);
or UO_1353 (O_1353,N_19579,N_19914);
nor UO_1354 (O_1354,N_19208,N_19989);
nand UO_1355 (O_1355,N_19526,N_19856);
xor UO_1356 (O_1356,N_19718,N_19205);
or UO_1357 (O_1357,N_19231,N_19585);
or UO_1358 (O_1358,N_19239,N_19721);
xnor UO_1359 (O_1359,N_19777,N_19345);
nor UO_1360 (O_1360,N_19852,N_19201);
or UO_1361 (O_1361,N_19588,N_19858);
or UO_1362 (O_1362,N_19551,N_19665);
nand UO_1363 (O_1363,N_19871,N_19545);
or UO_1364 (O_1364,N_19321,N_19963);
and UO_1365 (O_1365,N_19523,N_19330);
xnor UO_1366 (O_1366,N_19815,N_19849);
nand UO_1367 (O_1367,N_19243,N_19297);
nor UO_1368 (O_1368,N_19709,N_19258);
xnor UO_1369 (O_1369,N_19452,N_19708);
xor UO_1370 (O_1370,N_19808,N_19448);
nand UO_1371 (O_1371,N_19344,N_19745);
and UO_1372 (O_1372,N_19826,N_19636);
xnor UO_1373 (O_1373,N_19544,N_19397);
and UO_1374 (O_1374,N_19611,N_19459);
xnor UO_1375 (O_1375,N_19437,N_19713);
or UO_1376 (O_1376,N_19846,N_19517);
or UO_1377 (O_1377,N_19469,N_19304);
and UO_1378 (O_1378,N_19442,N_19436);
nor UO_1379 (O_1379,N_19839,N_19795);
xnor UO_1380 (O_1380,N_19572,N_19868);
nor UO_1381 (O_1381,N_19653,N_19612);
or UO_1382 (O_1382,N_19757,N_19521);
or UO_1383 (O_1383,N_19715,N_19788);
or UO_1384 (O_1384,N_19455,N_19696);
nor UO_1385 (O_1385,N_19398,N_19702);
xor UO_1386 (O_1386,N_19685,N_19444);
xnor UO_1387 (O_1387,N_19684,N_19665);
or UO_1388 (O_1388,N_19819,N_19481);
nor UO_1389 (O_1389,N_19451,N_19760);
nor UO_1390 (O_1390,N_19745,N_19814);
and UO_1391 (O_1391,N_19258,N_19289);
nand UO_1392 (O_1392,N_19313,N_19431);
or UO_1393 (O_1393,N_19796,N_19791);
nand UO_1394 (O_1394,N_19697,N_19287);
nor UO_1395 (O_1395,N_19725,N_19973);
or UO_1396 (O_1396,N_19927,N_19967);
nor UO_1397 (O_1397,N_19423,N_19680);
nand UO_1398 (O_1398,N_19232,N_19674);
nor UO_1399 (O_1399,N_19363,N_19364);
or UO_1400 (O_1400,N_19202,N_19335);
nand UO_1401 (O_1401,N_19880,N_19455);
nand UO_1402 (O_1402,N_19502,N_19564);
or UO_1403 (O_1403,N_19718,N_19367);
nor UO_1404 (O_1404,N_19412,N_19300);
nand UO_1405 (O_1405,N_19671,N_19337);
or UO_1406 (O_1406,N_19687,N_19915);
xnor UO_1407 (O_1407,N_19457,N_19595);
and UO_1408 (O_1408,N_19661,N_19360);
nand UO_1409 (O_1409,N_19528,N_19391);
nand UO_1410 (O_1410,N_19498,N_19208);
and UO_1411 (O_1411,N_19495,N_19535);
nand UO_1412 (O_1412,N_19931,N_19591);
nor UO_1413 (O_1413,N_19603,N_19799);
and UO_1414 (O_1414,N_19646,N_19359);
or UO_1415 (O_1415,N_19507,N_19433);
or UO_1416 (O_1416,N_19545,N_19681);
and UO_1417 (O_1417,N_19729,N_19404);
nor UO_1418 (O_1418,N_19631,N_19328);
nand UO_1419 (O_1419,N_19746,N_19341);
and UO_1420 (O_1420,N_19542,N_19422);
and UO_1421 (O_1421,N_19785,N_19323);
nand UO_1422 (O_1422,N_19929,N_19982);
nor UO_1423 (O_1423,N_19950,N_19425);
or UO_1424 (O_1424,N_19253,N_19884);
and UO_1425 (O_1425,N_19944,N_19806);
nor UO_1426 (O_1426,N_19641,N_19319);
nor UO_1427 (O_1427,N_19318,N_19431);
nor UO_1428 (O_1428,N_19411,N_19889);
nand UO_1429 (O_1429,N_19695,N_19828);
xnor UO_1430 (O_1430,N_19652,N_19219);
nor UO_1431 (O_1431,N_19992,N_19888);
nand UO_1432 (O_1432,N_19759,N_19480);
nand UO_1433 (O_1433,N_19700,N_19861);
or UO_1434 (O_1434,N_19799,N_19884);
xor UO_1435 (O_1435,N_19678,N_19343);
and UO_1436 (O_1436,N_19518,N_19749);
nand UO_1437 (O_1437,N_19613,N_19353);
and UO_1438 (O_1438,N_19846,N_19680);
or UO_1439 (O_1439,N_19640,N_19843);
and UO_1440 (O_1440,N_19540,N_19416);
or UO_1441 (O_1441,N_19913,N_19822);
nor UO_1442 (O_1442,N_19348,N_19552);
xor UO_1443 (O_1443,N_19450,N_19865);
xor UO_1444 (O_1444,N_19882,N_19240);
and UO_1445 (O_1445,N_19542,N_19612);
or UO_1446 (O_1446,N_19281,N_19250);
and UO_1447 (O_1447,N_19566,N_19509);
or UO_1448 (O_1448,N_19939,N_19682);
and UO_1449 (O_1449,N_19556,N_19435);
xnor UO_1450 (O_1450,N_19248,N_19775);
xor UO_1451 (O_1451,N_19615,N_19227);
nor UO_1452 (O_1452,N_19797,N_19896);
and UO_1453 (O_1453,N_19756,N_19233);
and UO_1454 (O_1454,N_19751,N_19250);
nand UO_1455 (O_1455,N_19300,N_19833);
nor UO_1456 (O_1456,N_19856,N_19732);
and UO_1457 (O_1457,N_19333,N_19447);
xnor UO_1458 (O_1458,N_19817,N_19993);
xor UO_1459 (O_1459,N_19258,N_19822);
xor UO_1460 (O_1460,N_19741,N_19370);
nor UO_1461 (O_1461,N_19572,N_19994);
nand UO_1462 (O_1462,N_19943,N_19968);
nor UO_1463 (O_1463,N_19525,N_19799);
nand UO_1464 (O_1464,N_19225,N_19412);
nor UO_1465 (O_1465,N_19727,N_19475);
or UO_1466 (O_1466,N_19209,N_19450);
nand UO_1467 (O_1467,N_19551,N_19480);
and UO_1468 (O_1468,N_19383,N_19754);
nand UO_1469 (O_1469,N_19801,N_19278);
nand UO_1470 (O_1470,N_19927,N_19660);
nor UO_1471 (O_1471,N_19529,N_19799);
nand UO_1472 (O_1472,N_19834,N_19457);
and UO_1473 (O_1473,N_19926,N_19502);
and UO_1474 (O_1474,N_19246,N_19704);
or UO_1475 (O_1475,N_19674,N_19671);
nor UO_1476 (O_1476,N_19284,N_19457);
and UO_1477 (O_1477,N_19230,N_19600);
or UO_1478 (O_1478,N_19528,N_19384);
nor UO_1479 (O_1479,N_19509,N_19976);
and UO_1480 (O_1480,N_19526,N_19805);
nand UO_1481 (O_1481,N_19950,N_19685);
xnor UO_1482 (O_1482,N_19656,N_19211);
and UO_1483 (O_1483,N_19759,N_19410);
nor UO_1484 (O_1484,N_19378,N_19284);
nor UO_1485 (O_1485,N_19708,N_19769);
nor UO_1486 (O_1486,N_19744,N_19976);
and UO_1487 (O_1487,N_19652,N_19701);
nor UO_1488 (O_1488,N_19304,N_19644);
xnor UO_1489 (O_1489,N_19348,N_19410);
or UO_1490 (O_1490,N_19752,N_19331);
xor UO_1491 (O_1491,N_19252,N_19728);
xor UO_1492 (O_1492,N_19332,N_19839);
or UO_1493 (O_1493,N_19219,N_19904);
or UO_1494 (O_1494,N_19383,N_19728);
or UO_1495 (O_1495,N_19697,N_19376);
and UO_1496 (O_1496,N_19316,N_19354);
nand UO_1497 (O_1497,N_19770,N_19812);
or UO_1498 (O_1498,N_19481,N_19252);
nor UO_1499 (O_1499,N_19924,N_19461);
or UO_1500 (O_1500,N_19367,N_19770);
nor UO_1501 (O_1501,N_19550,N_19774);
or UO_1502 (O_1502,N_19755,N_19217);
nand UO_1503 (O_1503,N_19910,N_19994);
or UO_1504 (O_1504,N_19831,N_19683);
nand UO_1505 (O_1505,N_19472,N_19260);
xor UO_1506 (O_1506,N_19356,N_19707);
and UO_1507 (O_1507,N_19229,N_19297);
or UO_1508 (O_1508,N_19477,N_19257);
xnor UO_1509 (O_1509,N_19717,N_19456);
and UO_1510 (O_1510,N_19452,N_19640);
and UO_1511 (O_1511,N_19344,N_19231);
nand UO_1512 (O_1512,N_19422,N_19837);
nor UO_1513 (O_1513,N_19475,N_19832);
nor UO_1514 (O_1514,N_19338,N_19568);
nand UO_1515 (O_1515,N_19849,N_19372);
xnor UO_1516 (O_1516,N_19790,N_19443);
or UO_1517 (O_1517,N_19562,N_19215);
or UO_1518 (O_1518,N_19804,N_19435);
nand UO_1519 (O_1519,N_19749,N_19855);
nor UO_1520 (O_1520,N_19669,N_19214);
xnor UO_1521 (O_1521,N_19267,N_19839);
nor UO_1522 (O_1522,N_19926,N_19887);
and UO_1523 (O_1523,N_19267,N_19944);
xor UO_1524 (O_1524,N_19231,N_19252);
or UO_1525 (O_1525,N_19893,N_19257);
or UO_1526 (O_1526,N_19737,N_19294);
nor UO_1527 (O_1527,N_19763,N_19674);
xor UO_1528 (O_1528,N_19226,N_19968);
or UO_1529 (O_1529,N_19347,N_19933);
or UO_1530 (O_1530,N_19866,N_19323);
or UO_1531 (O_1531,N_19571,N_19627);
nor UO_1532 (O_1532,N_19998,N_19470);
or UO_1533 (O_1533,N_19706,N_19283);
nor UO_1534 (O_1534,N_19431,N_19530);
xor UO_1535 (O_1535,N_19917,N_19224);
and UO_1536 (O_1536,N_19848,N_19869);
nand UO_1537 (O_1537,N_19646,N_19942);
nor UO_1538 (O_1538,N_19993,N_19766);
nor UO_1539 (O_1539,N_19550,N_19981);
or UO_1540 (O_1540,N_19271,N_19746);
nor UO_1541 (O_1541,N_19615,N_19610);
xnor UO_1542 (O_1542,N_19927,N_19216);
nor UO_1543 (O_1543,N_19422,N_19864);
or UO_1544 (O_1544,N_19477,N_19623);
and UO_1545 (O_1545,N_19989,N_19953);
and UO_1546 (O_1546,N_19549,N_19520);
nand UO_1547 (O_1547,N_19273,N_19271);
xnor UO_1548 (O_1548,N_19525,N_19625);
or UO_1549 (O_1549,N_19389,N_19782);
xnor UO_1550 (O_1550,N_19231,N_19283);
nor UO_1551 (O_1551,N_19721,N_19589);
or UO_1552 (O_1552,N_19345,N_19946);
nand UO_1553 (O_1553,N_19493,N_19283);
and UO_1554 (O_1554,N_19250,N_19361);
or UO_1555 (O_1555,N_19859,N_19268);
nor UO_1556 (O_1556,N_19915,N_19493);
xnor UO_1557 (O_1557,N_19226,N_19418);
or UO_1558 (O_1558,N_19579,N_19724);
or UO_1559 (O_1559,N_19880,N_19721);
xnor UO_1560 (O_1560,N_19279,N_19356);
or UO_1561 (O_1561,N_19865,N_19480);
or UO_1562 (O_1562,N_19907,N_19535);
xor UO_1563 (O_1563,N_19680,N_19984);
nor UO_1564 (O_1564,N_19520,N_19671);
xor UO_1565 (O_1565,N_19620,N_19285);
nand UO_1566 (O_1566,N_19933,N_19246);
or UO_1567 (O_1567,N_19942,N_19640);
nand UO_1568 (O_1568,N_19718,N_19900);
or UO_1569 (O_1569,N_19776,N_19493);
nor UO_1570 (O_1570,N_19286,N_19500);
and UO_1571 (O_1571,N_19936,N_19449);
or UO_1572 (O_1572,N_19565,N_19436);
or UO_1573 (O_1573,N_19881,N_19926);
nand UO_1574 (O_1574,N_19480,N_19931);
and UO_1575 (O_1575,N_19374,N_19706);
nand UO_1576 (O_1576,N_19703,N_19967);
xor UO_1577 (O_1577,N_19273,N_19263);
and UO_1578 (O_1578,N_19458,N_19793);
nand UO_1579 (O_1579,N_19385,N_19814);
xnor UO_1580 (O_1580,N_19823,N_19316);
nor UO_1581 (O_1581,N_19346,N_19301);
nand UO_1582 (O_1582,N_19354,N_19578);
or UO_1583 (O_1583,N_19861,N_19256);
or UO_1584 (O_1584,N_19782,N_19669);
nor UO_1585 (O_1585,N_19884,N_19737);
nand UO_1586 (O_1586,N_19855,N_19256);
nor UO_1587 (O_1587,N_19674,N_19311);
nand UO_1588 (O_1588,N_19924,N_19483);
nand UO_1589 (O_1589,N_19712,N_19840);
nand UO_1590 (O_1590,N_19708,N_19454);
nand UO_1591 (O_1591,N_19239,N_19597);
nand UO_1592 (O_1592,N_19869,N_19394);
or UO_1593 (O_1593,N_19836,N_19780);
and UO_1594 (O_1594,N_19973,N_19368);
nor UO_1595 (O_1595,N_19233,N_19660);
nor UO_1596 (O_1596,N_19450,N_19520);
or UO_1597 (O_1597,N_19416,N_19253);
nand UO_1598 (O_1598,N_19881,N_19274);
and UO_1599 (O_1599,N_19304,N_19648);
and UO_1600 (O_1600,N_19251,N_19760);
nor UO_1601 (O_1601,N_19387,N_19468);
nor UO_1602 (O_1602,N_19716,N_19594);
nand UO_1603 (O_1603,N_19799,N_19324);
nand UO_1604 (O_1604,N_19869,N_19912);
nor UO_1605 (O_1605,N_19434,N_19522);
nor UO_1606 (O_1606,N_19374,N_19442);
or UO_1607 (O_1607,N_19545,N_19339);
xor UO_1608 (O_1608,N_19270,N_19894);
nor UO_1609 (O_1609,N_19874,N_19940);
nand UO_1610 (O_1610,N_19833,N_19524);
xor UO_1611 (O_1611,N_19873,N_19349);
and UO_1612 (O_1612,N_19614,N_19917);
and UO_1613 (O_1613,N_19540,N_19760);
or UO_1614 (O_1614,N_19737,N_19684);
xnor UO_1615 (O_1615,N_19723,N_19648);
nand UO_1616 (O_1616,N_19924,N_19351);
nand UO_1617 (O_1617,N_19987,N_19456);
or UO_1618 (O_1618,N_19990,N_19711);
or UO_1619 (O_1619,N_19979,N_19965);
and UO_1620 (O_1620,N_19854,N_19775);
xor UO_1621 (O_1621,N_19978,N_19438);
nor UO_1622 (O_1622,N_19675,N_19894);
nor UO_1623 (O_1623,N_19772,N_19625);
xnor UO_1624 (O_1624,N_19419,N_19225);
or UO_1625 (O_1625,N_19760,N_19562);
xor UO_1626 (O_1626,N_19945,N_19290);
nor UO_1627 (O_1627,N_19961,N_19922);
nor UO_1628 (O_1628,N_19335,N_19249);
nor UO_1629 (O_1629,N_19644,N_19586);
xnor UO_1630 (O_1630,N_19597,N_19602);
nand UO_1631 (O_1631,N_19966,N_19874);
or UO_1632 (O_1632,N_19949,N_19716);
nand UO_1633 (O_1633,N_19964,N_19291);
nor UO_1634 (O_1634,N_19921,N_19247);
nand UO_1635 (O_1635,N_19468,N_19261);
xnor UO_1636 (O_1636,N_19467,N_19503);
xor UO_1637 (O_1637,N_19673,N_19628);
xor UO_1638 (O_1638,N_19853,N_19628);
nor UO_1639 (O_1639,N_19599,N_19814);
nand UO_1640 (O_1640,N_19743,N_19837);
nand UO_1641 (O_1641,N_19455,N_19827);
and UO_1642 (O_1642,N_19239,N_19905);
or UO_1643 (O_1643,N_19863,N_19248);
nor UO_1644 (O_1644,N_19292,N_19784);
nor UO_1645 (O_1645,N_19738,N_19875);
nand UO_1646 (O_1646,N_19269,N_19253);
nor UO_1647 (O_1647,N_19577,N_19671);
xnor UO_1648 (O_1648,N_19617,N_19524);
or UO_1649 (O_1649,N_19512,N_19389);
nor UO_1650 (O_1650,N_19655,N_19373);
and UO_1651 (O_1651,N_19718,N_19690);
and UO_1652 (O_1652,N_19575,N_19525);
and UO_1653 (O_1653,N_19542,N_19973);
and UO_1654 (O_1654,N_19782,N_19664);
and UO_1655 (O_1655,N_19857,N_19870);
nor UO_1656 (O_1656,N_19232,N_19716);
nand UO_1657 (O_1657,N_19920,N_19965);
nor UO_1658 (O_1658,N_19511,N_19309);
and UO_1659 (O_1659,N_19911,N_19939);
or UO_1660 (O_1660,N_19491,N_19384);
nor UO_1661 (O_1661,N_19772,N_19251);
xnor UO_1662 (O_1662,N_19880,N_19299);
nor UO_1663 (O_1663,N_19852,N_19411);
or UO_1664 (O_1664,N_19304,N_19442);
nor UO_1665 (O_1665,N_19325,N_19953);
nand UO_1666 (O_1666,N_19646,N_19793);
or UO_1667 (O_1667,N_19685,N_19563);
xor UO_1668 (O_1668,N_19494,N_19544);
xor UO_1669 (O_1669,N_19226,N_19507);
or UO_1670 (O_1670,N_19971,N_19867);
nand UO_1671 (O_1671,N_19397,N_19825);
and UO_1672 (O_1672,N_19931,N_19277);
nor UO_1673 (O_1673,N_19303,N_19340);
and UO_1674 (O_1674,N_19846,N_19455);
nand UO_1675 (O_1675,N_19413,N_19457);
xor UO_1676 (O_1676,N_19606,N_19417);
nand UO_1677 (O_1677,N_19952,N_19975);
or UO_1678 (O_1678,N_19340,N_19327);
nand UO_1679 (O_1679,N_19435,N_19584);
nand UO_1680 (O_1680,N_19638,N_19460);
nand UO_1681 (O_1681,N_19886,N_19682);
nor UO_1682 (O_1682,N_19233,N_19356);
nor UO_1683 (O_1683,N_19658,N_19626);
or UO_1684 (O_1684,N_19632,N_19290);
nand UO_1685 (O_1685,N_19349,N_19420);
nor UO_1686 (O_1686,N_19208,N_19693);
and UO_1687 (O_1687,N_19830,N_19955);
nand UO_1688 (O_1688,N_19644,N_19766);
nand UO_1689 (O_1689,N_19921,N_19203);
xnor UO_1690 (O_1690,N_19814,N_19818);
or UO_1691 (O_1691,N_19922,N_19464);
xnor UO_1692 (O_1692,N_19290,N_19983);
nand UO_1693 (O_1693,N_19914,N_19630);
nor UO_1694 (O_1694,N_19825,N_19472);
or UO_1695 (O_1695,N_19908,N_19524);
or UO_1696 (O_1696,N_19866,N_19748);
and UO_1697 (O_1697,N_19207,N_19921);
nor UO_1698 (O_1698,N_19223,N_19684);
or UO_1699 (O_1699,N_19885,N_19601);
and UO_1700 (O_1700,N_19509,N_19948);
or UO_1701 (O_1701,N_19848,N_19966);
xor UO_1702 (O_1702,N_19207,N_19504);
nor UO_1703 (O_1703,N_19808,N_19943);
nand UO_1704 (O_1704,N_19654,N_19559);
and UO_1705 (O_1705,N_19235,N_19472);
nor UO_1706 (O_1706,N_19969,N_19885);
nand UO_1707 (O_1707,N_19218,N_19819);
nand UO_1708 (O_1708,N_19967,N_19663);
nand UO_1709 (O_1709,N_19292,N_19758);
and UO_1710 (O_1710,N_19682,N_19258);
or UO_1711 (O_1711,N_19494,N_19599);
nand UO_1712 (O_1712,N_19622,N_19801);
nand UO_1713 (O_1713,N_19880,N_19651);
nand UO_1714 (O_1714,N_19255,N_19297);
nand UO_1715 (O_1715,N_19964,N_19990);
nor UO_1716 (O_1716,N_19293,N_19425);
nor UO_1717 (O_1717,N_19807,N_19818);
nor UO_1718 (O_1718,N_19745,N_19383);
or UO_1719 (O_1719,N_19851,N_19799);
and UO_1720 (O_1720,N_19847,N_19951);
nand UO_1721 (O_1721,N_19384,N_19671);
nand UO_1722 (O_1722,N_19765,N_19704);
and UO_1723 (O_1723,N_19208,N_19867);
and UO_1724 (O_1724,N_19299,N_19738);
xnor UO_1725 (O_1725,N_19635,N_19463);
nand UO_1726 (O_1726,N_19242,N_19225);
nor UO_1727 (O_1727,N_19926,N_19459);
nand UO_1728 (O_1728,N_19256,N_19871);
xor UO_1729 (O_1729,N_19887,N_19497);
and UO_1730 (O_1730,N_19205,N_19626);
xnor UO_1731 (O_1731,N_19418,N_19403);
nand UO_1732 (O_1732,N_19798,N_19874);
nor UO_1733 (O_1733,N_19976,N_19684);
nor UO_1734 (O_1734,N_19915,N_19565);
xnor UO_1735 (O_1735,N_19479,N_19543);
nand UO_1736 (O_1736,N_19382,N_19392);
or UO_1737 (O_1737,N_19936,N_19282);
and UO_1738 (O_1738,N_19353,N_19719);
or UO_1739 (O_1739,N_19746,N_19740);
and UO_1740 (O_1740,N_19847,N_19253);
or UO_1741 (O_1741,N_19979,N_19360);
nor UO_1742 (O_1742,N_19734,N_19263);
or UO_1743 (O_1743,N_19281,N_19480);
xnor UO_1744 (O_1744,N_19679,N_19672);
nor UO_1745 (O_1745,N_19233,N_19310);
xnor UO_1746 (O_1746,N_19510,N_19909);
xnor UO_1747 (O_1747,N_19957,N_19229);
and UO_1748 (O_1748,N_19961,N_19217);
nand UO_1749 (O_1749,N_19463,N_19348);
and UO_1750 (O_1750,N_19707,N_19216);
or UO_1751 (O_1751,N_19960,N_19435);
and UO_1752 (O_1752,N_19984,N_19400);
nor UO_1753 (O_1753,N_19734,N_19418);
xnor UO_1754 (O_1754,N_19218,N_19955);
or UO_1755 (O_1755,N_19836,N_19965);
nand UO_1756 (O_1756,N_19398,N_19981);
nand UO_1757 (O_1757,N_19898,N_19678);
nand UO_1758 (O_1758,N_19939,N_19981);
xnor UO_1759 (O_1759,N_19809,N_19707);
and UO_1760 (O_1760,N_19280,N_19512);
nand UO_1761 (O_1761,N_19200,N_19709);
nand UO_1762 (O_1762,N_19407,N_19231);
and UO_1763 (O_1763,N_19900,N_19745);
nand UO_1764 (O_1764,N_19505,N_19992);
nand UO_1765 (O_1765,N_19937,N_19947);
xor UO_1766 (O_1766,N_19741,N_19870);
and UO_1767 (O_1767,N_19606,N_19277);
nor UO_1768 (O_1768,N_19920,N_19891);
or UO_1769 (O_1769,N_19300,N_19653);
nor UO_1770 (O_1770,N_19211,N_19225);
xnor UO_1771 (O_1771,N_19869,N_19855);
nor UO_1772 (O_1772,N_19712,N_19721);
xor UO_1773 (O_1773,N_19753,N_19559);
or UO_1774 (O_1774,N_19667,N_19843);
and UO_1775 (O_1775,N_19943,N_19887);
nor UO_1776 (O_1776,N_19481,N_19412);
xor UO_1777 (O_1777,N_19628,N_19472);
nand UO_1778 (O_1778,N_19363,N_19836);
nand UO_1779 (O_1779,N_19919,N_19289);
and UO_1780 (O_1780,N_19480,N_19621);
nor UO_1781 (O_1781,N_19440,N_19961);
nor UO_1782 (O_1782,N_19551,N_19616);
or UO_1783 (O_1783,N_19582,N_19404);
and UO_1784 (O_1784,N_19341,N_19921);
nor UO_1785 (O_1785,N_19665,N_19849);
xor UO_1786 (O_1786,N_19930,N_19499);
nand UO_1787 (O_1787,N_19633,N_19465);
and UO_1788 (O_1788,N_19565,N_19259);
xnor UO_1789 (O_1789,N_19945,N_19970);
nor UO_1790 (O_1790,N_19701,N_19207);
and UO_1791 (O_1791,N_19492,N_19320);
nor UO_1792 (O_1792,N_19226,N_19491);
or UO_1793 (O_1793,N_19349,N_19964);
nand UO_1794 (O_1794,N_19777,N_19664);
xor UO_1795 (O_1795,N_19339,N_19857);
xor UO_1796 (O_1796,N_19433,N_19287);
xor UO_1797 (O_1797,N_19755,N_19917);
or UO_1798 (O_1798,N_19949,N_19475);
nor UO_1799 (O_1799,N_19887,N_19258);
nand UO_1800 (O_1800,N_19856,N_19938);
and UO_1801 (O_1801,N_19330,N_19426);
nor UO_1802 (O_1802,N_19801,N_19514);
nand UO_1803 (O_1803,N_19518,N_19604);
and UO_1804 (O_1804,N_19727,N_19532);
nand UO_1805 (O_1805,N_19369,N_19316);
xor UO_1806 (O_1806,N_19478,N_19968);
nor UO_1807 (O_1807,N_19467,N_19578);
nor UO_1808 (O_1808,N_19678,N_19945);
and UO_1809 (O_1809,N_19550,N_19985);
nor UO_1810 (O_1810,N_19437,N_19321);
nor UO_1811 (O_1811,N_19571,N_19523);
or UO_1812 (O_1812,N_19283,N_19707);
or UO_1813 (O_1813,N_19590,N_19200);
or UO_1814 (O_1814,N_19927,N_19250);
and UO_1815 (O_1815,N_19927,N_19485);
and UO_1816 (O_1816,N_19438,N_19522);
xor UO_1817 (O_1817,N_19675,N_19484);
xor UO_1818 (O_1818,N_19990,N_19524);
nand UO_1819 (O_1819,N_19795,N_19660);
xnor UO_1820 (O_1820,N_19467,N_19986);
xnor UO_1821 (O_1821,N_19942,N_19827);
nand UO_1822 (O_1822,N_19929,N_19354);
nor UO_1823 (O_1823,N_19655,N_19934);
nand UO_1824 (O_1824,N_19442,N_19786);
nand UO_1825 (O_1825,N_19566,N_19425);
nand UO_1826 (O_1826,N_19833,N_19665);
xnor UO_1827 (O_1827,N_19705,N_19412);
or UO_1828 (O_1828,N_19529,N_19622);
nor UO_1829 (O_1829,N_19374,N_19573);
or UO_1830 (O_1830,N_19991,N_19301);
and UO_1831 (O_1831,N_19555,N_19351);
nor UO_1832 (O_1832,N_19997,N_19246);
nor UO_1833 (O_1833,N_19465,N_19420);
or UO_1834 (O_1834,N_19679,N_19951);
nor UO_1835 (O_1835,N_19733,N_19619);
or UO_1836 (O_1836,N_19793,N_19493);
or UO_1837 (O_1837,N_19793,N_19677);
and UO_1838 (O_1838,N_19613,N_19967);
or UO_1839 (O_1839,N_19302,N_19386);
and UO_1840 (O_1840,N_19267,N_19673);
nor UO_1841 (O_1841,N_19453,N_19938);
or UO_1842 (O_1842,N_19916,N_19912);
nor UO_1843 (O_1843,N_19728,N_19632);
and UO_1844 (O_1844,N_19378,N_19774);
nand UO_1845 (O_1845,N_19699,N_19797);
xnor UO_1846 (O_1846,N_19486,N_19999);
nand UO_1847 (O_1847,N_19544,N_19427);
nand UO_1848 (O_1848,N_19491,N_19777);
nor UO_1849 (O_1849,N_19937,N_19528);
xnor UO_1850 (O_1850,N_19482,N_19224);
and UO_1851 (O_1851,N_19995,N_19318);
xor UO_1852 (O_1852,N_19633,N_19585);
xor UO_1853 (O_1853,N_19843,N_19385);
or UO_1854 (O_1854,N_19686,N_19254);
nor UO_1855 (O_1855,N_19888,N_19249);
and UO_1856 (O_1856,N_19942,N_19452);
or UO_1857 (O_1857,N_19260,N_19250);
nand UO_1858 (O_1858,N_19794,N_19738);
xor UO_1859 (O_1859,N_19314,N_19928);
or UO_1860 (O_1860,N_19488,N_19802);
nand UO_1861 (O_1861,N_19268,N_19851);
xnor UO_1862 (O_1862,N_19513,N_19914);
nand UO_1863 (O_1863,N_19674,N_19226);
nand UO_1864 (O_1864,N_19397,N_19482);
nor UO_1865 (O_1865,N_19452,N_19657);
or UO_1866 (O_1866,N_19811,N_19835);
nand UO_1867 (O_1867,N_19441,N_19482);
and UO_1868 (O_1868,N_19769,N_19776);
nor UO_1869 (O_1869,N_19847,N_19723);
xnor UO_1870 (O_1870,N_19274,N_19853);
nand UO_1871 (O_1871,N_19961,N_19615);
nand UO_1872 (O_1872,N_19634,N_19397);
nor UO_1873 (O_1873,N_19314,N_19941);
nand UO_1874 (O_1874,N_19992,N_19585);
xnor UO_1875 (O_1875,N_19507,N_19725);
or UO_1876 (O_1876,N_19627,N_19691);
nand UO_1877 (O_1877,N_19436,N_19605);
and UO_1878 (O_1878,N_19273,N_19788);
and UO_1879 (O_1879,N_19267,N_19871);
xor UO_1880 (O_1880,N_19876,N_19522);
nor UO_1881 (O_1881,N_19886,N_19429);
nand UO_1882 (O_1882,N_19594,N_19244);
xnor UO_1883 (O_1883,N_19313,N_19914);
or UO_1884 (O_1884,N_19402,N_19947);
nand UO_1885 (O_1885,N_19441,N_19940);
nand UO_1886 (O_1886,N_19432,N_19294);
nor UO_1887 (O_1887,N_19695,N_19977);
nor UO_1888 (O_1888,N_19583,N_19562);
nor UO_1889 (O_1889,N_19240,N_19616);
nor UO_1890 (O_1890,N_19565,N_19672);
and UO_1891 (O_1891,N_19836,N_19961);
xnor UO_1892 (O_1892,N_19723,N_19284);
xor UO_1893 (O_1893,N_19459,N_19661);
nand UO_1894 (O_1894,N_19377,N_19765);
xnor UO_1895 (O_1895,N_19309,N_19307);
and UO_1896 (O_1896,N_19451,N_19535);
xor UO_1897 (O_1897,N_19752,N_19576);
nor UO_1898 (O_1898,N_19569,N_19231);
and UO_1899 (O_1899,N_19847,N_19543);
and UO_1900 (O_1900,N_19512,N_19216);
nand UO_1901 (O_1901,N_19620,N_19866);
nor UO_1902 (O_1902,N_19407,N_19502);
nand UO_1903 (O_1903,N_19762,N_19268);
xnor UO_1904 (O_1904,N_19701,N_19534);
and UO_1905 (O_1905,N_19420,N_19672);
or UO_1906 (O_1906,N_19219,N_19310);
or UO_1907 (O_1907,N_19269,N_19926);
and UO_1908 (O_1908,N_19522,N_19933);
and UO_1909 (O_1909,N_19499,N_19344);
or UO_1910 (O_1910,N_19718,N_19446);
or UO_1911 (O_1911,N_19538,N_19230);
nor UO_1912 (O_1912,N_19522,N_19962);
nor UO_1913 (O_1913,N_19804,N_19537);
and UO_1914 (O_1914,N_19738,N_19372);
or UO_1915 (O_1915,N_19548,N_19544);
nand UO_1916 (O_1916,N_19515,N_19817);
or UO_1917 (O_1917,N_19304,N_19859);
nand UO_1918 (O_1918,N_19901,N_19382);
xnor UO_1919 (O_1919,N_19996,N_19811);
xnor UO_1920 (O_1920,N_19414,N_19992);
xor UO_1921 (O_1921,N_19371,N_19389);
nand UO_1922 (O_1922,N_19213,N_19878);
xor UO_1923 (O_1923,N_19649,N_19976);
nor UO_1924 (O_1924,N_19652,N_19595);
nor UO_1925 (O_1925,N_19273,N_19655);
xor UO_1926 (O_1926,N_19907,N_19874);
and UO_1927 (O_1927,N_19465,N_19284);
nor UO_1928 (O_1928,N_19825,N_19747);
nand UO_1929 (O_1929,N_19395,N_19408);
or UO_1930 (O_1930,N_19876,N_19449);
or UO_1931 (O_1931,N_19723,N_19247);
xnor UO_1932 (O_1932,N_19517,N_19552);
xnor UO_1933 (O_1933,N_19590,N_19899);
and UO_1934 (O_1934,N_19206,N_19622);
and UO_1935 (O_1935,N_19822,N_19624);
nor UO_1936 (O_1936,N_19912,N_19535);
and UO_1937 (O_1937,N_19822,N_19670);
and UO_1938 (O_1938,N_19765,N_19518);
and UO_1939 (O_1939,N_19870,N_19601);
or UO_1940 (O_1940,N_19763,N_19593);
nand UO_1941 (O_1941,N_19397,N_19383);
nand UO_1942 (O_1942,N_19232,N_19571);
xor UO_1943 (O_1943,N_19950,N_19910);
xnor UO_1944 (O_1944,N_19423,N_19448);
xnor UO_1945 (O_1945,N_19454,N_19768);
or UO_1946 (O_1946,N_19497,N_19293);
or UO_1947 (O_1947,N_19360,N_19395);
and UO_1948 (O_1948,N_19515,N_19942);
xor UO_1949 (O_1949,N_19384,N_19851);
nor UO_1950 (O_1950,N_19978,N_19510);
or UO_1951 (O_1951,N_19397,N_19882);
nand UO_1952 (O_1952,N_19892,N_19900);
xor UO_1953 (O_1953,N_19880,N_19371);
xor UO_1954 (O_1954,N_19236,N_19906);
xnor UO_1955 (O_1955,N_19393,N_19816);
and UO_1956 (O_1956,N_19478,N_19521);
nand UO_1957 (O_1957,N_19513,N_19620);
xnor UO_1958 (O_1958,N_19827,N_19462);
and UO_1959 (O_1959,N_19606,N_19211);
nor UO_1960 (O_1960,N_19518,N_19611);
xnor UO_1961 (O_1961,N_19850,N_19455);
nand UO_1962 (O_1962,N_19300,N_19401);
xor UO_1963 (O_1963,N_19674,N_19254);
xor UO_1964 (O_1964,N_19888,N_19237);
nor UO_1965 (O_1965,N_19323,N_19496);
or UO_1966 (O_1966,N_19447,N_19932);
nor UO_1967 (O_1967,N_19299,N_19385);
xnor UO_1968 (O_1968,N_19389,N_19785);
and UO_1969 (O_1969,N_19850,N_19703);
nand UO_1970 (O_1970,N_19294,N_19549);
or UO_1971 (O_1971,N_19844,N_19208);
xor UO_1972 (O_1972,N_19398,N_19558);
or UO_1973 (O_1973,N_19961,N_19523);
nand UO_1974 (O_1974,N_19359,N_19947);
or UO_1975 (O_1975,N_19847,N_19727);
nor UO_1976 (O_1976,N_19317,N_19260);
nor UO_1977 (O_1977,N_19561,N_19218);
nand UO_1978 (O_1978,N_19281,N_19538);
or UO_1979 (O_1979,N_19775,N_19830);
or UO_1980 (O_1980,N_19948,N_19434);
xnor UO_1981 (O_1981,N_19611,N_19495);
xnor UO_1982 (O_1982,N_19924,N_19304);
or UO_1983 (O_1983,N_19554,N_19814);
nand UO_1984 (O_1984,N_19912,N_19473);
and UO_1985 (O_1985,N_19723,N_19534);
xor UO_1986 (O_1986,N_19410,N_19321);
or UO_1987 (O_1987,N_19633,N_19416);
xor UO_1988 (O_1988,N_19772,N_19564);
xor UO_1989 (O_1989,N_19328,N_19837);
or UO_1990 (O_1990,N_19471,N_19979);
or UO_1991 (O_1991,N_19515,N_19395);
nor UO_1992 (O_1992,N_19786,N_19725);
nor UO_1993 (O_1993,N_19784,N_19649);
and UO_1994 (O_1994,N_19895,N_19827);
or UO_1995 (O_1995,N_19420,N_19813);
and UO_1996 (O_1996,N_19425,N_19345);
nor UO_1997 (O_1997,N_19412,N_19345);
nand UO_1998 (O_1998,N_19450,N_19806);
nand UO_1999 (O_1999,N_19935,N_19422);
nor UO_2000 (O_2000,N_19711,N_19909);
nor UO_2001 (O_2001,N_19814,N_19481);
nor UO_2002 (O_2002,N_19440,N_19858);
and UO_2003 (O_2003,N_19712,N_19803);
nand UO_2004 (O_2004,N_19618,N_19854);
xnor UO_2005 (O_2005,N_19828,N_19997);
or UO_2006 (O_2006,N_19744,N_19395);
nand UO_2007 (O_2007,N_19415,N_19898);
xnor UO_2008 (O_2008,N_19614,N_19691);
and UO_2009 (O_2009,N_19429,N_19841);
nand UO_2010 (O_2010,N_19900,N_19884);
or UO_2011 (O_2011,N_19402,N_19669);
nand UO_2012 (O_2012,N_19284,N_19476);
nand UO_2013 (O_2013,N_19348,N_19527);
xnor UO_2014 (O_2014,N_19371,N_19422);
xor UO_2015 (O_2015,N_19501,N_19530);
xnor UO_2016 (O_2016,N_19965,N_19733);
and UO_2017 (O_2017,N_19315,N_19386);
xor UO_2018 (O_2018,N_19971,N_19750);
and UO_2019 (O_2019,N_19594,N_19673);
nor UO_2020 (O_2020,N_19967,N_19815);
or UO_2021 (O_2021,N_19994,N_19697);
nand UO_2022 (O_2022,N_19518,N_19694);
nand UO_2023 (O_2023,N_19377,N_19240);
nor UO_2024 (O_2024,N_19239,N_19766);
and UO_2025 (O_2025,N_19251,N_19477);
and UO_2026 (O_2026,N_19513,N_19992);
and UO_2027 (O_2027,N_19939,N_19467);
xnor UO_2028 (O_2028,N_19489,N_19560);
nand UO_2029 (O_2029,N_19561,N_19259);
or UO_2030 (O_2030,N_19619,N_19411);
nor UO_2031 (O_2031,N_19988,N_19861);
and UO_2032 (O_2032,N_19812,N_19431);
and UO_2033 (O_2033,N_19448,N_19208);
xor UO_2034 (O_2034,N_19958,N_19758);
nor UO_2035 (O_2035,N_19422,N_19797);
nor UO_2036 (O_2036,N_19526,N_19310);
and UO_2037 (O_2037,N_19578,N_19561);
nand UO_2038 (O_2038,N_19491,N_19937);
nor UO_2039 (O_2039,N_19415,N_19821);
xor UO_2040 (O_2040,N_19425,N_19942);
or UO_2041 (O_2041,N_19936,N_19917);
nand UO_2042 (O_2042,N_19980,N_19637);
nand UO_2043 (O_2043,N_19356,N_19771);
or UO_2044 (O_2044,N_19498,N_19590);
xnor UO_2045 (O_2045,N_19686,N_19559);
or UO_2046 (O_2046,N_19759,N_19301);
nand UO_2047 (O_2047,N_19767,N_19984);
or UO_2048 (O_2048,N_19957,N_19277);
xnor UO_2049 (O_2049,N_19877,N_19919);
nor UO_2050 (O_2050,N_19245,N_19658);
nor UO_2051 (O_2051,N_19296,N_19533);
nand UO_2052 (O_2052,N_19460,N_19606);
or UO_2053 (O_2053,N_19263,N_19750);
nand UO_2054 (O_2054,N_19820,N_19755);
nand UO_2055 (O_2055,N_19865,N_19747);
nor UO_2056 (O_2056,N_19807,N_19484);
nor UO_2057 (O_2057,N_19350,N_19216);
nor UO_2058 (O_2058,N_19944,N_19947);
or UO_2059 (O_2059,N_19759,N_19292);
and UO_2060 (O_2060,N_19224,N_19504);
xor UO_2061 (O_2061,N_19741,N_19717);
nand UO_2062 (O_2062,N_19693,N_19717);
and UO_2063 (O_2063,N_19440,N_19569);
xnor UO_2064 (O_2064,N_19824,N_19908);
xnor UO_2065 (O_2065,N_19568,N_19920);
nand UO_2066 (O_2066,N_19269,N_19849);
xnor UO_2067 (O_2067,N_19826,N_19479);
nor UO_2068 (O_2068,N_19479,N_19848);
nand UO_2069 (O_2069,N_19677,N_19592);
xnor UO_2070 (O_2070,N_19385,N_19519);
nand UO_2071 (O_2071,N_19339,N_19746);
nand UO_2072 (O_2072,N_19292,N_19412);
xnor UO_2073 (O_2073,N_19789,N_19541);
nor UO_2074 (O_2074,N_19340,N_19857);
xor UO_2075 (O_2075,N_19884,N_19648);
nor UO_2076 (O_2076,N_19210,N_19697);
and UO_2077 (O_2077,N_19390,N_19585);
xor UO_2078 (O_2078,N_19626,N_19650);
and UO_2079 (O_2079,N_19283,N_19895);
nor UO_2080 (O_2080,N_19926,N_19596);
xnor UO_2081 (O_2081,N_19770,N_19919);
or UO_2082 (O_2082,N_19744,N_19839);
nand UO_2083 (O_2083,N_19303,N_19711);
or UO_2084 (O_2084,N_19603,N_19357);
nor UO_2085 (O_2085,N_19571,N_19328);
or UO_2086 (O_2086,N_19919,N_19245);
and UO_2087 (O_2087,N_19656,N_19276);
nand UO_2088 (O_2088,N_19699,N_19955);
nor UO_2089 (O_2089,N_19946,N_19514);
xnor UO_2090 (O_2090,N_19451,N_19820);
nor UO_2091 (O_2091,N_19465,N_19513);
nand UO_2092 (O_2092,N_19778,N_19919);
nor UO_2093 (O_2093,N_19771,N_19448);
or UO_2094 (O_2094,N_19383,N_19876);
and UO_2095 (O_2095,N_19317,N_19411);
xor UO_2096 (O_2096,N_19545,N_19467);
nand UO_2097 (O_2097,N_19929,N_19261);
xor UO_2098 (O_2098,N_19437,N_19753);
xor UO_2099 (O_2099,N_19416,N_19408);
or UO_2100 (O_2100,N_19644,N_19713);
nor UO_2101 (O_2101,N_19771,N_19772);
and UO_2102 (O_2102,N_19791,N_19343);
nor UO_2103 (O_2103,N_19996,N_19591);
nand UO_2104 (O_2104,N_19270,N_19217);
and UO_2105 (O_2105,N_19809,N_19641);
or UO_2106 (O_2106,N_19780,N_19666);
xor UO_2107 (O_2107,N_19743,N_19951);
and UO_2108 (O_2108,N_19791,N_19977);
xor UO_2109 (O_2109,N_19326,N_19344);
nor UO_2110 (O_2110,N_19704,N_19841);
nand UO_2111 (O_2111,N_19261,N_19722);
nand UO_2112 (O_2112,N_19818,N_19417);
xnor UO_2113 (O_2113,N_19926,N_19426);
or UO_2114 (O_2114,N_19210,N_19534);
xor UO_2115 (O_2115,N_19441,N_19862);
or UO_2116 (O_2116,N_19546,N_19470);
nand UO_2117 (O_2117,N_19349,N_19253);
nor UO_2118 (O_2118,N_19243,N_19338);
xor UO_2119 (O_2119,N_19417,N_19667);
nor UO_2120 (O_2120,N_19530,N_19744);
xnor UO_2121 (O_2121,N_19683,N_19989);
or UO_2122 (O_2122,N_19752,N_19269);
or UO_2123 (O_2123,N_19650,N_19957);
and UO_2124 (O_2124,N_19915,N_19826);
and UO_2125 (O_2125,N_19332,N_19485);
xor UO_2126 (O_2126,N_19623,N_19872);
xnor UO_2127 (O_2127,N_19419,N_19797);
nand UO_2128 (O_2128,N_19769,N_19575);
or UO_2129 (O_2129,N_19414,N_19618);
xor UO_2130 (O_2130,N_19792,N_19681);
and UO_2131 (O_2131,N_19750,N_19551);
and UO_2132 (O_2132,N_19727,N_19813);
or UO_2133 (O_2133,N_19220,N_19345);
nor UO_2134 (O_2134,N_19914,N_19524);
nand UO_2135 (O_2135,N_19476,N_19486);
nand UO_2136 (O_2136,N_19578,N_19731);
nand UO_2137 (O_2137,N_19974,N_19635);
nor UO_2138 (O_2138,N_19916,N_19201);
and UO_2139 (O_2139,N_19811,N_19965);
nand UO_2140 (O_2140,N_19916,N_19358);
nand UO_2141 (O_2141,N_19277,N_19413);
and UO_2142 (O_2142,N_19930,N_19450);
nor UO_2143 (O_2143,N_19241,N_19674);
and UO_2144 (O_2144,N_19491,N_19342);
nor UO_2145 (O_2145,N_19454,N_19985);
nor UO_2146 (O_2146,N_19450,N_19250);
nor UO_2147 (O_2147,N_19757,N_19687);
or UO_2148 (O_2148,N_19279,N_19621);
xor UO_2149 (O_2149,N_19263,N_19617);
nand UO_2150 (O_2150,N_19678,N_19846);
nor UO_2151 (O_2151,N_19387,N_19242);
nor UO_2152 (O_2152,N_19314,N_19814);
nand UO_2153 (O_2153,N_19252,N_19816);
nor UO_2154 (O_2154,N_19258,N_19652);
xor UO_2155 (O_2155,N_19635,N_19525);
or UO_2156 (O_2156,N_19950,N_19782);
nor UO_2157 (O_2157,N_19819,N_19798);
nand UO_2158 (O_2158,N_19276,N_19627);
nor UO_2159 (O_2159,N_19434,N_19657);
or UO_2160 (O_2160,N_19430,N_19697);
xnor UO_2161 (O_2161,N_19627,N_19950);
xor UO_2162 (O_2162,N_19275,N_19486);
nor UO_2163 (O_2163,N_19359,N_19236);
and UO_2164 (O_2164,N_19864,N_19638);
or UO_2165 (O_2165,N_19349,N_19756);
xor UO_2166 (O_2166,N_19841,N_19950);
and UO_2167 (O_2167,N_19710,N_19545);
or UO_2168 (O_2168,N_19385,N_19231);
nor UO_2169 (O_2169,N_19385,N_19506);
or UO_2170 (O_2170,N_19582,N_19823);
and UO_2171 (O_2171,N_19943,N_19518);
or UO_2172 (O_2172,N_19246,N_19689);
xor UO_2173 (O_2173,N_19586,N_19961);
and UO_2174 (O_2174,N_19843,N_19995);
xnor UO_2175 (O_2175,N_19845,N_19981);
nor UO_2176 (O_2176,N_19309,N_19302);
xnor UO_2177 (O_2177,N_19344,N_19653);
nor UO_2178 (O_2178,N_19970,N_19931);
xor UO_2179 (O_2179,N_19965,N_19878);
and UO_2180 (O_2180,N_19897,N_19270);
nand UO_2181 (O_2181,N_19572,N_19941);
or UO_2182 (O_2182,N_19925,N_19895);
or UO_2183 (O_2183,N_19892,N_19205);
xnor UO_2184 (O_2184,N_19745,N_19917);
or UO_2185 (O_2185,N_19424,N_19469);
xnor UO_2186 (O_2186,N_19732,N_19711);
nor UO_2187 (O_2187,N_19375,N_19785);
and UO_2188 (O_2188,N_19235,N_19229);
and UO_2189 (O_2189,N_19974,N_19647);
or UO_2190 (O_2190,N_19699,N_19513);
nand UO_2191 (O_2191,N_19730,N_19969);
or UO_2192 (O_2192,N_19678,N_19850);
or UO_2193 (O_2193,N_19422,N_19635);
nand UO_2194 (O_2194,N_19466,N_19672);
nor UO_2195 (O_2195,N_19292,N_19553);
and UO_2196 (O_2196,N_19730,N_19769);
nor UO_2197 (O_2197,N_19255,N_19263);
nand UO_2198 (O_2198,N_19670,N_19236);
and UO_2199 (O_2199,N_19333,N_19582);
nor UO_2200 (O_2200,N_19833,N_19467);
or UO_2201 (O_2201,N_19769,N_19242);
or UO_2202 (O_2202,N_19275,N_19465);
and UO_2203 (O_2203,N_19713,N_19534);
nand UO_2204 (O_2204,N_19453,N_19863);
or UO_2205 (O_2205,N_19355,N_19931);
and UO_2206 (O_2206,N_19691,N_19809);
nand UO_2207 (O_2207,N_19567,N_19795);
nand UO_2208 (O_2208,N_19642,N_19667);
nand UO_2209 (O_2209,N_19537,N_19494);
nor UO_2210 (O_2210,N_19438,N_19253);
or UO_2211 (O_2211,N_19700,N_19373);
or UO_2212 (O_2212,N_19308,N_19812);
and UO_2213 (O_2213,N_19904,N_19633);
xnor UO_2214 (O_2214,N_19415,N_19788);
nor UO_2215 (O_2215,N_19640,N_19625);
or UO_2216 (O_2216,N_19326,N_19429);
xor UO_2217 (O_2217,N_19280,N_19303);
nand UO_2218 (O_2218,N_19291,N_19281);
nor UO_2219 (O_2219,N_19892,N_19295);
nor UO_2220 (O_2220,N_19431,N_19638);
or UO_2221 (O_2221,N_19427,N_19672);
nor UO_2222 (O_2222,N_19657,N_19720);
nor UO_2223 (O_2223,N_19868,N_19462);
and UO_2224 (O_2224,N_19776,N_19283);
or UO_2225 (O_2225,N_19788,N_19309);
xnor UO_2226 (O_2226,N_19989,N_19347);
and UO_2227 (O_2227,N_19471,N_19818);
nand UO_2228 (O_2228,N_19204,N_19565);
xnor UO_2229 (O_2229,N_19784,N_19441);
nand UO_2230 (O_2230,N_19995,N_19725);
and UO_2231 (O_2231,N_19781,N_19642);
or UO_2232 (O_2232,N_19516,N_19462);
or UO_2233 (O_2233,N_19206,N_19680);
xnor UO_2234 (O_2234,N_19558,N_19621);
xnor UO_2235 (O_2235,N_19646,N_19795);
and UO_2236 (O_2236,N_19856,N_19476);
nand UO_2237 (O_2237,N_19391,N_19913);
xnor UO_2238 (O_2238,N_19515,N_19401);
xnor UO_2239 (O_2239,N_19892,N_19870);
nor UO_2240 (O_2240,N_19243,N_19679);
xnor UO_2241 (O_2241,N_19228,N_19771);
xnor UO_2242 (O_2242,N_19677,N_19657);
nor UO_2243 (O_2243,N_19250,N_19552);
nand UO_2244 (O_2244,N_19699,N_19963);
and UO_2245 (O_2245,N_19812,N_19409);
nor UO_2246 (O_2246,N_19723,N_19444);
xnor UO_2247 (O_2247,N_19401,N_19791);
nor UO_2248 (O_2248,N_19469,N_19868);
nand UO_2249 (O_2249,N_19422,N_19887);
nand UO_2250 (O_2250,N_19661,N_19414);
and UO_2251 (O_2251,N_19421,N_19319);
nand UO_2252 (O_2252,N_19287,N_19579);
nor UO_2253 (O_2253,N_19902,N_19245);
nor UO_2254 (O_2254,N_19998,N_19759);
xnor UO_2255 (O_2255,N_19768,N_19515);
xnor UO_2256 (O_2256,N_19295,N_19486);
nor UO_2257 (O_2257,N_19643,N_19558);
xor UO_2258 (O_2258,N_19775,N_19890);
xnor UO_2259 (O_2259,N_19770,N_19793);
or UO_2260 (O_2260,N_19600,N_19419);
xnor UO_2261 (O_2261,N_19609,N_19406);
and UO_2262 (O_2262,N_19237,N_19641);
nor UO_2263 (O_2263,N_19835,N_19800);
or UO_2264 (O_2264,N_19763,N_19482);
nor UO_2265 (O_2265,N_19693,N_19242);
nor UO_2266 (O_2266,N_19919,N_19405);
xnor UO_2267 (O_2267,N_19849,N_19405);
nand UO_2268 (O_2268,N_19604,N_19762);
or UO_2269 (O_2269,N_19873,N_19908);
and UO_2270 (O_2270,N_19808,N_19725);
nor UO_2271 (O_2271,N_19266,N_19470);
xnor UO_2272 (O_2272,N_19868,N_19309);
or UO_2273 (O_2273,N_19530,N_19495);
xnor UO_2274 (O_2274,N_19936,N_19227);
nand UO_2275 (O_2275,N_19654,N_19994);
xor UO_2276 (O_2276,N_19327,N_19706);
and UO_2277 (O_2277,N_19847,N_19632);
or UO_2278 (O_2278,N_19915,N_19936);
and UO_2279 (O_2279,N_19423,N_19932);
nand UO_2280 (O_2280,N_19897,N_19409);
and UO_2281 (O_2281,N_19401,N_19325);
and UO_2282 (O_2282,N_19533,N_19977);
nor UO_2283 (O_2283,N_19660,N_19877);
nand UO_2284 (O_2284,N_19211,N_19680);
nor UO_2285 (O_2285,N_19822,N_19588);
and UO_2286 (O_2286,N_19452,N_19594);
and UO_2287 (O_2287,N_19396,N_19310);
nand UO_2288 (O_2288,N_19639,N_19202);
or UO_2289 (O_2289,N_19561,N_19493);
or UO_2290 (O_2290,N_19348,N_19842);
xnor UO_2291 (O_2291,N_19962,N_19665);
or UO_2292 (O_2292,N_19853,N_19405);
and UO_2293 (O_2293,N_19694,N_19759);
or UO_2294 (O_2294,N_19255,N_19496);
xor UO_2295 (O_2295,N_19815,N_19825);
nand UO_2296 (O_2296,N_19315,N_19770);
xor UO_2297 (O_2297,N_19877,N_19420);
and UO_2298 (O_2298,N_19681,N_19720);
or UO_2299 (O_2299,N_19399,N_19593);
nand UO_2300 (O_2300,N_19333,N_19371);
and UO_2301 (O_2301,N_19698,N_19716);
nand UO_2302 (O_2302,N_19861,N_19978);
and UO_2303 (O_2303,N_19369,N_19651);
xor UO_2304 (O_2304,N_19413,N_19792);
nand UO_2305 (O_2305,N_19509,N_19951);
or UO_2306 (O_2306,N_19426,N_19811);
xor UO_2307 (O_2307,N_19547,N_19985);
nand UO_2308 (O_2308,N_19445,N_19645);
nor UO_2309 (O_2309,N_19586,N_19759);
or UO_2310 (O_2310,N_19466,N_19241);
xor UO_2311 (O_2311,N_19620,N_19332);
nor UO_2312 (O_2312,N_19709,N_19535);
and UO_2313 (O_2313,N_19524,N_19427);
and UO_2314 (O_2314,N_19271,N_19311);
or UO_2315 (O_2315,N_19269,N_19263);
nand UO_2316 (O_2316,N_19618,N_19862);
nand UO_2317 (O_2317,N_19673,N_19678);
nor UO_2318 (O_2318,N_19245,N_19874);
and UO_2319 (O_2319,N_19650,N_19765);
and UO_2320 (O_2320,N_19361,N_19242);
nor UO_2321 (O_2321,N_19204,N_19429);
and UO_2322 (O_2322,N_19233,N_19282);
nand UO_2323 (O_2323,N_19849,N_19710);
or UO_2324 (O_2324,N_19729,N_19252);
nor UO_2325 (O_2325,N_19549,N_19855);
and UO_2326 (O_2326,N_19925,N_19551);
nor UO_2327 (O_2327,N_19689,N_19418);
nand UO_2328 (O_2328,N_19541,N_19908);
nand UO_2329 (O_2329,N_19918,N_19832);
nand UO_2330 (O_2330,N_19866,N_19483);
nand UO_2331 (O_2331,N_19292,N_19546);
nand UO_2332 (O_2332,N_19729,N_19904);
and UO_2333 (O_2333,N_19786,N_19218);
or UO_2334 (O_2334,N_19452,N_19330);
xnor UO_2335 (O_2335,N_19227,N_19566);
or UO_2336 (O_2336,N_19487,N_19538);
or UO_2337 (O_2337,N_19446,N_19897);
xor UO_2338 (O_2338,N_19511,N_19946);
xnor UO_2339 (O_2339,N_19985,N_19945);
xor UO_2340 (O_2340,N_19527,N_19352);
nand UO_2341 (O_2341,N_19506,N_19723);
and UO_2342 (O_2342,N_19927,N_19317);
xor UO_2343 (O_2343,N_19391,N_19774);
nor UO_2344 (O_2344,N_19775,N_19465);
nand UO_2345 (O_2345,N_19540,N_19843);
nor UO_2346 (O_2346,N_19341,N_19632);
xor UO_2347 (O_2347,N_19977,N_19911);
xor UO_2348 (O_2348,N_19362,N_19921);
and UO_2349 (O_2349,N_19628,N_19831);
nor UO_2350 (O_2350,N_19700,N_19202);
or UO_2351 (O_2351,N_19468,N_19308);
nand UO_2352 (O_2352,N_19515,N_19535);
and UO_2353 (O_2353,N_19763,N_19455);
and UO_2354 (O_2354,N_19258,N_19673);
or UO_2355 (O_2355,N_19881,N_19824);
and UO_2356 (O_2356,N_19743,N_19540);
and UO_2357 (O_2357,N_19454,N_19276);
and UO_2358 (O_2358,N_19554,N_19990);
and UO_2359 (O_2359,N_19899,N_19646);
or UO_2360 (O_2360,N_19857,N_19216);
or UO_2361 (O_2361,N_19464,N_19466);
nand UO_2362 (O_2362,N_19776,N_19211);
nand UO_2363 (O_2363,N_19361,N_19625);
or UO_2364 (O_2364,N_19737,N_19676);
xor UO_2365 (O_2365,N_19732,N_19263);
nand UO_2366 (O_2366,N_19729,N_19817);
nor UO_2367 (O_2367,N_19931,N_19724);
and UO_2368 (O_2368,N_19714,N_19416);
nand UO_2369 (O_2369,N_19359,N_19976);
and UO_2370 (O_2370,N_19687,N_19745);
nor UO_2371 (O_2371,N_19740,N_19699);
or UO_2372 (O_2372,N_19218,N_19500);
nand UO_2373 (O_2373,N_19505,N_19430);
and UO_2374 (O_2374,N_19499,N_19221);
xnor UO_2375 (O_2375,N_19837,N_19767);
nand UO_2376 (O_2376,N_19489,N_19347);
nand UO_2377 (O_2377,N_19228,N_19674);
or UO_2378 (O_2378,N_19591,N_19828);
nand UO_2379 (O_2379,N_19561,N_19660);
xnor UO_2380 (O_2380,N_19592,N_19938);
nor UO_2381 (O_2381,N_19315,N_19498);
and UO_2382 (O_2382,N_19445,N_19828);
nor UO_2383 (O_2383,N_19940,N_19793);
nand UO_2384 (O_2384,N_19537,N_19945);
xor UO_2385 (O_2385,N_19584,N_19887);
nor UO_2386 (O_2386,N_19510,N_19590);
nand UO_2387 (O_2387,N_19563,N_19512);
and UO_2388 (O_2388,N_19733,N_19346);
or UO_2389 (O_2389,N_19649,N_19990);
or UO_2390 (O_2390,N_19729,N_19233);
xnor UO_2391 (O_2391,N_19463,N_19355);
xor UO_2392 (O_2392,N_19415,N_19995);
nand UO_2393 (O_2393,N_19400,N_19976);
nor UO_2394 (O_2394,N_19785,N_19253);
nand UO_2395 (O_2395,N_19516,N_19869);
nor UO_2396 (O_2396,N_19606,N_19740);
xnor UO_2397 (O_2397,N_19898,N_19977);
and UO_2398 (O_2398,N_19715,N_19208);
and UO_2399 (O_2399,N_19908,N_19367);
xor UO_2400 (O_2400,N_19747,N_19847);
nor UO_2401 (O_2401,N_19786,N_19230);
and UO_2402 (O_2402,N_19447,N_19236);
nor UO_2403 (O_2403,N_19880,N_19971);
and UO_2404 (O_2404,N_19858,N_19245);
or UO_2405 (O_2405,N_19958,N_19467);
nor UO_2406 (O_2406,N_19572,N_19301);
nand UO_2407 (O_2407,N_19557,N_19765);
or UO_2408 (O_2408,N_19937,N_19333);
and UO_2409 (O_2409,N_19358,N_19323);
nand UO_2410 (O_2410,N_19627,N_19768);
or UO_2411 (O_2411,N_19952,N_19918);
xor UO_2412 (O_2412,N_19878,N_19654);
nor UO_2413 (O_2413,N_19838,N_19227);
nand UO_2414 (O_2414,N_19822,N_19202);
nand UO_2415 (O_2415,N_19285,N_19743);
nor UO_2416 (O_2416,N_19964,N_19458);
nor UO_2417 (O_2417,N_19608,N_19845);
nand UO_2418 (O_2418,N_19740,N_19269);
or UO_2419 (O_2419,N_19389,N_19819);
or UO_2420 (O_2420,N_19694,N_19940);
nand UO_2421 (O_2421,N_19413,N_19681);
or UO_2422 (O_2422,N_19931,N_19613);
and UO_2423 (O_2423,N_19236,N_19312);
nor UO_2424 (O_2424,N_19866,N_19928);
and UO_2425 (O_2425,N_19375,N_19372);
nor UO_2426 (O_2426,N_19740,N_19796);
nor UO_2427 (O_2427,N_19428,N_19201);
xnor UO_2428 (O_2428,N_19532,N_19876);
nor UO_2429 (O_2429,N_19606,N_19271);
nor UO_2430 (O_2430,N_19831,N_19742);
xor UO_2431 (O_2431,N_19830,N_19917);
nor UO_2432 (O_2432,N_19330,N_19510);
or UO_2433 (O_2433,N_19556,N_19866);
and UO_2434 (O_2434,N_19304,N_19902);
xor UO_2435 (O_2435,N_19908,N_19298);
or UO_2436 (O_2436,N_19468,N_19846);
nor UO_2437 (O_2437,N_19264,N_19346);
nand UO_2438 (O_2438,N_19439,N_19642);
xnor UO_2439 (O_2439,N_19985,N_19225);
nor UO_2440 (O_2440,N_19721,N_19763);
or UO_2441 (O_2441,N_19551,N_19452);
xnor UO_2442 (O_2442,N_19329,N_19521);
xnor UO_2443 (O_2443,N_19365,N_19878);
nor UO_2444 (O_2444,N_19756,N_19591);
nor UO_2445 (O_2445,N_19993,N_19830);
nand UO_2446 (O_2446,N_19922,N_19862);
or UO_2447 (O_2447,N_19362,N_19599);
nor UO_2448 (O_2448,N_19862,N_19696);
nor UO_2449 (O_2449,N_19624,N_19550);
xor UO_2450 (O_2450,N_19339,N_19332);
nand UO_2451 (O_2451,N_19493,N_19871);
and UO_2452 (O_2452,N_19944,N_19802);
or UO_2453 (O_2453,N_19507,N_19932);
or UO_2454 (O_2454,N_19463,N_19399);
nor UO_2455 (O_2455,N_19790,N_19987);
or UO_2456 (O_2456,N_19979,N_19593);
nand UO_2457 (O_2457,N_19994,N_19831);
nand UO_2458 (O_2458,N_19423,N_19994);
nand UO_2459 (O_2459,N_19918,N_19577);
and UO_2460 (O_2460,N_19605,N_19699);
or UO_2461 (O_2461,N_19686,N_19211);
xnor UO_2462 (O_2462,N_19614,N_19777);
xnor UO_2463 (O_2463,N_19575,N_19970);
and UO_2464 (O_2464,N_19461,N_19935);
nand UO_2465 (O_2465,N_19880,N_19863);
nand UO_2466 (O_2466,N_19501,N_19280);
and UO_2467 (O_2467,N_19962,N_19533);
or UO_2468 (O_2468,N_19783,N_19606);
and UO_2469 (O_2469,N_19659,N_19887);
or UO_2470 (O_2470,N_19919,N_19606);
and UO_2471 (O_2471,N_19839,N_19253);
nand UO_2472 (O_2472,N_19218,N_19580);
and UO_2473 (O_2473,N_19211,N_19589);
and UO_2474 (O_2474,N_19902,N_19311);
or UO_2475 (O_2475,N_19888,N_19639);
or UO_2476 (O_2476,N_19382,N_19257);
or UO_2477 (O_2477,N_19860,N_19573);
and UO_2478 (O_2478,N_19503,N_19911);
nand UO_2479 (O_2479,N_19763,N_19552);
nand UO_2480 (O_2480,N_19852,N_19940);
or UO_2481 (O_2481,N_19564,N_19743);
and UO_2482 (O_2482,N_19214,N_19581);
nand UO_2483 (O_2483,N_19464,N_19222);
and UO_2484 (O_2484,N_19337,N_19240);
and UO_2485 (O_2485,N_19816,N_19417);
and UO_2486 (O_2486,N_19764,N_19786);
and UO_2487 (O_2487,N_19362,N_19774);
and UO_2488 (O_2488,N_19429,N_19868);
nor UO_2489 (O_2489,N_19889,N_19285);
xor UO_2490 (O_2490,N_19624,N_19726);
nand UO_2491 (O_2491,N_19438,N_19624);
nand UO_2492 (O_2492,N_19469,N_19498);
nand UO_2493 (O_2493,N_19836,N_19609);
nor UO_2494 (O_2494,N_19830,N_19294);
nor UO_2495 (O_2495,N_19636,N_19704);
nor UO_2496 (O_2496,N_19653,N_19680);
xor UO_2497 (O_2497,N_19968,N_19328);
nor UO_2498 (O_2498,N_19482,N_19834);
nor UO_2499 (O_2499,N_19560,N_19462);
endmodule