module basic_1500_15000_2000_100_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_507,In_92);
xor U1 (N_1,In_1254,In_306);
nor U2 (N_2,In_186,In_697);
nor U3 (N_3,In_836,In_1467);
nand U4 (N_4,In_925,In_530);
or U5 (N_5,In_1471,In_1237);
nand U6 (N_6,In_578,In_1178);
nand U7 (N_7,In_1084,In_377);
nand U8 (N_8,In_207,In_918);
or U9 (N_9,In_111,In_457);
or U10 (N_10,In_596,In_1223);
nor U11 (N_11,In_83,In_786);
and U12 (N_12,In_832,In_1034);
or U13 (N_13,In_282,In_78);
nor U14 (N_14,In_1390,In_843);
nand U15 (N_15,In_287,In_985);
and U16 (N_16,In_436,In_738);
and U17 (N_17,In_1456,In_588);
xnor U18 (N_18,In_120,In_12);
and U19 (N_19,In_568,In_945);
and U20 (N_20,In_1392,In_423);
and U21 (N_21,In_634,In_1410);
xor U22 (N_22,In_509,In_725);
nand U23 (N_23,In_67,In_651);
or U24 (N_24,In_1138,In_550);
or U25 (N_25,In_869,In_100);
or U26 (N_26,In_922,In_1062);
xnor U27 (N_27,In_890,In_1184);
xnor U28 (N_28,In_1336,In_876);
nand U29 (N_29,In_456,In_487);
nor U30 (N_30,In_52,In_1249);
and U31 (N_31,In_779,In_1337);
and U32 (N_32,In_212,In_899);
xor U33 (N_33,In_381,In_894);
and U34 (N_34,In_1141,In_424);
xnor U35 (N_35,In_956,In_136);
and U36 (N_36,In_1308,In_1204);
or U37 (N_37,In_965,In_1225);
nor U38 (N_38,In_1001,In_883);
nor U39 (N_39,In_1194,In_967);
and U40 (N_40,In_1380,In_388);
xor U41 (N_41,In_1140,In_574);
nor U42 (N_42,In_604,In_15);
nor U43 (N_43,In_1270,In_1195);
or U44 (N_44,In_1176,In_1170);
or U45 (N_45,In_1061,In_446);
xor U46 (N_46,In_122,In_13);
or U47 (N_47,In_1290,In_650);
nand U48 (N_48,In_1085,In_1401);
and U49 (N_49,In_1475,In_327);
and U50 (N_50,In_1422,In_426);
and U51 (N_51,In_1375,In_1257);
and U52 (N_52,In_379,In_102);
nor U53 (N_53,In_25,In_142);
nor U54 (N_54,In_368,In_1177);
nor U55 (N_55,In_514,In_587);
or U56 (N_56,In_1378,In_630);
xnor U57 (N_57,In_295,In_517);
nor U58 (N_58,In_953,In_230);
nor U59 (N_59,In_1108,In_1320);
nor U60 (N_60,In_1372,In_577);
or U61 (N_61,In_293,In_1165);
nand U62 (N_62,In_453,In_157);
xnor U63 (N_63,In_889,In_76);
and U64 (N_64,In_735,In_780);
and U65 (N_65,In_1027,In_320);
and U66 (N_66,In_93,In_104);
or U67 (N_67,In_1173,In_1368);
nand U68 (N_68,In_600,In_1030);
nand U69 (N_69,In_584,In_328);
nand U70 (N_70,In_661,In_5);
xnor U71 (N_71,In_1098,In_1388);
and U72 (N_72,In_940,In_752);
and U73 (N_73,In_916,In_1124);
xor U74 (N_74,In_713,In_166);
nor U75 (N_75,In_1384,In_97);
xnor U76 (N_76,In_1341,In_21);
and U77 (N_77,In_895,In_573);
nand U78 (N_78,In_1117,In_227);
and U79 (N_79,In_989,In_522);
and U80 (N_80,In_30,In_1219);
and U81 (N_81,In_810,In_515);
or U82 (N_82,In_1272,In_1258);
and U83 (N_83,In_422,In_1040);
or U84 (N_84,In_777,In_971);
xnor U85 (N_85,In_276,In_694);
nor U86 (N_86,In_891,In_586);
nand U87 (N_87,In_1322,In_837);
and U88 (N_88,In_109,In_753);
nor U89 (N_89,In_127,In_77);
or U90 (N_90,In_884,In_347);
nand U91 (N_91,In_937,In_490);
or U92 (N_92,In_265,In_94);
or U93 (N_93,In_1186,In_565);
nand U94 (N_94,In_299,In_66);
nor U95 (N_95,In_1492,In_405);
nand U96 (N_96,In_387,In_36);
or U97 (N_97,In_314,In_480);
xor U98 (N_98,In_110,In_666);
and U99 (N_99,In_1075,In_318);
and U100 (N_100,In_499,In_26);
and U101 (N_101,In_590,In_668);
or U102 (N_102,In_952,In_165);
nand U103 (N_103,In_1228,In_454);
nor U104 (N_104,In_244,In_1367);
nand U105 (N_105,In_1450,In_824);
nor U106 (N_106,In_1160,In_1215);
nor U107 (N_107,In_121,In_325);
and U108 (N_108,In_551,In_417);
and U109 (N_109,In_1139,In_1303);
or U110 (N_110,In_613,In_467);
nand U111 (N_111,In_1136,In_1291);
nand U112 (N_112,In_313,In_995);
nand U113 (N_113,In_431,In_1079);
or U114 (N_114,In_137,In_205);
or U115 (N_115,In_112,In_1469);
or U116 (N_116,In_776,In_1052);
and U117 (N_117,In_315,In_428);
or U118 (N_118,In_444,In_1312);
and U119 (N_119,In_1455,In_1196);
and U120 (N_120,In_385,In_1175);
and U121 (N_121,In_406,In_855);
and U122 (N_122,In_914,In_475);
and U123 (N_123,In_858,In_1025);
nand U124 (N_124,In_1042,In_1333);
or U125 (N_125,In_962,In_737);
and U126 (N_126,In_397,In_188);
or U127 (N_127,In_1125,In_1241);
nor U128 (N_128,In_116,In_744);
xnor U129 (N_129,In_1485,In_508);
xnor U130 (N_130,In_362,In_513);
and U131 (N_131,In_45,In_303);
nor U132 (N_132,In_1216,In_791);
xnor U133 (N_133,In_479,In_210);
and U134 (N_134,In_236,In_1438);
or U135 (N_135,In_1122,In_1360);
nand U136 (N_136,In_770,In_486);
and U137 (N_137,In_27,In_167);
and U138 (N_138,In_548,In_11);
xnor U139 (N_139,In_905,In_1123);
xor U140 (N_140,In_1484,In_1432);
nor U141 (N_141,In_881,In_250);
nor U142 (N_142,In_40,In_393);
nand U143 (N_143,In_168,In_699);
or U144 (N_144,In_1038,In_1202);
xor U145 (N_145,In_72,In_1399);
nand U146 (N_146,In_337,In_82);
or U147 (N_147,In_1444,In_35);
or U148 (N_148,In_1259,In_373);
and U149 (N_149,In_174,In_1406);
and U150 (N_150,In_353,In_346);
and U151 (N_151,In_656,In_723);
nand U152 (N_152,N_124,In_1442);
and U153 (N_153,In_612,In_7);
nand U154 (N_154,In_864,In_981);
and U155 (N_155,In_979,In_223);
nor U156 (N_156,In_321,In_1089);
xnor U157 (N_157,In_1120,In_1449);
and U158 (N_158,In_1073,In_118);
and U159 (N_159,In_1363,In_1376);
xor U160 (N_160,In_1133,N_45);
nand U161 (N_161,In_611,In_563);
xnor U162 (N_162,In_526,In_598);
and U163 (N_163,N_20,In_476);
nor U164 (N_164,In_156,In_255);
nor U165 (N_165,In_709,In_601);
and U166 (N_166,In_863,N_28);
nand U167 (N_167,In_710,In_1427);
xnor U168 (N_168,In_1226,In_1103);
or U169 (N_169,In_857,In_1386);
and U170 (N_170,In_284,In_196);
and U171 (N_171,In_660,In_736);
nand U172 (N_172,In_0,In_296);
xor U173 (N_173,In_1497,In_572);
xnor U174 (N_174,In_18,In_977);
nand U175 (N_175,In_835,In_705);
and U176 (N_176,In_474,In_1086);
or U177 (N_177,In_773,In_1113);
xnor U178 (N_178,In_462,In_22);
nand U179 (N_179,In_1131,In_1002);
or U180 (N_180,N_48,In_214);
nor U181 (N_181,In_412,In_1244);
and U182 (N_182,In_1317,In_1188);
nand U183 (N_183,In_286,N_11);
and U184 (N_184,In_1096,In_504);
nor U185 (N_185,In_1081,In_622);
nor U186 (N_186,In_473,In_1187);
nor U187 (N_187,In_481,In_242);
and U188 (N_188,In_1150,In_1477);
nand U189 (N_189,In_351,In_834);
nor U190 (N_190,In_759,In_825);
nand U191 (N_191,In_974,In_963);
nor U192 (N_192,In_65,In_542);
nor U193 (N_193,In_867,In_350);
or U194 (N_194,N_14,In_463);
nor U195 (N_195,N_89,In_966);
nor U196 (N_196,In_245,In_399);
xor U197 (N_197,In_620,In_1326);
nand U198 (N_198,In_332,In_363);
nand U199 (N_199,In_610,In_189);
and U200 (N_200,In_401,N_146);
and U201 (N_201,In_529,In_859);
nor U202 (N_202,In_947,In_781);
and U203 (N_203,N_64,In_460);
xor U204 (N_204,In_637,In_128);
and U205 (N_205,In_1354,In_430);
and U206 (N_206,In_1134,In_996);
nor U207 (N_207,In_1153,In_1301);
xor U208 (N_208,In_354,In_256);
nor U209 (N_209,In_1402,In_768);
nand U210 (N_210,In_1277,In_930);
xor U211 (N_211,In_264,In_224);
and U212 (N_212,In_570,In_1383);
nand U213 (N_213,In_980,In_356);
and U214 (N_214,N_63,In_410);
nor U215 (N_215,In_434,In_555);
nor U216 (N_216,N_55,In_557);
nor U217 (N_217,In_1049,In_689);
nand U218 (N_218,In_10,In_621);
or U219 (N_219,In_849,In_1221);
or U220 (N_220,In_144,In_1269);
nor U221 (N_221,In_263,In_1371);
nand U222 (N_222,N_106,In_202);
nor U223 (N_223,In_919,In_1035);
xor U224 (N_224,In_798,In_1490);
nor U225 (N_225,In_8,In_1071);
or U226 (N_226,In_1332,In_1126);
nand U227 (N_227,In_731,In_788);
or U228 (N_228,In_247,In_829);
or U229 (N_229,In_31,In_305);
nand U230 (N_230,In_783,In_1499);
nand U231 (N_231,In_1404,In_758);
and U232 (N_232,In_846,In_330);
nor U233 (N_233,In_1129,In_926);
and U234 (N_234,In_931,In_342);
or U235 (N_235,In_1200,In_969);
nand U236 (N_236,In_1026,In_1193);
or U237 (N_237,In_811,In_1130);
xnor U238 (N_238,In_1327,In_145);
nand U239 (N_239,In_1415,In_54);
xnor U240 (N_240,In_1171,In_349);
or U241 (N_241,In_1395,In_1099);
nor U242 (N_242,N_9,In_638);
and U243 (N_243,In_280,In_1053);
nand U244 (N_244,In_63,In_763);
xor U245 (N_245,In_690,In_856);
or U246 (N_246,In_813,In_98);
nor U247 (N_247,N_27,In_149);
nand U248 (N_248,In_1435,In_603);
nand U249 (N_249,In_334,In_179);
nand U250 (N_250,In_1345,N_145);
or U251 (N_251,In_1114,In_1447);
or U252 (N_252,In_643,In_1058);
and U253 (N_253,In_1431,In_975);
nor U254 (N_254,In_316,In_851);
and U255 (N_255,In_627,In_105);
nand U256 (N_256,In_564,In_1107);
and U257 (N_257,In_1016,In_283);
nand U258 (N_258,In_389,In_75);
xnor U259 (N_259,In_521,N_70);
xor U260 (N_260,In_964,In_1055);
nor U261 (N_261,In_1267,In_392);
nand U262 (N_262,In_701,In_1112);
nand U263 (N_263,N_149,In_614);
nand U264 (N_264,In_1292,In_271);
and U265 (N_265,In_1157,N_43);
nand U266 (N_266,In_103,In_1282);
xnor U267 (N_267,In_1210,In_942);
nor U268 (N_268,In_240,In_292);
or U269 (N_269,In_1095,In_1069);
or U270 (N_270,In_133,In_520);
nand U271 (N_271,N_41,In_175);
or U272 (N_272,In_148,In_41);
and U273 (N_273,In_19,In_1213);
nand U274 (N_274,In_1080,In_961);
or U275 (N_275,In_724,In_976);
or U276 (N_276,In_472,In_1146);
and U277 (N_277,In_88,In_1064);
or U278 (N_278,In_1247,In_1018);
xor U279 (N_279,In_57,In_743);
nor U280 (N_280,In_1393,In_277);
nor U281 (N_281,In_913,In_317);
or U282 (N_282,In_1032,N_84);
and U283 (N_283,In_567,In_1287);
nand U284 (N_284,N_127,In_23);
nor U285 (N_285,In_939,In_1208);
nor U286 (N_286,In_1305,In_579);
nand U287 (N_287,In_657,In_380);
xnor U288 (N_288,In_158,In_774);
or U289 (N_289,In_1232,In_172);
and U290 (N_290,In_1242,In_845);
nor U291 (N_291,In_1284,In_1077);
or U292 (N_292,In_1169,In_452);
nand U293 (N_293,In_132,In_445);
and U294 (N_294,In_421,In_1496);
and U295 (N_295,In_652,In_1364);
or U296 (N_296,N_88,In_853);
or U297 (N_297,In_478,In_441);
and U298 (N_298,In_635,In_1405);
nand U299 (N_299,N_87,In_451);
nor U300 (N_300,In_544,In_750);
or U301 (N_301,In_978,In_1275);
and U302 (N_302,N_144,In_1183);
or U303 (N_303,In_1295,In_807);
and U304 (N_304,In_778,In_512);
xnor U305 (N_305,In_806,N_167);
xnor U306 (N_306,In_669,In_532);
and U307 (N_307,In_273,In_1429);
or U308 (N_308,In_59,In_949);
or U309 (N_309,In_391,In_278);
nor U310 (N_310,In_1033,N_21);
nor U311 (N_311,In_360,In_48);
nand U312 (N_312,In_789,In_968);
nor U313 (N_313,In_345,N_57);
nor U314 (N_314,In_1464,In_184);
nor U315 (N_315,N_227,In_497);
xor U316 (N_316,In_1350,In_902);
nand U317 (N_317,N_36,N_40);
nor U318 (N_318,In_928,In_1201);
or U319 (N_319,In_695,In_1458);
nor U320 (N_320,In_1236,In_301);
nand U321 (N_321,In_866,In_576);
nand U322 (N_322,N_170,In_91);
nor U323 (N_323,In_231,In_169);
or U324 (N_324,N_134,In_1206);
and U325 (N_325,N_190,In_416);
or U326 (N_326,In_324,In_997);
nand U327 (N_327,In_691,In_496);
nor U328 (N_328,In_1211,N_39);
or U329 (N_329,In_617,In_1359);
xor U330 (N_330,In_907,In_17);
and U331 (N_331,In_1212,In_43);
nand U332 (N_332,In_192,In_193);
and U333 (N_333,In_1324,In_1209);
nor U334 (N_334,In_483,In_1421);
xor U335 (N_335,In_1065,In_1203);
nor U336 (N_336,In_1243,N_71);
nor U337 (N_337,In_470,In_1101);
nand U338 (N_338,In_1279,In_1022);
xnor U339 (N_339,In_782,In_817);
or U340 (N_340,In_801,In_455);
nand U341 (N_341,In_927,In_1423);
xor U342 (N_342,In_411,N_265);
or U343 (N_343,In_747,In_55);
nand U344 (N_344,In_527,In_1000);
nand U345 (N_345,In_983,In_716);
and U346 (N_346,In_1056,In_1274);
and U347 (N_347,N_102,In_1222);
nand U348 (N_348,In_646,In_672);
or U349 (N_349,In_352,In_1434);
xor U350 (N_350,In_1334,N_273);
nor U351 (N_351,In_402,In_1050);
xnor U352 (N_352,N_66,In_715);
or U353 (N_353,In_729,In_809);
nand U354 (N_354,In_1391,N_275);
nand U355 (N_355,In_734,In_663);
and U356 (N_356,In_331,In_870);
nor U357 (N_357,In_1381,N_139);
xnor U358 (N_358,In_90,In_1082);
nor U359 (N_359,N_100,In_221);
or U360 (N_360,N_161,N_44);
nand U361 (N_361,In_772,In_528);
and U362 (N_362,In_1309,In_1090);
or U363 (N_363,N_65,In_390);
nand U364 (N_364,In_685,In_2);
nand U365 (N_365,In_1009,In_921);
nor U366 (N_366,In_1044,In_1465);
or U367 (N_367,In_1362,In_254);
and U368 (N_368,In_6,In_123);
or U369 (N_369,In_1047,In_1088);
xor U370 (N_370,In_1468,In_712);
or U371 (N_371,In_260,In_270);
and U372 (N_372,In_429,In_1306);
or U373 (N_373,In_771,In_419);
and U374 (N_374,In_569,In_39);
or U375 (N_375,In_1298,In_1007);
nand U376 (N_376,In_1012,N_7);
nor U377 (N_377,In_746,In_1043);
nor U378 (N_378,N_51,In_1330);
nor U379 (N_379,N_142,In_131);
nand U380 (N_380,In_524,N_243);
xor U381 (N_381,In_721,N_19);
and U382 (N_382,In_593,In_1473);
nor U383 (N_383,In_450,In_225);
nand U384 (N_384,In_1351,N_268);
nor U385 (N_385,In_258,In_991);
and U386 (N_386,N_114,In_1266);
nand U387 (N_387,In_1297,In_992);
xor U388 (N_388,N_256,In_234);
xnor U389 (N_389,In_1460,In_289);
nor U390 (N_390,In_1353,In_203);
and U391 (N_391,In_1433,In_1036);
or U392 (N_392,N_199,N_181);
or U393 (N_393,In_369,In_176);
nand U394 (N_394,In_1229,In_639);
and U395 (N_395,N_203,N_165);
xor U396 (N_396,In_311,N_26);
or U397 (N_397,In_541,In_150);
nand U398 (N_398,In_605,N_175);
or U399 (N_399,In_1245,In_425);
and U400 (N_400,In_464,In_117);
and U401 (N_401,In_1239,In_233);
nand U402 (N_402,In_1425,In_631);
xnor U403 (N_403,In_1158,N_299);
or U404 (N_404,In_1394,In_1087);
xor U405 (N_405,N_220,In_711);
nand U406 (N_406,In_1357,In_1005);
nand U407 (N_407,In_181,In_970);
xnor U408 (N_408,In_1224,In_560);
and U409 (N_409,In_1299,In_687);
nand U410 (N_410,N_288,In_664);
xnor U411 (N_411,N_200,N_53);
nor U412 (N_412,In_885,In_850);
or U413 (N_413,In_262,In_1006);
nor U414 (N_414,N_115,N_221);
xor U415 (N_415,N_262,In_1358);
nand U416 (N_416,In_785,N_33);
or U417 (N_417,In_1121,N_193);
nor U418 (N_418,N_205,In_1255);
and U419 (N_419,In_153,In_183);
nand U420 (N_420,N_224,In_159);
or U421 (N_421,In_1028,In_440);
xor U422 (N_422,N_147,In_683);
nand U423 (N_423,In_396,In_1280);
and U424 (N_424,In_465,In_1314);
xor U425 (N_425,In_449,In_535);
nor U426 (N_426,N_245,N_185);
nor U427 (N_427,In_1066,In_1037);
nand U428 (N_428,In_547,In_340);
and U429 (N_429,In_1256,In_1181);
xor U430 (N_430,In_239,In_1168);
and U431 (N_431,In_364,In_365);
xnor U432 (N_432,In_1461,N_141);
nand U433 (N_433,In_336,In_162);
nor U434 (N_434,In_1179,In_190);
or U435 (N_435,In_519,In_173);
and U436 (N_436,In_491,In_1343);
xnor U437 (N_437,In_1057,N_110);
nor U438 (N_438,In_822,In_1109);
xor U439 (N_439,In_414,In_243);
xor U440 (N_440,In_272,In_1489);
or U441 (N_441,In_154,N_289);
or U442 (N_442,In_329,N_204);
xnor U443 (N_443,In_119,In_482);
and U444 (N_444,In_754,In_268);
and U445 (N_445,N_159,In_152);
xnor U446 (N_446,In_1106,N_156);
xnor U447 (N_447,In_862,In_727);
or U448 (N_448,In_823,In_1454);
xnor U449 (N_449,In_757,In_1340);
xnor U450 (N_450,In_717,N_314);
xor U451 (N_451,N_202,In_161);
nand U452 (N_452,In_987,In_1457);
or U453 (N_453,N_316,In_696);
nor U454 (N_454,N_178,In_787);
or U455 (N_455,N_397,In_197);
or U456 (N_456,In_1011,In_1338);
nand U457 (N_457,N_429,In_1);
xnor U458 (N_458,In_804,In_87);
or U459 (N_459,In_505,N_382);
or U460 (N_460,In_495,In_171);
xor U461 (N_461,N_92,In_248);
and U462 (N_462,In_554,In_1488);
nor U463 (N_463,In_552,In_1264);
and U464 (N_464,In_1355,N_123);
or U465 (N_465,In_488,N_404);
nor U466 (N_466,In_868,N_380);
nor U467 (N_467,In_1017,N_356);
nor U468 (N_468,N_361,In_510);
nand U469 (N_469,In_1142,N_189);
and U470 (N_470,N_8,In_427);
or U471 (N_471,In_1481,N_305);
or U472 (N_472,In_439,In_677);
and U473 (N_473,In_160,In_409);
or U474 (N_474,N_90,N_120);
and U475 (N_475,In_126,In_879);
nand U476 (N_476,In_1365,N_318);
nor U477 (N_477,In_714,In_1091);
nor U478 (N_478,In_629,In_917);
and U479 (N_479,N_283,N_341);
xor U480 (N_480,In_1104,N_422);
or U481 (N_481,In_933,In_582);
nand U482 (N_482,In_831,N_350);
nand U483 (N_483,In_14,In_115);
xnor U484 (N_484,In_108,N_136);
nor U485 (N_485,N_47,In_178);
nand U486 (N_486,In_85,In_218);
nor U487 (N_487,In_545,In_370);
xor U488 (N_488,In_900,In_415);
xnor U489 (N_489,In_493,In_944);
nand U490 (N_490,In_1143,In_537);
and U491 (N_491,In_335,In_1161);
or U492 (N_492,N_427,In_1278);
and U493 (N_493,N_98,In_733);
or U494 (N_494,In_594,N_436);
nor U495 (N_495,In_1311,N_81);
or U496 (N_496,N_386,In_794);
nor U497 (N_497,N_23,N_315);
nand U498 (N_498,In_177,In_766);
or U499 (N_499,In_1220,In_359);
xor U500 (N_500,In_348,In_1105);
and U501 (N_501,In_920,In_1408);
nand U502 (N_502,N_286,N_342);
nor U503 (N_503,In_732,N_187);
nor U504 (N_504,N_16,N_432);
xor U505 (N_505,In_816,In_1482);
nor U506 (N_506,N_56,N_254);
and U507 (N_507,N_329,N_135);
nand U508 (N_508,In_1293,In_1192);
and U509 (N_509,In_1054,In_659);
or U510 (N_510,N_3,In_322);
nand U511 (N_511,In_447,In_267);
or U512 (N_512,In_237,N_270);
and U513 (N_513,In_908,In_861);
or U514 (N_514,In_403,In_1452);
nand U515 (N_515,In_616,In_294);
nor U516 (N_516,In_297,N_169);
or U517 (N_517,In_655,In_799);
or U518 (N_518,N_425,N_259);
or U519 (N_519,In_703,In_1102);
nor U520 (N_520,In_1411,N_381);
or U521 (N_521,N_133,In_309);
nand U522 (N_522,In_1318,In_1361);
and U523 (N_523,In_226,N_137);
nor U524 (N_524,In_312,N_439);
nor U525 (N_525,In_1045,In_523);
xnor U526 (N_526,N_431,In_61);
xor U527 (N_527,In_1093,N_287);
xor U528 (N_528,In_125,N_118);
and U529 (N_529,N_339,In_675);
and U530 (N_530,In_880,In_418);
or U531 (N_531,In_138,N_168);
or U532 (N_532,In_892,In_503);
and U533 (N_533,In_95,In_673);
nor U534 (N_534,N_5,N_292);
xnor U535 (N_535,In_595,In_1483);
xnor U536 (N_536,In_633,N_163);
and U537 (N_537,N_4,In_187);
nor U538 (N_538,In_923,In_848);
xnor U539 (N_539,In_9,In_1167);
xor U540 (N_540,In_540,N_430);
nor U541 (N_541,In_1479,In_795);
nand U542 (N_542,In_707,In_602);
nand U543 (N_543,N_171,In_840);
nand U544 (N_544,In_1029,In_706);
nor U545 (N_545,In_625,In_1486);
nand U546 (N_546,In_1041,In_459);
nor U547 (N_547,In_874,In_762);
nand U548 (N_548,In_1190,In_338);
and U549 (N_549,N_17,N_362);
nor U550 (N_550,N_232,N_395);
nor U551 (N_551,In_198,N_277);
xnor U552 (N_552,In_1135,In_182);
xor U553 (N_553,N_151,N_296);
xnor U554 (N_554,In_143,In_1374);
xor U555 (N_555,In_1097,N_388);
or U556 (N_556,N_129,In_830);
nor U557 (N_557,N_35,In_761);
xnor U558 (N_558,N_34,In_1155);
xor U559 (N_559,In_489,In_339);
or U560 (N_560,N_210,N_411);
nand U561 (N_561,In_106,N_272);
xnor U562 (N_562,In_485,N_211);
xnor U563 (N_563,In_571,In_1466);
and U564 (N_564,N_101,In_1230);
and U565 (N_565,N_86,N_173);
and U566 (N_566,In_86,In_1480);
nand U567 (N_567,In_1231,In_1015);
xnor U568 (N_568,In_498,N_412);
nand U569 (N_569,In_626,In_1412);
xnor U570 (N_570,N_410,In_1413);
nor U571 (N_571,In_1416,In_395);
or U572 (N_572,In_534,N_400);
nand U573 (N_573,N_424,In_1352);
nand U574 (N_574,In_130,In_950);
xnor U575 (N_575,N_209,In_49);
or U576 (N_576,N_331,In_458);
nand U577 (N_577,In_1180,In_304);
nor U578 (N_578,N_192,In_222);
or U579 (N_579,In_827,N_72);
nor U580 (N_580,N_446,In_1377);
and U581 (N_581,In_812,In_366);
or U582 (N_582,N_330,N_284);
and U583 (N_583,N_1,In_1389);
nor U584 (N_584,In_838,N_417);
or U585 (N_585,In_982,In_1074);
xnor U586 (N_586,N_73,In_371);
xnor U587 (N_587,In_1248,In_1285);
nor U588 (N_588,In_1013,In_300);
and U589 (N_589,N_58,N_398);
or U590 (N_590,N_321,In_1470);
or U591 (N_591,N_182,N_208);
or U592 (N_592,N_311,In_704);
nand U593 (N_593,N_437,In_81);
or U594 (N_594,In_372,In_561);
xnor U595 (N_595,In_688,In_682);
or U596 (N_596,In_1072,In_671);
nand U597 (N_597,In_266,In_194);
or U598 (N_598,In_929,In_959);
nand U599 (N_599,In_1437,In_760);
or U600 (N_600,N_492,N_516);
and U601 (N_601,In_955,In_558);
xnor U602 (N_602,N_269,In_769);
and U603 (N_603,In_581,In_307);
and U604 (N_604,In_993,N_249);
or U605 (N_605,In_50,N_18);
xor U606 (N_606,In_1443,N_130);
or U607 (N_607,N_237,N_543);
or U608 (N_608,In_873,In_745);
nor U609 (N_609,In_860,In_1441);
or U610 (N_610,N_93,N_558);
and U611 (N_611,N_440,N_502);
nor U612 (N_612,N_183,N_217);
xnor U613 (N_613,In_559,N_393);
nand U614 (N_614,In_676,N_488);
nor U615 (N_615,N_500,N_477);
nand U616 (N_616,N_548,In_291);
nor U617 (N_617,In_341,In_1453);
and U618 (N_618,In_438,In_1164);
nand U619 (N_619,In_826,In_1302);
nor U620 (N_620,N_117,N_399);
or U621 (N_621,N_570,In_308);
or U622 (N_622,N_433,In_1260);
xor U623 (N_623,N_271,N_496);
xor U624 (N_624,N_459,N_153);
or U625 (N_625,In_1198,In_343);
nor U626 (N_626,In_803,N_461);
nand U627 (N_627,In_1403,In_793);
and U628 (N_628,N_94,In_279);
xnor U629 (N_629,In_1021,N_302);
xnor U630 (N_630,N_357,N_378);
nand U631 (N_631,In_1174,In_1092);
nor U632 (N_632,N_363,In_302);
or U633 (N_633,N_294,In_442);
nor U634 (N_634,N_248,N_239);
xor U635 (N_635,In_642,N_46);
or U636 (N_636,N_263,In_562);
nand U637 (N_637,N_367,N_463);
or U638 (N_638,In_1385,In_1116);
nand U639 (N_639,N_409,N_258);
and U640 (N_640,In_720,N_462);
nand U641 (N_641,In_47,In_1420);
and U642 (N_642,In_252,In_274);
nor U643 (N_643,In_323,N_423);
and U644 (N_644,In_1147,N_313);
and U645 (N_645,N_69,N_590);
nor U646 (N_646,N_74,In_238);
nor U647 (N_647,N_31,N_513);
xnor U648 (N_648,In_232,In_1024);
or U649 (N_649,N_253,In_1145);
nand U650 (N_650,In_654,N_534);
xor U651 (N_651,In_1235,In_893);
xor U652 (N_652,N_504,N_392);
xnor U653 (N_653,In_1476,In_546);
nor U654 (N_654,N_351,N_561);
nand U655 (N_655,In_201,In_139);
and U656 (N_656,N_6,N_125);
and U657 (N_657,N_352,N_498);
and U658 (N_658,In_1039,In_805);
nand U659 (N_659,In_24,N_402);
or U660 (N_660,In_1335,N_300);
nor U661 (N_661,In_1440,In_680);
xor U662 (N_662,In_319,In_180);
xor U663 (N_663,In_854,In_461);
nor U664 (N_664,In_1207,N_550);
xnor U665 (N_665,In_46,N_503);
nand U666 (N_666,N_520,In_1472);
or U667 (N_667,In_934,N_241);
xor U668 (N_668,N_585,In_797);
nor U669 (N_669,N_401,N_547);
xor U670 (N_670,N_415,In_935);
and U671 (N_671,In_326,In_1325);
and U672 (N_672,In_344,N_186);
or U673 (N_673,In_1307,N_379);
xnor U674 (N_674,In_585,N_335);
nor U675 (N_675,N_565,In_1078);
or U676 (N_676,N_99,In_468);
or U677 (N_677,N_279,N_317);
xnor U678 (N_678,In_994,N_68);
nand U679 (N_679,N_443,N_337);
or U680 (N_680,In_986,In_665);
or U681 (N_681,In_437,N_301);
or U682 (N_682,In_53,N_180);
and U683 (N_683,N_304,In_538);
nand U684 (N_684,In_722,In_51);
nand U685 (N_685,N_421,In_204);
xor U686 (N_686,N_128,In_151);
nor U687 (N_687,N_435,N_59);
nor U688 (N_688,N_107,In_549);
and U689 (N_689,N_230,In_742);
nand U690 (N_690,N_282,In_909);
nor U691 (N_691,N_238,N_291);
xnor U692 (N_692,In_62,N_80);
nand U693 (N_693,In_938,In_220);
nand U694 (N_694,N_479,N_177);
and U695 (N_695,N_236,In_719);
nand U696 (N_696,N_38,N_553);
nor U697 (N_697,N_428,N_15);
and U698 (N_698,N_491,In_200);
or U699 (N_699,In_1197,In_1424);
nand U700 (N_700,In_155,In_764);
nand U701 (N_701,N_261,In_1132);
and U702 (N_702,N_214,N_326);
or U703 (N_703,N_541,N_510);
xnor U704 (N_704,N_562,N_50);
xnor U705 (N_705,In_877,N_377);
xnor U706 (N_706,In_466,In_1346);
or U707 (N_707,N_372,In_1185);
nand U708 (N_708,N_581,N_226);
and U709 (N_709,N_371,N_111);
and U710 (N_710,In_833,In_960);
or U711 (N_711,N_387,N_348);
nor U712 (N_712,In_702,In_1100);
nand U713 (N_713,In_469,N_154);
or U714 (N_714,In_692,N_360);
or U715 (N_715,N_368,In_398);
nor U716 (N_716,N_176,N_460);
and U717 (N_717,In_249,In_1316);
or U718 (N_718,N_540,N_577);
and U719 (N_719,In_375,In_700);
nand U720 (N_720,In_1396,N_467);
nand U721 (N_721,In_80,N_96);
nor U722 (N_722,N_508,N_519);
or U723 (N_723,In_1014,N_524);
and U724 (N_724,N_408,N_472);
nand U725 (N_725,N_276,In_432);
or U726 (N_726,N_471,In_1119);
and U727 (N_727,N_438,N_567);
and U728 (N_728,In_1407,In_32);
xor U729 (N_729,N_242,N_246);
and U730 (N_730,In_1262,In_1289);
xor U731 (N_731,In_615,N_160);
nand U732 (N_732,In_257,In_79);
nand U733 (N_733,In_1323,In_1339);
nand U734 (N_734,In_84,In_649);
nand U735 (N_735,N_166,N_179);
nor U736 (N_736,In_382,In_141);
nor U737 (N_737,In_640,In_357);
xnor U738 (N_738,N_528,N_445);
and U739 (N_739,In_1268,N_201);
and U740 (N_740,N_599,In_275);
and U741 (N_741,N_507,In_670);
nand U742 (N_742,N_61,N_584);
xor U743 (N_743,In_448,N_105);
and U744 (N_744,In_1253,N_515);
xor U745 (N_745,N_546,In_539);
nor U746 (N_746,In_404,N_518);
or U747 (N_747,In_820,In_871);
nand U748 (N_748,N_589,In_89);
nand U749 (N_749,N_481,In_241);
nor U750 (N_750,In_828,In_74);
xor U751 (N_751,N_78,N_375);
nand U752 (N_752,N_686,In_674);
and U753 (N_753,In_872,N_158);
xor U754 (N_754,N_713,N_689);
nand U755 (N_755,N_613,N_434);
or U756 (N_756,N_307,N_555);
or U757 (N_757,In_1238,N_692);
or U758 (N_758,In_730,N_736);
nand U759 (N_759,In_69,In_839);
nor U760 (N_760,N_603,In_882);
nand U761 (N_761,In_841,N_624);
and U762 (N_762,In_998,In_1366);
and U763 (N_763,In_500,N_470);
nor U764 (N_764,N_523,N_654);
xnor U765 (N_765,In_1446,In_800);
or U766 (N_766,N_310,In_135);
and U767 (N_767,N_549,N_219);
and U768 (N_768,N_122,N_451);
nor U769 (N_769,In_678,N_582);
nor U770 (N_770,N_672,N_661);
or U771 (N_771,N_499,In_756);
xnor U772 (N_772,In_1451,N_24);
nand U773 (N_773,In_290,N_252);
nor U774 (N_774,N_490,N_740);
nor U775 (N_775,N_714,In_386);
or U776 (N_776,N_652,In_653);
nand U777 (N_777,N_116,N_629);
xor U778 (N_778,In_1349,In_1495);
or U779 (N_779,In_99,In_384);
xnor U780 (N_780,N_666,In_140);
nor U781 (N_781,N_625,N_630);
nand U782 (N_782,N_456,N_91);
xor U783 (N_783,N_207,In_16);
and U784 (N_784,N_669,In_814);
or U785 (N_785,N_675,N_349);
nand U786 (N_786,N_701,In_435);
nor U787 (N_787,N_578,In_1426);
and U788 (N_788,In_1273,N_697);
nand U789 (N_789,N_75,In_1217);
and U790 (N_790,N_525,In_628);
nor U791 (N_791,N_306,N_213);
and U792 (N_792,N_359,In_932);
or U793 (N_793,In_973,In_958);
or U794 (N_794,N_366,In_34);
nand U795 (N_795,N_728,N_643);
xor U796 (N_796,N_607,N_730);
nand U797 (N_797,N_468,N_685);
or U798 (N_798,N_702,In_897);
xnor U799 (N_799,In_1296,N_389);
or U800 (N_800,N_517,N_108);
nand U801 (N_801,N_679,N_483);
and U802 (N_802,N_484,In_209);
nand U803 (N_803,N_648,In_269);
or U804 (N_804,N_614,In_1162);
and U805 (N_805,In_1400,N_251);
nand U806 (N_806,N_396,In_477);
xnor U807 (N_807,In_1115,In_1369);
or U808 (N_808,N_152,In_1286);
and U809 (N_809,N_191,N_298);
or U810 (N_810,N_621,N_97);
nor U811 (N_811,N_267,N_698);
nor U812 (N_812,N_512,N_592);
and U813 (N_813,In_1059,In_1261);
xor U814 (N_814,N_343,N_234);
nor U815 (N_815,In_367,N_197);
nor U816 (N_816,N_601,N_580);
nand U817 (N_817,In_948,N_700);
nand U818 (N_818,In_1159,In_1128);
nor U819 (N_819,N_651,N_85);
nor U820 (N_820,N_391,N_83);
nor U821 (N_821,N_529,N_726);
nor U822 (N_822,In_259,N_662);
or U823 (N_823,In_64,N_29);
and U824 (N_824,N_478,In_943);
xnor U825 (N_825,N_257,N_67);
or U826 (N_826,N_95,In_20);
nor U827 (N_827,N_452,N_441);
xor U828 (N_828,N_667,In_591);
and U829 (N_829,N_636,N_450);
nand U830 (N_830,N_358,N_476);
nor U831 (N_831,In_1398,N_419);
xnor U832 (N_832,In_765,N_594);
nand U833 (N_833,N_143,In_1068);
nand U834 (N_834,N_526,N_568);
and U835 (N_835,N_413,In_1294);
xor U836 (N_836,N_748,In_1331);
nor U837 (N_837,In_728,N_223);
and U838 (N_838,N_537,N_355);
and U839 (N_839,N_749,In_1118);
and U840 (N_840,In_1191,N_196);
or U841 (N_841,N_655,N_328);
and U842 (N_842,In_58,N_574);
nor U843 (N_843,N_681,In_1397);
xnor U844 (N_844,In_1370,In_219);
and U845 (N_845,In_1003,In_553);
nor U846 (N_846,In_501,N_466);
nor U847 (N_847,In_1060,N_551);
and U848 (N_848,N_103,In_1265);
and U849 (N_849,N_712,N_708);
nand U850 (N_850,N_324,N_646);
or U851 (N_851,N_746,N_303);
or U852 (N_852,N_572,In_191);
and U853 (N_853,N_76,In_818);
nor U854 (N_854,N_593,N_416);
or U855 (N_855,N_140,In_533);
xor U856 (N_856,N_247,N_442);
xnor U857 (N_857,N_719,In_708);
or U858 (N_858,In_984,N_347);
or U859 (N_859,N_532,N_126);
xor U860 (N_860,N_340,N_737);
or U861 (N_861,In_1329,N_694);
nand U862 (N_862,In_1031,N_30);
or U863 (N_863,In_910,N_617);
xor U864 (N_864,N_742,N_42);
and U865 (N_865,In_215,N_738);
xnor U866 (N_866,In_358,In_1276);
nor U867 (N_867,N_619,In_1004);
or U868 (N_868,In_1205,N_79);
xnor U869 (N_869,N_721,N_618);
nand U870 (N_870,N_216,N_229);
and U871 (N_871,In_901,In_1347);
nor U872 (N_872,In_896,In_288);
nor U873 (N_873,In_681,N_215);
and U874 (N_874,N_622,N_673);
xnor U875 (N_875,In_56,N_13);
xnor U876 (N_876,N_627,N_49);
or U877 (N_877,In_1166,In_1094);
and U878 (N_878,In_886,N_22);
nand U879 (N_879,N_709,N_695);
xnor U880 (N_880,In_1373,N_720);
or U881 (N_881,N_255,In_1227);
nand U882 (N_882,N_545,N_383);
and U883 (N_883,N_119,In_1348);
nor U884 (N_884,In_1313,In_941);
or U885 (N_885,In_1310,N_486);
and U886 (N_886,N_725,N_290);
and U887 (N_887,In_107,N_597);
nand U888 (N_888,N_623,N_527);
xor U889 (N_889,N_370,In_206);
nand U890 (N_890,In_821,In_1023);
and U891 (N_891,N_744,N_650);
and U892 (N_892,N_683,N_113);
nand U893 (N_893,In_1382,In_990);
or U894 (N_894,In_333,N_374);
or U895 (N_895,In_1445,In_748);
nor U896 (N_896,N_678,N_390);
or U897 (N_897,In_531,N_676);
nand U898 (N_898,N_323,N_633);
nand U899 (N_899,In_211,N_162);
or U900 (N_900,N_474,In_253);
and U901 (N_901,N_787,In_589);
nor U902 (N_902,In_285,In_1067);
nor U903 (N_903,N_771,N_722);
nor U904 (N_904,In_1083,N_309);
nand U905 (N_905,In_1252,In_413);
xnor U906 (N_906,N_795,In_71);
nand U907 (N_907,N_588,N_691);
xnor U908 (N_908,In_420,N_121);
nor U909 (N_909,In_37,In_888);
nand U910 (N_910,N_826,In_1251);
nor U911 (N_911,N_864,N_631);
or U912 (N_912,In_679,In_543);
nand U913 (N_913,In_1462,N_354);
and U914 (N_914,N_858,In_815);
xnor U915 (N_915,N_586,In_693);
nor U916 (N_916,N_731,N_278);
nor U917 (N_917,N_734,N_754);
xnor U918 (N_918,N_505,N_325);
nor U919 (N_919,In_195,N_172);
or U920 (N_920,N_591,In_647);
nand U921 (N_921,In_556,N_554);
nor U922 (N_922,In_957,In_511);
nor U923 (N_923,N_878,N_839);
nor U924 (N_924,N_628,N_206);
nor U925 (N_925,In_251,N_418);
xor U926 (N_926,N_535,In_407);
or U927 (N_927,N_539,In_1234);
nand U928 (N_928,N_608,In_518);
and U929 (N_929,In_1288,In_924);
xnor U930 (N_930,In_624,N_816);
nor U931 (N_931,N_638,N_832);
nand U932 (N_932,N_52,N_705);
or U933 (N_933,N_863,In_146);
and U934 (N_934,N_222,In_310);
or U935 (N_935,N_319,N_148);
nor U936 (N_936,N_457,N_804);
or U937 (N_937,In_1218,N_752);
nor U938 (N_938,N_364,N_426);
and U939 (N_939,N_327,In_1214);
xor U940 (N_940,In_101,In_1010);
nor U941 (N_941,N_322,N_822);
nand U942 (N_942,In_502,In_1163);
or U943 (N_943,In_68,N_369);
or U944 (N_944,In_684,In_898);
or U945 (N_945,In_1240,N_333);
nor U946 (N_946,In_903,N_817);
nand U947 (N_947,In_383,In_1019);
xnor U948 (N_948,N_674,N_420);
xor U949 (N_949,N_658,In_775);
nor U950 (N_950,In_1474,In_525);
or U951 (N_951,In_374,In_619);
or U952 (N_952,N_757,N_764);
or U953 (N_953,In_583,N_869);
xnor U954 (N_954,N_716,N_807);
and U955 (N_955,N_810,In_1154);
nor U956 (N_956,N_865,In_199);
nor U957 (N_957,N_266,In_1156);
and U958 (N_958,In_662,N_198);
and U959 (N_959,N_642,N_250);
nor U960 (N_960,N_704,N_849);
and U961 (N_961,In_1127,N_521);
xnor U962 (N_962,N_768,N_373);
nor U963 (N_963,In_636,N_696);
nor U964 (N_964,In_1478,N_790);
xor U965 (N_965,In_972,In_819);
nor U966 (N_966,N_818,In_887);
xnor U967 (N_967,N_762,N_844);
xnor U968 (N_968,In_946,In_1491);
or U969 (N_969,N_855,N_583);
xor U970 (N_970,In_433,N_747);
xor U971 (N_971,In_912,In_951);
or U972 (N_972,N_264,N_464);
and U973 (N_973,In_784,In_645);
and U974 (N_974,N_659,N_827);
xor U975 (N_975,N_829,N_895);
and U976 (N_976,N_743,In_658);
or U977 (N_977,In_1271,In_1498);
xor U978 (N_978,N_727,N_406);
nand U979 (N_979,In_755,N_536);
or U980 (N_980,N_898,N_732);
nor U981 (N_981,N_711,N_260);
xor U982 (N_982,N_32,N_774);
nor U983 (N_983,N_334,In_216);
xnor U984 (N_984,N_814,N_893);
nand U985 (N_985,N_825,N_830);
nand U986 (N_986,N_852,N_12);
or U987 (N_987,N_766,N_109);
and U988 (N_988,N_861,N_723);
nand U989 (N_989,In_134,N_480);
xnor U990 (N_990,In_1417,N_285);
nor U991 (N_991,N_612,N_564);
and U992 (N_992,N_533,In_847);
and U993 (N_993,N_632,N_782);
xor U994 (N_994,N_575,In_208);
nand U995 (N_995,N_131,In_1304);
and U996 (N_996,N_493,In_1321);
or U997 (N_997,N_887,N_587);
or U998 (N_998,N_857,N_212);
xnor U999 (N_999,In_4,N_859);
nand U1000 (N_1000,N_854,N_596);
nand U1001 (N_1001,In_667,In_361);
xor U1002 (N_1002,N_338,In_802);
xor U1003 (N_1003,N_376,In_394);
nor U1004 (N_1004,N_530,In_686);
or U1005 (N_1005,In_96,N_218);
nand U1006 (N_1006,In_73,In_1182);
or U1007 (N_1007,N_559,N_332);
and U1008 (N_1008,In_516,In_163);
nand U1009 (N_1009,In_718,N_240);
and U1010 (N_1010,N_274,In_246);
nor U1011 (N_1011,N_866,N_640);
xor U1012 (N_1012,N_780,In_790);
nand U1013 (N_1013,N_756,N_792);
xnor U1014 (N_1014,N_407,In_471);
xnor U1015 (N_1015,N_458,N_888);
or U1016 (N_1016,N_62,N_751);
xor U1017 (N_1017,N_609,N_403);
xnor U1018 (N_1018,In_494,In_623);
and U1019 (N_1019,N_345,In_213);
nand U1020 (N_1020,In_44,In_3);
or U1021 (N_1021,N_293,N_10);
or U1022 (N_1022,In_484,In_33);
and U1023 (N_1023,N_602,N_563);
xnor U1024 (N_1024,N_794,N_693);
nand U1025 (N_1025,N_824,In_1148);
or U1026 (N_1026,N_860,N_644);
nor U1027 (N_1027,N_699,N_788);
and U1028 (N_1028,N_649,N_453);
nand U1029 (N_1029,N_786,N_600);
xor U1030 (N_1030,In_378,In_1463);
xnor U1031 (N_1031,N_772,In_1199);
nand U1032 (N_1032,In_443,In_740);
xor U1033 (N_1033,N_677,In_235);
xor U1034 (N_1034,In_1439,In_865);
or U1035 (N_1035,In_607,In_878);
nand U1036 (N_1036,N_544,N_556);
or U1037 (N_1037,N_891,N_781);
or U1038 (N_1038,N_706,N_784);
and U1039 (N_1039,N_885,In_129);
xor U1040 (N_1040,N_871,In_1414);
nor U1041 (N_1041,N_884,In_1063);
and U1042 (N_1042,N_802,N_174);
nor U1043 (N_1043,N_823,In_1430);
nand U1044 (N_1044,In_1137,In_1263);
or U1045 (N_1045,N_573,N_485);
xnor U1046 (N_1046,N_605,N_715);
nor U1047 (N_1047,In_400,N_465);
nand U1048 (N_1048,N_635,N_112);
xnor U1049 (N_1049,N_475,N_875);
and U1050 (N_1050,N_955,In_1448);
xor U1051 (N_1051,N_876,In_988);
nor U1052 (N_1052,N_988,N_923);
nand U1053 (N_1053,N_25,N_320);
or U1054 (N_1054,N_615,In_1151);
nor U1055 (N_1055,In_261,N_913);
or U1056 (N_1056,N_915,N_896);
nor U1057 (N_1057,In_1111,N_606);
or U1058 (N_1058,N_902,N_842);
xnor U1059 (N_1059,In_60,N_840);
nand U1060 (N_1060,N_710,N_910);
nand U1061 (N_1061,N_641,N_739);
xnor U1062 (N_1062,N_522,In_1046);
nor U1063 (N_1063,In_1493,N_281);
xnor U1064 (N_1064,N_184,N_899);
nand U1065 (N_1065,N_801,N_846);
xnor U1066 (N_1066,N_1003,In_1428);
or U1067 (N_1067,In_1172,N_971);
xnor U1068 (N_1068,N_610,N_783);
nor U1069 (N_1069,N_809,N_671);
and U1070 (N_1070,In_644,N_806);
and U1071 (N_1071,N_777,In_1459);
xnor U1072 (N_1072,N_886,N_194);
and U1073 (N_1073,N_837,N_741);
nor U1074 (N_1074,N_155,N_280);
and U1075 (N_1075,N_336,N_682);
or U1076 (N_1076,N_1044,In_29);
nand U1077 (N_1077,In_1149,N_912);
nand U1078 (N_1078,N_920,In_1233);
or U1079 (N_1079,N_538,In_408);
nor U1080 (N_1080,N_1022,In_536);
and U1081 (N_1081,N_803,N_932);
or U1082 (N_1082,N_60,N_835);
or U1083 (N_1083,N_948,N_983);
nand U1084 (N_1084,N_999,In_641);
nor U1085 (N_1085,In_1356,In_751);
nor U1086 (N_1086,N_1039,N_1032);
and U1087 (N_1087,In_580,N_813);
xor U1088 (N_1088,N_707,In_599);
xor U1089 (N_1089,N_892,N_1006);
nor U1090 (N_1090,N_244,N_365);
nand U1091 (N_1091,N_851,N_647);
or U1092 (N_1092,N_509,In_1344);
and U1093 (N_1093,N_1037,N_894);
nor U1094 (N_1094,N_964,N_1030);
or U1095 (N_1095,N_745,In_1300);
and U1096 (N_1096,N_1009,N_939);
or U1097 (N_1097,N_831,N_447);
nor U1098 (N_1098,N_872,In_904);
xnor U1099 (N_1099,N_940,In_618);
nand U1100 (N_1100,N_924,N_834);
nor U1101 (N_1101,N_560,N_501);
or U1102 (N_1102,N_960,N_850);
nand U1103 (N_1103,N_664,N_763);
and U1104 (N_1104,In_164,N_933);
nand U1105 (N_1105,N_946,N_938);
and U1106 (N_1106,N_922,In_875);
nor U1107 (N_1107,In_185,In_844);
nor U1108 (N_1108,In_1048,In_1008);
or U1109 (N_1109,N_506,N_576);
nor U1110 (N_1110,In_1070,In_113);
xnor U1111 (N_1111,N_921,N_856);
nor U1112 (N_1112,In_1076,N_965);
and U1113 (N_1113,In_1342,N_557);
nor U1114 (N_1114,N_847,N_845);
or U1115 (N_1115,N_970,N_1016);
nor U1116 (N_1116,N_755,N_966);
and U1117 (N_1117,N_495,N_799);
nor U1118 (N_1118,N_819,N_637);
nor U1119 (N_1119,N_930,N_1031);
or U1120 (N_1120,N_1021,N_639);
nor U1121 (N_1121,N_959,N_978);
or U1122 (N_1122,N_870,N_297);
or U1123 (N_1123,In_1409,N_634);
and U1124 (N_1124,In_1494,N_821);
nand U1125 (N_1125,N_980,N_779);
nand U1126 (N_1126,N_1035,In_147);
xor U1127 (N_1127,N_936,N_793);
or U1128 (N_1128,N_1026,N_308);
and U1129 (N_1129,N_668,N_903);
xnor U1130 (N_1130,N_684,N_1025);
nand U1131 (N_1131,N_982,N_473);
nor U1132 (N_1132,N_195,N_911);
nor U1133 (N_1133,N_974,N_941);
and U1134 (N_1134,N_405,N_680);
and U1135 (N_1135,N_947,N_665);
xnor U1136 (N_1136,In_936,N_949);
nand U1137 (N_1137,N_778,In_1144);
nor U1138 (N_1138,N_956,N_905);
or U1139 (N_1139,N_909,N_879);
xnor U1140 (N_1140,N_908,N_1043);
and U1141 (N_1141,N_164,N_616);
nand U1142 (N_1142,In_739,N_897);
or U1143 (N_1143,In_355,N_881);
and U1144 (N_1144,N_904,N_1024);
nand U1145 (N_1145,In_1387,In_1189);
and U1146 (N_1146,N_758,N_514);
nor U1147 (N_1147,N_935,N_989);
and U1148 (N_1148,N_566,In_767);
nand U1149 (N_1149,N_1046,N_918);
and U1150 (N_1150,N_917,N_901);
nor U1151 (N_1151,N_1019,N_957);
and U1152 (N_1152,N_653,N_934);
nand U1153 (N_1153,N_1010,N_765);
or U1154 (N_1154,In_1051,N_838);
nand U1155 (N_1155,N_1004,N_542);
or U1156 (N_1156,N_907,N_812);
or U1157 (N_1157,N_469,N_868);
and U1158 (N_1158,N_77,N_843);
nor U1159 (N_1159,N_511,In_1246);
or U1160 (N_1160,In_999,N_796);
or U1161 (N_1161,N_1023,N_703);
xnor U1162 (N_1162,In_749,N_1045);
or U1163 (N_1163,N_996,N_670);
xor U1164 (N_1164,N_995,N_811);
or U1165 (N_1165,N_494,N_384);
xnor U1166 (N_1166,In_906,N_1028);
xor U1167 (N_1167,N_1015,N_37);
xnor U1168 (N_1168,In_506,In_741);
nand U1169 (N_1169,N_984,N_138);
or U1170 (N_1170,N_225,N_950);
or U1171 (N_1171,N_1002,In_1283);
xor U1172 (N_1172,N_690,In_376);
nand U1173 (N_1173,N_900,N_235);
nor U1174 (N_1174,N_620,N_937);
nor U1175 (N_1175,N_945,N_497);
nor U1176 (N_1176,N_929,N_569);
nor U1177 (N_1177,N_836,N_853);
xor U1178 (N_1178,In_1328,N_1001);
xor U1179 (N_1179,N_954,N_54);
nand U1180 (N_1180,In_170,N_1008);
nor U1181 (N_1181,N_767,N_455);
nand U1182 (N_1182,N_188,N_1042);
nand U1183 (N_1183,In_1110,N_981);
or U1184 (N_1184,N_312,In_1436);
nand U1185 (N_1185,N_828,In_606);
nand U1186 (N_1186,N_928,N_353);
nand U1187 (N_1187,N_874,N_979);
nor U1188 (N_1188,N_953,N_394);
xnor U1189 (N_1189,N_985,N_961);
nor U1190 (N_1190,N_889,N_968);
xor U1191 (N_1191,In_698,N_993);
or U1192 (N_1192,In_124,N_798);
nor U1193 (N_1193,N_967,In_575);
xnor U1194 (N_1194,N_660,N_867);
or U1195 (N_1195,N_973,In_70);
nor U1196 (N_1196,N_1048,N_489);
and U1197 (N_1197,N_626,N_449);
or U1198 (N_1198,N_805,N_969);
or U1199 (N_1199,N_776,N_1005);
or U1200 (N_1200,N_1135,N_1117);
or U1201 (N_1201,N_882,In_1315);
and U1202 (N_1202,N_1171,N_1081);
or U1203 (N_1203,N_1186,N_992);
and U1204 (N_1204,N_1086,N_1192);
xnor U1205 (N_1205,N_1151,N_1071);
xor U1206 (N_1206,N_1125,N_1091);
or U1207 (N_1207,N_797,N_1085);
nand U1208 (N_1208,N_759,N_1185);
xor U1209 (N_1209,N_987,N_346);
nor U1210 (N_1210,N_1146,N_820);
nor U1211 (N_1211,N_1166,N_862);
and U1212 (N_1212,N_1112,N_1079);
or U1213 (N_1213,N_233,N_1173);
xor U1214 (N_1214,N_663,N_1142);
nand U1215 (N_1215,N_1182,In_608);
nand U1216 (N_1216,N_1111,N_1140);
nand U1217 (N_1217,In_1319,N_1180);
nand U1218 (N_1218,N_1056,N_1124);
and U1219 (N_1219,N_963,In_28);
nand U1220 (N_1220,N_1155,N_890);
or U1221 (N_1221,N_1114,N_1077);
xnor U1222 (N_1222,N_976,N_1109);
nor U1223 (N_1223,N_1167,N_448);
nor U1224 (N_1224,N_231,N_785);
nor U1225 (N_1225,N_1160,N_1165);
or U1226 (N_1226,N_1138,N_1104);
or U1227 (N_1227,N_1041,N_1148);
or U1228 (N_1228,In_911,N_228);
or U1229 (N_1229,N_735,In_42);
and U1230 (N_1230,N_1064,N_1070);
and U1231 (N_1231,In_1418,In_792);
and U1232 (N_1232,N_1115,N_733);
nor U1233 (N_1233,N_1059,N_1123);
and U1234 (N_1234,N_1051,N_552);
or U1235 (N_1235,N_1198,N_1100);
and U1236 (N_1236,N_927,N_1054);
or U1237 (N_1237,N_1020,N_1179);
and U1238 (N_1238,N_1122,N_1127);
and U1239 (N_1239,N_1121,N_1184);
or U1240 (N_1240,N_1027,N_611);
nand U1241 (N_1241,N_1000,N_1191);
and U1242 (N_1242,N_1156,N_1052);
or U1243 (N_1243,In_609,N_1069);
nor U1244 (N_1244,N_657,N_977);
xor U1245 (N_1245,N_1144,N_1065);
nand U1246 (N_1246,In_1487,N_1092);
nor U1247 (N_1247,N_760,N_1133);
or U1248 (N_1248,In_1250,N_1164);
or U1249 (N_1249,N_0,N_883);
nor U1250 (N_1250,In_217,N_962);
xnor U1251 (N_1251,N_753,N_1126);
nor U1252 (N_1252,N_1087,N_1088);
nand U1253 (N_1253,N_1187,N_1096);
nor U1254 (N_1254,In_298,N_931);
xor U1255 (N_1255,N_997,In_796);
and U1256 (N_1256,N_1047,N_656);
xor U1257 (N_1257,N_1060,N_994);
nand U1258 (N_1258,N_1113,N_1074);
and U1259 (N_1259,N_1188,N_385);
nand U1260 (N_1260,N_991,N_595);
xor U1261 (N_1261,N_943,N_1141);
nand U1262 (N_1262,N_775,In_592);
nor U1263 (N_1263,N_157,In_597);
nor U1264 (N_1264,N_1195,N_1145);
nor U1265 (N_1265,N_1116,N_880);
nor U1266 (N_1266,N_1034,N_916);
xnor U1267 (N_1267,N_1147,N_877);
and U1268 (N_1268,N_718,N_1062);
or U1269 (N_1269,In_492,N_1194);
or U1270 (N_1270,N_1018,N_729);
and U1271 (N_1271,N_815,N_1033);
or U1272 (N_1272,N_1101,N_1098);
nor U1273 (N_1273,N_1189,N_688);
and U1274 (N_1274,N_1097,N_1072);
xnor U1275 (N_1275,N_82,In_954);
nor U1276 (N_1276,N_1139,N_1061);
nand U1277 (N_1277,N_1108,N_1163);
or U1278 (N_1278,In_114,N_1093);
or U1279 (N_1279,N_848,N_972);
nor U1280 (N_1280,In_1379,In_842);
xnor U1281 (N_1281,N_914,N_1157);
nor U1282 (N_1282,N_808,N_687);
nand U1283 (N_1283,N_1110,N_1149);
and U1284 (N_1284,In_808,N_919);
or U1285 (N_1285,In_632,N_1129);
and U1286 (N_1286,N_1153,N_1181);
xnor U1287 (N_1287,N_1036,N_833);
or U1288 (N_1288,N_717,N_1178);
and U1289 (N_1289,N_295,N_1068);
nor U1290 (N_1290,N_926,N_1103);
and U1291 (N_1291,N_1134,N_1067);
or U1292 (N_1292,N_769,N_454);
xor U1293 (N_1293,N_1076,In_1419);
nor U1294 (N_1294,N_1128,N_1075);
or U1295 (N_1295,N_1174,N_604);
nand U1296 (N_1296,N_1199,N_344);
nor U1297 (N_1297,N_1050,In_1281);
nand U1298 (N_1298,N_414,N_1130);
nor U1299 (N_1299,N_925,In_852);
nor U1300 (N_1300,N_1082,N_1177);
nor U1301 (N_1301,In_648,In_915);
nor U1302 (N_1302,N_1162,N_1172);
nand U1303 (N_1303,N_1106,N_1066);
nor U1304 (N_1304,N_1038,N_958);
or U1305 (N_1305,N_1159,N_1058);
nand U1306 (N_1306,N_1095,N_724);
xnor U1307 (N_1307,N_1143,N_789);
nand U1308 (N_1308,N_773,N_1169);
and U1309 (N_1309,N_1132,N_1136);
xor U1310 (N_1310,N_1055,N_906);
or U1311 (N_1311,N_1154,N_645);
nor U1312 (N_1312,N_1131,In_726);
and U1313 (N_1313,N_150,In_229);
and U1314 (N_1314,N_1099,N_1161);
or U1315 (N_1315,N_1083,N_132);
or U1316 (N_1316,N_1190,N_951);
nand U1317 (N_1317,N_444,N_1089);
nand U1318 (N_1318,N_1080,N_1120);
xor U1319 (N_1319,N_1073,N_1152);
nand U1320 (N_1320,N_1057,N_579);
xnor U1321 (N_1321,N_1040,N_1102);
or U1322 (N_1322,N_1078,N_1049);
nand U1323 (N_1323,N_1183,N_944);
and U1324 (N_1324,In_566,N_104);
or U1325 (N_1325,N_531,In_1152);
and U1326 (N_1326,N_2,N_873);
nor U1327 (N_1327,N_1150,N_1014);
xor U1328 (N_1328,N_750,N_800);
nand U1329 (N_1329,N_770,N_841);
or U1330 (N_1330,N_1193,N_1090);
nor U1331 (N_1331,N_1029,N_998);
or U1332 (N_1332,N_1053,N_1119);
and U1333 (N_1333,N_791,N_1137);
nor U1334 (N_1334,N_1175,N_1012);
or U1335 (N_1335,N_1094,In_281);
nor U1336 (N_1336,In_1020,N_1011);
xnor U1337 (N_1337,N_990,N_986);
xnor U1338 (N_1338,N_571,In_228);
nor U1339 (N_1339,N_1176,N_942);
or U1340 (N_1340,N_1063,N_1158);
xor U1341 (N_1341,N_952,N_1168);
or U1342 (N_1342,N_975,N_1105);
or U1343 (N_1343,N_761,N_1017);
or U1344 (N_1344,N_1118,N_1197);
nand U1345 (N_1345,N_1196,N_482);
nor U1346 (N_1346,In_38,N_598);
and U1347 (N_1347,N_1107,N_1007);
xor U1348 (N_1348,N_487,N_1084);
nor U1349 (N_1349,N_1170,N_1013);
nor U1350 (N_1350,N_1340,N_1254);
and U1351 (N_1351,N_1307,N_1313);
and U1352 (N_1352,N_1237,N_1322);
xnor U1353 (N_1353,N_1293,N_1258);
xor U1354 (N_1354,N_1251,N_1305);
and U1355 (N_1355,N_1252,N_1270);
xor U1356 (N_1356,N_1288,N_1223);
or U1357 (N_1357,N_1284,N_1343);
nor U1358 (N_1358,N_1285,N_1204);
nand U1359 (N_1359,N_1331,N_1294);
and U1360 (N_1360,N_1300,N_1325);
and U1361 (N_1361,N_1346,N_1334);
xor U1362 (N_1362,N_1231,N_1221);
nor U1363 (N_1363,N_1224,N_1215);
and U1364 (N_1364,N_1276,N_1347);
nand U1365 (N_1365,N_1228,N_1281);
xor U1366 (N_1366,N_1292,N_1262);
and U1367 (N_1367,N_1314,N_1326);
xor U1368 (N_1368,N_1213,N_1210);
or U1369 (N_1369,N_1220,N_1286);
nor U1370 (N_1370,N_1219,N_1304);
or U1371 (N_1371,N_1238,N_1225);
or U1372 (N_1372,N_1207,N_1266);
nand U1373 (N_1373,N_1310,N_1247);
xnor U1374 (N_1374,N_1250,N_1202);
nand U1375 (N_1375,N_1261,N_1277);
and U1376 (N_1376,N_1200,N_1249);
nand U1377 (N_1377,N_1203,N_1315);
xor U1378 (N_1378,N_1243,N_1302);
xnor U1379 (N_1379,N_1218,N_1268);
xor U1380 (N_1380,N_1248,N_1312);
or U1381 (N_1381,N_1338,N_1235);
nor U1382 (N_1382,N_1308,N_1341);
and U1383 (N_1383,N_1299,N_1280);
or U1384 (N_1384,N_1208,N_1269);
xnor U1385 (N_1385,N_1232,N_1241);
xnor U1386 (N_1386,N_1318,N_1216);
nor U1387 (N_1387,N_1255,N_1327);
or U1388 (N_1388,N_1244,N_1283);
or U1389 (N_1389,N_1201,N_1265);
and U1390 (N_1390,N_1306,N_1212);
or U1391 (N_1391,N_1298,N_1301);
and U1392 (N_1392,N_1287,N_1316);
nand U1393 (N_1393,N_1339,N_1209);
nor U1394 (N_1394,N_1336,N_1332);
xor U1395 (N_1395,N_1321,N_1227);
or U1396 (N_1396,N_1329,N_1289);
and U1397 (N_1397,N_1328,N_1337);
or U1398 (N_1398,N_1240,N_1279);
nand U1399 (N_1399,N_1282,N_1273);
nand U1400 (N_1400,N_1317,N_1217);
or U1401 (N_1401,N_1236,N_1330);
or U1402 (N_1402,N_1349,N_1275);
nand U1403 (N_1403,N_1271,N_1263);
and U1404 (N_1404,N_1206,N_1256);
xor U1405 (N_1405,N_1259,N_1260);
nand U1406 (N_1406,N_1272,N_1296);
xor U1407 (N_1407,N_1233,N_1274);
or U1408 (N_1408,N_1345,N_1246);
and U1409 (N_1409,N_1226,N_1319);
xnor U1410 (N_1410,N_1264,N_1229);
xor U1411 (N_1411,N_1278,N_1245);
nor U1412 (N_1412,N_1344,N_1335);
or U1413 (N_1413,N_1348,N_1214);
nor U1414 (N_1414,N_1297,N_1230);
and U1415 (N_1415,N_1291,N_1211);
and U1416 (N_1416,N_1333,N_1239);
nand U1417 (N_1417,N_1234,N_1267);
nor U1418 (N_1418,N_1303,N_1320);
nand U1419 (N_1419,N_1205,N_1222);
or U1420 (N_1420,N_1311,N_1342);
or U1421 (N_1421,N_1290,N_1323);
and U1422 (N_1422,N_1253,N_1324);
and U1423 (N_1423,N_1257,N_1242);
and U1424 (N_1424,N_1309,N_1295);
or U1425 (N_1425,N_1303,N_1214);
or U1426 (N_1426,N_1331,N_1240);
nand U1427 (N_1427,N_1325,N_1218);
and U1428 (N_1428,N_1226,N_1254);
xnor U1429 (N_1429,N_1250,N_1204);
nand U1430 (N_1430,N_1214,N_1347);
and U1431 (N_1431,N_1212,N_1329);
or U1432 (N_1432,N_1210,N_1307);
xnor U1433 (N_1433,N_1332,N_1208);
nor U1434 (N_1434,N_1291,N_1329);
and U1435 (N_1435,N_1298,N_1346);
xor U1436 (N_1436,N_1347,N_1282);
nand U1437 (N_1437,N_1281,N_1233);
and U1438 (N_1438,N_1302,N_1285);
nor U1439 (N_1439,N_1266,N_1303);
xor U1440 (N_1440,N_1282,N_1287);
and U1441 (N_1441,N_1267,N_1342);
nor U1442 (N_1442,N_1223,N_1330);
and U1443 (N_1443,N_1314,N_1282);
nand U1444 (N_1444,N_1322,N_1256);
nor U1445 (N_1445,N_1300,N_1210);
nor U1446 (N_1446,N_1200,N_1283);
nand U1447 (N_1447,N_1276,N_1290);
xnor U1448 (N_1448,N_1231,N_1233);
nand U1449 (N_1449,N_1261,N_1248);
nand U1450 (N_1450,N_1268,N_1243);
and U1451 (N_1451,N_1325,N_1312);
nand U1452 (N_1452,N_1291,N_1203);
xnor U1453 (N_1453,N_1232,N_1220);
nand U1454 (N_1454,N_1202,N_1303);
nand U1455 (N_1455,N_1209,N_1303);
or U1456 (N_1456,N_1328,N_1287);
and U1457 (N_1457,N_1293,N_1345);
nand U1458 (N_1458,N_1208,N_1279);
xor U1459 (N_1459,N_1257,N_1203);
nand U1460 (N_1460,N_1241,N_1211);
xnor U1461 (N_1461,N_1239,N_1250);
xor U1462 (N_1462,N_1289,N_1211);
xnor U1463 (N_1463,N_1292,N_1349);
nor U1464 (N_1464,N_1294,N_1202);
nand U1465 (N_1465,N_1247,N_1255);
xnor U1466 (N_1466,N_1330,N_1217);
xnor U1467 (N_1467,N_1202,N_1230);
and U1468 (N_1468,N_1323,N_1320);
nand U1469 (N_1469,N_1275,N_1309);
xor U1470 (N_1470,N_1262,N_1313);
xnor U1471 (N_1471,N_1289,N_1214);
nor U1472 (N_1472,N_1212,N_1266);
or U1473 (N_1473,N_1329,N_1230);
nor U1474 (N_1474,N_1225,N_1236);
and U1475 (N_1475,N_1348,N_1326);
xor U1476 (N_1476,N_1300,N_1219);
nand U1477 (N_1477,N_1286,N_1273);
xnor U1478 (N_1478,N_1242,N_1245);
and U1479 (N_1479,N_1206,N_1301);
nand U1480 (N_1480,N_1270,N_1260);
xnor U1481 (N_1481,N_1297,N_1272);
or U1482 (N_1482,N_1255,N_1331);
and U1483 (N_1483,N_1210,N_1257);
xnor U1484 (N_1484,N_1239,N_1349);
xor U1485 (N_1485,N_1251,N_1285);
and U1486 (N_1486,N_1228,N_1225);
xnor U1487 (N_1487,N_1271,N_1276);
or U1488 (N_1488,N_1315,N_1284);
or U1489 (N_1489,N_1273,N_1292);
nor U1490 (N_1490,N_1243,N_1301);
nor U1491 (N_1491,N_1211,N_1262);
nand U1492 (N_1492,N_1225,N_1254);
nand U1493 (N_1493,N_1274,N_1286);
and U1494 (N_1494,N_1299,N_1262);
nor U1495 (N_1495,N_1319,N_1294);
or U1496 (N_1496,N_1246,N_1262);
nor U1497 (N_1497,N_1275,N_1310);
nor U1498 (N_1498,N_1220,N_1208);
xnor U1499 (N_1499,N_1298,N_1320);
xor U1500 (N_1500,N_1382,N_1362);
nor U1501 (N_1501,N_1494,N_1496);
or U1502 (N_1502,N_1453,N_1482);
nand U1503 (N_1503,N_1465,N_1407);
and U1504 (N_1504,N_1446,N_1434);
nand U1505 (N_1505,N_1397,N_1406);
nand U1506 (N_1506,N_1416,N_1438);
xor U1507 (N_1507,N_1352,N_1387);
xnor U1508 (N_1508,N_1363,N_1464);
nand U1509 (N_1509,N_1450,N_1492);
nand U1510 (N_1510,N_1399,N_1460);
or U1511 (N_1511,N_1415,N_1481);
nor U1512 (N_1512,N_1400,N_1371);
xnor U1513 (N_1513,N_1489,N_1471);
and U1514 (N_1514,N_1467,N_1451);
and U1515 (N_1515,N_1404,N_1497);
or U1516 (N_1516,N_1487,N_1355);
or U1517 (N_1517,N_1479,N_1385);
nand U1518 (N_1518,N_1475,N_1380);
xor U1519 (N_1519,N_1490,N_1364);
and U1520 (N_1520,N_1486,N_1377);
nor U1521 (N_1521,N_1441,N_1393);
and U1522 (N_1522,N_1356,N_1498);
or U1523 (N_1523,N_1493,N_1459);
nor U1524 (N_1524,N_1436,N_1414);
nor U1525 (N_1525,N_1366,N_1373);
or U1526 (N_1526,N_1369,N_1430);
and U1527 (N_1527,N_1367,N_1383);
nor U1528 (N_1528,N_1432,N_1395);
nand U1529 (N_1529,N_1403,N_1483);
or U1530 (N_1530,N_1427,N_1463);
nand U1531 (N_1531,N_1480,N_1444);
nor U1532 (N_1532,N_1412,N_1445);
or U1533 (N_1533,N_1431,N_1388);
or U1534 (N_1534,N_1474,N_1370);
xnor U1535 (N_1535,N_1386,N_1372);
nor U1536 (N_1536,N_1457,N_1358);
or U1537 (N_1537,N_1449,N_1476);
nor U1538 (N_1538,N_1433,N_1376);
or U1539 (N_1539,N_1409,N_1439);
or U1540 (N_1540,N_1477,N_1423);
xor U1541 (N_1541,N_1421,N_1405);
nor U1542 (N_1542,N_1428,N_1417);
xnor U1543 (N_1543,N_1359,N_1375);
xnor U1544 (N_1544,N_1411,N_1485);
xor U1545 (N_1545,N_1473,N_1442);
nand U1546 (N_1546,N_1499,N_1437);
or U1547 (N_1547,N_1461,N_1422);
and U1548 (N_1548,N_1484,N_1455);
xnor U1549 (N_1549,N_1396,N_1491);
nor U1550 (N_1550,N_1454,N_1470);
or U1551 (N_1551,N_1389,N_1447);
or U1552 (N_1552,N_1435,N_1448);
nor U1553 (N_1553,N_1360,N_1468);
and U1554 (N_1554,N_1425,N_1354);
or U1555 (N_1555,N_1478,N_1424);
xnor U1556 (N_1556,N_1401,N_1353);
and U1557 (N_1557,N_1452,N_1419);
or U1558 (N_1558,N_1378,N_1374);
nand U1559 (N_1559,N_1410,N_1420);
nor U1560 (N_1560,N_1413,N_1429);
nor U1561 (N_1561,N_1381,N_1394);
xor U1562 (N_1562,N_1462,N_1443);
nor U1563 (N_1563,N_1469,N_1495);
or U1564 (N_1564,N_1384,N_1458);
nand U1565 (N_1565,N_1357,N_1392);
xnor U1566 (N_1566,N_1402,N_1472);
nand U1567 (N_1567,N_1390,N_1398);
xor U1568 (N_1568,N_1365,N_1408);
xor U1569 (N_1569,N_1361,N_1426);
or U1570 (N_1570,N_1379,N_1456);
or U1571 (N_1571,N_1488,N_1351);
nand U1572 (N_1572,N_1418,N_1466);
or U1573 (N_1573,N_1391,N_1440);
nor U1574 (N_1574,N_1350,N_1368);
and U1575 (N_1575,N_1404,N_1388);
and U1576 (N_1576,N_1496,N_1378);
and U1577 (N_1577,N_1386,N_1403);
and U1578 (N_1578,N_1374,N_1411);
nand U1579 (N_1579,N_1353,N_1467);
nor U1580 (N_1580,N_1412,N_1405);
and U1581 (N_1581,N_1498,N_1477);
nand U1582 (N_1582,N_1400,N_1490);
and U1583 (N_1583,N_1426,N_1459);
nor U1584 (N_1584,N_1499,N_1482);
xor U1585 (N_1585,N_1487,N_1489);
or U1586 (N_1586,N_1461,N_1363);
xor U1587 (N_1587,N_1357,N_1411);
and U1588 (N_1588,N_1489,N_1438);
and U1589 (N_1589,N_1420,N_1475);
nor U1590 (N_1590,N_1395,N_1463);
nand U1591 (N_1591,N_1352,N_1467);
or U1592 (N_1592,N_1442,N_1432);
xor U1593 (N_1593,N_1403,N_1378);
nand U1594 (N_1594,N_1470,N_1411);
xor U1595 (N_1595,N_1463,N_1384);
and U1596 (N_1596,N_1403,N_1407);
nand U1597 (N_1597,N_1386,N_1384);
and U1598 (N_1598,N_1487,N_1433);
and U1599 (N_1599,N_1411,N_1462);
xnor U1600 (N_1600,N_1460,N_1443);
or U1601 (N_1601,N_1451,N_1382);
or U1602 (N_1602,N_1424,N_1487);
nor U1603 (N_1603,N_1477,N_1428);
nor U1604 (N_1604,N_1450,N_1374);
and U1605 (N_1605,N_1358,N_1437);
nand U1606 (N_1606,N_1474,N_1390);
and U1607 (N_1607,N_1436,N_1482);
nor U1608 (N_1608,N_1365,N_1392);
nand U1609 (N_1609,N_1446,N_1380);
nor U1610 (N_1610,N_1407,N_1470);
or U1611 (N_1611,N_1359,N_1354);
or U1612 (N_1612,N_1363,N_1408);
and U1613 (N_1613,N_1411,N_1435);
and U1614 (N_1614,N_1440,N_1379);
xor U1615 (N_1615,N_1418,N_1358);
xnor U1616 (N_1616,N_1378,N_1445);
nand U1617 (N_1617,N_1457,N_1424);
nand U1618 (N_1618,N_1371,N_1465);
and U1619 (N_1619,N_1366,N_1426);
xnor U1620 (N_1620,N_1366,N_1441);
nand U1621 (N_1621,N_1382,N_1459);
or U1622 (N_1622,N_1447,N_1485);
nor U1623 (N_1623,N_1400,N_1406);
nand U1624 (N_1624,N_1498,N_1388);
or U1625 (N_1625,N_1350,N_1492);
nor U1626 (N_1626,N_1430,N_1444);
xnor U1627 (N_1627,N_1451,N_1367);
nand U1628 (N_1628,N_1450,N_1421);
nor U1629 (N_1629,N_1409,N_1443);
nand U1630 (N_1630,N_1367,N_1493);
and U1631 (N_1631,N_1489,N_1407);
or U1632 (N_1632,N_1492,N_1461);
xnor U1633 (N_1633,N_1413,N_1439);
xnor U1634 (N_1634,N_1376,N_1429);
nand U1635 (N_1635,N_1490,N_1495);
xor U1636 (N_1636,N_1372,N_1473);
and U1637 (N_1637,N_1455,N_1490);
or U1638 (N_1638,N_1442,N_1380);
or U1639 (N_1639,N_1380,N_1467);
and U1640 (N_1640,N_1461,N_1471);
and U1641 (N_1641,N_1414,N_1474);
xnor U1642 (N_1642,N_1477,N_1476);
and U1643 (N_1643,N_1431,N_1437);
xnor U1644 (N_1644,N_1429,N_1436);
or U1645 (N_1645,N_1378,N_1432);
nor U1646 (N_1646,N_1426,N_1454);
nor U1647 (N_1647,N_1414,N_1368);
nor U1648 (N_1648,N_1423,N_1427);
and U1649 (N_1649,N_1407,N_1474);
xor U1650 (N_1650,N_1507,N_1623);
or U1651 (N_1651,N_1520,N_1625);
and U1652 (N_1652,N_1552,N_1615);
nand U1653 (N_1653,N_1647,N_1621);
nand U1654 (N_1654,N_1540,N_1572);
nand U1655 (N_1655,N_1579,N_1606);
nand U1656 (N_1656,N_1521,N_1557);
xor U1657 (N_1657,N_1523,N_1586);
or U1658 (N_1658,N_1614,N_1644);
or U1659 (N_1659,N_1519,N_1533);
and U1660 (N_1660,N_1584,N_1575);
xnor U1661 (N_1661,N_1600,N_1541);
xor U1662 (N_1662,N_1649,N_1610);
nor U1663 (N_1663,N_1555,N_1568);
or U1664 (N_1664,N_1554,N_1510);
nand U1665 (N_1665,N_1642,N_1609);
and U1666 (N_1666,N_1622,N_1641);
or U1667 (N_1667,N_1602,N_1538);
xnor U1668 (N_1668,N_1593,N_1603);
nor U1669 (N_1669,N_1578,N_1545);
xor U1670 (N_1670,N_1503,N_1558);
or U1671 (N_1671,N_1619,N_1516);
nor U1672 (N_1672,N_1639,N_1501);
nor U1673 (N_1673,N_1601,N_1630);
or U1674 (N_1674,N_1645,N_1574);
xor U1675 (N_1675,N_1515,N_1536);
xor U1676 (N_1676,N_1635,N_1620);
and U1677 (N_1677,N_1522,N_1542);
nand U1678 (N_1678,N_1599,N_1583);
nand U1679 (N_1679,N_1532,N_1548);
xnor U1680 (N_1680,N_1513,N_1627);
and U1681 (N_1681,N_1518,N_1544);
nand U1682 (N_1682,N_1556,N_1570);
nand U1683 (N_1683,N_1514,N_1592);
xor U1684 (N_1684,N_1616,N_1626);
nor U1685 (N_1685,N_1581,N_1508);
nand U1686 (N_1686,N_1631,N_1607);
nor U1687 (N_1687,N_1543,N_1524);
or U1688 (N_1688,N_1563,N_1577);
xnor U1689 (N_1689,N_1505,N_1559);
and U1690 (N_1690,N_1638,N_1608);
and U1691 (N_1691,N_1596,N_1560);
nor U1692 (N_1692,N_1643,N_1640);
and U1693 (N_1693,N_1509,N_1605);
nor U1694 (N_1694,N_1594,N_1589);
nor U1695 (N_1695,N_1613,N_1636);
xnor U1696 (N_1696,N_1550,N_1502);
and U1697 (N_1697,N_1504,N_1565);
nor U1698 (N_1698,N_1646,N_1597);
or U1699 (N_1699,N_1534,N_1537);
and U1700 (N_1700,N_1648,N_1585);
or U1701 (N_1701,N_1618,N_1611);
and U1702 (N_1702,N_1569,N_1629);
and U1703 (N_1703,N_1562,N_1531);
and U1704 (N_1704,N_1528,N_1500);
xnor U1705 (N_1705,N_1595,N_1590);
xnor U1706 (N_1706,N_1549,N_1527);
nor U1707 (N_1707,N_1612,N_1529);
and U1708 (N_1708,N_1547,N_1580);
xnor U1709 (N_1709,N_1564,N_1566);
nor U1710 (N_1710,N_1546,N_1591);
nor U1711 (N_1711,N_1588,N_1637);
xnor U1712 (N_1712,N_1624,N_1604);
xor U1713 (N_1713,N_1573,N_1617);
xor U1714 (N_1714,N_1535,N_1567);
xnor U1715 (N_1715,N_1632,N_1525);
and U1716 (N_1716,N_1526,N_1511);
xnor U1717 (N_1717,N_1587,N_1634);
nor U1718 (N_1718,N_1561,N_1517);
nand U1719 (N_1719,N_1553,N_1598);
xnor U1720 (N_1720,N_1530,N_1576);
nand U1721 (N_1721,N_1633,N_1539);
nand U1722 (N_1722,N_1512,N_1582);
or U1723 (N_1723,N_1506,N_1551);
nand U1724 (N_1724,N_1571,N_1628);
xnor U1725 (N_1725,N_1531,N_1507);
nand U1726 (N_1726,N_1552,N_1643);
nor U1727 (N_1727,N_1528,N_1561);
nand U1728 (N_1728,N_1566,N_1582);
or U1729 (N_1729,N_1570,N_1511);
xnor U1730 (N_1730,N_1575,N_1607);
or U1731 (N_1731,N_1589,N_1631);
nor U1732 (N_1732,N_1614,N_1605);
xor U1733 (N_1733,N_1538,N_1617);
or U1734 (N_1734,N_1509,N_1517);
or U1735 (N_1735,N_1591,N_1612);
nor U1736 (N_1736,N_1594,N_1542);
nor U1737 (N_1737,N_1567,N_1542);
nor U1738 (N_1738,N_1548,N_1554);
or U1739 (N_1739,N_1596,N_1551);
or U1740 (N_1740,N_1519,N_1527);
nand U1741 (N_1741,N_1603,N_1591);
or U1742 (N_1742,N_1620,N_1567);
nand U1743 (N_1743,N_1545,N_1573);
nor U1744 (N_1744,N_1611,N_1645);
nand U1745 (N_1745,N_1559,N_1611);
or U1746 (N_1746,N_1603,N_1634);
or U1747 (N_1747,N_1561,N_1581);
nor U1748 (N_1748,N_1551,N_1609);
nand U1749 (N_1749,N_1567,N_1557);
or U1750 (N_1750,N_1544,N_1627);
nor U1751 (N_1751,N_1518,N_1638);
or U1752 (N_1752,N_1527,N_1505);
xor U1753 (N_1753,N_1598,N_1575);
nor U1754 (N_1754,N_1533,N_1617);
xor U1755 (N_1755,N_1522,N_1629);
nand U1756 (N_1756,N_1636,N_1624);
nor U1757 (N_1757,N_1622,N_1565);
nand U1758 (N_1758,N_1616,N_1596);
or U1759 (N_1759,N_1566,N_1559);
or U1760 (N_1760,N_1526,N_1552);
nor U1761 (N_1761,N_1613,N_1648);
and U1762 (N_1762,N_1530,N_1590);
nand U1763 (N_1763,N_1500,N_1516);
and U1764 (N_1764,N_1533,N_1590);
or U1765 (N_1765,N_1574,N_1540);
nand U1766 (N_1766,N_1563,N_1535);
nand U1767 (N_1767,N_1593,N_1646);
xnor U1768 (N_1768,N_1628,N_1502);
xor U1769 (N_1769,N_1553,N_1534);
xnor U1770 (N_1770,N_1571,N_1595);
and U1771 (N_1771,N_1611,N_1561);
xor U1772 (N_1772,N_1552,N_1645);
or U1773 (N_1773,N_1502,N_1510);
nand U1774 (N_1774,N_1598,N_1534);
nand U1775 (N_1775,N_1537,N_1572);
or U1776 (N_1776,N_1532,N_1646);
or U1777 (N_1777,N_1598,N_1529);
and U1778 (N_1778,N_1543,N_1640);
nand U1779 (N_1779,N_1639,N_1572);
and U1780 (N_1780,N_1539,N_1568);
xnor U1781 (N_1781,N_1600,N_1524);
nor U1782 (N_1782,N_1585,N_1511);
or U1783 (N_1783,N_1534,N_1563);
or U1784 (N_1784,N_1642,N_1615);
or U1785 (N_1785,N_1615,N_1532);
nor U1786 (N_1786,N_1562,N_1577);
or U1787 (N_1787,N_1613,N_1577);
nand U1788 (N_1788,N_1547,N_1558);
or U1789 (N_1789,N_1550,N_1514);
nor U1790 (N_1790,N_1502,N_1647);
or U1791 (N_1791,N_1634,N_1614);
xnor U1792 (N_1792,N_1615,N_1521);
xor U1793 (N_1793,N_1531,N_1630);
or U1794 (N_1794,N_1627,N_1525);
nor U1795 (N_1795,N_1538,N_1511);
and U1796 (N_1796,N_1513,N_1527);
and U1797 (N_1797,N_1644,N_1637);
and U1798 (N_1798,N_1617,N_1535);
xor U1799 (N_1799,N_1500,N_1581);
or U1800 (N_1800,N_1750,N_1699);
and U1801 (N_1801,N_1777,N_1779);
or U1802 (N_1802,N_1761,N_1690);
nor U1803 (N_1803,N_1653,N_1687);
and U1804 (N_1804,N_1788,N_1717);
nand U1805 (N_1805,N_1658,N_1725);
xor U1806 (N_1806,N_1766,N_1710);
and U1807 (N_1807,N_1714,N_1659);
and U1808 (N_1808,N_1774,N_1666);
or U1809 (N_1809,N_1764,N_1726);
and U1810 (N_1810,N_1753,N_1684);
xnor U1811 (N_1811,N_1702,N_1707);
and U1812 (N_1812,N_1731,N_1694);
xor U1813 (N_1813,N_1770,N_1723);
and U1814 (N_1814,N_1744,N_1675);
xor U1815 (N_1815,N_1718,N_1679);
xor U1816 (N_1816,N_1660,N_1654);
or U1817 (N_1817,N_1734,N_1746);
or U1818 (N_1818,N_1719,N_1754);
xnor U1819 (N_1819,N_1745,N_1672);
nor U1820 (N_1820,N_1790,N_1676);
xor U1821 (N_1821,N_1767,N_1737);
or U1822 (N_1822,N_1792,N_1677);
nand U1823 (N_1823,N_1681,N_1652);
or U1824 (N_1824,N_1655,N_1784);
nand U1825 (N_1825,N_1757,N_1693);
nor U1826 (N_1826,N_1711,N_1782);
or U1827 (N_1827,N_1682,N_1789);
and U1828 (N_1828,N_1667,N_1722);
xor U1829 (N_1829,N_1650,N_1793);
xor U1830 (N_1830,N_1748,N_1662);
and U1831 (N_1831,N_1794,N_1771);
nand U1832 (N_1832,N_1747,N_1712);
and U1833 (N_1833,N_1716,N_1729);
nor U1834 (N_1834,N_1760,N_1697);
or U1835 (N_1835,N_1698,N_1673);
nand U1836 (N_1836,N_1786,N_1688);
and U1837 (N_1837,N_1683,N_1778);
xor U1838 (N_1838,N_1674,N_1678);
nand U1839 (N_1839,N_1759,N_1663);
nand U1840 (N_1840,N_1765,N_1705);
and U1841 (N_1841,N_1724,N_1772);
xnor U1842 (N_1842,N_1689,N_1708);
nand U1843 (N_1843,N_1691,N_1735);
or U1844 (N_1844,N_1739,N_1670);
xor U1845 (N_1845,N_1721,N_1709);
nand U1846 (N_1846,N_1657,N_1661);
or U1847 (N_1847,N_1756,N_1651);
xor U1848 (N_1848,N_1799,N_1776);
nand U1849 (N_1849,N_1781,N_1785);
xor U1850 (N_1850,N_1783,N_1686);
nand U1851 (N_1851,N_1692,N_1743);
nand U1852 (N_1852,N_1740,N_1704);
nor U1853 (N_1853,N_1669,N_1796);
and U1854 (N_1854,N_1762,N_1780);
xnor U1855 (N_1855,N_1668,N_1749);
xor U1856 (N_1856,N_1727,N_1787);
or U1857 (N_1857,N_1755,N_1713);
xor U1858 (N_1858,N_1733,N_1732);
or U1859 (N_1859,N_1706,N_1696);
xnor U1860 (N_1860,N_1664,N_1752);
or U1861 (N_1861,N_1741,N_1720);
and U1862 (N_1862,N_1730,N_1685);
or U1863 (N_1863,N_1795,N_1695);
and U1864 (N_1864,N_1728,N_1700);
and U1865 (N_1865,N_1768,N_1798);
nor U1866 (N_1866,N_1736,N_1656);
nor U1867 (N_1867,N_1742,N_1797);
nand U1868 (N_1868,N_1758,N_1680);
xor U1869 (N_1869,N_1775,N_1715);
and U1870 (N_1870,N_1703,N_1671);
xnor U1871 (N_1871,N_1773,N_1763);
and U1872 (N_1872,N_1791,N_1769);
or U1873 (N_1873,N_1751,N_1738);
nand U1874 (N_1874,N_1701,N_1665);
and U1875 (N_1875,N_1667,N_1663);
and U1876 (N_1876,N_1655,N_1776);
or U1877 (N_1877,N_1740,N_1793);
and U1878 (N_1878,N_1701,N_1755);
and U1879 (N_1879,N_1660,N_1664);
nor U1880 (N_1880,N_1772,N_1661);
xor U1881 (N_1881,N_1705,N_1777);
and U1882 (N_1882,N_1714,N_1705);
nor U1883 (N_1883,N_1678,N_1733);
xnor U1884 (N_1884,N_1663,N_1733);
nand U1885 (N_1885,N_1768,N_1761);
nor U1886 (N_1886,N_1722,N_1760);
xor U1887 (N_1887,N_1724,N_1659);
nand U1888 (N_1888,N_1767,N_1687);
nor U1889 (N_1889,N_1770,N_1778);
nand U1890 (N_1890,N_1671,N_1731);
nor U1891 (N_1891,N_1711,N_1767);
and U1892 (N_1892,N_1655,N_1749);
xor U1893 (N_1893,N_1783,N_1662);
or U1894 (N_1894,N_1672,N_1711);
and U1895 (N_1895,N_1780,N_1670);
xnor U1896 (N_1896,N_1772,N_1748);
nor U1897 (N_1897,N_1700,N_1683);
or U1898 (N_1898,N_1727,N_1660);
nor U1899 (N_1899,N_1669,N_1772);
and U1900 (N_1900,N_1781,N_1757);
or U1901 (N_1901,N_1698,N_1701);
nand U1902 (N_1902,N_1794,N_1744);
or U1903 (N_1903,N_1736,N_1724);
nor U1904 (N_1904,N_1650,N_1698);
nand U1905 (N_1905,N_1762,N_1689);
or U1906 (N_1906,N_1782,N_1702);
nand U1907 (N_1907,N_1655,N_1723);
nand U1908 (N_1908,N_1734,N_1785);
nor U1909 (N_1909,N_1789,N_1659);
nand U1910 (N_1910,N_1691,N_1757);
xor U1911 (N_1911,N_1658,N_1796);
nand U1912 (N_1912,N_1743,N_1776);
xnor U1913 (N_1913,N_1750,N_1695);
nor U1914 (N_1914,N_1698,N_1737);
nor U1915 (N_1915,N_1769,N_1681);
nand U1916 (N_1916,N_1774,N_1665);
or U1917 (N_1917,N_1673,N_1760);
xnor U1918 (N_1918,N_1706,N_1794);
or U1919 (N_1919,N_1757,N_1793);
nor U1920 (N_1920,N_1797,N_1695);
nand U1921 (N_1921,N_1696,N_1652);
and U1922 (N_1922,N_1693,N_1682);
and U1923 (N_1923,N_1794,N_1738);
and U1924 (N_1924,N_1664,N_1670);
nand U1925 (N_1925,N_1757,N_1664);
xnor U1926 (N_1926,N_1736,N_1679);
xor U1927 (N_1927,N_1762,N_1766);
and U1928 (N_1928,N_1761,N_1665);
or U1929 (N_1929,N_1778,N_1695);
and U1930 (N_1930,N_1675,N_1692);
nand U1931 (N_1931,N_1693,N_1707);
nor U1932 (N_1932,N_1732,N_1765);
and U1933 (N_1933,N_1706,N_1683);
or U1934 (N_1934,N_1745,N_1655);
nand U1935 (N_1935,N_1681,N_1717);
xnor U1936 (N_1936,N_1738,N_1688);
or U1937 (N_1937,N_1664,N_1792);
nor U1938 (N_1938,N_1661,N_1673);
or U1939 (N_1939,N_1799,N_1777);
and U1940 (N_1940,N_1728,N_1705);
and U1941 (N_1941,N_1791,N_1669);
or U1942 (N_1942,N_1667,N_1686);
xnor U1943 (N_1943,N_1716,N_1690);
xor U1944 (N_1944,N_1747,N_1674);
nor U1945 (N_1945,N_1728,N_1673);
or U1946 (N_1946,N_1701,N_1783);
nor U1947 (N_1947,N_1729,N_1747);
or U1948 (N_1948,N_1790,N_1788);
nor U1949 (N_1949,N_1740,N_1738);
nand U1950 (N_1950,N_1853,N_1890);
nor U1951 (N_1951,N_1816,N_1857);
and U1952 (N_1952,N_1948,N_1834);
xnor U1953 (N_1953,N_1880,N_1810);
nor U1954 (N_1954,N_1870,N_1926);
nor U1955 (N_1955,N_1862,N_1815);
and U1956 (N_1956,N_1932,N_1920);
or U1957 (N_1957,N_1827,N_1824);
nand U1958 (N_1958,N_1947,N_1944);
or U1959 (N_1959,N_1930,N_1937);
and U1960 (N_1960,N_1836,N_1900);
xor U1961 (N_1961,N_1917,N_1883);
and U1962 (N_1962,N_1822,N_1925);
and U1963 (N_1963,N_1929,N_1909);
xor U1964 (N_1964,N_1907,N_1935);
nand U1965 (N_1965,N_1820,N_1833);
and U1966 (N_1966,N_1840,N_1844);
nor U1967 (N_1967,N_1855,N_1941);
and U1968 (N_1968,N_1848,N_1913);
or U1969 (N_1969,N_1901,N_1832);
and U1970 (N_1970,N_1878,N_1921);
or U1971 (N_1971,N_1928,N_1940);
xor U1972 (N_1972,N_1851,N_1875);
and U1973 (N_1973,N_1897,N_1846);
or U1974 (N_1974,N_1854,N_1885);
nand U1975 (N_1975,N_1889,N_1893);
and U1976 (N_1976,N_1879,N_1830);
nor U1977 (N_1977,N_1887,N_1821);
xnor U1978 (N_1978,N_1871,N_1835);
and U1979 (N_1979,N_1868,N_1945);
nand U1980 (N_1980,N_1805,N_1807);
xnor U1981 (N_1981,N_1906,N_1946);
nor U1982 (N_1982,N_1873,N_1852);
nand U1983 (N_1983,N_1892,N_1899);
or U1984 (N_1984,N_1841,N_1902);
nor U1985 (N_1985,N_1933,N_1813);
xor U1986 (N_1986,N_1860,N_1812);
nand U1987 (N_1987,N_1886,N_1837);
nand U1988 (N_1988,N_1914,N_1845);
or U1989 (N_1989,N_1898,N_1814);
nand U1990 (N_1990,N_1839,N_1884);
or U1991 (N_1991,N_1842,N_1936);
and U1992 (N_1992,N_1924,N_1918);
and U1993 (N_1993,N_1874,N_1904);
or U1994 (N_1994,N_1934,N_1804);
and U1995 (N_1995,N_1865,N_1801);
nor U1996 (N_1996,N_1927,N_1903);
xor U1997 (N_1997,N_1912,N_1919);
xnor U1998 (N_1998,N_1877,N_1911);
and U1999 (N_1999,N_1803,N_1872);
nor U2000 (N_2000,N_1847,N_1876);
xor U2001 (N_2001,N_1866,N_1838);
and U2002 (N_2002,N_1881,N_1861);
and U2003 (N_2003,N_1811,N_1819);
or U2004 (N_2004,N_1905,N_1888);
nor U2005 (N_2005,N_1843,N_1910);
xor U2006 (N_2006,N_1923,N_1850);
nor U2007 (N_2007,N_1915,N_1939);
or U2008 (N_2008,N_1931,N_1825);
nand U2009 (N_2009,N_1943,N_1891);
and U2010 (N_2010,N_1922,N_1858);
and U2011 (N_2011,N_1949,N_1869);
nor U2012 (N_2012,N_1800,N_1863);
nand U2013 (N_2013,N_1882,N_1818);
or U2014 (N_2014,N_1859,N_1896);
xnor U2015 (N_2015,N_1806,N_1867);
nor U2016 (N_2016,N_1826,N_1829);
nor U2017 (N_2017,N_1849,N_1864);
nand U2018 (N_2018,N_1908,N_1894);
and U2019 (N_2019,N_1938,N_1802);
and U2020 (N_2020,N_1808,N_1895);
nor U2021 (N_2021,N_1828,N_1942);
nand U2022 (N_2022,N_1823,N_1856);
and U2023 (N_2023,N_1831,N_1817);
nor U2024 (N_2024,N_1809,N_1916);
and U2025 (N_2025,N_1825,N_1892);
nor U2026 (N_2026,N_1928,N_1882);
nand U2027 (N_2027,N_1835,N_1810);
and U2028 (N_2028,N_1898,N_1879);
xnor U2029 (N_2029,N_1847,N_1947);
or U2030 (N_2030,N_1831,N_1858);
nand U2031 (N_2031,N_1897,N_1913);
xnor U2032 (N_2032,N_1869,N_1918);
xor U2033 (N_2033,N_1870,N_1860);
xnor U2034 (N_2034,N_1806,N_1826);
and U2035 (N_2035,N_1908,N_1862);
xnor U2036 (N_2036,N_1807,N_1818);
xor U2037 (N_2037,N_1818,N_1933);
or U2038 (N_2038,N_1870,N_1884);
nor U2039 (N_2039,N_1933,N_1896);
and U2040 (N_2040,N_1866,N_1904);
nand U2041 (N_2041,N_1929,N_1890);
nand U2042 (N_2042,N_1836,N_1819);
xor U2043 (N_2043,N_1943,N_1933);
nor U2044 (N_2044,N_1911,N_1891);
and U2045 (N_2045,N_1882,N_1844);
nor U2046 (N_2046,N_1884,N_1804);
nand U2047 (N_2047,N_1896,N_1865);
or U2048 (N_2048,N_1901,N_1862);
or U2049 (N_2049,N_1829,N_1843);
nand U2050 (N_2050,N_1935,N_1905);
and U2051 (N_2051,N_1939,N_1937);
nand U2052 (N_2052,N_1821,N_1851);
and U2053 (N_2053,N_1907,N_1903);
and U2054 (N_2054,N_1949,N_1914);
and U2055 (N_2055,N_1861,N_1918);
nand U2056 (N_2056,N_1946,N_1826);
or U2057 (N_2057,N_1871,N_1891);
nand U2058 (N_2058,N_1893,N_1880);
nand U2059 (N_2059,N_1840,N_1936);
or U2060 (N_2060,N_1891,N_1821);
xor U2061 (N_2061,N_1848,N_1843);
nand U2062 (N_2062,N_1875,N_1862);
or U2063 (N_2063,N_1808,N_1911);
and U2064 (N_2064,N_1938,N_1867);
xnor U2065 (N_2065,N_1946,N_1932);
and U2066 (N_2066,N_1944,N_1817);
or U2067 (N_2067,N_1829,N_1840);
nand U2068 (N_2068,N_1921,N_1902);
and U2069 (N_2069,N_1904,N_1895);
or U2070 (N_2070,N_1903,N_1825);
nor U2071 (N_2071,N_1888,N_1879);
nor U2072 (N_2072,N_1939,N_1930);
nor U2073 (N_2073,N_1883,N_1895);
nand U2074 (N_2074,N_1868,N_1879);
and U2075 (N_2075,N_1900,N_1819);
and U2076 (N_2076,N_1847,N_1815);
or U2077 (N_2077,N_1812,N_1811);
nand U2078 (N_2078,N_1879,N_1931);
or U2079 (N_2079,N_1850,N_1916);
and U2080 (N_2080,N_1811,N_1806);
nand U2081 (N_2081,N_1924,N_1863);
nor U2082 (N_2082,N_1940,N_1888);
xor U2083 (N_2083,N_1815,N_1849);
xnor U2084 (N_2084,N_1944,N_1886);
nand U2085 (N_2085,N_1908,N_1835);
xnor U2086 (N_2086,N_1861,N_1886);
xnor U2087 (N_2087,N_1945,N_1835);
and U2088 (N_2088,N_1848,N_1849);
or U2089 (N_2089,N_1856,N_1884);
xor U2090 (N_2090,N_1921,N_1867);
and U2091 (N_2091,N_1847,N_1878);
xnor U2092 (N_2092,N_1874,N_1928);
and U2093 (N_2093,N_1801,N_1896);
nand U2094 (N_2094,N_1910,N_1875);
nand U2095 (N_2095,N_1891,N_1886);
xor U2096 (N_2096,N_1888,N_1891);
nand U2097 (N_2097,N_1920,N_1847);
nand U2098 (N_2098,N_1945,N_1905);
or U2099 (N_2099,N_1820,N_1889);
nor U2100 (N_2100,N_2015,N_2073);
xor U2101 (N_2101,N_2006,N_2010);
nand U2102 (N_2102,N_2025,N_2081);
or U2103 (N_2103,N_2092,N_2083);
nor U2104 (N_2104,N_2000,N_2078);
nand U2105 (N_2105,N_2020,N_1979);
xnor U2106 (N_2106,N_2035,N_1997);
xor U2107 (N_2107,N_1950,N_1985);
xor U2108 (N_2108,N_2008,N_1959);
nor U2109 (N_2109,N_1972,N_2028);
and U2110 (N_2110,N_2065,N_2087);
or U2111 (N_2111,N_2039,N_2053);
or U2112 (N_2112,N_2096,N_1967);
xor U2113 (N_2113,N_2002,N_1983);
or U2114 (N_2114,N_2062,N_1951);
nor U2115 (N_2115,N_2068,N_1984);
and U2116 (N_2116,N_1999,N_2012);
nor U2117 (N_2117,N_2057,N_2085);
xnor U2118 (N_2118,N_1953,N_2097);
nand U2119 (N_2119,N_1955,N_2038);
or U2120 (N_2120,N_1978,N_1971);
nor U2121 (N_2121,N_1995,N_2029);
and U2122 (N_2122,N_1977,N_2009);
nand U2123 (N_2123,N_2059,N_1980);
xor U2124 (N_2124,N_2089,N_2060);
or U2125 (N_2125,N_2032,N_1988);
nor U2126 (N_2126,N_2041,N_2023);
or U2127 (N_2127,N_2033,N_2050);
nand U2128 (N_2128,N_2088,N_2095);
nand U2129 (N_2129,N_1989,N_2086);
and U2130 (N_2130,N_2036,N_2007);
nand U2131 (N_2131,N_2055,N_2013);
and U2132 (N_2132,N_2063,N_2045);
and U2133 (N_2133,N_2044,N_2070);
nand U2134 (N_2134,N_2051,N_1961);
or U2135 (N_2135,N_2071,N_2034);
or U2136 (N_2136,N_2042,N_1954);
or U2137 (N_2137,N_1975,N_2075);
and U2138 (N_2138,N_1976,N_1969);
nor U2139 (N_2139,N_1996,N_2003);
and U2140 (N_2140,N_2001,N_2084);
or U2141 (N_2141,N_1966,N_1965);
nand U2142 (N_2142,N_2047,N_2019);
xnor U2143 (N_2143,N_1963,N_2080);
xor U2144 (N_2144,N_1991,N_1992);
xnor U2145 (N_2145,N_2018,N_2016);
or U2146 (N_2146,N_2077,N_2021);
nand U2147 (N_2147,N_2082,N_2011);
xor U2148 (N_2148,N_2076,N_2026);
nor U2149 (N_2149,N_1960,N_2030);
nor U2150 (N_2150,N_2052,N_2005);
nor U2151 (N_2151,N_1956,N_2064);
xor U2152 (N_2152,N_1974,N_2093);
nor U2153 (N_2153,N_2056,N_2024);
xor U2154 (N_2154,N_2054,N_2058);
xor U2155 (N_2155,N_2067,N_2072);
nor U2156 (N_2156,N_2091,N_2048);
nand U2157 (N_2157,N_2066,N_1981);
nor U2158 (N_2158,N_2043,N_2061);
and U2159 (N_2159,N_2040,N_1964);
and U2160 (N_2160,N_1962,N_2098);
or U2161 (N_2161,N_2090,N_2004);
xor U2162 (N_2162,N_2046,N_2014);
nand U2163 (N_2163,N_2099,N_2094);
and U2164 (N_2164,N_1994,N_2027);
or U2165 (N_2165,N_1958,N_2037);
xnor U2166 (N_2166,N_2031,N_1987);
nor U2167 (N_2167,N_1957,N_2079);
xor U2168 (N_2168,N_2049,N_1982);
or U2169 (N_2169,N_2022,N_1973);
and U2170 (N_2170,N_1986,N_1990);
nand U2171 (N_2171,N_1970,N_2074);
xnor U2172 (N_2172,N_2017,N_2069);
nand U2173 (N_2173,N_1998,N_1952);
and U2174 (N_2174,N_1993,N_1968);
or U2175 (N_2175,N_2052,N_2012);
xnor U2176 (N_2176,N_2032,N_2077);
or U2177 (N_2177,N_2024,N_2093);
and U2178 (N_2178,N_2097,N_2030);
or U2179 (N_2179,N_1970,N_2029);
nand U2180 (N_2180,N_2093,N_2027);
nand U2181 (N_2181,N_1977,N_2001);
or U2182 (N_2182,N_2002,N_2000);
or U2183 (N_2183,N_2073,N_1961);
xnor U2184 (N_2184,N_2033,N_2097);
nor U2185 (N_2185,N_2038,N_2093);
or U2186 (N_2186,N_1997,N_2017);
nor U2187 (N_2187,N_2010,N_2042);
nand U2188 (N_2188,N_2030,N_2074);
xnor U2189 (N_2189,N_1987,N_1960);
nor U2190 (N_2190,N_1997,N_1965);
xor U2191 (N_2191,N_2022,N_2036);
nor U2192 (N_2192,N_1972,N_2053);
or U2193 (N_2193,N_2035,N_2047);
or U2194 (N_2194,N_2050,N_2085);
nor U2195 (N_2195,N_1975,N_1995);
nor U2196 (N_2196,N_2066,N_2096);
nand U2197 (N_2197,N_2039,N_2001);
nand U2198 (N_2198,N_2085,N_2014);
or U2199 (N_2199,N_1968,N_1958);
xnor U2200 (N_2200,N_1963,N_2051);
nor U2201 (N_2201,N_2071,N_2008);
nand U2202 (N_2202,N_2016,N_2042);
and U2203 (N_2203,N_2065,N_2053);
nand U2204 (N_2204,N_1997,N_2065);
xnor U2205 (N_2205,N_2025,N_2072);
and U2206 (N_2206,N_2073,N_2084);
or U2207 (N_2207,N_1996,N_1985);
and U2208 (N_2208,N_2022,N_2032);
or U2209 (N_2209,N_1992,N_1988);
nor U2210 (N_2210,N_1950,N_1966);
nor U2211 (N_2211,N_1993,N_2014);
nand U2212 (N_2212,N_2035,N_2057);
xor U2213 (N_2213,N_1958,N_1992);
xnor U2214 (N_2214,N_2043,N_2013);
xnor U2215 (N_2215,N_2057,N_2082);
nand U2216 (N_2216,N_1976,N_1950);
nand U2217 (N_2217,N_2076,N_2029);
nor U2218 (N_2218,N_2084,N_2091);
nand U2219 (N_2219,N_2010,N_2018);
nor U2220 (N_2220,N_2030,N_2059);
nor U2221 (N_2221,N_2047,N_2007);
nor U2222 (N_2222,N_2091,N_2075);
and U2223 (N_2223,N_2017,N_2066);
or U2224 (N_2224,N_2086,N_1969);
nand U2225 (N_2225,N_2026,N_2019);
and U2226 (N_2226,N_2057,N_1973);
xnor U2227 (N_2227,N_2082,N_1965);
xnor U2228 (N_2228,N_1985,N_2097);
or U2229 (N_2229,N_1979,N_1975);
and U2230 (N_2230,N_2089,N_2046);
or U2231 (N_2231,N_2077,N_2011);
nor U2232 (N_2232,N_2013,N_2078);
nor U2233 (N_2233,N_2005,N_2054);
or U2234 (N_2234,N_2046,N_2011);
and U2235 (N_2235,N_2095,N_2055);
and U2236 (N_2236,N_2004,N_2011);
and U2237 (N_2237,N_2009,N_2081);
nand U2238 (N_2238,N_1950,N_2037);
xnor U2239 (N_2239,N_2013,N_2095);
or U2240 (N_2240,N_2091,N_1998);
nand U2241 (N_2241,N_1964,N_2058);
nor U2242 (N_2242,N_1996,N_2017);
or U2243 (N_2243,N_1980,N_2009);
xnor U2244 (N_2244,N_1961,N_1968);
nor U2245 (N_2245,N_1967,N_2027);
nor U2246 (N_2246,N_2026,N_1963);
nand U2247 (N_2247,N_2010,N_2038);
xnor U2248 (N_2248,N_2027,N_1966);
nand U2249 (N_2249,N_1982,N_1996);
or U2250 (N_2250,N_2143,N_2102);
and U2251 (N_2251,N_2182,N_2214);
nor U2252 (N_2252,N_2124,N_2222);
or U2253 (N_2253,N_2239,N_2204);
nand U2254 (N_2254,N_2186,N_2174);
nor U2255 (N_2255,N_2135,N_2201);
and U2256 (N_2256,N_2205,N_2152);
and U2257 (N_2257,N_2199,N_2147);
nand U2258 (N_2258,N_2206,N_2232);
and U2259 (N_2259,N_2118,N_2101);
nor U2260 (N_2260,N_2168,N_2244);
nand U2261 (N_2261,N_2234,N_2129);
xor U2262 (N_2262,N_2200,N_2188);
nand U2263 (N_2263,N_2228,N_2242);
nand U2264 (N_2264,N_2149,N_2105);
xnor U2265 (N_2265,N_2133,N_2218);
or U2266 (N_2266,N_2187,N_2181);
or U2267 (N_2267,N_2245,N_2126);
xnor U2268 (N_2268,N_2190,N_2219);
and U2269 (N_2269,N_2236,N_2213);
nand U2270 (N_2270,N_2194,N_2158);
and U2271 (N_2271,N_2111,N_2211);
nand U2272 (N_2272,N_2137,N_2166);
and U2273 (N_2273,N_2109,N_2120);
nand U2274 (N_2274,N_2249,N_2134);
and U2275 (N_2275,N_2198,N_2170);
nor U2276 (N_2276,N_2171,N_2238);
xnor U2277 (N_2277,N_2131,N_2221);
and U2278 (N_2278,N_2121,N_2172);
and U2279 (N_2279,N_2145,N_2140);
or U2280 (N_2280,N_2155,N_2193);
nor U2281 (N_2281,N_2130,N_2144);
xor U2282 (N_2282,N_2136,N_2164);
or U2283 (N_2283,N_2165,N_2233);
xor U2284 (N_2284,N_2248,N_2151);
or U2285 (N_2285,N_2196,N_2108);
nand U2286 (N_2286,N_2104,N_2119);
or U2287 (N_2287,N_2107,N_2113);
or U2288 (N_2288,N_2192,N_2180);
nor U2289 (N_2289,N_2128,N_2235);
or U2290 (N_2290,N_2202,N_2173);
nor U2291 (N_2291,N_2197,N_2243);
and U2292 (N_2292,N_2210,N_2115);
and U2293 (N_2293,N_2241,N_2220);
nand U2294 (N_2294,N_2162,N_2106);
and U2295 (N_2295,N_2231,N_2150);
and U2296 (N_2296,N_2195,N_2125);
nor U2297 (N_2297,N_2161,N_2215);
xnor U2298 (N_2298,N_2229,N_2157);
nor U2299 (N_2299,N_2189,N_2226);
nor U2300 (N_2300,N_2225,N_2114);
nor U2301 (N_2301,N_2240,N_2224);
xor U2302 (N_2302,N_2223,N_2127);
nor U2303 (N_2303,N_2217,N_2167);
nor U2304 (N_2304,N_2156,N_2141);
nor U2305 (N_2305,N_2179,N_2246);
nand U2306 (N_2306,N_2176,N_2146);
and U2307 (N_2307,N_2191,N_2183);
nor U2308 (N_2308,N_2100,N_2153);
and U2309 (N_2309,N_2154,N_2178);
and U2310 (N_2310,N_2142,N_2184);
xnor U2311 (N_2311,N_2110,N_2123);
and U2312 (N_2312,N_2230,N_2103);
and U2313 (N_2313,N_2132,N_2138);
and U2314 (N_2314,N_2209,N_2175);
xnor U2315 (N_2315,N_2116,N_2169);
xnor U2316 (N_2316,N_2203,N_2160);
nand U2317 (N_2317,N_2117,N_2227);
xnor U2318 (N_2318,N_2159,N_2148);
and U2319 (N_2319,N_2208,N_2185);
nor U2320 (N_2320,N_2212,N_2139);
or U2321 (N_2321,N_2177,N_2163);
xor U2322 (N_2322,N_2207,N_2247);
nand U2323 (N_2323,N_2112,N_2237);
and U2324 (N_2324,N_2216,N_2122);
and U2325 (N_2325,N_2148,N_2203);
and U2326 (N_2326,N_2235,N_2111);
nand U2327 (N_2327,N_2124,N_2171);
nand U2328 (N_2328,N_2216,N_2133);
or U2329 (N_2329,N_2137,N_2233);
and U2330 (N_2330,N_2243,N_2224);
or U2331 (N_2331,N_2166,N_2131);
or U2332 (N_2332,N_2173,N_2130);
or U2333 (N_2333,N_2177,N_2157);
nand U2334 (N_2334,N_2226,N_2149);
nor U2335 (N_2335,N_2109,N_2191);
or U2336 (N_2336,N_2203,N_2195);
nand U2337 (N_2337,N_2121,N_2138);
nor U2338 (N_2338,N_2116,N_2142);
xor U2339 (N_2339,N_2249,N_2209);
xor U2340 (N_2340,N_2142,N_2171);
nand U2341 (N_2341,N_2150,N_2138);
nor U2342 (N_2342,N_2135,N_2114);
or U2343 (N_2343,N_2105,N_2156);
xnor U2344 (N_2344,N_2120,N_2196);
nor U2345 (N_2345,N_2156,N_2158);
xnor U2346 (N_2346,N_2196,N_2123);
or U2347 (N_2347,N_2108,N_2163);
xnor U2348 (N_2348,N_2117,N_2103);
and U2349 (N_2349,N_2188,N_2242);
and U2350 (N_2350,N_2213,N_2247);
xnor U2351 (N_2351,N_2188,N_2124);
nand U2352 (N_2352,N_2155,N_2148);
xor U2353 (N_2353,N_2127,N_2241);
and U2354 (N_2354,N_2188,N_2233);
nor U2355 (N_2355,N_2207,N_2229);
and U2356 (N_2356,N_2222,N_2176);
nand U2357 (N_2357,N_2173,N_2234);
or U2358 (N_2358,N_2104,N_2165);
nor U2359 (N_2359,N_2115,N_2172);
or U2360 (N_2360,N_2120,N_2241);
nor U2361 (N_2361,N_2134,N_2175);
or U2362 (N_2362,N_2204,N_2197);
xnor U2363 (N_2363,N_2149,N_2240);
xor U2364 (N_2364,N_2147,N_2103);
and U2365 (N_2365,N_2174,N_2133);
xor U2366 (N_2366,N_2223,N_2143);
nor U2367 (N_2367,N_2147,N_2108);
xnor U2368 (N_2368,N_2174,N_2200);
xnor U2369 (N_2369,N_2134,N_2246);
nand U2370 (N_2370,N_2224,N_2119);
xnor U2371 (N_2371,N_2191,N_2142);
xor U2372 (N_2372,N_2225,N_2132);
nand U2373 (N_2373,N_2133,N_2195);
xor U2374 (N_2374,N_2118,N_2125);
xor U2375 (N_2375,N_2237,N_2119);
xnor U2376 (N_2376,N_2118,N_2131);
nand U2377 (N_2377,N_2143,N_2165);
nor U2378 (N_2378,N_2152,N_2145);
nand U2379 (N_2379,N_2173,N_2183);
nand U2380 (N_2380,N_2224,N_2128);
and U2381 (N_2381,N_2182,N_2211);
nor U2382 (N_2382,N_2223,N_2179);
and U2383 (N_2383,N_2117,N_2191);
and U2384 (N_2384,N_2149,N_2215);
nand U2385 (N_2385,N_2213,N_2142);
xnor U2386 (N_2386,N_2198,N_2241);
xnor U2387 (N_2387,N_2225,N_2150);
nand U2388 (N_2388,N_2103,N_2237);
and U2389 (N_2389,N_2202,N_2203);
xnor U2390 (N_2390,N_2188,N_2199);
xor U2391 (N_2391,N_2199,N_2154);
or U2392 (N_2392,N_2235,N_2209);
xnor U2393 (N_2393,N_2238,N_2203);
nor U2394 (N_2394,N_2181,N_2231);
or U2395 (N_2395,N_2239,N_2162);
nand U2396 (N_2396,N_2156,N_2192);
nand U2397 (N_2397,N_2122,N_2244);
or U2398 (N_2398,N_2246,N_2170);
xnor U2399 (N_2399,N_2110,N_2196);
or U2400 (N_2400,N_2390,N_2304);
or U2401 (N_2401,N_2334,N_2250);
nor U2402 (N_2402,N_2279,N_2309);
or U2403 (N_2403,N_2264,N_2362);
and U2404 (N_2404,N_2267,N_2252);
nand U2405 (N_2405,N_2271,N_2317);
nor U2406 (N_2406,N_2367,N_2262);
nor U2407 (N_2407,N_2310,N_2280);
xnor U2408 (N_2408,N_2260,N_2360);
nand U2409 (N_2409,N_2303,N_2361);
nor U2410 (N_2410,N_2290,N_2278);
nor U2411 (N_2411,N_2393,N_2327);
nand U2412 (N_2412,N_2286,N_2266);
nor U2413 (N_2413,N_2268,N_2296);
and U2414 (N_2414,N_2275,N_2381);
nand U2415 (N_2415,N_2373,N_2337);
or U2416 (N_2416,N_2340,N_2265);
and U2417 (N_2417,N_2282,N_2394);
xor U2418 (N_2418,N_2272,N_2354);
and U2419 (N_2419,N_2289,N_2295);
nor U2420 (N_2420,N_2395,N_2342);
or U2421 (N_2421,N_2294,N_2325);
nor U2422 (N_2422,N_2357,N_2297);
and U2423 (N_2423,N_2256,N_2356);
and U2424 (N_2424,N_2391,N_2348);
or U2425 (N_2425,N_2322,N_2253);
xnor U2426 (N_2426,N_2321,N_2331);
nor U2427 (N_2427,N_2378,N_2397);
nor U2428 (N_2428,N_2336,N_2349);
or U2429 (N_2429,N_2270,N_2314);
or U2430 (N_2430,N_2254,N_2351);
nor U2431 (N_2431,N_2287,N_2399);
nand U2432 (N_2432,N_2383,N_2338);
xor U2433 (N_2433,N_2341,N_2323);
nand U2434 (N_2434,N_2277,N_2259);
xnor U2435 (N_2435,N_2311,N_2333);
or U2436 (N_2436,N_2330,N_2358);
nor U2437 (N_2437,N_2308,N_2380);
nor U2438 (N_2438,N_2344,N_2258);
nand U2439 (N_2439,N_2305,N_2350);
and U2440 (N_2440,N_2285,N_2276);
xnor U2441 (N_2441,N_2298,N_2257);
xnor U2442 (N_2442,N_2332,N_2307);
and U2443 (N_2443,N_2335,N_2251);
nor U2444 (N_2444,N_2386,N_2316);
nor U2445 (N_2445,N_2369,N_2320);
or U2446 (N_2446,N_2384,N_2387);
and U2447 (N_2447,N_2346,N_2388);
or U2448 (N_2448,N_2375,N_2283);
or U2449 (N_2449,N_2299,N_2364);
xor U2450 (N_2450,N_2263,N_2255);
nor U2451 (N_2451,N_2365,N_2398);
and U2452 (N_2452,N_2345,N_2302);
and U2453 (N_2453,N_2352,N_2372);
nand U2454 (N_2454,N_2261,N_2371);
nand U2455 (N_2455,N_2291,N_2392);
and U2456 (N_2456,N_2319,N_2269);
nor U2457 (N_2457,N_2293,N_2281);
nor U2458 (N_2458,N_2273,N_2315);
xor U2459 (N_2459,N_2347,N_2382);
or U2460 (N_2460,N_2306,N_2292);
xnor U2461 (N_2461,N_2363,N_2284);
and U2462 (N_2462,N_2374,N_2368);
nor U2463 (N_2463,N_2313,N_2329);
nor U2464 (N_2464,N_2326,N_2377);
xnor U2465 (N_2465,N_2376,N_2312);
nand U2466 (N_2466,N_2389,N_2396);
or U2467 (N_2467,N_2385,N_2353);
xnor U2468 (N_2468,N_2318,N_2355);
or U2469 (N_2469,N_2301,N_2370);
nand U2470 (N_2470,N_2324,N_2366);
nand U2471 (N_2471,N_2343,N_2339);
nor U2472 (N_2472,N_2288,N_2379);
nor U2473 (N_2473,N_2300,N_2328);
nand U2474 (N_2474,N_2274,N_2359);
xnor U2475 (N_2475,N_2346,N_2338);
xor U2476 (N_2476,N_2275,N_2319);
nand U2477 (N_2477,N_2277,N_2294);
xor U2478 (N_2478,N_2293,N_2317);
or U2479 (N_2479,N_2297,N_2312);
nor U2480 (N_2480,N_2291,N_2332);
xnor U2481 (N_2481,N_2331,N_2305);
xor U2482 (N_2482,N_2354,N_2274);
and U2483 (N_2483,N_2303,N_2280);
and U2484 (N_2484,N_2347,N_2308);
xnor U2485 (N_2485,N_2332,N_2357);
xnor U2486 (N_2486,N_2314,N_2344);
xnor U2487 (N_2487,N_2343,N_2277);
xor U2488 (N_2488,N_2268,N_2398);
xnor U2489 (N_2489,N_2253,N_2372);
nand U2490 (N_2490,N_2276,N_2256);
and U2491 (N_2491,N_2377,N_2373);
or U2492 (N_2492,N_2299,N_2311);
and U2493 (N_2493,N_2355,N_2384);
or U2494 (N_2494,N_2392,N_2398);
or U2495 (N_2495,N_2350,N_2292);
and U2496 (N_2496,N_2364,N_2334);
and U2497 (N_2497,N_2321,N_2357);
or U2498 (N_2498,N_2304,N_2383);
or U2499 (N_2499,N_2299,N_2334);
and U2500 (N_2500,N_2314,N_2267);
xor U2501 (N_2501,N_2340,N_2319);
nand U2502 (N_2502,N_2394,N_2324);
nand U2503 (N_2503,N_2376,N_2386);
nand U2504 (N_2504,N_2301,N_2369);
nor U2505 (N_2505,N_2321,N_2308);
nor U2506 (N_2506,N_2331,N_2368);
nor U2507 (N_2507,N_2328,N_2310);
nand U2508 (N_2508,N_2349,N_2271);
nand U2509 (N_2509,N_2356,N_2347);
nor U2510 (N_2510,N_2316,N_2288);
or U2511 (N_2511,N_2376,N_2369);
nand U2512 (N_2512,N_2376,N_2274);
and U2513 (N_2513,N_2390,N_2316);
and U2514 (N_2514,N_2320,N_2313);
nand U2515 (N_2515,N_2332,N_2382);
or U2516 (N_2516,N_2281,N_2384);
nor U2517 (N_2517,N_2352,N_2391);
nor U2518 (N_2518,N_2281,N_2347);
and U2519 (N_2519,N_2320,N_2311);
xor U2520 (N_2520,N_2333,N_2390);
or U2521 (N_2521,N_2370,N_2260);
nand U2522 (N_2522,N_2386,N_2300);
or U2523 (N_2523,N_2290,N_2266);
xor U2524 (N_2524,N_2356,N_2325);
xnor U2525 (N_2525,N_2273,N_2369);
and U2526 (N_2526,N_2256,N_2384);
and U2527 (N_2527,N_2295,N_2291);
and U2528 (N_2528,N_2337,N_2301);
or U2529 (N_2529,N_2299,N_2362);
xor U2530 (N_2530,N_2356,N_2273);
nor U2531 (N_2531,N_2386,N_2352);
nand U2532 (N_2532,N_2328,N_2277);
nor U2533 (N_2533,N_2287,N_2298);
or U2534 (N_2534,N_2332,N_2282);
and U2535 (N_2535,N_2266,N_2399);
and U2536 (N_2536,N_2254,N_2305);
xnor U2537 (N_2537,N_2360,N_2297);
and U2538 (N_2538,N_2380,N_2315);
or U2539 (N_2539,N_2336,N_2255);
xor U2540 (N_2540,N_2284,N_2397);
nor U2541 (N_2541,N_2364,N_2323);
nand U2542 (N_2542,N_2306,N_2371);
and U2543 (N_2543,N_2394,N_2267);
nor U2544 (N_2544,N_2375,N_2398);
nor U2545 (N_2545,N_2288,N_2259);
xor U2546 (N_2546,N_2342,N_2344);
nor U2547 (N_2547,N_2366,N_2287);
or U2548 (N_2548,N_2352,N_2382);
and U2549 (N_2549,N_2361,N_2257);
nor U2550 (N_2550,N_2434,N_2546);
nor U2551 (N_2551,N_2411,N_2444);
nand U2552 (N_2552,N_2548,N_2495);
and U2553 (N_2553,N_2538,N_2506);
nand U2554 (N_2554,N_2504,N_2440);
and U2555 (N_2555,N_2472,N_2484);
or U2556 (N_2556,N_2507,N_2425);
xnor U2557 (N_2557,N_2417,N_2456);
or U2558 (N_2558,N_2403,N_2547);
nand U2559 (N_2559,N_2458,N_2463);
xor U2560 (N_2560,N_2493,N_2497);
nor U2561 (N_2561,N_2470,N_2525);
and U2562 (N_2562,N_2457,N_2537);
or U2563 (N_2563,N_2449,N_2503);
xor U2564 (N_2564,N_2433,N_2439);
nand U2565 (N_2565,N_2467,N_2448);
nor U2566 (N_2566,N_2476,N_2531);
and U2567 (N_2567,N_2475,N_2438);
xnor U2568 (N_2568,N_2435,N_2533);
and U2569 (N_2569,N_2481,N_2514);
and U2570 (N_2570,N_2446,N_2541);
xor U2571 (N_2571,N_2494,N_2492);
or U2572 (N_2572,N_2509,N_2469);
xnor U2573 (N_2573,N_2518,N_2498);
nor U2574 (N_2574,N_2523,N_2487);
and U2575 (N_2575,N_2404,N_2445);
nand U2576 (N_2576,N_2510,N_2473);
nor U2577 (N_2577,N_2406,N_2480);
xnor U2578 (N_2578,N_2521,N_2464);
xor U2579 (N_2579,N_2419,N_2505);
xnor U2580 (N_2580,N_2465,N_2474);
and U2581 (N_2581,N_2401,N_2413);
or U2582 (N_2582,N_2522,N_2530);
xor U2583 (N_2583,N_2544,N_2549);
nand U2584 (N_2584,N_2526,N_2532);
and U2585 (N_2585,N_2441,N_2415);
or U2586 (N_2586,N_2428,N_2426);
or U2587 (N_2587,N_2519,N_2462);
nand U2588 (N_2588,N_2491,N_2418);
nand U2589 (N_2589,N_2460,N_2432);
xor U2590 (N_2590,N_2517,N_2408);
and U2591 (N_2591,N_2468,N_2452);
xnor U2592 (N_2592,N_2430,N_2500);
and U2593 (N_2593,N_2423,N_2486);
nand U2594 (N_2594,N_2443,N_2429);
xor U2595 (N_2595,N_2454,N_2499);
nand U2596 (N_2596,N_2453,N_2516);
nand U2597 (N_2597,N_2402,N_2529);
or U2598 (N_2598,N_2539,N_2501);
nor U2599 (N_2599,N_2407,N_2515);
nand U2600 (N_2600,N_2485,N_2540);
nor U2601 (N_2601,N_2461,N_2412);
and U2602 (N_2602,N_2508,N_2524);
nand U2603 (N_2603,N_2450,N_2421);
and U2604 (N_2604,N_2534,N_2488);
xor U2605 (N_2605,N_2427,N_2442);
nand U2606 (N_2606,N_2490,N_2471);
or U2607 (N_2607,N_2542,N_2400);
xnor U2608 (N_2608,N_2528,N_2422);
and U2609 (N_2609,N_2527,N_2424);
nand U2610 (N_2610,N_2502,N_2479);
nand U2611 (N_2611,N_2511,N_2477);
nor U2612 (N_2612,N_2405,N_2520);
or U2613 (N_2613,N_2483,N_2447);
nand U2614 (N_2614,N_2414,N_2416);
and U2615 (N_2615,N_2512,N_2478);
xor U2616 (N_2616,N_2437,N_2536);
nor U2617 (N_2617,N_2513,N_2496);
nand U2618 (N_2618,N_2489,N_2535);
nand U2619 (N_2619,N_2409,N_2466);
nand U2620 (N_2620,N_2455,N_2459);
and U2621 (N_2621,N_2543,N_2420);
or U2622 (N_2622,N_2410,N_2451);
nand U2623 (N_2623,N_2431,N_2545);
xor U2624 (N_2624,N_2482,N_2436);
and U2625 (N_2625,N_2439,N_2477);
xor U2626 (N_2626,N_2458,N_2533);
or U2627 (N_2627,N_2517,N_2511);
xnor U2628 (N_2628,N_2416,N_2546);
nor U2629 (N_2629,N_2514,N_2509);
xor U2630 (N_2630,N_2421,N_2500);
nand U2631 (N_2631,N_2415,N_2522);
nand U2632 (N_2632,N_2494,N_2425);
and U2633 (N_2633,N_2447,N_2466);
nand U2634 (N_2634,N_2498,N_2546);
nor U2635 (N_2635,N_2501,N_2426);
or U2636 (N_2636,N_2535,N_2430);
and U2637 (N_2637,N_2512,N_2483);
nor U2638 (N_2638,N_2542,N_2500);
or U2639 (N_2639,N_2400,N_2519);
and U2640 (N_2640,N_2483,N_2418);
nand U2641 (N_2641,N_2528,N_2461);
and U2642 (N_2642,N_2517,N_2528);
and U2643 (N_2643,N_2530,N_2508);
xor U2644 (N_2644,N_2490,N_2462);
or U2645 (N_2645,N_2443,N_2455);
xnor U2646 (N_2646,N_2404,N_2539);
or U2647 (N_2647,N_2429,N_2442);
nand U2648 (N_2648,N_2523,N_2470);
nor U2649 (N_2649,N_2455,N_2463);
and U2650 (N_2650,N_2503,N_2542);
xor U2651 (N_2651,N_2438,N_2494);
xor U2652 (N_2652,N_2488,N_2503);
nand U2653 (N_2653,N_2408,N_2418);
nor U2654 (N_2654,N_2401,N_2423);
or U2655 (N_2655,N_2418,N_2433);
nor U2656 (N_2656,N_2473,N_2463);
xnor U2657 (N_2657,N_2418,N_2498);
and U2658 (N_2658,N_2542,N_2539);
nand U2659 (N_2659,N_2443,N_2413);
xnor U2660 (N_2660,N_2464,N_2493);
nor U2661 (N_2661,N_2485,N_2503);
nor U2662 (N_2662,N_2535,N_2525);
xor U2663 (N_2663,N_2415,N_2518);
and U2664 (N_2664,N_2524,N_2537);
and U2665 (N_2665,N_2417,N_2429);
nand U2666 (N_2666,N_2415,N_2455);
and U2667 (N_2667,N_2415,N_2479);
and U2668 (N_2668,N_2468,N_2501);
xor U2669 (N_2669,N_2432,N_2446);
and U2670 (N_2670,N_2401,N_2527);
xnor U2671 (N_2671,N_2403,N_2500);
nand U2672 (N_2672,N_2448,N_2462);
and U2673 (N_2673,N_2457,N_2486);
nand U2674 (N_2674,N_2401,N_2475);
xnor U2675 (N_2675,N_2493,N_2475);
xnor U2676 (N_2676,N_2448,N_2530);
and U2677 (N_2677,N_2537,N_2508);
nand U2678 (N_2678,N_2533,N_2447);
xor U2679 (N_2679,N_2479,N_2463);
xnor U2680 (N_2680,N_2415,N_2516);
xor U2681 (N_2681,N_2442,N_2528);
nand U2682 (N_2682,N_2436,N_2470);
nor U2683 (N_2683,N_2445,N_2535);
nor U2684 (N_2684,N_2463,N_2509);
nand U2685 (N_2685,N_2488,N_2413);
nor U2686 (N_2686,N_2442,N_2498);
nor U2687 (N_2687,N_2469,N_2415);
nand U2688 (N_2688,N_2481,N_2427);
nand U2689 (N_2689,N_2528,N_2515);
xnor U2690 (N_2690,N_2463,N_2522);
and U2691 (N_2691,N_2493,N_2512);
nand U2692 (N_2692,N_2536,N_2470);
xnor U2693 (N_2693,N_2401,N_2421);
nor U2694 (N_2694,N_2477,N_2540);
xor U2695 (N_2695,N_2413,N_2495);
and U2696 (N_2696,N_2535,N_2456);
or U2697 (N_2697,N_2450,N_2469);
or U2698 (N_2698,N_2524,N_2400);
xor U2699 (N_2699,N_2433,N_2461);
xnor U2700 (N_2700,N_2598,N_2641);
or U2701 (N_2701,N_2583,N_2678);
and U2702 (N_2702,N_2624,N_2653);
or U2703 (N_2703,N_2627,N_2589);
or U2704 (N_2704,N_2600,N_2669);
or U2705 (N_2705,N_2637,N_2675);
nand U2706 (N_2706,N_2585,N_2689);
xnor U2707 (N_2707,N_2683,N_2552);
nand U2708 (N_2708,N_2558,N_2607);
xnor U2709 (N_2709,N_2658,N_2693);
xor U2710 (N_2710,N_2599,N_2622);
nor U2711 (N_2711,N_2605,N_2659);
xor U2712 (N_2712,N_2666,N_2566);
or U2713 (N_2713,N_2628,N_2630);
xnor U2714 (N_2714,N_2632,N_2651);
nand U2715 (N_2715,N_2640,N_2676);
nand U2716 (N_2716,N_2602,N_2687);
and U2717 (N_2717,N_2686,N_2684);
or U2718 (N_2718,N_2579,N_2673);
nor U2719 (N_2719,N_2642,N_2612);
nand U2720 (N_2720,N_2633,N_2577);
or U2721 (N_2721,N_2679,N_2616);
xnor U2722 (N_2722,N_2575,N_2587);
or U2723 (N_2723,N_2643,N_2674);
xor U2724 (N_2724,N_2609,N_2681);
and U2725 (N_2725,N_2672,N_2621);
nor U2726 (N_2726,N_2625,N_2608);
nor U2727 (N_2727,N_2593,N_2650);
nand U2728 (N_2728,N_2578,N_2572);
xor U2729 (N_2729,N_2570,N_2574);
nor U2730 (N_2730,N_2644,N_2638);
nand U2731 (N_2731,N_2639,N_2680);
nor U2732 (N_2732,N_2648,N_2554);
xor U2733 (N_2733,N_2576,N_2594);
and U2734 (N_2734,N_2565,N_2614);
xor U2735 (N_2735,N_2569,N_2584);
xnor U2736 (N_2736,N_2571,N_2695);
or U2737 (N_2737,N_2677,N_2664);
nand U2738 (N_2738,N_2610,N_2655);
and U2739 (N_2739,N_2634,N_2645);
and U2740 (N_2740,N_2568,N_2690);
nor U2741 (N_2741,N_2604,N_2567);
or U2742 (N_2742,N_2652,N_2699);
nor U2743 (N_2743,N_2619,N_2596);
nor U2744 (N_2744,N_2635,N_2682);
xor U2745 (N_2745,N_2557,N_2691);
nor U2746 (N_2746,N_2620,N_2559);
xor U2747 (N_2747,N_2564,N_2696);
or U2748 (N_2748,N_2671,N_2629);
or U2749 (N_2749,N_2623,N_2586);
and U2750 (N_2750,N_2603,N_2626);
xnor U2751 (N_2751,N_2560,N_2592);
xor U2752 (N_2752,N_2646,N_2551);
or U2753 (N_2753,N_2606,N_2697);
and U2754 (N_2754,N_2556,N_2661);
and U2755 (N_2755,N_2688,N_2694);
and U2756 (N_2756,N_2662,N_2670);
nand U2757 (N_2757,N_2663,N_2657);
and U2758 (N_2758,N_2555,N_2647);
xor U2759 (N_2759,N_2582,N_2563);
and U2760 (N_2760,N_2668,N_2562);
and U2761 (N_2761,N_2580,N_2692);
or U2762 (N_2762,N_2611,N_2581);
nand U2763 (N_2763,N_2595,N_2597);
and U2764 (N_2764,N_2590,N_2685);
and U2765 (N_2765,N_2617,N_2660);
xnor U2766 (N_2766,N_2553,N_2631);
and U2767 (N_2767,N_2591,N_2656);
and U2768 (N_2768,N_2601,N_2588);
and U2769 (N_2769,N_2550,N_2613);
xor U2770 (N_2770,N_2561,N_2698);
and U2771 (N_2771,N_2649,N_2573);
nand U2772 (N_2772,N_2618,N_2615);
nand U2773 (N_2773,N_2665,N_2654);
nor U2774 (N_2774,N_2636,N_2667);
xor U2775 (N_2775,N_2596,N_2663);
nor U2776 (N_2776,N_2634,N_2687);
and U2777 (N_2777,N_2603,N_2580);
and U2778 (N_2778,N_2687,N_2589);
and U2779 (N_2779,N_2586,N_2660);
nor U2780 (N_2780,N_2630,N_2681);
nor U2781 (N_2781,N_2568,N_2660);
nor U2782 (N_2782,N_2649,N_2577);
or U2783 (N_2783,N_2552,N_2640);
xor U2784 (N_2784,N_2648,N_2697);
or U2785 (N_2785,N_2662,N_2604);
xor U2786 (N_2786,N_2640,N_2576);
nor U2787 (N_2787,N_2624,N_2603);
xnor U2788 (N_2788,N_2608,N_2670);
or U2789 (N_2789,N_2687,N_2618);
and U2790 (N_2790,N_2611,N_2665);
or U2791 (N_2791,N_2657,N_2618);
xor U2792 (N_2792,N_2684,N_2587);
and U2793 (N_2793,N_2633,N_2611);
nor U2794 (N_2794,N_2553,N_2665);
and U2795 (N_2795,N_2650,N_2673);
xor U2796 (N_2796,N_2666,N_2670);
and U2797 (N_2797,N_2580,N_2605);
and U2798 (N_2798,N_2599,N_2621);
or U2799 (N_2799,N_2658,N_2578);
nor U2800 (N_2800,N_2617,N_2678);
and U2801 (N_2801,N_2617,N_2644);
xor U2802 (N_2802,N_2694,N_2591);
nand U2803 (N_2803,N_2674,N_2605);
xor U2804 (N_2804,N_2627,N_2587);
nor U2805 (N_2805,N_2551,N_2690);
or U2806 (N_2806,N_2603,N_2630);
or U2807 (N_2807,N_2588,N_2589);
nor U2808 (N_2808,N_2648,N_2571);
nor U2809 (N_2809,N_2581,N_2642);
and U2810 (N_2810,N_2658,N_2640);
nor U2811 (N_2811,N_2699,N_2600);
xnor U2812 (N_2812,N_2596,N_2599);
nand U2813 (N_2813,N_2597,N_2638);
xor U2814 (N_2814,N_2579,N_2555);
nand U2815 (N_2815,N_2599,N_2697);
xor U2816 (N_2816,N_2677,N_2565);
or U2817 (N_2817,N_2697,N_2605);
nand U2818 (N_2818,N_2684,N_2582);
and U2819 (N_2819,N_2688,N_2568);
nor U2820 (N_2820,N_2562,N_2568);
nand U2821 (N_2821,N_2593,N_2665);
nand U2822 (N_2822,N_2640,N_2568);
nor U2823 (N_2823,N_2609,N_2670);
and U2824 (N_2824,N_2625,N_2558);
and U2825 (N_2825,N_2600,N_2685);
xor U2826 (N_2826,N_2589,N_2621);
nor U2827 (N_2827,N_2672,N_2642);
or U2828 (N_2828,N_2558,N_2594);
nor U2829 (N_2829,N_2550,N_2666);
and U2830 (N_2830,N_2656,N_2586);
xnor U2831 (N_2831,N_2550,N_2608);
nor U2832 (N_2832,N_2642,N_2636);
nand U2833 (N_2833,N_2676,N_2687);
xnor U2834 (N_2834,N_2607,N_2677);
nor U2835 (N_2835,N_2604,N_2574);
or U2836 (N_2836,N_2593,N_2616);
or U2837 (N_2837,N_2638,N_2680);
and U2838 (N_2838,N_2577,N_2586);
nand U2839 (N_2839,N_2596,N_2623);
nand U2840 (N_2840,N_2564,N_2620);
nor U2841 (N_2841,N_2642,N_2626);
xnor U2842 (N_2842,N_2552,N_2568);
nand U2843 (N_2843,N_2632,N_2681);
nor U2844 (N_2844,N_2597,N_2683);
or U2845 (N_2845,N_2659,N_2693);
nor U2846 (N_2846,N_2591,N_2633);
nand U2847 (N_2847,N_2621,N_2603);
nor U2848 (N_2848,N_2675,N_2609);
xnor U2849 (N_2849,N_2653,N_2576);
and U2850 (N_2850,N_2713,N_2825);
and U2851 (N_2851,N_2775,N_2815);
nor U2852 (N_2852,N_2723,N_2780);
xor U2853 (N_2853,N_2833,N_2757);
and U2854 (N_2854,N_2779,N_2834);
nor U2855 (N_2855,N_2786,N_2846);
nand U2856 (N_2856,N_2738,N_2734);
and U2857 (N_2857,N_2709,N_2719);
nor U2858 (N_2858,N_2704,N_2816);
and U2859 (N_2859,N_2739,N_2756);
and U2860 (N_2860,N_2839,N_2819);
or U2861 (N_2861,N_2826,N_2702);
or U2862 (N_2862,N_2761,N_2740);
and U2863 (N_2863,N_2751,N_2804);
xor U2864 (N_2864,N_2706,N_2812);
xnor U2865 (N_2865,N_2749,N_2727);
nor U2866 (N_2866,N_2799,N_2722);
nand U2867 (N_2867,N_2845,N_2712);
and U2868 (N_2868,N_2837,N_2800);
nand U2869 (N_2869,N_2742,N_2741);
and U2870 (N_2870,N_2755,N_2790);
nor U2871 (N_2871,N_2758,N_2848);
or U2872 (N_2872,N_2787,N_2847);
or U2873 (N_2873,N_2822,N_2827);
nor U2874 (N_2874,N_2817,N_2836);
or U2875 (N_2875,N_2809,N_2746);
nor U2876 (N_2876,N_2745,N_2841);
or U2877 (N_2877,N_2724,N_2744);
nand U2878 (N_2878,N_2801,N_2843);
nor U2879 (N_2879,N_2732,N_2705);
and U2880 (N_2880,N_2830,N_2820);
and U2881 (N_2881,N_2823,N_2838);
or U2882 (N_2882,N_2793,N_2776);
and U2883 (N_2883,N_2835,N_2710);
xor U2884 (N_2884,N_2729,N_2849);
or U2885 (N_2885,N_2720,N_2763);
or U2886 (N_2886,N_2764,N_2728);
and U2887 (N_2887,N_2831,N_2700);
xnor U2888 (N_2888,N_2777,N_2708);
or U2889 (N_2889,N_2802,N_2767);
nand U2890 (N_2890,N_2731,N_2736);
xor U2891 (N_2891,N_2721,N_2711);
nand U2892 (N_2892,N_2785,N_2759);
nand U2893 (N_2893,N_2806,N_2791);
or U2894 (N_2894,N_2789,N_2842);
nor U2895 (N_2895,N_2753,N_2718);
nand U2896 (N_2896,N_2768,N_2730);
nor U2897 (N_2897,N_2784,N_2829);
or U2898 (N_2898,N_2807,N_2707);
xnor U2899 (N_2899,N_2778,N_2725);
nand U2900 (N_2900,N_2840,N_2781);
or U2901 (N_2901,N_2714,N_2716);
or U2902 (N_2902,N_2792,N_2743);
and U2903 (N_2903,N_2797,N_2828);
xnor U2904 (N_2904,N_2765,N_2798);
xnor U2905 (N_2905,N_2821,N_2747);
and U2906 (N_2906,N_2783,N_2771);
nand U2907 (N_2907,N_2774,N_2818);
and U2908 (N_2908,N_2769,N_2773);
nor U2909 (N_2909,N_2752,N_2770);
xor U2910 (N_2910,N_2788,N_2795);
or U2911 (N_2911,N_2803,N_2735);
or U2912 (N_2912,N_2844,N_2808);
nand U2913 (N_2913,N_2810,N_2717);
nor U2914 (N_2914,N_2796,N_2715);
xor U2915 (N_2915,N_2703,N_2754);
nor U2916 (N_2916,N_2766,N_2824);
xnor U2917 (N_2917,N_2772,N_2750);
nor U2918 (N_2918,N_2794,N_2782);
xnor U2919 (N_2919,N_2726,N_2748);
or U2920 (N_2920,N_2737,N_2813);
and U2921 (N_2921,N_2762,N_2811);
and U2922 (N_2922,N_2814,N_2760);
xor U2923 (N_2923,N_2701,N_2805);
and U2924 (N_2924,N_2733,N_2832);
or U2925 (N_2925,N_2782,N_2793);
nor U2926 (N_2926,N_2725,N_2732);
nor U2927 (N_2927,N_2789,N_2746);
and U2928 (N_2928,N_2805,N_2773);
xor U2929 (N_2929,N_2806,N_2837);
or U2930 (N_2930,N_2720,N_2833);
or U2931 (N_2931,N_2756,N_2785);
nor U2932 (N_2932,N_2757,N_2714);
nand U2933 (N_2933,N_2792,N_2754);
nor U2934 (N_2934,N_2826,N_2742);
nand U2935 (N_2935,N_2788,N_2742);
and U2936 (N_2936,N_2763,N_2840);
nand U2937 (N_2937,N_2809,N_2808);
and U2938 (N_2938,N_2844,N_2764);
and U2939 (N_2939,N_2723,N_2823);
and U2940 (N_2940,N_2762,N_2775);
xnor U2941 (N_2941,N_2739,N_2791);
or U2942 (N_2942,N_2778,N_2703);
xor U2943 (N_2943,N_2775,N_2821);
xor U2944 (N_2944,N_2812,N_2787);
xnor U2945 (N_2945,N_2705,N_2832);
or U2946 (N_2946,N_2759,N_2717);
or U2947 (N_2947,N_2777,N_2808);
or U2948 (N_2948,N_2724,N_2834);
and U2949 (N_2949,N_2718,N_2777);
or U2950 (N_2950,N_2718,N_2801);
and U2951 (N_2951,N_2721,N_2777);
and U2952 (N_2952,N_2713,N_2727);
nor U2953 (N_2953,N_2785,N_2832);
xnor U2954 (N_2954,N_2712,N_2817);
xor U2955 (N_2955,N_2717,N_2706);
xor U2956 (N_2956,N_2784,N_2758);
and U2957 (N_2957,N_2722,N_2797);
or U2958 (N_2958,N_2736,N_2828);
or U2959 (N_2959,N_2772,N_2757);
xor U2960 (N_2960,N_2835,N_2765);
or U2961 (N_2961,N_2769,N_2810);
or U2962 (N_2962,N_2752,N_2775);
and U2963 (N_2963,N_2802,N_2822);
xor U2964 (N_2964,N_2804,N_2797);
nor U2965 (N_2965,N_2705,N_2723);
nor U2966 (N_2966,N_2823,N_2718);
and U2967 (N_2967,N_2704,N_2745);
xnor U2968 (N_2968,N_2708,N_2768);
nand U2969 (N_2969,N_2719,N_2809);
and U2970 (N_2970,N_2736,N_2797);
nor U2971 (N_2971,N_2757,N_2762);
xor U2972 (N_2972,N_2796,N_2746);
or U2973 (N_2973,N_2739,N_2714);
nor U2974 (N_2974,N_2743,N_2744);
nand U2975 (N_2975,N_2702,N_2822);
nand U2976 (N_2976,N_2820,N_2793);
xnor U2977 (N_2977,N_2846,N_2845);
or U2978 (N_2978,N_2844,N_2813);
nand U2979 (N_2979,N_2848,N_2718);
and U2980 (N_2980,N_2815,N_2723);
nor U2981 (N_2981,N_2766,N_2775);
or U2982 (N_2982,N_2817,N_2830);
nand U2983 (N_2983,N_2726,N_2761);
or U2984 (N_2984,N_2823,N_2707);
and U2985 (N_2985,N_2720,N_2761);
nor U2986 (N_2986,N_2797,N_2765);
or U2987 (N_2987,N_2749,N_2778);
nor U2988 (N_2988,N_2711,N_2829);
or U2989 (N_2989,N_2845,N_2758);
nand U2990 (N_2990,N_2733,N_2767);
nor U2991 (N_2991,N_2787,N_2833);
or U2992 (N_2992,N_2787,N_2700);
nor U2993 (N_2993,N_2848,N_2721);
nand U2994 (N_2994,N_2787,N_2805);
xor U2995 (N_2995,N_2807,N_2784);
and U2996 (N_2996,N_2825,N_2835);
xnor U2997 (N_2997,N_2780,N_2796);
nor U2998 (N_2998,N_2794,N_2846);
or U2999 (N_2999,N_2776,N_2742);
xor U3000 (N_3000,N_2886,N_2935);
nor U3001 (N_3001,N_2961,N_2869);
xnor U3002 (N_3002,N_2968,N_2911);
or U3003 (N_3003,N_2972,N_2983);
nand U3004 (N_3004,N_2970,N_2898);
nand U3005 (N_3005,N_2978,N_2964);
xnor U3006 (N_3006,N_2969,N_2884);
nor U3007 (N_3007,N_2854,N_2872);
or U3008 (N_3008,N_2913,N_2953);
nor U3009 (N_3009,N_2862,N_2954);
or U3010 (N_3010,N_2988,N_2867);
or U3011 (N_3011,N_2910,N_2918);
nand U3012 (N_3012,N_2891,N_2896);
or U3013 (N_3013,N_2981,N_2966);
nor U3014 (N_3014,N_2903,N_2945);
nor U3015 (N_3015,N_2979,N_2864);
nand U3016 (N_3016,N_2925,N_2990);
and U3017 (N_3017,N_2857,N_2874);
or U3018 (N_3018,N_2938,N_2985);
nand U3019 (N_3019,N_2955,N_2996);
or U3020 (N_3020,N_2951,N_2971);
xnor U3021 (N_3021,N_2948,N_2940);
nor U3022 (N_3022,N_2957,N_2958);
or U3023 (N_3023,N_2899,N_2924);
and U3024 (N_3024,N_2930,N_2851);
xnor U3025 (N_3025,N_2998,N_2895);
nand U3026 (N_3026,N_2859,N_2976);
nand U3027 (N_3027,N_2991,N_2977);
xnor U3028 (N_3028,N_2893,N_2926);
and U3029 (N_3029,N_2865,N_2875);
nor U3030 (N_3030,N_2878,N_2931);
nand U3031 (N_3031,N_2959,N_2944);
nand U3032 (N_3032,N_2897,N_2919);
and U3033 (N_3033,N_2852,N_2994);
xor U3034 (N_3034,N_2863,N_2912);
nand U3035 (N_3035,N_2923,N_2889);
nand U3036 (N_3036,N_2853,N_2965);
xor U3037 (N_3037,N_2992,N_2892);
xnor U3038 (N_3038,N_2933,N_2932);
nand U3039 (N_3039,N_2902,N_2962);
nand U3040 (N_3040,N_2984,N_2974);
nor U3041 (N_3041,N_2942,N_2937);
xor U3042 (N_3042,N_2963,N_2861);
or U3043 (N_3043,N_2997,N_2900);
or U3044 (N_3044,N_2880,N_2989);
nand U3045 (N_3045,N_2882,N_2927);
nor U3046 (N_3046,N_2905,N_2890);
nand U3047 (N_3047,N_2855,N_2995);
nand U3048 (N_3048,N_2916,N_2894);
xnor U3049 (N_3049,N_2941,N_2947);
and U3050 (N_3050,N_2879,N_2939);
and U3051 (N_3051,N_2888,N_2936);
xnor U3052 (N_3052,N_2856,N_2858);
and U3053 (N_3053,N_2887,N_2904);
xor U3054 (N_3054,N_2866,N_2908);
xor U3055 (N_3055,N_2914,N_2986);
and U3056 (N_3056,N_2973,N_2956);
xnor U3057 (N_3057,N_2920,N_2876);
nand U3058 (N_3058,N_2883,N_2917);
nor U3059 (N_3059,N_2885,N_2949);
or U3060 (N_3060,N_2928,N_2934);
xnor U3061 (N_3061,N_2987,N_2946);
or U3062 (N_3062,N_2980,N_2943);
nor U3063 (N_3063,N_2921,N_2860);
and U3064 (N_3064,N_2952,N_2915);
and U3065 (N_3065,N_2960,N_2922);
xor U3066 (N_3066,N_2907,N_2850);
or U3067 (N_3067,N_2870,N_2909);
nor U3068 (N_3068,N_2873,N_2993);
and U3069 (N_3069,N_2906,N_2881);
xnor U3070 (N_3070,N_2982,N_2929);
and U3071 (N_3071,N_2999,N_2868);
xnor U3072 (N_3072,N_2877,N_2871);
or U3073 (N_3073,N_2950,N_2975);
xor U3074 (N_3074,N_2901,N_2967);
nand U3075 (N_3075,N_2870,N_2861);
nor U3076 (N_3076,N_2993,N_2972);
nand U3077 (N_3077,N_2902,N_2908);
nand U3078 (N_3078,N_2870,N_2941);
and U3079 (N_3079,N_2911,N_2895);
xor U3080 (N_3080,N_2897,N_2879);
xor U3081 (N_3081,N_2918,N_2886);
nor U3082 (N_3082,N_2866,N_2915);
or U3083 (N_3083,N_2866,N_2882);
and U3084 (N_3084,N_2953,N_2921);
or U3085 (N_3085,N_2978,N_2899);
xor U3086 (N_3086,N_2862,N_2989);
nand U3087 (N_3087,N_2934,N_2904);
nor U3088 (N_3088,N_2850,N_2864);
nor U3089 (N_3089,N_2892,N_2931);
and U3090 (N_3090,N_2863,N_2991);
and U3091 (N_3091,N_2888,N_2900);
and U3092 (N_3092,N_2937,N_2995);
and U3093 (N_3093,N_2891,N_2899);
xnor U3094 (N_3094,N_2913,N_2886);
or U3095 (N_3095,N_2949,N_2971);
and U3096 (N_3096,N_2894,N_2936);
xor U3097 (N_3097,N_2893,N_2954);
nand U3098 (N_3098,N_2959,N_2899);
nor U3099 (N_3099,N_2885,N_2901);
xor U3100 (N_3100,N_2965,N_2980);
and U3101 (N_3101,N_2943,N_2959);
nand U3102 (N_3102,N_2898,N_2855);
xnor U3103 (N_3103,N_2886,N_2961);
or U3104 (N_3104,N_2991,N_2981);
and U3105 (N_3105,N_2969,N_2939);
xnor U3106 (N_3106,N_2877,N_2969);
or U3107 (N_3107,N_2893,N_2941);
nand U3108 (N_3108,N_2861,N_2943);
nor U3109 (N_3109,N_2908,N_2869);
and U3110 (N_3110,N_2893,N_2990);
or U3111 (N_3111,N_2936,N_2982);
and U3112 (N_3112,N_2856,N_2932);
or U3113 (N_3113,N_2951,N_2924);
nor U3114 (N_3114,N_2973,N_2915);
nand U3115 (N_3115,N_2987,N_2962);
nor U3116 (N_3116,N_2890,N_2897);
nor U3117 (N_3117,N_2903,N_2894);
nor U3118 (N_3118,N_2933,N_2882);
and U3119 (N_3119,N_2852,N_2931);
nand U3120 (N_3120,N_2920,N_2928);
or U3121 (N_3121,N_2933,N_2911);
xnor U3122 (N_3122,N_2946,N_2979);
nand U3123 (N_3123,N_2920,N_2997);
and U3124 (N_3124,N_2875,N_2950);
xor U3125 (N_3125,N_2936,N_2903);
xor U3126 (N_3126,N_2874,N_2930);
and U3127 (N_3127,N_2859,N_2897);
or U3128 (N_3128,N_2962,N_2999);
xnor U3129 (N_3129,N_2928,N_2935);
nor U3130 (N_3130,N_2937,N_2863);
or U3131 (N_3131,N_2870,N_2995);
xnor U3132 (N_3132,N_2965,N_2916);
xor U3133 (N_3133,N_2927,N_2984);
or U3134 (N_3134,N_2950,N_2856);
nor U3135 (N_3135,N_2893,N_2946);
xor U3136 (N_3136,N_2965,N_2935);
and U3137 (N_3137,N_2888,N_2850);
nand U3138 (N_3138,N_2903,N_2955);
nand U3139 (N_3139,N_2853,N_2874);
nand U3140 (N_3140,N_2890,N_2867);
and U3141 (N_3141,N_2976,N_2866);
nor U3142 (N_3142,N_2917,N_2882);
or U3143 (N_3143,N_2914,N_2941);
xnor U3144 (N_3144,N_2890,N_2864);
xnor U3145 (N_3145,N_2934,N_2946);
nand U3146 (N_3146,N_2957,N_2924);
nand U3147 (N_3147,N_2921,N_2923);
nand U3148 (N_3148,N_2886,N_2916);
nor U3149 (N_3149,N_2882,N_2964);
nand U3150 (N_3150,N_3109,N_3075);
nor U3151 (N_3151,N_3094,N_3099);
or U3152 (N_3152,N_3124,N_3015);
xnor U3153 (N_3153,N_3062,N_3056);
nor U3154 (N_3154,N_3043,N_3106);
nor U3155 (N_3155,N_3126,N_3129);
nor U3156 (N_3156,N_3070,N_3082);
nand U3157 (N_3157,N_3083,N_3141);
nor U3158 (N_3158,N_3093,N_3134);
nor U3159 (N_3159,N_3088,N_3135);
nor U3160 (N_3160,N_3024,N_3001);
and U3161 (N_3161,N_3107,N_3097);
nand U3162 (N_3162,N_3013,N_3098);
xor U3163 (N_3163,N_3038,N_3022);
xnor U3164 (N_3164,N_3058,N_3104);
xor U3165 (N_3165,N_3128,N_3130);
xnor U3166 (N_3166,N_3139,N_3054);
xor U3167 (N_3167,N_3017,N_3089);
or U3168 (N_3168,N_3047,N_3048);
nand U3169 (N_3169,N_3080,N_3147);
xor U3170 (N_3170,N_3084,N_3050);
and U3171 (N_3171,N_3142,N_3076);
nand U3172 (N_3172,N_3121,N_3049);
nand U3173 (N_3173,N_3133,N_3005);
nand U3174 (N_3174,N_3060,N_3132);
nor U3175 (N_3175,N_3012,N_3113);
xor U3176 (N_3176,N_3127,N_3009);
nor U3177 (N_3177,N_3023,N_3105);
nor U3178 (N_3178,N_3069,N_3136);
nand U3179 (N_3179,N_3042,N_3125);
or U3180 (N_3180,N_3033,N_3149);
and U3181 (N_3181,N_3072,N_3111);
and U3182 (N_3182,N_3085,N_3031);
and U3183 (N_3183,N_3041,N_3006);
nor U3184 (N_3184,N_3144,N_3091);
xor U3185 (N_3185,N_3067,N_3077);
and U3186 (N_3186,N_3131,N_3010);
xor U3187 (N_3187,N_3074,N_3008);
and U3188 (N_3188,N_3143,N_3137);
xnor U3189 (N_3189,N_3071,N_3061);
nand U3190 (N_3190,N_3039,N_3028);
nor U3191 (N_3191,N_3035,N_3102);
or U3192 (N_3192,N_3020,N_3116);
or U3193 (N_3193,N_3115,N_3087);
or U3194 (N_3194,N_3016,N_3000);
and U3195 (N_3195,N_3003,N_3034);
and U3196 (N_3196,N_3138,N_3073);
and U3197 (N_3197,N_3146,N_3140);
nand U3198 (N_3198,N_3051,N_3103);
nor U3199 (N_3199,N_3118,N_3078);
and U3200 (N_3200,N_3100,N_3057);
nand U3201 (N_3201,N_3002,N_3026);
xor U3202 (N_3202,N_3110,N_3108);
and U3203 (N_3203,N_3081,N_3025);
xor U3204 (N_3204,N_3066,N_3119);
and U3205 (N_3205,N_3032,N_3052);
and U3206 (N_3206,N_3092,N_3007);
nor U3207 (N_3207,N_3086,N_3059);
or U3208 (N_3208,N_3055,N_3029);
nor U3209 (N_3209,N_3004,N_3011);
nand U3210 (N_3210,N_3037,N_3120);
xnor U3211 (N_3211,N_3019,N_3021);
and U3212 (N_3212,N_3046,N_3018);
and U3213 (N_3213,N_3040,N_3063);
or U3214 (N_3214,N_3145,N_3095);
nor U3215 (N_3215,N_3090,N_3079);
nand U3216 (N_3216,N_3027,N_3065);
xnor U3217 (N_3217,N_3101,N_3068);
or U3218 (N_3218,N_3117,N_3044);
xnor U3219 (N_3219,N_3030,N_3148);
nor U3220 (N_3220,N_3096,N_3122);
xnor U3221 (N_3221,N_3123,N_3036);
nand U3222 (N_3222,N_3045,N_3114);
or U3223 (N_3223,N_3112,N_3064);
xor U3224 (N_3224,N_3014,N_3053);
and U3225 (N_3225,N_3141,N_3099);
and U3226 (N_3226,N_3113,N_3125);
or U3227 (N_3227,N_3050,N_3137);
xnor U3228 (N_3228,N_3138,N_3102);
nand U3229 (N_3229,N_3078,N_3072);
xor U3230 (N_3230,N_3142,N_3107);
nand U3231 (N_3231,N_3039,N_3105);
nand U3232 (N_3232,N_3085,N_3088);
or U3233 (N_3233,N_3059,N_3072);
nor U3234 (N_3234,N_3027,N_3087);
nor U3235 (N_3235,N_3130,N_3017);
and U3236 (N_3236,N_3067,N_3074);
and U3237 (N_3237,N_3068,N_3059);
nor U3238 (N_3238,N_3049,N_3096);
or U3239 (N_3239,N_3023,N_3132);
or U3240 (N_3240,N_3014,N_3133);
nor U3241 (N_3241,N_3066,N_3131);
and U3242 (N_3242,N_3115,N_3041);
and U3243 (N_3243,N_3055,N_3058);
or U3244 (N_3244,N_3147,N_3111);
nand U3245 (N_3245,N_3067,N_3091);
xnor U3246 (N_3246,N_3045,N_3030);
or U3247 (N_3247,N_3023,N_3021);
xnor U3248 (N_3248,N_3009,N_3097);
or U3249 (N_3249,N_3103,N_3134);
xor U3250 (N_3250,N_3131,N_3052);
nor U3251 (N_3251,N_3062,N_3112);
and U3252 (N_3252,N_3119,N_3148);
xnor U3253 (N_3253,N_3028,N_3097);
nor U3254 (N_3254,N_3056,N_3125);
and U3255 (N_3255,N_3089,N_3064);
and U3256 (N_3256,N_3067,N_3096);
or U3257 (N_3257,N_3148,N_3073);
nand U3258 (N_3258,N_3069,N_3037);
nand U3259 (N_3259,N_3021,N_3123);
and U3260 (N_3260,N_3084,N_3063);
nor U3261 (N_3261,N_3083,N_3000);
nand U3262 (N_3262,N_3018,N_3109);
or U3263 (N_3263,N_3082,N_3073);
xnor U3264 (N_3264,N_3032,N_3126);
or U3265 (N_3265,N_3112,N_3087);
nor U3266 (N_3266,N_3109,N_3061);
nor U3267 (N_3267,N_3014,N_3076);
or U3268 (N_3268,N_3149,N_3050);
or U3269 (N_3269,N_3130,N_3051);
or U3270 (N_3270,N_3019,N_3001);
or U3271 (N_3271,N_3029,N_3120);
and U3272 (N_3272,N_3126,N_3102);
or U3273 (N_3273,N_3001,N_3138);
nor U3274 (N_3274,N_3068,N_3022);
nor U3275 (N_3275,N_3022,N_3118);
xnor U3276 (N_3276,N_3109,N_3147);
nor U3277 (N_3277,N_3035,N_3062);
or U3278 (N_3278,N_3100,N_3074);
and U3279 (N_3279,N_3107,N_3006);
and U3280 (N_3280,N_3027,N_3044);
xor U3281 (N_3281,N_3045,N_3060);
nor U3282 (N_3282,N_3111,N_3122);
nor U3283 (N_3283,N_3037,N_3026);
xnor U3284 (N_3284,N_3097,N_3126);
or U3285 (N_3285,N_3090,N_3122);
xor U3286 (N_3286,N_3134,N_3034);
nand U3287 (N_3287,N_3097,N_3006);
and U3288 (N_3288,N_3047,N_3051);
and U3289 (N_3289,N_3017,N_3109);
and U3290 (N_3290,N_3059,N_3095);
nor U3291 (N_3291,N_3105,N_3148);
nor U3292 (N_3292,N_3015,N_3107);
nor U3293 (N_3293,N_3110,N_3044);
nand U3294 (N_3294,N_3058,N_3080);
and U3295 (N_3295,N_3047,N_3083);
xnor U3296 (N_3296,N_3081,N_3111);
and U3297 (N_3297,N_3088,N_3030);
xnor U3298 (N_3298,N_3140,N_3108);
nor U3299 (N_3299,N_3145,N_3123);
nand U3300 (N_3300,N_3177,N_3163);
or U3301 (N_3301,N_3186,N_3222);
nand U3302 (N_3302,N_3249,N_3285);
nor U3303 (N_3303,N_3245,N_3180);
nand U3304 (N_3304,N_3255,N_3184);
or U3305 (N_3305,N_3251,N_3195);
and U3306 (N_3306,N_3232,N_3275);
xnor U3307 (N_3307,N_3281,N_3240);
or U3308 (N_3308,N_3233,N_3223);
and U3309 (N_3309,N_3253,N_3261);
xnor U3310 (N_3310,N_3269,N_3214);
or U3311 (N_3311,N_3264,N_3297);
nor U3312 (N_3312,N_3156,N_3162);
xnor U3313 (N_3313,N_3262,N_3290);
nor U3314 (N_3314,N_3260,N_3203);
and U3315 (N_3315,N_3234,N_3194);
xnor U3316 (N_3316,N_3287,N_3244);
nand U3317 (N_3317,N_3252,N_3207);
nand U3318 (N_3318,N_3173,N_3201);
xor U3319 (N_3319,N_3196,N_3190);
or U3320 (N_3320,N_3272,N_3289);
xnor U3321 (N_3321,N_3217,N_3288);
nand U3322 (N_3322,N_3200,N_3158);
nand U3323 (N_3323,N_3185,N_3270);
xnor U3324 (N_3324,N_3182,N_3266);
xor U3325 (N_3325,N_3188,N_3208);
nor U3326 (N_3326,N_3284,N_3237);
or U3327 (N_3327,N_3229,N_3187);
nand U3328 (N_3328,N_3176,N_3226);
nor U3329 (N_3329,N_3213,N_3283);
nand U3330 (N_3330,N_3206,N_3204);
xor U3331 (N_3331,N_3227,N_3299);
nand U3332 (N_3332,N_3168,N_3157);
xor U3333 (N_3333,N_3220,N_3216);
nand U3334 (N_3334,N_3164,N_3265);
or U3335 (N_3335,N_3174,N_3243);
nor U3336 (N_3336,N_3155,N_3293);
or U3337 (N_3337,N_3179,N_3231);
nor U3338 (N_3338,N_3193,N_3254);
xnor U3339 (N_3339,N_3211,N_3246);
nand U3340 (N_3340,N_3171,N_3292);
or U3341 (N_3341,N_3271,N_3259);
nor U3342 (N_3342,N_3242,N_3170);
or U3343 (N_3343,N_3236,N_3250);
nor U3344 (N_3344,N_3181,N_3276);
or U3345 (N_3345,N_3169,N_3152);
or U3346 (N_3346,N_3159,N_3202);
or U3347 (N_3347,N_3298,N_3280);
and U3348 (N_3348,N_3192,N_3215);
and U3349 (N_3349,N_3224,N_3268);
nand U3350 (N_3350,N_3175,N_3278);
and U3351 (N_3351,N_3256,N_3277);
or U3352 (N_3352,N_3228,N_3166);
or U3353 (N_3353,N_3221,N_3153);
nor U3354 (N_3354,N_3219,N_3257);
nor U3355 (N_3355,N_3183,N_3274);
xor U3356 (N_3356,N_3178,N_3151);
xor U3357 (N_3357,N_3209,N_3225);
xnor U3358 (N_3358,N_3279,N_3248);
nand U3359 (N_3359,N_3197,N_3161);
xnor U3360 (N_3360,N_3286,N_3172);
or U3361 (N_3361,N_3198,N_3258);
and U3362 (N_3362,N_3165,N_3296);
xor U3363 (N_3363,N_3160,N_3238);
nor U3364 (N_3364,N_3212,N_3294);
and U3365 (N_3365,N_3189,N_3218);
xnor U3366 (N_3366,N_3150,N_3205);
nand U3367 (N_3367,N_3241,N_3273);
nor U3368 (N_3368,N_3295,N_3154);
and U3369 (N_3369,N_3167,N_3263);
or U3370 (N_3370,N_3191,N_3239);
nor U3371 (N_3371,N_3235,N_3230);
and U3372 (N_3372,N_3282,N_3291);
or U3373 (N_3373,N_3210,N_3267);
nand U3374 (N_3374,N_3247,N_3199);
and U3375 (N_3375,N_3265,N_3226);
and U3376 (N_3376,N_3152,N_3175);
and U3377 (N_3377,N_3206,N_3162);
nand U3378 (N_3378,N_3288,N_3286);
xnor U3379 (N_3379,N_3197,N_3165);
and U3380 (N_3380,N_3279,N_3261);
nand U3381 (N_3381,N_3215,N_3207);
nor U3382 (N_3382,N_3182,N_3299);
or U3383 (N_3383,N_3258,N_3154);
and U3384 (N_3384,N_3164,N_3199);
or U3385 (N_3385,N_3192,N_3160);
and U3386 (N_3386,N_3212,N_3218);
and U3387 (N_3387,N_3195,N_3167);
nor U3388 (N_3388,N_3190,N_3270);
xor U3389 (N_3389,N_3286,N_3217);
nor U3390 (N_3390,N_3177,N_3228);
nand U3391 (N_3391,N_3236,N_3209);
or U3392 (N_3392,N_3199,N_3223);
or U3393 (N_3393,N_3274,N_3291);
nor U3394 (N_3394,N_3224,N_3156);
nor U3395 (N_3395,N_3157,N_3287);
nor U3396 (N_3396,N_3196,N_3213);
xor U3397 (N_3397,N_3253,N_3170);
nor U3398 (N_3398,N_3176,N_3211);
or U3399 (N_3399,N_3277,N_3209);
and U3400 (N_3400,N_3180,N_3172);
nand U3401 (N_3401,N_3176,N_3294);
or U3402 (N_3402,N_3230,N_3234);
nand U3403 (N_3403,N_3199,N_3237);
or U3404 (N_3404,N_3250,N_3185);
nor U3405 (N_3405,N_3238,N_3184);
or U3406 (N_3406,N_3280,N_3196);
xor U3407 (N_3407,N_3192,N_3231);
nor U3408 (N_3408,N_3202,N_3297);
xnor U3409 (N_3409,N_3159,N_3231);
and U3410 (N_3410,N_3237,N_3154);
xnor U3411 (N_3411,N_3258,N_3260);
xor U3412 (N_3412,N_3170,N_3153);
nand U3413 (N_3413,N_3263,N_3243);
nand U3414 (N_3414,N_3288,N_3176);
nor U3415 (N_3415,N_3184,N_3156);
xnor U3416 (N_3416,N_3207,N_3238);
nand U3417 (N_3417,N_3292,N_3261);
nand U3418 (N_3418,N_3153,N_3242);
or U3419 (N_3419,N_3245,N_3151);
xnor U3420 (N_3420,N_3232,N_3201);
and U3421 (N_3421,N_3224,N_3259);
xor U3422 (N_3422,N_3204,N_3260);
and U3423 (N_3423,N_3230,N_3295);
nor U3424 (N_3424,N_3253,N_3173);
nand U3425 (N_3425,N_3238,N_3208);
or U3426 (N_3426,N_3238,N_3162);
and U3427 (N_3427,N_3290,N_3282);
xor U3428 (N_3428,N_3209,N_3178);
nor U3429 (N_3429,N_3164,N_3207);
and U3430 (N_3430,N_3249,N_3186);
nand U3431 (N_3431,N_3236,N_3237);
or U3432 (N_3432,N_3197,N_3254);
nand U3433 (N_3433,N_3243,N_3162);
nor U3434 (N_3434,N_3266,N_3184);
nor U3435 (N_3435,N_3211,N_3240);
xnor U3436 (N_3436,N_3184,N_3191);
nand U3437 (N_3437,N_3164,N_3216);
nand U3438 (N_3438,N_3198,N_3248);
xor U3439 (N_3439,N_3190,N_3208);
and U3440 (N_3440,N_3296,N_3243);
or U3441 (N_3441,N_3194,N_3237);
and U3442 (N_3442,N_3263,N_3230);
or U3443 (N_3443,N_3229,N_3236);
xnor U3444 (N_3444,N_3192,N_3269);
nor U3445 (N_3445,N_3282,N_3199);
nand U3446 (N_3446,N_3286,N_3254);
or U3447 (N_3447,N_3208,N_3203);
nand U3448 (N_3448,N_3268,N_3231);
and U3449 (N_3449,N_3189,N_3238);
xor U3450 (N_3450,N_3339,N_3378);
xnor U3451 (N_3451,N_3344,N_3418);
nand U3452 (N_3452,N_3317,N_3333);
nor U3453 (N_3453,N_3314,N_3323);
nor U3454 (N_3454,N_3365,N_3332);
xnor U3455 (N_3455,N_3316,N_3373);
nor U3456 (N_3456,N_3442,N_3381);
xnor U3457 (N_3457,N_3355,N_3393);
nand U3458 (N_3458,N_3440,N_3385);
or U3459 (N_3459,N_3307,N_3356);
and U3460 (N_3460,N_3380,N_3342);
and U3461 (N_3461,N_3387,N_3347);
xor U3462 (N_3462,N_3375,N_3384);
or U3463 (N_3463,N_3352,N_3383);
nor U3464 (N_3464,N_3345,N_3376);
nor U3465 (N_3465,N_3422,N_3372);
and U3466 (N_3466,N_3327,N_3358);
and U3467 (N_3467,N_3368,N_3382);
and U3468 (N_3468,N_3338,N_3424);
nor U3469 (N_3469,N_3444,N_3417);
xor U3470 (N_3470,N_3340,N_3407);
xor U3471 (N_3471,N_3438,N_3366);
nor U3472 (N_3472,N_3404,N_3349);
nand U3473 (N_3473,N_3426,N_3441);
or U3474 (N_3474,N_3446,N_3421);
and U3475 (N_3475,N_3405,N_3392);
or U3476 (N_3476,N_3434,N_3359);
nor U3477 (N_3477,N_3389,N_3377);
xnor U3478 (N_3478,N_3348,N_3374);
xor U3479 (N_3479,N_3411,N_3361);
xnor U3480 (N_3480,N_3413,N_3300);
and U3481 (N_3481,N_3394,N_3326);
and U3482 (N_3482,N_3341,N_3427);
and U3483 (N_3483,N_3335,N_3325);
nand U3484 (N_3484,N_3319,N_3329);
and U3485 (N_3485,N_3312,N_3390);
nor U3486 (N_3486,N_3334,N_3437);
and U3487 (N_3487,N_3448,N_3363);
nor U3488 (N_3488,N_3430,N_3410);
nand U3489 (N_3489,N_3449,N_3397);
nor U3490 (N_3490,N_3400,N_3406);
or U3491 (N_3491,N_3416,N_3306);
nand U3492 (N_3492,N_3310,N_3414);
nor U3493 (N_3493,N_3425,N_3360);
nand U3494 (N_3494,N_3346,N_3354);
xor U3495 (N_3495,N_3353,N_3433);
nand U3496 (N_3496,N_3403,N_3322);
xnor U3497 (N_3497,N_3315,N_3402);
nand U3498 (N_3498,N_3398,N_3313);
nor U3499 (N_3499,N_3370,N_3304);
nor U3500 (N_3500,N_3367,N_3409);
nand U3501 (N_3501,N_3431,N_3330);
nand U3502 (N_3502,N_3399,N_3324);
or U3503 (N_3503,N_3337,N_3331);
nor U3504 (N_3504,N_3302,N_3351);
nand U3505 (N_3505,N_3412,N_3321);
nand U3506 (N_3506,N_3320,N_3308);
xnor U3507 (N_3507,N_3391,N_3386);
nor U3508 (N_3508,N_3305,N_3379);
and U3509 (N_3509,N_3309,N_3439);
nand U3510 (N_3510,N_3364,N_3369);
nand U3511 (N_3511,N_3318,N_3362);
or U3512 (N_3512,N_3357,N_3336);
nor U3513 (N_3513,N_3447,N_3388);
nor U3514 (N_3514,N_3328,N_3350);
nand U3515 (N_3515,N_3428,N_3423);
and U3516 (N_3516,N_3445,N_3415);
and U3517 (N_3517,N_3420,N_3301);
nand U3518 (N_3518,N_3343,N_3371);
nor U3519 (N_3519,N_3395,N_3408);
nor U3520 (N_3520,N_3401,N_3396);
xnor U3521 (N_3521,N_3419,N_3443);
or U3522 (N_3522,N_3429,N_3435);
nor U3523 (N_3523,N_3311,N_3303);
nor U3524 (N_3524,N_3436,N_3432);
xor U3525 (N_3525,N_3404,N_3378);
nor U3526 (N_3526,N_3326,N_3360);
and U3527 (N_3527,N_3415,N_3303);
or U3528 (N_3528,N_3424,N_3405);
nor U3529 (N_3529,N_3441,N_3408);
nor U3530 (N_3530,N_3432,N_3376);
and U3531 (N_3531,N_3362,N_3321);
and U3532 (N_3532,N_3405,N_3301);
and U3533 (N_3533,N_3362,N_3342);
xnor U3534 (N_3534,N_3394,N_3351);
and U3535 (N_3535,N_3315,N_3380);
nand U3536 (N_3536,N_3436,N_3413);
nor U3537 (N_3537,N_3419,N_3368);
nand U3538 (N_3538,N_3338,N_3445);
nand U3539 (N_3539,N_3329,N_3348);
xnor U3540 (N_3540,N_3440,N_3334);
nor U3541 (N_3541,N_3435,N_3352);
and U3542 (N_3542,N_3379,N_3427);
xnor U3543 (N_3543,N_3446,N_3365);
and U3544 (N_3544,N_3413,N_3349);
or U3545 (N_3545,N_3336,N_3416);
and U3546 (N_3546,N_3353,N_3356);
or U3547 (N_3547,N_3334,N_3434);
or U3548 (N_3548,N_3318,N_3338);
nor U3549 (N_3549,N_3410,N_3355);
xor U3550 (N_3550,N_3400,N_3446);
or U3551 (N_3551,N_3395,N_3387);
xor U3552 (N_3552,N_3438,N_3374);
and U3553 (N_3553,N_3410,N_3307);
xnor U3554 (N_3554,N_3427,N_3355);
nand U3555 (N_3555,N_3437,N_3424);
xnor U3556 (N_3556,N_3449,N_3344);
xor U3557 (N_3557,N_3313,N_3354);
or U3558 (N_3558,N_3393,N_3339);
or U3559 (N_3559,N_3363,N_3379);
xor U3560 (N_3560,N_3437,N_3341);
and U3561 (N_3561,N_3377,N_3353);
or U3562 (N_3562,N_3446,N_3420);
nand U3563 (N_3563,N_3380,N_3339);
or U3564 (N_3564,N_3315,N_3379);
nand U3565 (N_3565,N_3403,N_3423);
and U3566 (N_3566,N_3344,N_3423);
and U3567 (N_3567,N_3373,N_3412);
xnor U3568 (N_3568,N_3397,N_3385);
and U3569 (N_3569,N_3408,N_3442);
and U3570 (N_3570,N_3390,N_3446);
or U3571 (N_3571,N_3374,N_3419);
or U3572 (N_3572,N_3329,N_3386);
or U3573 (N_3573,N_3338,N_3392);
or U3574 (N_3574,N_3389,N_3384);
xnor U3575 (N_3575,N_3319,N_3306);
nor U3576 (N_3576,N_3319,N_3322);
nor U3577 (N_3577,N_3300,N_3379);
xor U3578 (N_3578,N_3391,N_3323);
nand U3579 (N_3579,N_3379,N_3401);
nor U3580 (N_3580,N_3301,N_3423);
nand U3581 (N_3581,N_3442,N_3430);
nor U3582 (N_3582,N_3358,N_3396);
nor U3583 (N_3583,N_3344,N_3374);
nor U3584 (N_3584,N_3413,N_3380);
nor U3585 (N_3585,N_3403,N_3323);
and U3586 (N_3586,N_3301,N_3422);
or U3587 (N_3587,N_3363,N_3384);
or U3588 (N_3588,N_3397,N_3446);
and U3589 (N_3589,N_3330,N_3415);
nand U3590 (N_3590,N_3384,N_3369);
nand U3591 (N_3591,N_3313,N_3342);
nor U3592 (N_3592,N_3307,N_3350);
and U3593 (N_3593,N_3316,N_3411);
nor U3594 (N_3594,N_3407,N_3424);
or U3595 (N_3595,N_3405,N_3428);
and U3596 (N_3596,N_3304,N_3346);
and U3597 (N_3597,N_3356,N_3434);
or U3598 (N_3598,N_3303,N_3302);
and U3599 (N_3599,N_3428,N_3418);
xnor U3600 (N_3600,N_3497,N_3489);
nand U3601 (N_3601,N_3468,N_3453);
or U3602 (N_3602,N_3533,N_3562);
and U3603 (N_3603,N_3558,N_3572);
xnor U3604 (N_3604,N_3554,N_3561);
nand U3605 (N_3605,N_3485,N_3538);
or U3606 (N_3606,N_3487,N_3596);
nand U3607 (N_3607,N_3503,N_3512);
or U3608 (N_3608,N_3593,N_3484);
nor U3609 (N_3609,N_3551,N_3535);
xnor U3610 (N_3610,N_3482,N_3595);
nor U3611 (N_3611,N_3496,N_3478);
or U3612 (N_3612,N_3576,N_3462);
nand U3613 (N_3613,N_3521,N_3454);
xnor U3614 (N_3614,N_3455,N_3559);
or U3615 (N_3615,N_3479,N_3466);
and U3616 (N_3616,N_3560,N_3520);
nor U3617 (N_3617,N_3569,N_3540);
nand U3618 (N_3618,N_3575,N_3529);
xor U3619 (N_3619,N_3473,N_3506);
xnor U3620 (N_3620,N_3480,N_3567);
and U3621 (N_3621,N_3470,N_3579);
or U3622 (N_3622,N_3458,N_3452);
xnor U3623 (N_3623,N_3585,N_3501);
xor U3624 (N_3624,N_3451,N_3543);
xor U3625 (N_3625,N_3589,N_3588);
and U3626 (N_3626,N_3481,N_3528);
nor U3627 (N_3627,N_3460,N_3536);
nor U3628 (N_3628,N_3517,N_3518);
or U3629 (N_3629,N_3499,N_3465);
nand U3630 (N_3630,N_3586,N_3582);
nand U3631 (N_3631,N_3508,N_3553);
xor U3632 (N_3632,N_3594,N_3461);
nand U3633 (N_3633,N_3568,N_3564);
nand U3634 (N_3634,N_3534,N_3515);
xor U3635 (N_3635,N_3587,N_3477);
nor U3636 (N_3636,N_3527,N_3495);
xnor U3637 (N_3637,N_3548,N_3549);
and U3638 (N_3638,N_3504,N_3476);
xnor U3639 (N_3639,N_3519,N_3581);
or U3640 (N_3640,N_3571,N_3463);
xnor U3641 (N_3641,N_3577,N_3511);
and U3642 (N_3642,N_3509,N_3552);
xor U3643 (N_3643,N_3513,N_3598);
nand U3644 (N_3644,N_3486,N_3464);
nand U3645 (N_3645,N_3471,N_3532);
and U3646 (N_3646,N_3524,N_3541);
nand U3647 (N_3647,N_3469,N_3474);
or U3648 (N_3648,N_3556,N_3578);
xor U3649 (N_3649,N_3597,N_3494);
nor U3650 (N_3650,N_3592,N_3502);
nand U3651 (N_3651,N_3491,N_3514);
nand U3652 (N_3652,N_3459,N_3584);
and U3653 (N_3653,N_3545,N_3555);
xnor U3654 (N_3654,N_3590,N_3542);
nor U3655 (N_3655,N_3537,N_3550);
or U3656 (N_3656,N_3450,N_3547);
and U3657 (N_3657,N_3483,N_3526);
nand U3658 (N_3658,N_3488,N_3544);
nor U3659 (N_3659,N_3500,N_3472);
and U3660 (N_3660,N_3583,N_3591);
and U3661 (N_3661,N_3498,N_3507);
and U3662 (N_3662,N_3539,N_3493);
nand U3663 (N_3663,N_3457,N_3599);
nor U3664 (N_3664,N_3565,N_3475);
nor U3665 (N_3665,N_3505,N_3490);
or U3666 (N_3666,N_3563,N_3492);
and U3667 (N_3667,N_3516,N_3523);
nor U3668 (N_3668,N_3566,N_3510);
nor U3669 (N_3669,N_3531,N_3522);
or U3670 (N_3670,N_3570,N_3546);
and U3671 (N_3671,N_3456,N_3573);
nor U3672 (N_3672,N_3574,N_3530);
nor U3673 (N_3673,N_3467,N_3525);
and U3674 (N_3674,N_3580,N_3557);
xnor U3675 (N_3675,N_3591,N_3483);
nor U3676 (N_3676,N_3548,N_3577);
and U3677 (N_3677,N_3471,N_3583);
and U3678 (N_3678,N_3555,N_3508);
nand U3679 (N_3679,N_3452,N_3590);
nand U3680 (N_3680,N_3453,N_3481);
xnor U3681 (N_3681,N_3542,N_3547);
or U3682 (N_3682,N_3451,N_3539);
nand U3683 (N_3683,N_3565,N_3480);
nand U3684 (N_3684,N_3475,N_3599);
or U3685 (N_3685,N_3501,N_3595);
or U3686 (N_3686,N_3466,N_3477);
nand U3687 (N_3687,N_3595,N_3525);
nand U3688 (N_3688,N_3510,N_3527);
nor U3689 (N_3689,N_3471,N_3509);
or U3690 (N_3690,N_3457,N_3451);
nor U3691 (N_3691,N_3546,N_3485);
xnor U3692 (N_3692,N_3469,N_3477);
nand U3693 (N_3693,N_3510,N_3578);
nand U3694 (N_3694,N_3502,N_3555);
and U3695 (N_3695,N_3456,N_3586);
nor U3696 (N_3696,N_3453,N_3465);
xor U3697 (N_3697,N_3560,N_3598);
xnor U3698 (N_3698,N_3555,N_3463);
xor U3699 (N_3699,N_3553,N_3450);
xnor U3700 (N_3700,N_3588,N_3466);
or U3701 (N_3701,N_3593,N_3552);
nand U3702 (N_3702,N_3506,N_3593);
or U3703 (N_3703,N_3480,N_3595);
or U3704 (N_3704,N_3488,N_3489);
and U3705 (N_3705,N_3453,N_3578);
nor U3706 (N_3706,N_3576,N_3469);
nand U3707 (N_3707,N_3548,N_3455);
nor U3708 (N_3708,N_3583,N_3563);
and U3709 (N_3709,N_3500,N_3590);
nand U3710 (N_3710,N_3552,N_3530);
or U3711 (N_3711,N_3599,N_3580);
and U3712 (N_3712,N_3484,N_3526);
and U3713 (N_3713,N_3497,N_3491);
or U3714 (N_3714,N_3459,N_3494);
nand U3715 (N_3715,N_3560,N_3592);
and U3716 (N_3716,N_3538,N_3541);
nand U3717 (N_3717,N_3535,N_3489);
xor U3718 (N_3718,N_3515,N_3461);
and U3719 (N_3719,N_3471,N_3523);
nor U3720 (N_3720,N_3519,N_3511);
and U3721 (N_3721,N_3562,N_3591);
or U3722 (N_3722,N_3549,N_3595);
xnor U3723 (N_3723,N_3477,N_3513);
or U3724 (N_3724,N_3478,N_3539);
and U3725 (N_3725,N_3523,N_3464);
nor U3726 (N_3726,N_3591,N_3581);
nor U3727 (N_3727,N_3560,N_3588);
xor U3728 (N_3728,N_3560,N_3480);
and U3729 (N_3729,N_3568,N_3582);
xor U3730 (N_3730,N_3500,N_3501);
nand U3731 (N_3731,N_3569,N_3537);
or U3732 (N_3732,N_3548,N_3596);
or U3733 (N_3733,N_3584,N_3496);
nand U3734 (N_3734,N_3583,N_3492);
and U3735 (N_3735,N_3552,N_3482);
and U3736 (N_3736,N_3584,N_3559);
nand U3737 (N_3737,N_3489,N_3578);
xor U3738 (N_3738,N_3529,N_3577);
nand U3739 (N_3739,N_3510,N_3564);
and U3740 (N_3740,N_3554,N_3494);
xnor U3741 (N_3741,N_3528,N_3482);
nor U3742 (N_3742,N_3457,N_3467);
or U3743 (N_3743,N_3578,N_3467);
nor U3744 (N_3744,N_3588,N_3579);
nand U3745 (N_3745,N_3512,N_3504);
or U3746 (N_3746,N_3492,N_3479);
nor U3747 (N_3747,N_3565,N_3548);
and U3748 (N_3748,N_3486,N_3450);
nor U3749 (N_3749,N_3563,N_3541);
and U3750 (N_3750,N_3624,N_3601);
nand U3751 (N_3751,N_3659,N_3635);
and U3752 (N_3752,N_3608,N_3676);
nor U3753 (N_3753,N_3725,N_3696);
xnor U3754 (N_3754,N_3654,N_3611);
nand U3755 (N_3755,N_3678,N_3629);
nand U3756 (N_3756,N_3721,N_3717);
and U3757 (N_3757,N_3685,N_3726);
nand U3758 (N_3758,N_3609,N_3620);
xnor U3759 (N_3759,N_3748,N_3680);
or U3760 (N_3760,N_3708,N_3677);
nand U3761 (N_3761,N_3715,N_3667);
xnor U3762 (N_3762,N_3714,N_3710);
or U3763 (N_3763,N_3622,N_3655);
or U3764 (N_3764,N_3692,N_3687);
xnor U3765 (N_3765,N_3604,N_3602);
nand U3766 (N_3766,N_3630,N_3631);
xnor U3767 (N_3767,N_3665,N_3746);
and U3768 (N_3768,N_3724,N_3691);
or U3769 (N_3769,N_3645,N_3713);
nor U3770 (N_3770,N_3640,N_3606);
nor U3771 (N_3771,N_3628,N_3623);
or U3772 (N_3772,N_3730,N_3682);
xor U3773 (N_3773,N_3657,N_3658);
and U3774 (N_3774,N_3668,N_3605);
and U3775 (N_3775,N_3613,N_3743);
nand U3776 (N_3776,N_3663,N_3625);
or U3777 (N_3777,N_3664,N_3650);
and U3778 (N_3778,N_3643,N_3616);
nor U3779 (N_3779,N_3637,N_3711);
or U3780 (N_3780,N_3626,N_3722);
or U3781 (N_3781,N_3669,N_3690);
xnor U3782 (N_3782,N_3614,N_3633);
or U3783 (N_3783,N_3706,N_3653);
nor U3784 (N_3784,N_3749,N_3707);
and U3785 (N_3785,N_3673,N_3745);
xnor U3786 (N_3786,N_3694,N_3652);
nor U3787 (N_3787,N_3686,N_3612);
and U3788 (N_3788,N_3693,N_3709);
and U3789 (N_3789,N_3732,N_3720);
and U3790 (N_3790,N_3660,N_3747);
nor U3791 (N_3791,N_3716,N_3639);
nand U3792 (N_3792,N_3671,N_3644);
nor U3793 (N_3793,N_3619,N_3674);
xor U3794 (N_3794,N_3675,N_3603);
or U3795 (N_3795,N_3649,N_3607);
and U3796 (N_3796,N_3742,N_3723);
or U3797 (N_3797,N_3627,N_3734);
xnor U3798 (N_3798,N_3684,N_3672);
nand U3799 (N_3799,N_3615,N_3646);
or U3800 (N_3800,N_3700,N_3718);
nor U3801 (N_3801,N_3728,N_3698);
and U3802 (N_3802,N_3704,N_3705);
nand U3803 (N_3803,N_3648,N_3699);
nand U3804 (N_3804,N_3632,N_3712);
and U3805 (N_3805,N_3679,N_3642);
nand U3806 (N_3806,N_3736,N_3670);
or U3807 (N_3807,N_3727,N_3740);
or U3808 (N_3808,N_3610,N_3731);
xor U3809 (N_3809,N_3733,N_3738);
xnor U3810 (N_3810,N_3741,N_3737);
or U3811 (N_3811,N_3636,N_3600);
xnor U3812 (N_3812,N_3617,N_3621);
nor U3813 (N_3813,N_3744,N_3647);
and U3814 (N_3814,N_3662,N_3735);
nor U3815 (N_3815,N_3651,N_3666);
or U3816 (N_3816,N_3702,N_3634);
nor U3817 (N_3817,N_3681,N_3701);
nor U3818 (N_3818,N_3739,N_3641);
or U3819 (N_3819,N_3688,N_3689);
nand U3820 (N_3820,N_3683,N_3656);
and U3821 (N_3821,N_3719,N_3661);
xnor U3822 (N_3822,N_3618,N_3695);
nor U3823 (N_3823,N_3729,N_3703);
xnor U3824 (N_3824,N_3638,N_3697);
nor U3825 (N_3825,N_3718,N_3665);
nand U3826 (N_3826,N_3636,N_3604);
and U3827 (N_3827,N_3733,N_3647);
and U3828 (N_3828,N_3605,N_3661);
nand U3829 (N_3829,N_3674,N_3606);
or U3830 (N_3830,N_3714,N_3729);
nand U3831 (N_3831,N_3666,N_3715);
and U3832 (N_3832,N_3673,N_3699);
nor U3833 (N_3833,N_3605,N_3601);
nor U3834 (N_3834,N_3682,N_3697);
or U3835 (N_3835,N_3662,N_3701);
and U3836 (N_3836,N_3729,N_3682);
nor U3837 (N_3837,N_3661,N_3705);
and U3838 (N_3838,N_3606,N_3727);
nand U3839 (N_3839,N_3688,N_3666);
or U3840 (N_3840,N_3612,N_3658);
and U3841 (N_3841,N_3710,N_3630);
or U3842 (N_3842,N_3619,N_3616);
and U3843 (N_3843,N_3735,N_3695);
xor U3844 (N_3844,N_3699,N_3608);
nor U3845 (N_3845,N_3646,N_3634);
or U3846 (N_3846,N_3700,N_3652);
nand U3847 (N_3847,N_3641,N_3658);
and U3848 (N_3848,N_3615,N_3696);
and U3849 (N_3849,N_3644,N_3725);
xnor U3850 (N_3850,N_3684,N_3627);
nor U3851 (N_3851,N_3679,N_3688);
nand U3852 (N_3852,N_3671,N_3652);
xnor U3853 (N_3853,N_3747,N_3693);
nor U3854 (N_3854,N_3702,N_3612);
nand U3855 (N_3855,N_3662,N_3697);
nand U3856 (N_3856,N_3689,N_3707);
xor U3857 (N_3857,N_3740,N_3688);
or U3858 (N_3858,N_3741,N_3605);
xor U3859 (N_3859,N_3605,N_3720);
xor U3860 (N_3860,N_3645,N_3718);
nand U3861 (N_3861,N_3632,N_3635);
and U3862 (N_3862,N_3740,N_3665);
xnor U3863 (N_3863,N_3739,N_3639);
or U3864 (N_3864,N_3647,N_3644);
and U3865 (N_3865,N_3684,N_3660);
nor U3866 (N_3866,N_3646,N_3719);
or U3867 (N_3867,N_3657,N_3616);
and U3868 (N_3868,N_3706,N_3723);
nor U3869 (N_3869,N_3697,N_3725);
and U3870 (N_3870,N_3653,N_3690);
and U3871 (N_3871,N_3685,N_3612);
and U3872 (N_3872,N_3735,N_3671);
and U3873 (N_3873,N_3681,N_3678);
nor U3874 (N_3874,N_3614,N_3680);
xnor U3875 (N_3875,N_3657,N_3738);
and U3876 (N_3876,N_3610,N_3694);
and U3877 (N_3877,N_3688,N_3746);
and U3878 (N_3878,N_3605,N_3637);
xnor U3879 (N_3879,N_3689,N_3645);
nor U3880 (N_3880,N_3641,N_3616);
and U3881 (N_3881,N_3602,N_3601);
nand U3882 (N_3882,N_3707,N_3634);
xnor U3883 (N_3883,N_3652,N_3609);
nand U3884 (N_3884,N_3612,N_3735);
xnor U3885 (N_3885,N_3638,N_3635);
and U3886 (N_3886,N_3700,N_3645);
or U3887 (N_3887,N_3721,N_3697);
nor U3888 (N_3888,N_3622,N_3709);
or U3889 (N_3889,N_3670,N_3649);
xor U3890 (N_3890,N_3655,N_3680);
or U3891 (N_3891,N_3648,N_3743);
and U3892 (N_3892,N_3642,N_3601);
nand U3893 (N_3893,N_3718,N_3671);
or U3894 (N_3894,N_3749,N_3647);
nand U3895 (N_3895,N_3646,N_3675);
or U3896 (N_3896,N_3674,N_3657);
or U3897 (N_3897,N_3628,N_3690);
xor U3898 (N_3898,N_3728,N_3615);
nor U3899 (N_3899,N_3704,N_3659);
or U3900 (N_3900,N_3861,N_3863);
and U3901 (N_3901,N_3871,N_3896);
or U3902 (N_3902,N_3857,N_3840);
xor U3903 (N_3903,N_3800,N_3845);
nand U3904 (N_3904,N_3773,N_3842);
and U3905 (N_3905,N_3819,N_3843);
or U3906 (N_3906,N_3841,N_3855);
and U3907 (N_3907,N_3898,N_3897);
or U3908 (N_3908,N_3880,N_3883);
xnor U3909 (N_3909,N_3776,N_3766);
or U3910 (N_3910,N_3762,N_3849);
nand U3911 (N_3911,N_3780,N_3879);
xor U3912 (N_3912,N_3852,N_3866);
nor U3913 (N_3913,N_3836,N_3789);
nor U3914 (N_3914,N_3752,N_3761);
nor U3915 (N_3915,N_3893,N_3763);
and U3916 (N_3916,N_3755,N_3760);
xor U3917 (N_3917,N_3796,N_3869);
nor U3918 (N_3918,N_3881,N_3826);
or U3919 (N_3919,N_3811,N_3782);
or U3920 (N_3920,N_3794,N_3848);
and U3921 (N_3921,N_3859,N_3805);
nor U3922 (N_3922,N_3781,N_3793);
nand U3923 (N_3923,N_3851,N_3778);
xnor U3924 (N_3924,N_3830,N_3885);
and U3925 (N_3925,N_3801,N_3816);
nand U3926 (N_3926,N_3838,N_3821);
and U3927 (N_3927,N_3825,N_3813);
and U3928 (N_3928,N_3812,N_3783);
nand U3929 (N_3929,N_3798,N_3853);
nand U3930 (N_3930,N_3847,N_3768);
xor U3931 (N_3931,N_3809,N_3831);
nand U3932 (N_3932,N_3772,N_3829);
or U3933 (N_3933,N_3788,N_3799);
nand U3934 (N_3934,N_3784,N_3822);
nor U3935 (N_3935,N_3758,N_3786);
nand U3936 (N_3936,N_3834,N_3878);
or U3937 (N_3937,N_3876,N_3790);
nor U3938 (N_3938,N_3895,N_3894);
or U3939 (N_3939,N_3808,N_3804);
and U3940 (N_3940,N_3774,N_3815);
or U3941 (N_3941,N_3820,N_3806);
nor U3942 (N_3942,N_3884,N_3846);
or U3943 (N_3943,N_3810,N_3817);
nor U3944 (N_3944,N_3889,N_3890);
xnor U3945 (N_3945,N_3888,N_3837);
or U3946 (N_3946,N_3899,N_3814);
or U3947 (N_3947,N_3870,N_3865);
and U3948 (N_3948,N_3795,N_3751);
xnor U3949 (N_3949,N_3777,N_3892);
or U3950 (N_3950,N_3860,N_3858);
or U3951 (N_3951,N_3791,N_3792);
xor U3952 (N_3952,N_3854,N_3770);
nor U3953 (N_3953,N_3807,N_3891);
xnor U3954 (N_3954,N_3864,N_3818);
nor U3955 (N_3955,N_3824,N_3832);
xnor U3956 (N_3956,N_3839,N_3756);
or U3957 (N_3957,N_3844,N_3887);
and U3958 (N_3958,N_3771,N_3872);
and U3959 (N_3959,N_3750,N_3764);
nand U3960 (N_3960,N_3875,N_3850);
nor U3961 (N_3961,N_3828,N_3787);
nand U3962 (N_3962,N_3874,N_3797);
nand U3963 (N_3963,N_3779,N_3823);
and U3964 (N_3964,N_3868,N_3856);
nand U3965 (N_3965,N_3757,N_3882);
nand U3966 (N_3966,N_3886,N_3862);
nand U3967 (N_3967,N_3785,N_3867);
nand U3968 (N_3968,N_3775,N_3759);
or U3969 (N_3969,N_3753,N_3754);
nor U3970 (N_3970,N_3835,N_3769);
and U3971 (N_3971,N_3803,N_3833);
nand U3972 (N_3972,N_3767,N_3802);
and U3973 (N_3973,N_3877,N_3873);
nor U3974 (N_3974,N_3827,N_3765);
and U3975 (N_3975,N_3794,N_3837);
or U3976 (N_3976,N_3821,N_3812);
or U3977 (N_3977,N_3752,N_3807);
nand U3978 (N_3978,N_3896,N_3899);
or U3979 (N_3979,N_3799,N_3839);
or U3980 (N_3980,N_3849,N_3876);
nand U3981 (N_3981,N_3793,N_3792);
and U3982 (N_3982,N_3898,N_3769);
and U3983 (N_3983,N_3890,N_3836);
xor U3984 (N_3984,N_3835,N_3813);
xnor U3985 (N_3985,N_3856,N_3870);
nor U3986 (N_3986,N_3782,N_3898);
nand U3987 (N_3987,N_3825,N_3839);
nand U3988 (N_3988,N_3824,N_3884);
xnor U3989 (N_3989,N_3880,N_3806);
xnor U3990 (N_3990,N_3804,N_3793);
and U3991 (N_3991,N_3886,N_3870);
or U3992 (N_3992,N_3805,N_3754);
or U3993 (N_3993,N_3862,N_3813);
xor U3994 (N_3994,N_3819,N_3800);
xnor U3995 (N_3995,N_3776,N_3774);
and U3996 (N_3996,N_3786,N_3800);
and U3997 (N_3997,N_3809,N_3846);
or U3998 (N_3998,N_3884,N_3803);
and U3999 (N_3999,N_3897,N_3886);
and U4000 (N_4000,N_3857,N_3873);
nand U4001 (N_4001,N_3898,N_3873);
nor U4002 (N_4002,N_3759,N_3895);
nor U4003 (N_4003,N_3863,N_3784);
nor U4004 (N_4004,N_3798,N_3780);
nand U4005 (N_4005,N_3860,N_3816);
xnor U4006 (N_4006,N_3759,N_3879);
nor U4007 (N_4007,N_3833,N_3812);
and U4008 (N_4008,N_3798,N_3808);
nand U4009 (N_4009,N_3832,N_3780);
xnor U4010 (N_4010,N_3774,N_3809);
or U4011 (N_4011,N_3841,N_3879);
nand U4012 (N_4012,N_3823,N_3887);
nand U4013 (N_4013,N_3872,N_3750);
nor U4014 (N_4014,N_3794,N_3858);
or U4015 (N_4015,N_3789,N_3870);
xor U4016 (N_4016,N_3796,N_3772);
nand U4017 (N_4017,N_3835,N_3782);
or U4018 (N_4018,N_3842,N_3881);
and U4019 (N_4019,N_3789,N_3883);
xnor U4020 (N_4020,N_3804,N_3882);
and U4021 (N_4021,N_3773,N_3752);
or U4022 (N_4022,N_3750,N_3893);
nand U4023 (N_4023,N_3782,N_3874);
nor U4024 (N_4024,N_3858,N_3799);
and U4025 (N_4025,N_3884,N_3856);
xnor U4026 (N_4026,N_3813,N_3778);
or U4027 (N_4027,N_3770,N_3845);
or U4028 (N_4028,N_3843,N_3875);
and U4029 (N_4029,N_3820,N_3772);
and U4030 (N_4030,N_3889,N_3851);
and U4031 (N_4031,N_3856,N_3887);
nor U4032 (N_4032,N_3770,N_3844);
nor U4033 (N_4033,N_3769,N_3863);
and U4034 (N_4034,N_3764,N_3766);
and U4035 (N_4035,N_3899,N_3877);
or U4036 (N_4036,N_3877,N_3897);
or U4037 (N_4037,N_3782,N_3880);
nor U4038 (N_4038,N_3751,N_3808);
nand U4039 (N_4039,N_3886,N_3765);
nand U4040 (N_4040,N_3761,N_3791);
nand U4041 (N_4041,N_3887,N_3795);
nand U4042 (N_4042,N_3764,N_3790);
xor U4043 (N_4043,N_3875,N_3837);
or U4044 (N_4044,N_3760,N_3859);
xnor U4045 (N_4045,N_3820,N_3777);
or U4046 (N_4046,N_3827,N_3866);
nand U4047 (N_4047,N_3851,N_3818);
xor U4048 (N_4048,N_3856,N_3753);
xor U4049 (N_4049,N_3774,N_3800);
nor U4050 (N_4050,N_3950,N_3983);
nand U4051 (N_4051,N_4025,N_4017);
xor U4052 (N_4052,N_3997,N_3968);
and U4053 (N_4053,N_4028,N_3921);
xnor U4054 (N_4054,N_3916,N_4000);
nand U4055 (N_4055,N_4019,N_4034);
nor U4056 (N_4056,N_4032,N_3977);
and U4057 (N_4057,N_4040,N_3938);
nand U4058 (N_4058,N_3984,N_3973);
or U4059 (N_4059,N_3939,N_3962);
or U4060 (N_4060,N_3904,N_4003);
xor U4061 (N_4061,N_3918,N_3937);
xnor U4062 (N_4062,N_3985,N_3947);
nor U4063 (N_4063,N_3945,N_4024);
or U4064 (N_4064,N_4033,N_3948);
or U4065 (N_4065,N_4011,N_3999);
xor U4066 (N_4066,N_3978,N_3920);
xor U4067 (N_4067,N_3987,N_3993);
nor U4068 (N_4068,N_3908,N_3955);
nand U4069 (N_4069,N_4037,N_3942);
nand U4070 (N_4070,N_3946,N_3956);
nor U4071 (N_4071,N_4029,N_3917);
nand U4072 (N_4072,N_3992,N_3923);
nor U4073 (N_4073,N_3924,N_3915);
or U4074 (N_4074,N_3912,N_3965);
and U4075 (N_4075,N_4031,N_4016);
and U4076 (N_4076,N_3951,N_3905);
nand U4077 (N_4077,N_4012,N_4046);
nand U4078 (N_4078,N_4022,N_4035);
nand U4079 (N_4079,N_3922,N_3909);
or U4080 (N_4080,N_4018,N_3961);
xor U4081 (N_4081,N_3996,N_3903);
nor U4082 (N_4082,N_3925,N_4036);
xnor U4083 (N_4083,N_3991,N_3998);
or U4084 (N_4084,N_3927,N_4030);
nor U4085 (N_4085,N_4044,N_4045);
or U4086 (N_4086,N_3953,N_3960);
or U4087 (N_4087,N_3952,N_4013);
nand U4088 (N_4088,N_3976,N_3926);
xor U4089 (N_4089,N_3994,N_4047);
xor U4090 (N_4090,N_3936,N_4038);
nor U4091 (N_4091,N_3981,N_3906);
nand U4092 (N_4092,N_3974,N_3967);
and U4093 (N_4093,N_3958,N_3929);
and U4094 (N_4094,N_3910,N_3944);
xor U4095 (N_4095,N_4004,N_3982);
nor U4096 (N_4096,N_4001,N_3986);
and U4097 (N_4097,N_3988,N_4014);
nand U4098 (N_4098,N_3959,N_4015);
nand U4099 (N_4099,N_4042,N_3954);
or U4100 (N_4100,N_3930,N_3932);
nor U4101 (N_4101,N_3995,N_4002);
nand U4102 (N_4102,N_4005,N_4007);
or U4103 (N_4103,N_3949,N_3931);
nor U4104 (N_4104,N_4023,N_4041);
and U4105 (N_4105,N_3940,N_3919);
nor U4106 (N_4106,N_3941,N_3902);
and U4107 (N_4107,N_3989,N_4048);
xor U4108 (N_4108,N_3911,N_4039);
or U4109 (N_4109,N_3900,N_3966);
and U4110 (N_4110,N_3934,N_3907);
xnor U4111 (N_4111,N_3971,N_3933);
nand U4112 (N_4112,N_4010,N_3980);
and U4113 (N_4113,N_4021,N_3970);
or U4114 (N_4114,N_4043,N_4026);
nand U4115 (N_4115,N_3979,N_4020);
xnor U4116 (N_4116,N_3969,N_3914);
nand U4117 (N_4117,N_3957,N_4009);
nand U4118 (N_4118,N_4049,N_3935);
nand U4119 (N_4119,N_3943,N_4006);
nor U4120 (N_4120,N_3928,N_3964);
nor U4121 (N_4121,N_3913,N_4008);
nor U4122 (N_4122,N_3901,N_4027);
xor U4123 (N_4123,N_3990,N_3975);
or U4124 (N_4124,N_3972,N_3963);
and U4125 (N_4125,N_3970,N_3944);
and U4126 (N_4126,N_3960,N_3989);
nor U4127 (N_4127,N_3953,N_3904);
nand U4128 (N_4128,N_3912,N_4023);
nor U4129 (N_4129,N_4021,N_3975);
nand U4130 (N_4130,N_3914,N_3965);
nand U4131 (N_4131,N_3907,N_3953);
nand U4132 (N_4132,N_3940,N_4031);
xor U4133 (N_4133,N_3976,N_3984);
and U4134 (N_4134,N_4002,N_3913);
xor U4135 (N_4135,N_3907,N_3984);
or U4136 (N_4136,N_3972,N_3993);
nand U4137 (N_4137,N_3947,N_4034);
nor U4138 (N_4138,N_3966,N_3983);
or U4139 (N_4139,N_3945,N_4002);
nand U4140 (N_4140,N_3929,N_3959);
and U4141 (N_4141,N_4037,N_3922);
nand U4142 (N_4142,N_4039,N_3998);
nand U4143 (N_4143,N_3943,N_3945);
xnor U4144 (N_4144,N_3973,N_4003);
nand U4145 (N_4145,N_4013,N_3973);
and U4146 (N_4146,N_3958,N_3902);
and U4147 (N_4147,N_3950,N_3951);
nand U4148 (N_4148,N_3916,N_3993);
xor U4149 (N_4149,N_3915,N_3906);
or U4150 (N_4150,N_3967,N_3919);
xor U4151 (N_4151,N_3995,N_3964);
nor U4152 (N_4152,N_4002,N_3977);
nand U4153 (N_4153,N_4033,N_3966);
nand U4154 (N_4154,N_3925,N_4021);
nand U4155 (N_4155,N_4004,N_3988);
nand U4156 (N_4156,N_3956,N_4011);
xor U4157 (N_4157,N_4032,N_4033);
nand U4158 (N_4158,N_3973,N_3930);
or U4159 (N_4159,N_3946,N_3943);
nor U4160 (N_4160,N_4036,N_3996);
nand U4161 (N_4161,N_3920,N_3935);
or U4162 (N_4162,N_3983,N_4029);
or U4163 (N_4163,N_3973,N_3913);
nor U4164 (N_4164,N_4027,N_4029);
xnor U4165 (N_4165,N_3911,N_3978);
xnor U4166 (N_4166,N_4027,N_3955);
and U4167 (N_4167,N_3973,N_4025);
nand U4168 (N_4168,N_4027,N_3919);
nand U4169 (N_4169,N_3999,N_4012);
and U4170 (N_4170,N_3940,N_3929);
or U4171 (N_4171,N_4007,N_3997);
xor U4172 (N_4172,N_3996,N_4009);
or U4173 (N_4173,N_3988,N_3993);
nor U4174 (N_4174,N_4019,N_3912);
xor U4175 (N_4175,N_3982,N_3992);
xnor U4176 (N_4176,N_3905,N_3910);
nand U4177 (N_4177,N_3997,N_3907);
and U4178 (N_4178,N_4044,N_4010);
nand U4179 (N_4179,N_3911,N_3970);
or U4180 (N_4180,N_3908,N_3978);
xnor U4181 (N_4181,N_3931,N_4004);
and U4182 (N_4182,N_3992,N_4025);
or U4183 (N_4183,N_4026,N_3920);
xnor U4184 (N_4184,N_4007,N_4041);
and U4185 (N_4185,N_3910,N_3929);
nor U4186 (N_4186,N_3946,N_3986);
nor U4187 (N_4187,N_4029,N_3902);
and U4188 (N_4188,N_4048,N_3905);
and U4189 (N_4189,N_3967,N_3938);
or U4190 (N_4190,N_4031,N_3984);
nor U4191 (N_4191,N_3941,N_3904);
and U4192 (N_4192,N_4043,N_4012);
nor U4193 (N_4193,N_3974,N_3928);
nand U4194 (N_4194,N_4008,N_3910);
nor U4195 (N_4195,N_3951,N_3988);
and U4196 (N_4196,N_3935,N_4018);
nand U4197 (N_4197,N_3980,N_3945);
or U4198 (N_4198,N_3979,N_3941);
nor U4199 (N_4199,N_4015,N_4008);
or U4200 (N_4200,N_4120,N_4054);
or U4201 (N_4201,N_4177,N_4088);
nand U4202 (N_4202,N_4076,N_4194);
nand U4203 (N_4203,N_4119,N_4132);
and U4204 (N_4204,N_4199,N_4189);
nand U4205 (N_4205,N_4158,N_4106);
nor U4206 (N_4206,N_4184,N_4197);
or U4207 (N_4207,N_4053,N_4138);
and U4208 (N_4208,N_4107,N_4142);
or U4209 (N_4209,N_4080,N_4090);
nand U4210 (N_4210,N_4069,N_4172);
and U4211 (N_4211,N_4055,N_4061);
xnor U4212 (N_4212,N_4124,N_4081);
xor U4213 (N_4213,N_4178,N_4133);
xor U4214 (N_4214,N_4166,N_4185);
nand U4215 (N_4215,N_4131,N_4195);
nand U4216 (N_4216,N_4099,N_4072);
xnor U4217 (N_4217,N_4078,N_4058);
or U4218 (N_4218,N_4174,N_4187);
nor U4219 (N_4219,N_4112,N_4063);
nand U4220 (N_4220,N_4176,N_4074);
nor U4221 (N_4221,N_4051,N_4162);
nand U4222 (N_4222,N_4159,N_4192);
nand U4223 (N_4223,N_4102,N_4059);
or U4224 (N_4224,N_4136,N_4079);
or U4225 (N_4225,N_4151,N_4121);
or U4226 (N_4226,N_4156,N_4104);
nand U4227 (N_4227,N_4070,N_4164);
and U4228 (N_4228,N_4165,N_4064);
and U4229 (N_4229,N_4157,N_4052);
and U4230 (N_4230,N_4186,N_4170);
nand U4231 (N_4231,N_4116,N_4188);
and U4232 (N_4232,N_4193,N_4179);
or U4233 (N_4233,N_4180,N_4089);
nor U4234 (N_4234,N_4075,N_4113);
or U4235 (N_4235,N_4163,N_4128);
or U4236 (N_4236,N_4153,N_4182);
xnor U4237 (N_4237,N_4095,N_4082);
nor U4238 (N_4238,N_4169,N_4139);
nor U4239 (N_4239,N_4065,N_4160);
nand U4240 (N_4240,N_4198,N_4145);
nor U4241 (N_4241,N_4127,N_4083);
nand U4242 (N_4242,N_4050,N_4130);
or U4243 (N_4243,N_4115,N_4111);
and U4244 (N_4244,N_4126,N_4062);
xor U4245 (N_4245,N_4068,N_4161);
nand U4246 (N_4246,N_4150,N_4167);
xor U4247 (N_4247,N_4143,N_4109);
xnor U4248 (N_4248,N_4141,N_4093);
nor U4249 (N_4249,N_4097,N_4190);
or U4250 (N_4250,N_4085,N_4096);
and U4251 (N_4251,N_4173,N_4129);
xnor U4252 (N_4252,N_4086,N_4066);
or U4253 (N_4253,N_4149,N_4117);
nand U4254 (N_4254,N_4137,N_4060);
nor U4255 (N_4255,N_4110,N_4168);
nand U4256 (N_4256,N_4057,N_4123);
or U4257 (N_4257,N_4100,N_4067);
nand U4258 (N_4258,N_4144,N_4175);
nor U4259 (N_4259,N_4071,N_4148);
xnor U4260 (N_4260,N_4098,N_4125);
nor U4261 (N_4261,N_4103,N_4114);
nor U4262 (N_4262,N_4118,N_4140);
xnor U4263 (N_4263,N_4108,N_4101);
and U4264 (N_4264,N_4147,N_4196);
nand U4265 (N_4265,N_4171,N_4084);
nor U4266 (N_4266,N_4154,N_4094);
or U4267 (N_4267,N_4073,N_4092);
xor U4268 (N_4268,N_4155,N_4105);
nor U4269 (N_4269,N_4191,N_4087);
xnor U4270 (N_4270,N_4056,N_4181);
xnor U4271 (N_4271,N_4091,N_4077);
and U4272 (N_4272,N_4183,N_4146);
nand U4273 (N_4273,N_4134,N_4135);
nand U4274 (N_4274,N_4122,N_4152);
nor U4275 (N_4275,N_4092,N_4170);
nand U4276 (N_4276,N_4062,N_4089);
nand U4277 (N_4277,N_4148,N_4194);
or U4278 (N_4278,N_4196,N_4158);
nand U4279 (N_4279,N_4173,N_4150);
or U4280 (N_4280,N_4060,N_4124);
or U4281 (N_4281,N_4123,N_4175);
xor U4282 (N_4282,N_4084,N_4132);
and U4283 (N_4283,N_4102,N_4161);
or U4284 (N_4284,N_4178,N_4082);
xnor U4285 (N_4285,N_4086,N_4160);
xor U4286 (N_4286,N_4174,N_4135);
nand U4287 (N_4287,N_4136,N_4174);
nor U4288 (N_4288,N_4160,N_4087);
nand U4289 (N_4289,N_4189,N_4050);
and U4290 (N_4290,N_4191,N_4193);
nor U4291 (N_4291,N_4181,N_4176);
or U4292 (N_4292,N_4084,N_4193);
nor U4293 (N_4293,N_4185,N_4190);
or U4294 (N_4294,N_4177,N_4073);
xnor U4295 (N_4295,N_4064,N_4118);
nor U4296 (N_4296,N_4126,N_4079);
xor U4297 (N_4297,N_4084,N_4074);
nand U4298 (N_4298,N_4163,N_4132);
nor U4299 (N_4299,N_4101,N_4122);
and U4300 (N_4300,N_4179,N_4078);
or U4301 (N_4301,N_4146,N_4191);
nand U4302 (N_4302,N_4196,N_4095);
or U4303 (N_4303,N_4107,N_4191);
or U4304 (N_4304,N_4138,N_4142);
nor U4305 (N_4305,N_4056,N_4053);
nand U4306 (N_4306,N_4118,N_4090);
nand U4307 (N_4307,N_4169,N_4140);
nand U4308 (N_4308,N_4113,N_4157);
nor U4309 (N_4309,N_4085,N_4174);
nor U4310 (N_4310,N_4109,N_4089);
nand U4311 (N_4311,N_4100,N_4098);
xor U4312 (N_4312,N_4165,N_4166);
nand U4313 (N_4313,N_4187,N_4150);
nor U4314 (N_4314,N_4083,N_4163);
and U4315 (N_4315,N_4076,N_4147);
nand U4316 (N_4316,N_4131,N_4079);
nand U4317 (N_4317,N_4076,N_4173);
xnor U4318 (N_4318,N_4162,N_4083);
and U4319 (N_4319,N_4169,N_4160);
xnor U4320 (N_4320,N_4159,N_4058);
xor U4321 (N_4321,N_4185,N_4088);
or U4322 (N_4322,N_4195,N_4156);
and U4323 (N_4323,N_4074,N_4101);
nand U4324 (N_4324,N_4050,N_4112);
nand U4325 (N_4325,N_4106,N_4097);
nor U4326 (N_4326,N_4184,N_4088);
or U4327 (N_4327,N_4066,N_4181);
or U4328 (N_4328,N_4171,N_4102);
or U4329 (N_4329,N_4150,N_4102);
or U4330 (N_4330,N_4069,N_4174);
nand U4331 (N_4331,N_4150,N_4125);
nand U4332 (N_4332,N_4156,N_4105);
nand U4333 (N_4333,N_4068,N_4073);
xnor U4334 (N_4334,N_4064,N_4147);
nor U4335 (N_4335,N_4186,N_4177);
xor U4336 (N_4336,N_4070,N_4191);
and U4337 (N_4337,N_4191,N_4109);
nand U4338 (N_4338,N_4141,N_4106);
or U4339 (N_4339,N_4115,N_4127);
or U4340 (N_4340,N_4076,N_4050);
xor U4341 (N_4341,N_4055,N_4181);
and U4342 (N_4342,N_4126,N_4113);
nor U4343 (N_4343,N_4161,N_4058);
nand U4344 (N_4344,N_4085,N_4067);
nor U4345 (N_4345,N_4179,N_4124);
xnor U4346 (N_4346,N_4146,N_4156);
and U4347 (N_4347,N_4104,N_4077);
or U4348 (N_4348,N_4127,N_4186);
or U4349 (N_4349,N_4105,N_4107);
xor U4350 (N_4350,N_4218,N_4217);
and U4351 (N_4351,N_4283,N_4289);
nor U4352 (N_4352,N_4339,N_4298);
or U4353 (N_4353,N_4277,N_4315);
xnor U4354 (N_4354,N_4320,N_4331);
nor U4355 (N_4355,N_4286,N_4343);
xor U4356 (N_4356,N_4338,N_4318);
nor U4357 (N_4357,N_4221,N_4346);
nor U4358 (N_4358,N_4275,N_4208);
and U4359 (N_4359,N_4235,N_4348);
and U4360 (N_4360,N_4322,N_4333);
xnor U4361 (N_4361,N_4269,N_4266);
nor U4362 (N_4362,N_4213,N_4259);
and U4363 (N_4363,N_4291,N_4206);
and U4364 (N_4364,N_4345,N_4327);
or U4365 (N_4365,N_4223,N_4272);
nor U4366 (N_4366,N_4230,N_4232);
or U4367 (N_4367,N_4287,N_4212);
nand U4368 (N_4368,N_4281,N_4317);
xnor U4369 (N_4369,N_4246,N_4226);
nand U4370 (N_4370,N_4216,N_4313);
xnor U4371 (N_4371,N_4279,N_4271);
nor U4372 (N_4372,N_4285,N_4200);
or U4373 (N_4373,N_4202,N_4326);
nor U4374 (N_4374,N_4300,N_4260);
and U4375 (N_4375,N_4311,N_4301);
nor U4376 (N_4376,N_4342,N_4314);
or U4377 (N_4377,N_4270,N_4236);
xnor U4378 (N_4378,N_4328,N_4267);
or U4379 (N_4379,N_4250,N_4316);
xor U4380 (N_4380,N_4253,N_4290);
nor U4381 (N_4381,N_4214,N_4280);
nand U4382 (N_4382,N_4302,N_4288);
or U4383 (N_4383,N_4325,N_4274);
nor U4384 (N_4384,N_4305,N_4349);
nand U4385 (N_4385,N_4244,N_4263);
nor U4386 (N_4386,N_4207,N_4304);
and U4387 (N_4387,N_4215,N_4347);
nand U4388 (N_4388,N_4310,N_4340);
nor U4389 (N_4389,N_4255,N_4324);
nor U4390 (N_4390,N_4257,N_4252);
xnor U4391 (N_4391,N_4262,N_4341);
or U4392 (N_4392,N_4224,N_4335);
nand U4393 (N_4393,N_4323,N_4231);
and U4394 (N_4394,N_4222,N_4303);
nand U4395 (N_4395,N_4309,N_4306);
nor U4396 (N_4396,N_4233,N_4220);
or U4397 (N_4397,N_4241,N_4209);
and U4398 (N_4398,N_4293,N_4243);
or U4399 (N_4399,N_4295,N_4261);
nand U4400 (N_4400,N_4312,N_4227);
or U4401 (N_4401,N_4219,N_4268);
xnor U4402 (N_4402,N_4332,N_4296);
and U4403 (N_4403,N_4211,N_4284);
nand U4404 (N_4404,N_4204,N_4201);
xor U4405 (N_4405,N_4264,N_4245);
xnor U4406 (N_4406,N_4321,N_4234);
nor U4407 (N_4407,N_4247,N_4334);
or U4408 (N_4408,N_4308,N_4265);
xnor U4409 (N_4409,N_4210,N_4344);
xor U4410 (N_4410,N_4249,N_4251);
nand U4411 (N_4411,N_4254,N_4242);
and U4412 (N_4412,N_4239,N_4237);
and U4413 (N_4413,N_4276,N_4278);
xnor U4414 (N_4414,N_4225,N_4299);
and U4415 (N_4415,N_4248,N_4297);
xnor U4416 (N_4416,N_4336,N_4329);
or U4417 (N_4417,N_4228,N_4238);
nand U4418 (N_4418,N_4203,N_4292);
nand U4419 (N_4419,N_4273,N_4337);
xnor U4420 (N_4420,N_4282,N_4307);
xor U4421 (N_4421,N_4205,N_4229);
nor U4422 (N_4422,N_4319,N_4330);
nor U4423 (N_4423,N_4258,N_4256);
nand U4424 (N_4424,N_4240,N_4294);
or U4425 (N_4425,N_4271,N_4319);
nand U4426 (N_4426,N_4237,N_4235);
or U4427 (N_4427,N_4342,N_4209);
or U4428 (N_4428,N_4213,N_4338);
and U4429 (N_4429,N_4313,N_4270);
nor U4430 (N_4430,N_4263,N_4333);
and U4431 (N_4431,N_4220,N_4329);
nand U4432 (N_4432,N_4247,N_4327);
and U4433 (N_4433,N_4243,N_4227);
nand U4434 (N_4434,N_4347,N_4283);
xor U4435 (N_4435,N_4296,N_4333);
and U4436 (N_4436,N_4239,N_4215);
nor U4437 (N_4437,N_4329,N_4240);
or U4438 (N_4438,N_4342,N_4302);
and U4439 (N_4439,N_4342,N_4250);
xor U4440 (N_4440,N_4345,N_4263);
xnor U4441 (N_4441,N_4292,N_4334);
and U4442 (N_4442,N_4237,N_4260);
or U4443 (N_4443,N_4216,N_4314);
and U4444 (N_4444,N_4290,N_4339);
xor U4445 (N_4445,N_4257,N_4304);
and U4446 (N_4446,N_4216,N_4291);
nand U4447 (N_4447,N_4252,N_4344);
and U4448 (N_4448,N_4332,N_4343);
xor U4449 (N_4449,N_4241,N_4240);
and U4450 (N_4450,N_4340,N_4255);
nor U4451 (N_4451,N_4201,N_4299);
nor U4452 (N_4452,N_4225,N_4342);
xnor U4453 (N_4453,N_4329,N_4303);
xor U4454 (N_4454,N_4313,N_4294);
nand U4455 (N_4455,N_4247,N_4314);
nor U4456 (N_4456,N_4231,N_4311);
or U4457 (N_4457,N_4306,N_4335);
nor U4458 (N_4458,N_4247,N_4218);
and U4459 (N_4459,N_4225,N_4270);
or U4460 (N_4460,N_4283,N_4284);
xor U4461 (N_4461,N_4247,N_4240);
or U4462 (N_4462,N_4347,N_4336);
nand U4463 (N_4463,N_4300,N_4201);
or U4464 (N_4464,N_4213,N_4264);
nand U4465 (N_4465,N_4307,N_4206);
or U4466 (N_4466,N_4340,N_4267);
nand U4467 (N_4467,N_4300,N_4307);
nor U4468 (N_4468,N_4259,N_4238);
and U4469 (N_4469,N_4231,N_4349);
and U4470 (N_4470,N_4309,N_4259);
nor U4471 (N_4471,N_4316,N_4212);
and U4472 (N_4472,N_4221,N_4236);
nor U4473 (N_4473,N_4267,N_4310);
xnor U4474 (N_4474,N_4204,N_4249);
or U4475 (N_4475,N_4262,N_4243);
and U4476 (N_4476,N_4333,N_4349);
nand U4477 (N_4477,N_4346,N_4250);
nor U4478 (N_4478,N_4238,N_4287);
xnor U4479 (N_4479,N_4300,N_4322);
or U4480 (N_4480,N_4203,N_4324);
nand U4481 (N_4481,N_4294,N_4284);
or U4482 (N_4482,N_4329,N_4278);
or U4483 (N_4483,N_4303,N_4348);
nand U4484 (N_4484,N_4282,N_4252);
and U4485 (N_4485,N_4301,N_4334);
or U4486 (N_4486,N_4287,N_4233);
nand U4487 (N_4487,N_4275,N_4332);
nor U4488 (N_4488,N_4274,N_4238);
nor U4489 (N_4489,N_4261,N_4344);
nand U4490 (N_4490,N_4226,N_4277);
nand U4491 (N_4491,N_4275,N_4273);
or U4492 (N_4492,N_4241,N_4298);
nand U4493 (N_4493,N_4206,N_4293);
or U4494 (N_4494,N_4314,N_4313);
and U4495 (N_4495,N_4328,N_4322);
xnor U4496 (N_4496,N_4326,N_4308);
nand U4497 (N_4497,N_4316,N_4246);
and U4498 (N_4498,N_4248,N_4226);
nand U4499 (N_4499,N_4346,N_4306);
nor U4500 (N_4500,N_4412,N_4473);
or U4501 (N_4501,N_4486,N_4383);
nand U4502 (N_4502,N_4494,N_4453);
nand U4503 (N_4503,N_4462,N_4372);
nor U4504 (N_4504,N_4454,N_4392);
nor U4505 (N_4505,N_4360,N_4418);
and U4506 (N_4506,N_4489,N_4482);
xnor U4507 (N_4507,N_4370,N_4463);
or U4508 (N_4508,N_4409,N_4407);
nor U4509 (N_4509,N_4378,N_4417);
nand U4510 (N_4510,N_4406,N_4468);
or U4511 (N_4511,N_4426,N_4404);
or U4512 (N_4512,N_4456,N_4476);
and U4513 (N_4513,N_4386,N_4359);
nor U4514 (N_4514,N_4403,N_4373);
xnor U4515 (N_4515,N_4495,N_4355);
nand U4516 (N_4516,N_4379,N_4371);
or U4517 (N_4517,N_4375,N_4430);
nor U4518 (N_4518,N_4433,N_4479);
and U4519 (N_4519,N_4483,N_4429);
xnor U4520 (N_4520,N_4437,N_4465);
nor U4521 (N_4521,N_4478,N_4408);
and U4522 (N_4522,N_4496,N_4410);
xnor U4523 (N_4523,N_4491,N_4405);
nand U4524 (N_4524,N_4461,N_4424);
xnor U4525 (N_4525,N_4364,N_4469);
or U4526 (N_4526,N_4385,N_4438);
and U4527 (N_4527,N_4369,N_4449);
or U4528 (N_4528,N_4363,N_4365);
nand U4529 (N_4529,N_4415,N_4466);
nand U4530 (N_4530,N_4451,N_4395);
and U4531 (N_4531,N_4450,N_4354);
or U4532 (N_4532,N_4487,N_4377);
nor U4533 (N_4533,N_4401,N_4477);
and U4534 (N_4534,N_4423,N_4380);
xor U4535 (N_4535,N_4366,N_4356);
nor U4536 (N_4536,N_4400,N_4436);
xor U4537 (N_4537,N_4367,N_4471);
xor U4538 (N_4538,N_4414,N_4499);
or U4539 (N_4539,N_4493,N_4381);
and U4540 (N_4540,N_4484,N_4445);
and U4541 (N_4541,N_4472,N_4458);
nor U4542 (N_4542,N_4441,N_4442);
nand U4543 (N_4543,N_4455,N_4419);
nand U4544 (N_4544,N_4498,N_4431);
xnor U4545 (N_4545,N_4402,N_4420);
nor U4546 (N_4546,N_4439,N_4452);
nor U4547 (N_4547,N_4459,N_4413);
and U4548 (N_4548,N_4432,N_4362);
and U4549 (N_4549,N_4434,N_4368);
nor U4550 (N_4550,N_4464,N_4447);
nor U4551 (N_4551,N_4352,N_4384);
or U4552 (N_4552,N_4394,N_4376);
or U4553 (N_4553,N_4391,N_4492);
or U4554 (N_4554,N_4353,N_4422);
xnor U4555 (N_4555,N_4397,N_4443);
or U4556 (N_4556,N_4399,N_4448);
nor U4557 (N_4557,N_4393,N_4350);
or U4558 (N_4558,N_4440,N_4382);
nand U4559 (N_4559,N_4390,N_4374);
nand U4560 (N_4560,N_4435,N_4388);
nand U4561 (N_4561,N_4389,N_4396);
or U4562 (N_4562,N_4481,N_4497);
nand U4563 (N_4563,N_4444,N_4416);
nor U4564 (N_4564,N_4357,N_4361);
xnor U4565 (N_4565,N_4398,N_4490);
xnor U4566 (N_4566,N_4480,N_4460);
nand U4567 (N_4567,N_4488,N_4411);
nor U4568 (N_4568,N_4387,N_4457);
or U4569 (N_4569,N_4421,N_4446);
and U4570 (N_4570,N_4358,N_4351);
or U4571 (N_4571,N_4475,N_4428);
nor U4572 (N_4572,N_4470,N_4425);
xnor U4573 (N_4573,N_4474,N_4427);
or U4574 (N_4574,N_4467,N_4485);
and U4575 (N_4575,N_4494,N_4411);
nor U4576 (N_4576,N_4471,N_4494);
nand U4577 (N_4577,N_4486,N_4373);
nor U4578 (N_4578,N_4353,N_4360);
nand U4579 (N_4579,N_4420,N_4437);
or U4580 (N_4580,N_4372,N_4367);
nand U4581 (N_4581,N_4422,N_4374);
nor U4582 (N_4582,N_4434,N_4461);
or U4583 (N_4583,N_4387,N_4421);
or U4584 (N_4584,N_4481,N_4357);
nor U4585 (N_4585,N_4409,N_4351);
xnor U4586 (N_4586,N_4486,N_4445);
nor U4587 (N_4587,N_4352,N_4357);
xnor U4588 (N_4588,N_4447,N_4492);
or U4589 (N_4589,N_4352,N_4481);
or U4590 (N_4590,N_4365,N_4369);
nand U4591 (N_4591,N_4463,N_4458);
nor U4592 (N_4592,N_4386,N_4420);
nand U4593 (N_4593,N_4449,N_4370);
xor U4594 (N_4594,N_4428,N_4427);
nand U4595 (N_4595,N_4485,N_4474);
or U4596 (N_4596,N_4382,N_4468);
nand U4597 (N_4597,N_4426,N_4408);
xor U4598 (N_4598,N_4358,N_4448);
nor U4599 (N_4599,N_4468,N_4461);
and U4600 (N_4600,N_4408,N_4437);
nor U4601 (N_4601,N_4459,N_4468);
and U4602 (N_4602,N_4442,N_4368);
xnor U4603 (N_4603,N_4491,N_4457);
nor U4604 (N_4604,N_4358,N_4393);
and U4605 (N_4605,N_4452,N_4454);
and U4606 (N_4606,N_4490,N_4374);
xnor U4607 (N_4607,N_4396,N_4351);
or U4608 (N_4608,N_4367,N_4485);
and U4609 (N_4609,N_4433,N_4467);
xor U4610 (N_4610,N_4425,N_4406);
or U4611 (N_4611,N_4493,N_4477);
xor U4612 (N_4612,N_4444,N_4466);
nand U4613 (N_4613,N_4392,N_4446);
or U4614 (N_4614,N_4401,N_4449);
nand U4615 (N_4615,N_4402,N_4477);
and U4616 (N_4616,N_4467,N_4475);
xnor U4617 (N_4617,N_4461,N_4394);
and U4618 (N_4618,N_4374,N_4426);
nor U4619 (N_4619,N_4380,N_4405);
xor U4620 (N_4620,N_4357,N_4461);
xor U4621 (N_4621,N_4387,N_4473);
nand U4622 (N_4622,N_4392,N_4495);
nor U4623 (N_4623,N_4353,N_4412);
and U4624 (N_4624,N_4432,N_4451);
and U4625 (N_4625,N_4461,N_4489);
nor U4626 (N_4626,N_4452,N_4469);
nand U4627 (N_4627,N_4411,N_4424);
and U4628 (N_4628,N_4490,N_4481);
nor U4629 (N_4629,N_4383,N_4366);
and U4630 (N_4630,N_4483,N_4375);
xnor U4631 (N_4631,N_4351,N_4462);
and U4632 (N_4632,N_4489,N_4398);
xnor U4633 (N_4633,N_4447,N_4363);
nor U4634 (N_4634,N_4439,N_4413);
nand U4635 (N_4635,N_4486,N_4479);
xor U4636 (N_4636,N_4454,N_4389);
xnor U4637 (N_4637,N_4436,N_4482);
and U4638 (N_4638,N_4399,N_4379);
and U4639 (N_4639,N_4352,N_4412);
nor U4640 (N_4640,N_4493,N_4357);
nand U4641 (N_4641,N_4498,N_4452);
nor U4642 (N_4642,N_4413,N_4464);
nor U4643 (N_4643,N_4413,N_4367);
or U4644 (N_4644,N_4406,N_4379);
nor U4645 (N_4645,N_4408,N_4397);
or U4646 (N_4646,N_4383,N_4442);
nor U4647 (N_4647,N_4418,N_4405);
or U4648 (N_4648,N_4448,N_4384);
xnor U4649 (N_4649,N_4458,N_4350);
nor U4650 (N_4650,N_4611,N_4605);
xnor U4651 (N_4651,N_4609,N_4520);
xnor U4652 (N_4652,N_4563,N_4649);
and U4653 (N_4653,N_4573,N_4562);
or U4654 (N_4654,N_4642,N_4510);
nand U4655 (N_4655,N_4637,N_4513);
and U4656 (N_4656,N_4534,N_4557);
nand U4657 (N_4657,N_4623,N_4554);
and U4658 (N_4658,N_4645,N_4580);
nand U4659 (N_4659,N_4505,N_4618);
nand U4660 (N_4660,N_4641,N_4561);
or U4661 (N_4661,N_4575,N_4526);
or U4662 (N_4662,N_4521,N_4643);
nor U4663 (N_4663,N_4548,N_4558);
nor U4664 (N_4664,N_4602,N_4585);
nand U4665 (N_4665,N_4604,N_4582);
nand U4666 (N_4666,N_4509,N_4572);
and U4667 (N_4667,N_4647,N_4535);
and U4668 (N_4668,N_4538,N_4570);
or U4669 (N_4669,N_4587,N_4595);
and U4670 (N_4670,N_4626,N_4593);
and U4671 (N_4671,N_4567,N_4581);
nand U4672 (N_4672,N_4603,N_4512);
and U4673 (N_4673,N_4627,N_4571);
nor U4674 (N_4674,N_4615,N_4516);
or U4675 (N_4675,N_4519,N_4569);
xnor U4676 (N_4676,N_4613,N_4524);
xor U4677 (N_4677,N_4583,N_4619);
nand U4678 (N_4678,N_4547,N_4511);
nor U4679 (N_4679,N_4636,N_4523);
xor U4680 (N_4680,N_4531,N_4500);
xor U4681 (N_4681,N_4638,N_4617);
nand U4682 (N_4682,N_4600,N_4622);
nand U4683 (N_4683,N_4527,N_4525);
xnor U4684 (N_4684,N_4620,N_4586);
xnor U4685 (N_4685,N_4514,N_4559);
xor U4686 (N_4686,N_4579,N_4560);
nand U4687 (N_4687,N_4503,N_4549);
nand U4688 (N_4688,N_4553,N_4644);
nor U4689 (N_4689,N_4590,N_4536);
or U4690 (N_4690,N_4631,N_4608);
nor U4691 (N_4691,N_4634,N_4610);
and U4692 (N_4692,N_4614,N_4566);
or U4693 (N_4693,N_4628,N_4541);
xor U4694 (N_4694,N_4506,N_4597);
and U4695 (N_4695,N_4630,N_4598);
nand U4696 (N_4696,N_4577,N_4594);
nor U4697 (N_4697,N_4621,N_4502);
nand U4698 (N_4698,N_4550,N_4545);
nand U4699 (N_4699,N_4646,N_4522);
nor U4700 (N_4700,N_4625,N_4504);
nor U4701 (N_4701,N_4635,N_4543);
and U4702 (N_4702,N_4515,N_4529);
or U4703 (N_4703,N_4624,N_4546);
xnor U4704 (N_4704,N_4599,N_4539);
nor U4705 (N_4705,N_4556,N_4612);
nand U4706 (N_4706,N_4639,N_4508);
xnor U4707 (N_4707,N_4640,N_4540);
and U4708 (N_4708,N_4584,N_4578);
nand U4709 (N_4709,N_4537,N_4530);
xor U4710 (N_4710,N_4633,N_4596);
or U4711 (N_4711,N_4607,N_4565);
or U4712 (N_4712,N_4589,N_4532);
nor U4713 (N_4713,N_4501,N_4588);
xor U4714 (N_4714,N_4544,N_4518);
or U4715 (N_4715,N_4632,N_4528);
and U4716 (N_4716,N_4648,N_4564);
or U4717 (N_4717,N_4517,N_4629);
nand U4718 (N_4718,N_4574,N_4507);
and U4719 (N_4719,N_4616,N_4542);
nor U4720 (N_4720,N_4552,N_4568);
nand U4721 (N_4721,N_4606,N_4555);
nor U4722 (N_4722,N_4551,N_4601);
nor U4723 (N_4723,N_4533,N_4592);
nor U4724 (N_4724,N_4591,N_4576);
nor U4725 (N_4725,N_4566,N_4539);
xnor U4726 (N_4726,N_4533,N_4637);
or U4727 (N_4727,N_4583,N_4646);
nor U4728 (N_4728,N_4620,N_4563);
or U4729 (N_4729,N_4503,N_4563);
nand U4730 (N_4730,N_4629,N_4508);
nand U4731 (N_4731,N_4567,N_4625);
nand U4732 (N_4732,N_4596,N_4511);
nor U4733 (N_4733,N_4647,N_4643);
and U4734 (N_4734,N_4588,N_4608);
nor U4735 (N_4735,N_4573,N_4526);
nor U4736 (N_4736,N_4522,N_4550);
and U4737 (N_4737,N_4598,N_4508);
nor U4738 (N_4738,N_4579,N_4531);
nand U4739 (N_4739,N_4625,N_4586);
and U4740 (N_4740,N_4647,N_4624);
nor U4741 (N_4741,N_4582,N_4544);
nand U4742 (N_4742,N_4545,N_4629);
xor U4743 (N_4743,N_4549,N_4640);
nand U4744 (N_4744,N_4555,N_4629);
xor U4745 (N_4745,N_4619,N_4566);
xor U4746 (N_4746,N_4529,N_4639);
nand U4747 (N_4747,N_4613,N_4614);
and U4748 (N_4748,N_4629,N_4643);
nor U4749 (N_4749,N_4534,N_4501);
nor U4750 (N_4750,N_4629,N_4564);
and U4751 (N_4751,N_4525,N_4639);
xnor U4752 (N_4752,N_4555,N_4526);
nor U4753 (N_4753,N_4606,N_4550);
nand U4754 (N_4754,N_4615,N_4509);
and U4755 (N_4755,N_4568,N_4621);
nor U4756 (N_4756,N_4542,N_4523);
nand U4757 (N_4757,N_4587,N_4513);
nor U4758 (N_4758,N_4580,N_4619);
xor U4759 (N_4759,N_4583,N_4591);
or U4760 (N_4760,N_4539,N_4569);
nand U4761 (N_4761,N_4558,N_4594);
or U4762 (N_4762,N_4573,N_4599);
nand U4763 (N_4763,N_4583,N_4576);
nand U4764 (N_4764,N_4585,N_4579);
xnor U4765 (N_4765,N_4602,N_4632);
nor U4766 (N_4766,N_4547,N_4593);
nor U4767 (N_4767,N_4635,N_4518);
nor U4768 (N_4768,N_4554,N_4612);
nor U4769 (N_4769,N_4548,N_4586);
xor U4770 (N_4770,N_4511,N_4530);
nand U4771 (N_4771,N_4570,N_4577);
or U4772 (N_4772,N_4504,N_4554);
nor U4773 (N_4773,N_4531,N_4569);
and U4774 (N_4774,N_4567,N_4632);
nand U4775 (N_4775,N_4619,N_4501);
or U4776 (N_4776,N_4581,N_4516);
and U4777 (N_4777,N_4568,N_4531);
or U4778 (N_4778,N_4545,N_4605);
or U4779 (N_4779,N_4534,N_4559);
or U4780 (N_4780,N_4612,N_4632);
or U4781 (N_4781,N_4597,N_4548);
and U4782 (N_4782,N_4556,N_4563);
nand U4783 (N_4783,N_4642,N_4632);
nor U4784 (N_4784,N_4577,N_4534);
nor U4785 (N_4785,N_4583,N_4605);
nor U4786 (N_4786,N_4515,N_4635);
nand U4787 (N_4787,N_4629,N_4500);
or U4788 (N_4788,N_4610,N_4588);
or U4789 (N_4789,N_4620,N_4597);
and U4790 (N_4790,N_4623,N_4642);
or U4791 (N_4791,N_4578,N_4594);
nor U4792 (N_4792,N_4543,N_4630);
and U4793 (N_4793,N_4541,N_4554);
nand U4794 (N_4794,N_4623,N_4601);
xnor U4795 (N_4795,N_4643,N_4520);
nor U4796 (N_4796,N_4510,N_4596);
nand U4797 (N_4797,N_4531,N_4586);
and U4798 (N_4798,N_4569,N_4566);
or U4799 (N_4799,N_4525,N_4503);
nand U4800 (N_4800,N_4681,N_4791);
nand U4801 (N_4801,N_4798,N_4771);
nand U4802 (N_4802,N_4678,N_4754);
nor U4803 (N_4803,N_4714,N_4783);
xor U4804 (N_4804,N_4677,N_4658);
xnor U4805 (N_4805,N_4661,N_4653);
or U4806 (N_4806,N_4762,N_4696);
and U4807 (N_4807,N_4724,N_4730);
xor U4808 (N_4808,N_4773,N_4682);
nor U4809 (N_4809,N_4794,N_4704);
nor U4810 (N_4810,N_4793,N_4728);
nand U4811 (N_4811,N_4721,N_4778);
and U4812 (N_4812,N_4756,N_4675);
nand U4813 (N_4813,N_4715,N_4680);
and U4814 (N_4814,N_4779,N_4750);
nor U4815 (N_4815,N_4748,N_4781);
or U4816 (N_4816,N_4753,N_4763);
and U4817 (N_4817,N_4692,N_4788);
nand U4818 (N_4818,N_4786,N_4743);
nor U4819 (N_4819,N_4709,N_4796);
and U4820 (N_4820,N_4758,N_4686);
nand U4821 (N_4821,N_4745,N_4711);
nor U4822 (N_4822,N_4747,N_4736);
nand U4823 (N_4823,N_4738,N_4760);
nand U4824 (N_4824,N_4701,N_4734);
nand U4825 (N_4825,N_4713,N_4703);
xor U4826 (N_4826,N_4782,N_4769);
nor U4827 (N_4827,N_4690,N_4666);
and U4828 (N_4828,N_4770,N_4664);
nand U4829 (N_4829,N_4797,N_4685);
nand U4830 (N_4830,N_4732,N_4751);
nand U4831 (N_4831,N_4670,N_4727);
or U4832 (N_4832,N_4710,N_4722);
nand U4833 (N_4833,N_4651,N_4687);
nand U4834 (N_4834,N_4777,N_4699);
or U4835 (N_4835,N_4739,N_4667);
nand U4836 (N_4836,N_4659,N_4707);
and U4837 (N_4837,N_4656,N_4723);
nand U4838 (N_4838,N_4652,N_4671);
nor U4839 (N_4839,N_4761,N_4700);
and U4840 (N_4840,N_4705,N_4755);
xor U4841 (N_4841,N_4650,N_4749);
xnor U4842 (N_4842,N_4717,N_4683);
nand U4843 (N_4843,N_4662,N_4708);
nor U4844 (N_4844,N_4746,N_4772);
and U4845 (N_4845,N_4693,N_4785);
xor U4846 (N_4846,N_4716,N_4698);
nand U4847 (N_4847,N_4684,N_4688);
xor U4848 (N_4848,N_4689,N_4695);
or U4849 (N_4849,N_4702,N_4737);
or U4850 (N_4850,N_4726,N_4789);
and U4851 (N_4851,N_4764,N_4733);
xor U4852 (N_4852,N_4691,N_4757);
nand U4853 (N_4853,N_4694,N_4657);
nand U4854 (N_4854,N_4731,N_4655);
nor U4855 (N_4855,N_4741,N_4742);
nand U4856 (N_4856,N_4676,N_4792);
and U4857 (N_4857,N_4766,N_4799);
or U4858 (N_4858,N_4725,N_4776);
nor U4859 (N_4859,N_4679,N_4744);
nand U4860 (N_4860,N_4654,N_4706);
xnor U4861 (N_4861,N_4787,N_4719);
and U4862 (N_4862,N_4668,N_4669);
nand U4863 (N_4863,N_4740,N_4663);
or U4864 (N_4864,N_4674,N_4673);
xnor U4865 (N_4865,N_4795,N_4759);
and U4866 (N_4866,N_4774,N_4735);
nor U4867 (N_4867,N_4718,N_4790);
and U4868 (N_4868,N_4729,N_4767);
and U4869 (N_4869,N_4665,N_4784);
and U4870 (N_4870,N_4660,N_4712);
xnor U4871 (N_4871,N_4780,N_4720);
xnor U4872 (N_4872,N_4768,N_4775);
and U4873 (N_4873,N_4765,N_4752);
or U4874 (N_4874,N_4672,N_4697);
nand U4875 (N_4875,N_4738,N_4791);
nor U4876 (N_4876,N_4767,N_4679);
nand U4877 (N_4877,N_4779,N_4695);
or U4878 (N_4878,N_4740,N_4709);
nand U4879 (N_4879,N_4776,N_4678);
nand U4880 (N_4880,N_4655,N_4756);
nand U4881 (N_4881,N_4743,N_4746);
and U4882 (N_4882,N_4670,N_4722);
and U4883 (N_4883,N_4730,N_4725);
or U4884 (N_4884,N_4707,N_4763);
xor U4885 (N_4885,N_4771,N_4736);
or U4886 (N_4886,N_4761,N_4687);
nand U4887 (N_4887,N_4715,N_4728);
xor U4888 (N_4888,N_4771,N_4670);
and U4889 (N_4889,N_4744,N_4663);
nor U4890 (N_4890,N_4795,N_4722);
xnor U4891 (N_4891,N_4715,N_4655);
and U4892 (N_4892,N_4792,N_4795);
and U4893 (N_4893,N_4676,N_4777);
nor U4894 (N_4894,N_4776,N_4773);
xnor U4895 (N_4895,N_4726,N_4740);
nand U4896 (N_4896,N_4691,N_4793);
or U4897 (N_4897,N_4667,N_4735);
nand U4898 (N_4898,N_4654,N_4650);
or U4899 (N_4899,N_4747,N_4690);
or U4900 (N_4900,N_4732,N_4782);
and U4901 (N_4901,N_4656,N_4764);
or U4902 (N_4902,N_4742,N_4711);
xor U4903 (N_4903,N_4762,N_4687);
or U4904 (N_4904,N_4731,N_4658);
xor U4905 (N_4905,N_4700,N_4695);
nand U4906 (N_4906,N_4754,N_4782);
nor U4907 (N_4907,N_4699,N_4692);
xor U4908 (N_4908,N_4731,N_4676);
nand U4909 (N_4909,N_4666,N_4695);
or U4910 (N_4910,N_4686,N_4796);
or U4911 (N_4911,N_4699,N_4723);
nor U4912 (N_4912,N_4661,N_4797);
nor U4913 (N_4913,N_4717,N_4714);
and U4914 (N_4914,N_4717,N_4712);
xnor U4915 (N_4915,N_4702,N_4713);
or U4916 (N_4916,N_4706,N_4788);
nand U4917 (N_4917,N_4657,N_4720);
and U4918 (N_4918,N_4735,N_4744);
nand U4919 (N_4919,N_4682,N_4772);
and U4920 (N_4920,N_4752,N_4776);
nand U4921 (N_4921,N_4681,N_4742);
nand U4922 (N_4922,N_4767,N_4794);
nor U4923 (N_4923,N_4732,N_4785);
or U4924 (N_4924,N_4655,N_4722);
or U4925 (N_4925,N_4797,N_4741);
xnor U4926 (N_4926,N_4740,N_4756);
or U4927 (N_4927,N_4740,N_4755);
and U4928 (N_4928,N_4701,N_4708);
or U4929 (N_4929,N_4745,N_4781);
nor U4930 (N_4930,N_4694,N_4717);
and U4931 (N_4931,N_4709,N_4654);
nor U4932 (N_4932,N_4753,N_4718);
or U4933 (N_4933,N_4670,N_4764);
nor U4934 (N_4934,N_4677,N_4792);
and U4935 (N_4935,N_4712,N_4750);
xnor U4936 (N_4936,N_4735,N_4787);
xnor U4937 (N_4937,N_4712,N_4665);
nand U4938 (N_4938,N_4728,N_4683);
or U4939 (N_4939,N_4741,N_4767);
nor U4940 (N_4940,N_4794,N_4751);
xnor U4941 (N_4941,N_4667,N_4707);
nand U4942 (N_4942,N_4666,N_4722);
or U4943 (N_4943,N_4664,N_4653);
nand U4944 (N_4944,N_4651,N_4670);
xor U4945 (N_4945,N_4680,N_4659);
or U4946 (N_4946,N_4719,N_4791);
nor U4947 (N_4947,N_4658,N_4661);
nand U4948 (N_4948,N_4769,N_4714);
nand U4949 (N_4949,N_4685,N_4735);
nor U4950 (N_4950,N_4811,N_4935);
xnor U4951 (N_4951,N_4858,N_4844);
xor U4952 (N_4952,N_4940,N_4913);
or U4953 (N_4953,N_4944,N_4895);
and U4954 (N_4954,N_4828,N_4800);
xor U4955 (N_4955,N_4904,N_4856);
and U4956 (N_4956,N_4901,N_4910);
nand U4957 (N_4957,N_4946,N_4863);
nor U4958 (N_4958,N_4880,N_4833);
nor U4959 (N_4959,N_4902,N_4877);
or U4960 (N_4960,N_4889,N_4825);
nand U4961 (N_4961,N_4906,N_4829);
and U4962 (N_4962,N_4948,N_4941);
or U4963 (N_4963,N_4843,N_4879);
nand U4964 (N_4964,N_4848,N_4839);
and U4965 (N_4965,N_4882,N_4868);
nand U4966 (N_4966,N_4846,N_4900);
or U4967 (N_4967,N_4893,N_4857);
xor U4968 (N_4968,N_4938,N_4826);
xor U4969 (N_4969,N_4860,N_4908);
or U4970 (N_4970,N_4914,N_4830);
xnor U4971 (N_4971,N_4907,N_4928);
and U4972 (N_4972,N_4850,N_4849);
or U4973 (N_4973,N_4945,N_4929);
nor U4974 (N_4974,N_4834,N_4947);
nor U4975 (N_4975,N_4837,N_4869);
nand U4976 (N_4976,N_4832,N_4836);
nand U4977 (N_4977,N_4864,N_4911);
nor U4978 (N_4978,N_4896,N_4930);
and U4979 (N_4979,N_4861,N_4926);
and U4980 (N_4980,N_4912,N_4892);
and U4981 (N_4981,N_4862,N_4899);
nand U4982 (N_4982,N_4838,N_4887);
and U4983 (N_4983,N_4949,N_4924);
and U4984 (N_4984,N_4805,N_4808);
nor U4985 (N_4985,N_4865,N_4890);
or U4986 (N_4986,N_4927,N_4853);
or U4987 (N_4987,N_4898,N_4883);
or U4988 (N_4988,N_4822,N_4866);
and U4989 (N_4989,N_4814,N_4842);
nor U4990 (N_4990,N_4859,N_4937);
or U4991 (N_4991,N_4855,N_4897);
and U4992 (N_4992,N_4824,N_4820);
xor U4993 (N_4993,N_4806,N_4886);
xnor U4994 (N_4994,N_4835,N_4871);
nor U4995 (N_4995,N_4942,N_4810);
and U4996 (N_4996,N_4872,N_4867);
nor U4997 (N_4997,N_4801,N_4919);
and U4998 (N_4998,N_4870,N_4813);
nor U4999 (N_4999,N_4809,N_4921);
or U5000 (N_5000,N_4854,N_4816);
nor U5001 (N_5001,N_4888,N_4873);
or U5002 (N_5002,N_4934,N_4920);
or U5003 (N_5003,N_4922,N_4812);
or U5004 (N_5004,N_4841,N_4909);
nor U5005 (N_5005,N_4851,N_4821);
and U5006 (N_5006,N_4894,N_4933);
and U5007 (N_5007,N_4905,N_4807);
and U5008 (N_5008,N_4923,N_4823);
nor U5009 (N_5009,N_4916,N_4847);
nand U5010 (N_5010,N_4891,N_4818);
nand U5011 (N_5011,N_4915,N_4875);
xnor U5012 (N_5012,N_4943,N_4936);
nand U5013 (N_5013,N_4840,N_4852);
and U5014 (N_5014,N_4881,N_4931);
and U5015 (N_5015,N_4903,N_4878);
and U5016 (N_5016,N_4885,N_4815);
and U5017 (N_5017,N_4939,N_4932);
xor U5018 (N_5018,N_4884,N_4918);
or U5019 (N_5019,N_4845,N_4917);
or U5020 (N_5020,N_4803,N_4817);
nand U5021 (N_5021,N_4876,N_4874);
nand U5022 (N_5022,N_4819,N_4802);
xor U5023 (N_5023,N_4925,N_4804);
nand U5024 (N_5024,N_4831,N_4827);
and U5025 (N_5025,N_4865,N_4882);
nor U5026 (N_5026,N_4828,N_4821);
nor U5027 (N_5027,N_4926,N_4895);
and U5028 (N_5028,N_4924,N_4851);
or U5029 (N_5029,N_4801,N_4912);
and U5030 (N_5030,N_4817,N_4913);
and U5031 (N_5031,N_4851,N_4839);
nor U5032 (N_5032,N_4869,N_4948);
and U5033 (N_5033,N_4920,N_4848);
nor U5034 (N_5034,N_4872,N_4838);
or U5035 (N_5035,N_4937,N_4837);
and U5036 (N_5036,N_4842,N_4833);
xnor U5037 (N_5037,N_4807,N_4874);
or U5038 (N_5038,N_4918,N_4816);
xnor U5039 (N_5039,N_4877,N_4843);
xor U5040 (N_5040,N_4866,N_4855);
nor U5041 (N_5041,N_4800,N_4875);
or U5042 (N_5042,N_4935,N_4914);
xnor U5043 (N_5043,N_4908,N_4843);
nor U5044 (N_5044,N_4876,N_4870);
xnor U5045 (N_5045,N_4827,N_4873);
and U5046 (N_5046,N_4827,N_4921);
xnor U5047 (N_5047,N_4928,N_4940);
nand U5048 (N_5048,N_4948,N_4879);
and U5049 (N_5049,N_4805,N_4830);
nor U5050 (N_5050,N_4910,N_4832);
and U5051 (N_5051,N_4858,N_4939);
and U5052 (N_5052,N_4841,N_4807);
nand U5053 (N_5053,N_4896,N_4802);
and U5054 (N_5054,N_4826,N_4944);
nand U5055 (N_5055,N_4890,N_4884);
and U5056 (N_5056,N_4841,N_4876);
and U5057 (N_5057,N_4863,N_4853);
xnor U5058 (N_5058,N_4943,N_4836);
or U5059 (N_5059,N_4862,N_4931);
or U5060 (N_5060,N_4933,N_4819);
xor U5061 (N_5061,N_4910,N_4919);
or U5062 (N_5062,N_4904,N_4838);
or U5063 (N_5063,N_4915,N_4943);
xor U5064 (N_5064,N_4909,N_4824);
nand U5065 (N_5065,N_4893,N_4912);
nor U5066 (N_5066,N_4884,N_4932);
nand U5067 (N_5067,N_4928,N_4827);
xnor U5068 (N_5068,N_4824,N_4830);
xor U5069 (N_5069,N_4846,N_4813);
and U5070 (N_5070,N_4879,N_4947);
or U5071 (N_5071,N_4840,N_4890);
nand U5072 (N_5072,N_4870,N_4895);
and U5073 (N_5073,N_4887,N_4868);
and U5074 (N_5074,N_4854,N_4869);
nand U5075 (N_5075,N_4887,N_4863);
or U5076 (N_5076,N_4868,N_4838);
nor U5077 (N_5077,N_4862,N_4940);
xor U5078 (N_5078,N_4807,N_4931);
nor U5079 (N_5079,N_4916,N_4863);
nor U5080 (N_5080,N_4873,N_4947);
and U5081 (N_5081,N_4855,N_4869);
xor U5082 (N_5082,N_4871,N_4931);
or U5083 (N_5083,N_4921,N_4867);
and U5084 (N_5084,N_4897,N_4842);
xor U5085 (N_5085,N_4933,N_4843);
nand U5086 (N_5086,N_4864,N_4858);
nand U5087 (N_5087,N_4806,N_4919);
and U5088 (N_5088,N_4802,N_4858);
nor U5089 (N_5089,N_4850,N_4903);
nand U5090 (N_5090,N_4832,N_4884);
nor U5091 (N_5091,N_4927,N_4864);
and U5092 (N_5092,N_4932,N_4807);
nand U5093 (N_5093,N_4905,N_4948);
nand U5094 (N_5094,N_4874,N_4912);
xnor U5095 (N_5095,N_4876,N_4832);
xnor U5096 (N_5096,N_4819,N_4939);
xor U5097 (N_5097,N_4908,N_4857);
nor U5098 (N_5098,N_4818,N_4839);
nor U5099 (N_5099,N_4851,N_4864);
nand U5100 (N_5100,N_5067,N_5006);
and U5101 (N_5101,N_4983,N_4980);
nor U5102 (N_5102,N_5047,N_4998);
and U5103 (N_5103,N_5005,N_5083);
nor U5104 (N_5104,N_4972,N_5072);
or U5105 (N_5105,N_5073,N_4963);
nand U5106 (N_5106,N_4953,N_5063);
and U5107 (N_5107,N_5029,N_5008);
nand U5108 (N_5108,N_5015,N_4986);
or U5109 (N_5109,N_5041,N_4952);
and U5110 (N_5110,N_5070,N_5040);
nand U5111 (N_5111,N_5039,N_5016);
and U5112 (N_5112,N_5060,N_5032);
nand U5113 (N_5113,N_4993,N_5010);
and U5114 (N_5114,N_4988,N_5004);
or U5115 (N_5115,N_5075,N_4959);
nand U5116 (N_5116,N_5024,N_4954);
and U5117 (N_5117,N_5023,N_5019);
or U5118 (N_5118,N_5002,N_5077);
and U5119 (N_5119,N_5052,N_5020);
or U5120 (N_5120,N_4982,N_5093);
xor U5121 (N_5121,N_4964,N_4961);
and U5122 (N_5122,N_4978,N_4973);
and U5123 (N_5123,N_5097,N_5034);
nor U5124 (N_5124,N_4991,N_5076);
and U5125 (N_5125,N_5090,N_4957);
and U5126 (N_5126,N_5055,N_5095);
and U5127 (N_5127,N_5058,N_5053);
or U5128 (N_5128,N_4979,N_5089);
xor U5129 (N_5129,N_4984,N_5009);
and U5130 (N_5130,N_5081,N_5001);
nor U5131 (N_5131,N_5098,N_5013);
nand U5132 (N_5132,N_4962,N_4974);
xnor U5133 (N_5133,N_4950,N_5078);
nand U5134 (N_5134,N_5003,N_5022);
and U5135 (N_5135,N_4969,N_4977);
nand U5136 (N_5136,N_5031,N_4971);
and U5137 (N_5137,N_5045,N_5017);
and U5138 (N_5138,N_5085,N_5014);
nor U5139 (N_5139,N_4956,N_5092);
or U5140 (N_5140,N_5042,N_5071);
or U5141 (N_5141,N_4955,N_4985);
or U5142 (N_5142,N_4996,N_4995);
and U5143 (N_5143,N_5080,N_4966);
or U5144 (N_5144,N_5064,N_5021);
xor U5145 (N_5145,N_5059,N_4994);
nor U5146 (N_5146,N_5056,N_5050);
or U5147 (N_5147,N_5043,N_4989);
and U5148 (N_5148,N_5065,N_5057);
and U5149 (N_5149,N_4990,N_4967);
or U5150 (N_5150,N_4997,N_5086);
xor U5151 (N_5151,N_4987,N_5061);
nor U5152 (N_5152,N_4999,N_5037);
or U5153 (N_5153,N_4960,N_5000);
xor U5154 (N_5154,N_5033,N_5038);
and U5155 (N_5155,N_5011,N_5027);
and U5156 (N_5156,N_5066,N_5087);
nand U5157 (N_5157,N_5030,N_4975);
nand U5158 (N_5158,N_5049,N_5026);
nand U5159 (N_5159,N_4958,N_5048);
xor U5160 (N_5160,N_5074,N_5091);
nand U5161 (N_5161,N_5012,N_5062);
nor U5162 (N_5162,N_4951,N_4965);
and U5163 (N_5163,N_4981,N_5018);
or U5164 (N_5164,N_5036,N_4976);
or U5165 (N_5165,N_5007,N_4992);
xor U5166 (N_5166,N_5088,N_5028);
nand U5167 (N_5167,N_4970,N_5054);
and U5168 (N_5168,N_5082,N_5051);
and U5169 (N_5169,N_5044,N_5084);
nand U5170 (N_5170,N_4968,N_5094);
or U5171 (N_5171,N_5079,N_5099);
or U5172 (N_5172,N_5046,N_5068);
and U5173 (N_5173,N_5069,N_5025);
nand U5174 (N_5174,N_5035,N_5096);
nor U5175 (N_5175,N_5071,N_5068);
or U5176 (N_5176,N_5033,N_4981);
and U5177 (N_5177,N_5001,N_5040);
xnor U5178 (N_5178,N_4957,N_4960);
or U5179 (N_5179,N_5039,N_5047);
or U5180 (N_5180,N_5093,N_4963);
nand U5181 (N_5181,N_5020,N_5023);
or U5182 (N_5182,N_5085,N_5053);
nand U5183 (N_5183,N_4995,N_4963);
or U5184 (N_5184,N_5010,N_5048);
or U5185 (N_5185,N_4964,N_5041);
or U5186 (N_5186,N_5058,N_5070);
nand U5187 (N_5187,N_4964,N_5056);
and U5188 (N_5188,N_4978,N_4980);
xnor U5189 (N_5189,N_4997,N_5035);
or U5190 (N_5190,N_4986,N_5097);
or U5191 (N_5191,N_5045,N_5080);
nor U5192 (N_5192,N_5028,N_5020);
xnor U5193 (N_5193,N_5054,N_5073);
xnor U5194 (N_5194,N_5068,N_5021);
or U5195 (N_5195,N_5084,N_4967);
nand U5196 (N_5196,N_5052,N_5039);
and U5197 (N_5197,N_5042,N_5095);
xor U5198 (N_5198,N_5028,N_4980);
nor U5199 (N_5199,N_5088,N_5071);
nand U5200 (N_5200,N_4969,N_5081);
or U5201 (N_5201,N_5075,N_5048);
nor U5202 (N_5202,N_5088,N_5070);
and U5203 (N_5203,N_5017,N_5038);
xnor U5204 (N_5204,N_5087,N_5052);
nand U5205 (N_5205,N_5034,N_4965);
or U5206 (N_5206,N_4996,N_5080);
xor U5207 (N_5207,N_4964,N_5053);
or U5208 (N_5208,N_4963,N_5006);
nand U5209 (N_5209,N_4972,N_5064);
and U5210 (N_5210,N_4976,N_5099);
xor U5211 (N_5211,N_5029,N_4972);
nor U5212 (N_5212,N_4988,N_5007);
xnor U5213 (N_5213,N_5038,N_5025);
nor U5214 (N_5214,N_5039,N_5003);
or U5215 (N_5215,N_4957,N_4972);
nor U5216 (N_5216,N_5047,N_5061);
xor U5217 (N_5217,N_4998,N_4994);
or U5218 (N_5218,N_4984,N_5074);
nor U5219 (N_5219,N_4952,N_5000);
xor U5220 (N_5220,N_5099,N_4992);
nor U5221 (N_5221,N_5063,N_5025);
nand U5222 (N_5222,N_5017,N_5095);
and U5223 (N_5223,N_5010,N_4991);
and U5224 (N_5224,N_5021,N_5033);
nor U5225 (N_5225,N_5037,N_5070);
or U5226 (N_5226,N_4983,N_5084);
nand U5227 (N_5227,N_4986,N_4953);
or U5228 (N_5228,N_5083,N_4951);
or U5229 (N_5229,N_5089,N_5054);
and U5230 (N_5230,N_4965,N_5051);
and U5231 (N_5231,N_5044,N_5054);
nor U5232 (N_5232,N_5064,N_5068);
and U5233 (N_5233,N_4987,N_5029);
and U5234 (N_5234,N_5027,N_4962);
nand U5235 (N_5235,N_5013,N_5000);
and U5236 (N_5236,N_5095,N_5032);
nand U5237 (N_5237,N_4960,N_5097);
nand U5238 (N_5238,N_4953,N_5093);
nand U5239 (N_5239,N_5067,N_5014);
nand U5240 (N_5240,N_5024,N_4982);
or U5241 (N_5241,N_5089,N_5065);
or U5242 (N_5242,N_5092,N_5084);
and U5243 (N_5243,N_5050,N_5003);
nor U5244 (N_5244,N_5051,N_5034);
nand U5245 (N_5245,N_5026,N_4973);
nor U5246 (N_5246,N_4979,N_5048);
nand U5247 (N_5247,N_5087,N_5099);
or U5248 (N_5248,N_5069,N_5088);
and U5249 (N_5249,N_5083,N_4989);
nand U5250 (N_5250,N_5247,N_5119);
or U5251 (N_5251,N_5193,N_5186);
or U5252 (N_5252,N_5127,N_5242);
or U5253 (N_5253,N_5101,N_5149);
nor U5254 (N_5254,N_5156,N_5103);
xor U5255 (N_5255,N_5126,N_5150);
nand U5256 (N_5256,N_5217,N_5215);
and U5257 (N_5257,N_5225,N_5134);
nor U5258 (N_5258,N_5209,N_5138);
and U5259 (N_5259,N_5113,N_5195);
and U5260 (N_5260,N_5108,N_5173);
and U5261 (N_5261,N_5184,N_5190);
xor U5262 (N_5262,N_5171,N_5216);
nor U5263 (N_5263,N_5107,N_5191);
xor U5264 (N_5264,N_5109,N_5223);
or U5265 (N_5265,N_5131,N_5221);
and U5266 (N_5266,N_5220,N_5144);
or U5267 (N_5267,N_5181,N_5233);
or U5268 (N_5268,N_5231,N_5129);
and U5269 (N_5269,N_5100,N_5140);
or U5270 (N_5270,N_5204,N_5199);
or U5271 (N_5271,N_5122,N_5170);
xnor U5272 (N_5272,N_5174,N_5192);
or U5273 (N_5273,N_5178,N_5194);
nand U5274 (N_5274,N_5137,N_5118);
xnor U5275 (N_5275,N_5154,N_5133);
or U5276 (N_5276,N_5239,N_5185);
xnor U5277 (N_5277,N_5224,N_5197);
nand U5278 (N_5278,N_5219,N_5106);
and U5279 (N_5279,N_5240,N_5172);
nand U5280 (N_5280,N_5228,N_5214);
nand U5281 (N_5281,N_5164,N_5165);
xnor U5282 (N_5282,N_5182,N_5167);
and U5283 (N_5283,N_5222,N_5203);
xor U5284 (N_5284,N_5143,N_5176);
and U5285 (N_5285,N_5128,N_5160);
nor U5286 (N_5286,N_5115,N_5230);
or U5287 (N_5287,N_5177,N_5152);
nand U5288 (N_5288,N_5227,N_5237);
and U5289 (N_5289,N_5201,N_5147);
xnor U5290 (N_5290,N_5166,N_5207);
nand U5291 (N_5291,N_5168,N_5141);
xnor U5292 (N_5292,N_5132,N_5198);
xor U5293 (N_5293,N_5120,N_5187);
nor U5294 (N_5294,N_5111,N_5241);
and U5295 (N_5295,N_5145,N_5124);
and U5296 (N_5296,N_5236,N_5249);
nor U5297 (N_5297,N_5246,N_5169);
nor U5298 (N_5298,N_5206,N_5205);
xor U5299 (N_5299,N_5202,N_5235);
nor U5300 (N_5300,N_5123,N_5229);
nor U5301 (N_5301,N_5200,N_5148);
nand U5302 (N_5302,N_5157,N_5125);
and U5303 (N_5303,N_5155,N_5175);
nand U5304 (N_5304,N_5248,N_5116);
nor U5305 (N_5305,N_5189,N_5243);
or U5306 (N_5306,N_5180,N_5121);
nand U5307 (N_5307,N_5151,N_5211);
and U5308 (N_5308,N_5104,N_5210);
nor U5309 (N_5309,N_5196,N_5158);
and U5310 (N_5310,N_5244,N_5110);
nand U5311 (N_5311,N_5212,N_5153);
nand U5312 (N_5312,N_5117,N_5226);
nor U5313 (N_5313,N_5102,N_5232);
xnor U5314 (N_5314,N_5159,N_5162);
and U5315 (N_5315,N_5179,N_5234);
or U5316 (N_5316,N_5146,N_5163);
nand U5317 (N_5317,N_5161,N_5135);
nand U5318 (N_5318,N_5114,N_5183);
nand U5319 (N_5319,N_5112,N_5136);
and U5320 (N_5320,N_5142,N_5218);
nand U5321 (N_5321,N_5188,N_5130);
nand U5322 (N_5322,N_5213,N_5245);
nand U5323 (N_5323,N_5208,N_5105);
nand U5324 (N_5324,N_5238,N_5139);
or U5325 (N_5325,N_5236,N_5146);
xor U5326 (N_5326,N_5162,N_5212);
or U5327 (N_5327,N_5199,N_5110);
nor U5328 (N_5328,N_5171,N_5181);
or U5329 (N_5329,N_5205,N_5110);
or U5330 (N_5330,N_5195,N_5248);
and U5331 (N_5331,N_5195,N_5234);
nor U5332 (N_5332,N_5194,N_5139);
nand U5333 (N_5333,N_5203,N_5105);
xor U5334 (N_5334,N_5245,N_5179);
and U5335 (N_5335,N_5135,N_5185);
and U5336 (N_5336,N_5131,N_5180);
or U5337 (N_5337,N_5220,N_5200);
nand U5338 (N_5338,N_5134,N_5161);
or U5339 (N_5339,N_5135,N_5192);
nor U5340 (N_5340,N_5108,N_5117);
and U5341 (N_5341,N_5203,N_5226);
nand U5342 (N_5342,N_5150,N_5237);
or U5343 (N_5343,N_5131,N_5106);
nor U5344 (N_5344,N_5205,N_5100);
and U5345 (N_5345,N_5206,N_5193);
nand U5346 (N_5346,N_5142,N_5220);
or U5347 (N_5347,N_5169,N_5100);
xnor U5348 (N_5348,N_5199,N_5173);
or U5349 (N_5349,N_5168,N_5142);
and U5350 (N_5350,N_5190,N_5162);
nor U5351 (N_5351,N_5134,N_5242);
nor U5352 (N_5352,N_5128,N_5224);
nor U5353 (N_5353,N_5223,N_5243);
nor U5354 (N_5354,N_5157,N_5140);
and U5355 (N_5355,N_5104,N_5162);
and U5356 (N_5356,N_5169,N_5121);
nand U5357 (N_5357,N_5215,N_5127);
xor U5358 (N_5358,N_5130,N_5125);
nor U5359 (N_5359,N_5197,N_5228);
nand U5360 (N_5360,N_5224,N_5248);
nor U5361 (N_5361,N_5241,N_5116);
nand U5362 (N_5362,N_5221,N_5187);
nand U5363 (N_5363,N_5222,N_5119);
and U5364 (N_5364,N_5209,N_5169);
or U5365 (N_5365,N_5134,N_5193);
nand U5366 (N_5366,N_5249,N_5168);
or U5367 (N_5367,N_5140,N_5101);
nor U5368 (N_5368,N_5109,N_5112);
and U5369 (N_5369,N_5161,N_5180);
nand U5370 (N_5370,N_5231,N_5112);
or U5371 (N_5371,N_5191,N_5242);
or U5372 (N_5372,N_5112,N_5181);
or U5373 (N_5373,N_5198,N_5226);
and U5374 (N_5374,N_5189,N_5237);
nor U5375 (N_5375,N_5224,N_5131);
xnor U5376 (N_5376,N_5148,N_5101);
xor U5377 (N_5377,N_5192,N_5142);
xor U5378 (N_5378,N_5159,N_5153);
and U5379 (N_5379,N_5183,N_5246);
xor U5380 (N_5380,N_5131,N_5209);
and U5381 (N_5381,N_5223,N_5202);
nor U5382 (N_5382,N_5178,N_5195);
nor U5383 (N_5383,N_5152,N_5195);
xor U5384 (N_5384,N_5185,N_5232);
nand U5385 (N_5385,N_5241,N_5203);
nand U5386 (N_5386,N_5229,N_5126);
nor U5387 (N_5387,N_5211,N_5153);
or U5388 (N_5388,N_5224,N_5225);
nor U5389 (N_5389,N_5177,N_5102);
xnor U5390 (N_5390,N_5202,N_5144);
xnor U5391 (N_5391,N_5206,N_5176);
nor U5392 (N_5392,N_5131,N_5146);
or U5393 (N_5393,N_5161,N_5100);
xnor U5394 (N_5394,N_5116,N_5104);
nand U5395 (N_5395,N_5199,N_5240);
or U5396 (N_5396,N_5153,N_5201);
xor U5397 (N_5397,N_5170,N_5131);
or U5398 (N_5398,N_5123,N_5137);
nor U5399 (N_5399,N_5203,N_5245);
or U5400 (N_5400,N_5250,N_5341);
nor U5401 (N_5401,N_5292,N_5373);
xnor U5402 (N_5402,N_5327,N_5375);
nor U5403 (N_5403,N_5371,N_5272);
nor U5404 (N_5404,N_5259,N_5304);
or U5405 (N_5405,N_5367,N_5344);
and U5406 (N_5406,N_5377,N_5286);
nand U5407 (N_5407,N_5325,N_5295);
and U5408 (N_5408,N_5326,N_5294);
or U5409 (N_5409,N_5330,N_5346);
nand U5410 (N_5410,N_5310,N_5253);
and U5411 (N_5411,N_5313,N_5334);
xnor U5412 (N_5412,N_5335,N_5254);
nand U5413 (N_5413,N_5372,N_5279);
or U5414 (N_5414,N_5257,N_5343);
or U5415 (N_5415,N_5391,N_5317);
and U5416 (N_5416,N_5303,N_5350);
xor U5417 (N_5417,N_5278,N_5352);
or U5418 (N_5418,N_5287,N_5368);
or U5419 (N_5419,N_5282,N_5338);
nand U5420 (N_5420,N_5263,N_5379);
xnor U5421 (N_5421,N_5289,N_5293);
and U5422 (N_5422,N_5322,N_5308);
nor U5423 (N_5423,N_5386,N_5385);
nor U5424 (N_5424,N_5388,N_5281);
nor U5425 (N_5425,N_5273,N_5331);
and U5426 (N_5426,N_5268,N_5356);
xnor U5427 (N_5427,N_5347,N_5353);
nand U5428 (N_5428,N_5261,N_5363);
or U5429 (N_5429,N_5298,N_5328);
nand U5430 (N_5430,N_5323,N_5351);
and U5431 (N_5431,N_5291,N_5258);
and U5432 (N_5432,N_5396,N_5296);
nor U5433 (N_5433,N_5364,N_5290);
xor U5434 (N_5434,N_5288,N_5264);
and U5435 (N_5435,N_5309,N_5321);
nand U5436 (N_5436,N_5384,N_5271);
and U5437 (N_5437,N_5333,N_5398);
xnor U5438 (N_5438,N_5387,N_5252);
nor U5439 (N_5439,N_5359,N_5393);
or U5440 (N_5440,N_5340,N_5284);
nand U5441 (N_5441,N_5262,N_5299);
nor U5442 (N_5442,N_5378,N_5357);
xor U5443 (N_5443,N_5365,N_5280);
and U5444 (N_5444,N_5318,N_5332);
nor U5445 (N_5445,N_5305,N_5306);
nor U5446 (N_5446,N_5320,N_5329);
xor U5447 (N_5447,N_5361,N_5256);
nor U5448 (N_5448,N_5297,N_5337);
nand U5449 (N_5449,N_5369,N_5397);
nor U5450 (N_5450,N_5383,N_5362);
nand U5451 (N_5451,N_5319,N_5349);
nand U5452 (N_5452,N_5266,N_5301);
xor U5453 (N_5453,N_5307,N_5345);
and U5454 (N_5454,N_5392,N_5265);
nand U5455 (N_5455,N_5342,N_5267);
nor U5456 (N_5456,N_5380,N_5390);
and U5457 (N_5457,N_5339,N_5382);
xor U5458 (N_5458,N_5395,N_5389);
and U5459 (N_5459,N_5274,N_5358);
and U5460 (N_5460,N_5314,N_5355);
xnor U5461 (N_5461,N_5366,N_5270);
nor U5462 (N_5462,N_5251,N_5311);
nor U5463 (N_5463,N_5374,N_5285);
and U5464 (N_5464,N_5276,N_5269);
nand U5465 (N_5465,N_5283,N_5277);
nand U5466 (N_5466,N_5399,N_5324);
and U5467 (N_5467,N_5312,N_5302);
or U5468 (N_5468,N_5376,N_5255);
and U5469 (N_5469,N_5336,N_5381);
nor U5470 (N_5470,N_5348,N_5315);
and U5471 (N_5471,N_5316,N_5260);
nand U5472 (N_5472,N_5360,N_5354);
or U5473 (N_5473,N_5275,N_5370);
or U5474 (N_5474,N_5300,N_5394);
or U5475 (N_5475,N_5310,N_5355);
nand U5476 (N_5476,N_5378,N_5262);
and U5477 (N_5477,N_5348,N_5387);
xor U5478 (N_5478,N_5382,N_5254);
or U5479 (N_5479,N_5377,N_5307);
nor U5480 (N_5480,N_5389,N_5263);
and U5481 (N_5481,N_5308,N_5330);
and U5482 (N_5482,N_5382,N_5375);
and U5483 (N_5483,N_5327,N_5293);
nor U5484 (N_5484,N_5358,N_5353);
nor U5485 (N_5485,N_5253,N_5252);
nor U5486 (N_5486,N_5376,N_5377);
nor U5487 (N_5487,N_5362,N_5391);
xnor U5488 (N_5488,N_5398,N_5282);
nand U5489 (N_5489,N_5392,N_5386);
xnor U5490 (N_5490,N_5368,N_5292);
xor U5491 (N_5491,N_5389,N_5281);
nor U5492 (N_5492,N_5335,N_5391);
nand U5493 (N_5493,N_5310,N_5283);
nand U5494 (N_5494,N_5276,N_5302);
nor U5495 (N_5495,N_5394,N_5296);
nor U5496 (N_5496,N_5304,N_5324);
and U5497 (N_5497,N_5266,N_5393);
nor U5498 (N_5498,N_5385,N_5336);
and U5499 (N_5499,N_5288,N_5305);
nor U5500 (N_5500,N_5318,N_5341);
nand U5501 (N_5501,N_5337,N_5280);
xor U5502 (N_5502,N_5371,N_5364);
xor U5503 (N_5503,N_5350,N_5379);
or U5504 (N_5504,N_5375,N_5271);
nor U5505 (N_5505,N_5395,N_5343);
or U5506 (N_5506,N_5384,N_5286);
or U5507 (N_5507,N_5293,N_5254);
nand U5508 (N_5508,N_5280,N_5383);
and U5509 (N_5509,N_5365,N_5326);
and U5510 (N_5510,N_5272,N_5335);
nand U5511 (N_5511,N_5328,N_5349);
nor U5512 (N_5512,N_5251,N_5396);
and U5513 (N_5513,N_5388,N_5293);
nor U5514 (N_5514,N_5362,N_5364);
xnor U5515 (N_5515,N_5365,N_5334);
nor U5516 (N_5516,N_5289,N_5256);
nor U5517 (N_5517,N_5348,N_5304);
or U5518 (N_5518,N_5307,N_5258);
and U5519 (N_5519,N_5313,N_5250);
nor U5520 (N_5520,N_5376,N_5328);
nand U5521 (N_5521,N_5259,N_5359);
xnor U5522 (N_5522,N_5374,N_5328);
nor U5523 (N_5523,N_5298,N_5276);
or U5524 (N_5524,N_5380,N_5372);
and U5525 (N_5525,N_5389,N_5335);
or U5526 (N_5526,N_5387,N_5382);
nand U5527 (N_5527,N_5282,N_5290);
xnor U5528 (N_5528,N_5346,N_5277);
xor U5529 (N_5529,N_5290,N_5373);
nor U5530 (N_5530,N_5363,N_5368);
nand U5531 (N_5531,N_5281,N_5362);
nand U5532 (N_5532,N_5355,N_5335);
nand U5533 (N_5533,N_5265,N_5294);
or U5534 (N_5534,N_5359,N_5374);
nor U5535 (N_5535,N_5333,N_5261);
and U5536 (N_5536,N_5273,N_5377);
or U5537 (N_5537,N_5351,N_5326);
and U5538 (N_5538,N_5267,N_5268);
xnor U5539 (N_5539,N_5267,N_5337);
nor U5540 (N_5540,N_5302,N_5315);
nand U5541 (N_5541,N_5265,N_5326);
nand U5542 (N_5542,N_5259,N_5338);
xor U5543 (N_5543,N_5353,N_5386);
or U5544 (N_5544,N_5250,N_5397);
or U5545 (N_5545,N_5373,N_5309);
or U5546 (N_5546,N_5314,N_5300);
nor U5547 (N_5547,N_5365,N_5277);
xnor U5548 (N_5548,N_5323,N_5287);
or U5549 (N_5549,N_5272,N_5268);
or U5550 (N_5550,N_5486,N_5428);
xnor U5551 (N_5551,N_5535,N_5460);
or U5552 (N_5552,N_5512,N_5465);
nor U5553 (N_5553,N_5422,N_5418);
xor U5554 (N_5554,N_5541,N_5425);
nor U5555 (N_5555,N_5544,N_5493);
nand U5556 (N_5556,N_5522,N_5520);
xor U5557 (N_5557,N_5506,N_5417);
and U5558 (N_5558,N_5497,N_5476);
and U5559 (N_5559,N_5434,N_5549);
nand U5560 (N_5560,N_5433,N_5401);
or U5561 (N_5561,N_5537,N_5431);
and U5562 (N_5562,N_5446,N_5450);
nor U5563 (N_5563,N_5546,N_5441);
and U5564 (N_5564,N_5454,N_5402);
nor U5565 (N_5565,N_5403,N_5490);
nand U5566 (N_5566,N_5468,N_5479);
xor U5567 (N_5567,N_5459,N_5455);
nor U5568 (N_5568,N_5429,N_5464);
nand U5569 (N_5569,N_5426,N_5525);
xnor U5570 (N_5570,N_5534,N_5487);
nor U5571 (N_5571,N_5496,N_5437);
nand U5572 (N_5572,N_5410,N_5444);
nand U5573 (N_5573,N_5538,N_5474);
nor U5574 (N_5574,N_5472,N_5438);
nand U5575 (N_5575,N_5475,N_5469);
or U5576 (N_5576,N_5420,N_5529);
xor U5577 (N_5577,N_5443,N_5415);
xnor U5578 (N_5578,N_5533,N_5408);
and U5579 (N_5579,N_5463,N_5423);
or U5580 (N_5580,N_5482,N_5526);
nor U5581 (N_5581,N_5511,N_5416);
or U5582 (N_5582,N_5405,N_5532);
nand U5583 (N_5583,N_5519,N_5499);
nor U5584 (N_5584,N_5518,N_5409);
nand U5585 (N_5585,N_5500,N_5439);
nor U5586 (N_5586,N_5400,N_5435);
and U5587 (N_5587,N_5461,N_5510);
nor U5588 (N_5588,N_5427,N_5412);
nor U5589 (N_5589,N_5456,N_5473);
and U5590 (N_5590,N_5527,N_5515);
nand U5591 (N_5591,N_5492,N_5502);
nand U5592 (N_5592,N_5507,N_5501);
nor U5593 (N_5593,N_5452,N_5514);
nand U5594 (N_5594,N_5407,N_5543);
and U5595 (N_5595,N_5498,N_5466);
xor U5596 (N_5596,N_5458,N_5489);
xor U5597 (N_5597,N_5513,N_5547);
xnor U5598 (N_5598,N_5545,N_5536);
and U5599 (N_5599,N_5548,N_5508);
xnor U5600 (N_5600,N_5540,N_5424);
or U5601 (N_5601,N_5457,N_5447);
or U5602 (N_5602,N_5503,N_5421);
nand U5603 (N_5603,N_5542,N_5539);
and U5604 (N_5604,N_5523,N_5445);
and U5605 (N_5605,N_5478,N_5432);
nand U5606 (N_5606,N_5430,N_5524);
nand U5607 (N_5607,N_5494,N_5462);
or U5608 (N_5608,N_5521,N_5491);
nand U5609 (N_5609,N_5495,N_5449);
xnor U5610 (N_5610,N_5467,N_5477);
or U5611 (N_5611,N_5436,N_5406);
xor U5612 (N_5612,N_5481,N_5411);
nand U5613 (N_5613,N_5404,N_5470);
and U5614 (N_5614,N_5483,N_5451);
or U5615 (N_5615,N_5517,N_5442);
nand U5616 (N_5616,N_5528,N_5413);
nand U5617 (N_5617,N_5531,N_5480);
nand U5618 (N_5618,N_5530,N_5504);
or U5619 (N_5619,N_5516,N_5505);
nor U5620 (N_5620,N_5440,N_5448);
xor U5621 (N_5621,N_5488,N_5471);
and U5622 (N_5622,N_5414,N_5509);
and U5623 (N_5623,N_5485,N_5453);
or U5624 (N_5624,N_5419,N_5484);
and U5625 (N_5625,N_5425,N_5495);
or U5626 (N_5626,N_5443,N_5525);
and U5627 (N_5627,N_5505,N_5476);
and U5628 (N_5628,N_5498,N_5531);
xnor U5629 (N_5629,N_5414,N_5484);
xor U5630 (N_5630,N_5495,N_5527);
xnor U5631 (N_5631,N_5442,N_5505);
nor U5632 (N_5632,N_5418,N_5466);
xor U5633 (N_5633,N_5465,N_5403);
nand U5634 (N_5634,N_5421,N_5416);
nand U5635 (N_5635,N_5481,N_5488);
or U5636 (N_5636,N_5434,N_5409);
and U5637 (N_5637,N_5476,N_5464);
nand U5638 (N_5638,N_5507,N_5544);
or U5639 (N_5639,N_5534,N_5478);
xor U5640 (N_5640,N_5498,N_5543);
xor U5641 (N_5641,N_5445,N_5415);
nand U5642 (N_5642,N_5545,N_5494);
xor U5643 (N_5643,N_5435,N_5494);
xor U5644 (N_5644,N_5493,N_5425);
xor U5645 (N_5645,N_5521,N_5421);
or U5646 (N_5646,N_5490,N_5458);
and U5647 (N_5647,N_5513,N_5480);
and U5648 (N_5648,N_5538,N_5439);
or U5649 (N_5649,N_5504,N_5435);
and U5650 (N_5650,N_5491,N_5526);
nand U5651 (N_5651,N_5425,N_5481);
xor U5652 (N_5652,N_5542,N_5471);
xnor U5653 (N_5653,N_5508,N_5443);
nand U5654 (N_5654,N_5428,N_5489);
xor U5655 (N_5655,N_5444,N_5503);
xor U5656 (N_5656,N_5408,N_5427);
nor U5657 (N_5657,N_5454,N_5439);
nor U5658 (N_5658,N_5461,N_5408);
nand U5659 (N_5659,N_5489,N_5440);
nor U5660 (N_5660,N_5413,N_5495);
nor U5661 (N_5661,N_5524,N_5538);
or U5662 (N_5662,N_5443,N_5493);
and U5663 (N_5663,N_5465,N_5470);
nor U5664 (N_5664,N_5521,N_5447);
nor U5665 (N_5665,N_5432,N_5450);
or U5666 (N_5666,N_5451,N_5434);
and U5667 (N_5667,N_5469,N_5514);
and U5668 (N_5668,N_5444,N_5431);
nor U5669 (N_5669,N_5417,N_5504);
xnor U5670 (N_5670,N_5405,N_5461);
nand U5671 (N_5671,N_5503,N_5526);
and U5672 (N_5672,N_5468,N_5417);
or U5673 (N_5673,N_5509,N_5517);
or U5674 (N_5674,N_5484,N_5412);
or U5675 (N_5675,N_5442,N_5532);
or U5676 (N_5676,N_5484,N_5430);
or U5677 (N_5677,N_5480,N_5534);
xor U5678 (N_5678,N_5464,N_5462);
xnor U5679 (N_5679,N_5430,N_5450);
nor U5680 (N_5680,N_5478,N_5449);
nor U5681 (N_5681,N_5417,N_5421);
nor U5682 (N_5682,N_5514,N_5543);
or U5683 (N_5683,N_5433,N_5471);
nor U5684 (N_5684,N_5495,N_5544);
or U5685 (N_5685,N_5414,N_5453);
or U5686 (N_5686,N_5460,N_5541);
or U5687 (N_5687,N_5460,N_5441);
or U5688 (N_5688,N_5459,N_5442);
and U5689 (N_5689,N_5433,N_5462);
and U5690 (N_5690,N_5538,N_5500);
nand U5691 (N_5691,N_5484,N_5425);
xor U5692 (N_5692,N_5474,N_5419);
nand U5693 (N_5693,N_5487,N_5432);
nor U5694 (N_5694,N_5538,N_5433);
nor U5695 (N_5695,N_5449,N_5447);
and U5696 (N_5696,N_5488,N_5420);
xnor U5697 (N_5697,N_5480,N_5475);
and U5698 (N_5698,N_5502,N_5432);
nand U5699 (N_5699,N_5483,N_5518);
or U5700 (N_5700,N_5603,N_5660);
xnor U5701 (N_5701,N_5612,N_5601);
nand U5702 (N_5702,N_5652,N_5676);
xnor U5703 (N_5703,N_5677,N_5688);
or U5704 (N_5704,N_5646,N_5566);
and U5705 (N_5705,N_5574,N_5699);
nand U5706 (N_5706,N_5620,N_5696);
and U5707 (N_5707,N_5551,N_5568);
xnor U5708 (N_5708,N_5619,N_5599);
or U5709 (N_5709,N_5689,N_5608);
and U5710 (N_5710,N_5559,N_5591);
nand U5711 (N_5711,N_5665,N_5633);
and U5712 (N_5712,N_5658,N_5655);
nand U5713 (N_5713,N_5663,N_5570);
and U5714 (N_5714,N_5583,N_5640);
and U5715 (N_5715,N_5651,N_5563);
nor U5716 (N_5716,N_5674,N_5616);
nand U5717 (N_5717,N_5664,N_5595);
nor U5718 (N_5718,N_5680,N_5589);
xnor U5719 (N_5719,N_5550,N_5587);
xnor U5720 (N_5720,N_5592,N_5602);
nand U5721 (N_5721,N_5572,N_5683);
or U5722 (N_5722,N_5690,N_5594);
and U5723 (N_5723,N_5637,N_5684);
nand U5724 (N_5724,N_5626,N_5562);
nand U5725 (N_5725,N_5631,N_5695);
or U5726 (N_5726,N_5615,N_5569);
nand U5727 (N_5727,N_5600,N_5634);
and U5728 (N_5728,N_5630,N_5613);
nand U5729 (N_5729,N_5628,N_5649);
xor U5730 (N_5730,N_5596,N_5672);
nand U5731 (N_5731,N_5573,N_5698);
and U5732 (N_5732,N_5641,N_5668);
and U5733 (N_5733,N_5565,N_5555);
and U5734 (N_5734,N_5697,N_5582);
or U5735 (N_5735,N_5597,N_5560);
nand U5736 (N_5736,N_5667,N_5632);
nand U5737 (N_5737,N_5564,N_5686);
nor U5738 (N_5738,N_5627,N_5653);
nand U5739 (N_5739,N_5584,N_5693);
nor U5740 (N_5740,N_5561,N_5575);
and U5741 (N_5741,N_5650,N_5580);
xor U5742 (N_5742,N_5638,N_5687);
xnor U5743 (N_5743,N_5648,N_5553);
and U5744 (N_5744,N_5669,N_5557);
xor U5745 (N_5745,N_5656,N_5552);
nand U5746 (N_5746,N_5643,N_5675);
nand U5747 (N_5747,N_5678,N_5579);
and U5748 (N_5748,N_5654,N_5625);
and U5749 (N_5749,N_5585,N_5621);
nor U5750 (N_5750,N_5682,N_5618);
nor U5751 (N_5751,N_5586,N_5614);
xnor U5752 (N_5752,N_5681,N_5610);
nor U5753 (N_5753,N_5666,N_5611);
and U5754 (N_5754,N_5662,N_5581);
and U5755 (N_5755,N_5644,N_5607);
or U5756 (N_5756,N_5558,N_5685);
nand U5757 (N_5757,N_5571,N_5598);
or U5758 (N_5758,N_5694,N_5673);
xnor U5759 (N_5759,N_5661,N_5554);
or U5760 (N_5760,N_5593,N_5606);
or U5761 (N_5761,N_5636,N_5576);
nand U5762 (N_5762,N_5567,N_5657);
or U5763 (N_5763,N_5556,N_5692);
and U5764 (N_5764,N_5605,N_5691);
and U5765 (N_5765,N_5629,N_5647);
nand U5766 (N_5766,N_5588,N_5671);
and U5767 (N_5767,N_5577,N_5624);
and U5768 (N_5768,N_5622,N_5609);
or U5769 (N_5769,N_5639,N_5659);
xor U5770 (N_5770,N_5617,N_5604);
xnor U5771 (N_5771,N_5578,N_5645);
xor U5772 (N_5772,N_5679,N_5642);
and U5773 (N_5773,N_5590,N_5635);
nor U5774 (N_5774,N_5670,N_5623);
nor U5775 (N_5775,N_5661,N_5572);
and U5776 (N_5776,N_5558,N_5676);
or U5777 (N_5777,N_5685,N_5561);
or U5778 (N_5778,N_5636,N_5607);
or U5779 (N_5779,N_5578,N_5671);
nand U5780 (N_5780,N_5607,N_5551);
and U5781 (N_5781,N_5573,N_5586);
xor U5782 (N_5782,N_5660,N_5611);
and U5783 (N_5783,N_5565,N_5590);
and U5784 (N_5784,N_5694,N_5578);
and U5785 (N_5785,N_5589,N_5553);
nand U5786 (N_5786,N_5584,N_5624);
and U5787 (N_5787,N_5591,N_5628);
xnor U5788 (N_5788,N_5602,N_5614);
xnor U5789 (N_5789,N_5648,N_5666);
or U5790 (N_5790,N_5645,N_5592);
or U5791 (N_5791,N_5674,N_5554);
nand U5792 (N_5792,N_5685,N_5643);
xor U5793 (N_5793,N_5646,N_5619);
nor U5794 (N_5794,N_5591,N_5696);
nor U5795 (N_5795,N_5681,N_5663);
nor U5796 (N_5796,N_5605,N_5648);
or U5797 (N_5797,N_5627,N_5699);
nand U5798 (N_5798,N_5560,N_5624);
and U5799 (N_5799,N_5632,N_5685);
or U5800 (N_5800,N_5629,N_5630);
or U5801 (N_5801,N_5551,N_5682);
xnor U5802 (N_5802,N_5570,N_5696);
nor U5803 (N_5803,N_5697,N_5579);
nor U5804 (N_5804,N_5646,N_5588);
or U5805 (N_5805,N_5565,N_5662);
nor U5806 (N_5806,N_5586,N_5650);
and U5807 (N_5807,N_5698,N_5612);
and U5808 (N_5808,N_5575,N_5674);
and U5809 (N_5809,N_5634,N_5550);
xor U5810 (N_5810,N_5577,N_5696);
nor U5811 (N_5811,N_5651,N_5622);
nor U5812 (N_5812,N_5688,N_5654);
xor U5813 (N_5813,N_5602,N_5604);
or U5814 (N_5814,N_5663,N_5566);
xor U5815 (N_5815,N_5681,N_5568);
nand U5816 (N_5816,N_5614,N_5653);
and U5817 (N_5817,N_5582,N_5656);
or U5818 (N_5818,N_5658,N_5649);
nor U5819 (N_5819,N_5663,N_5632);
nor U5820 (N_5820,N_5563,N_5673);
nor U5821 (N_5821,N_5690,N_5557);
or U5822 (N_5822,N_5561,N_5627);
xnor U5823 (N_5823,N_5681,N_5692);
and U5824 (N_5824,N_5552,N_5604);
xnor U5825 (N_5825,N_5642,N_5581);
xor U5826 (N_5826,N_5697,N_5688);
nand U5827 (N_5827,N_5627,N_5564);
nor U5828 (N_5828,N_5689,N_5682);
and U5829 (N_5829,N_5641,N_5634);
nor U5830 (N_5830,N_5613,N_5632);
nand U5831 (N_5831,N_5603,N_5580);
xor U5832 (N_5832,N_5643,N_5647);
and U5833 (N_5833,N_5666,N_5579);
xnor U5834 (N_5834,N_5659,N_5677);
or U5835 (N_5835,N_5662,N_5558);
or U5836 (N_5836,N_5662,N_5631);
or U5837 (N_5837,N_5649,N_5699);
or U5838 (N_5838,N_5627,N_5698);
or U5839 (N_5839,N_5628,N_5695);
or U5840 (N_5840,N_5615,N_5584);
nor U5841 (N_5841,N_5615,N_5638);
nand U5842 (N_5842,N_5571,N_5639);
nand U5843 (N_5843,N_5601,N_5577);
nor U5844 (N_5844,N_5698,N_5681);
xor U5845 (N_5845,N_5593,N_5579);
or U5846 (N_5846,N_5661,N_5609);
or U5847 (N_5847,N_5556,N_5590);
or U5848 (N_5848,N_5688,N_5683);
xnor U5849 (N_5849,N_5669,N_5698);
nor U5850 (N_5850,N_5767,N_5816);
nor U5851 (N_5851,N_5808,N_5706);
nand U5852 (N_5852,N_5712,N_5805);
and U5853 (N_5853,N_5792,N_5727);
nor U5854 (N_5854,N_5766,N_5705);
nor U5855 (N_5855,N_5783,N_5701);
and U5856 (N_5856,N_5804,N_5787);
nand U5857 (N_5857,N_5715,N_5829);
and U5858 (N_5858,N_5822,N_5745);
and U5859 (N_5859,N_5785,N_5809);
xor U5860 (N_5860,N_5841,N_5832);
xor U5861 (N_5861,N_5790,N_5834);
nor U5862 (N_5862,N_5759,N_5702);
or U5863 (N_5863,N_5716,N_5728);
or U5864 (N_5864,N_5771,N_5833);
and U5865 (N_5865,N_5704,N_5796);
or U5866 (N_5866,N_5773,N_5847);
nor U5867 (N_5867,N_5752,N_5818);
nor U5868 (N_5868,N_5776,N_5733);
and U5869 (N_5869,N_5844,N_5801);
nand U5870 (N_5870,N_5718,N_5837);
and U5871 (N_5871,N_5813,N_5746);
and U5872 (N_5872,N_5772,N_5838);
xnor U5873 (N_5873,N_5764,N_5730);
xnor U5874 (N_5874,N_5800,N_5775);
nor U5875 (N_5875,N_5774,N_5793);
nand U5876 (N_5876,N_5724,N_5794);
and U5877 (N_5877,N_5843,N_5779);
and U5878 (N_5878,N_5781,N_5731);
nor U5879 (N_5879,N_5842,N_5812);
and U5880 (N_5880,N_5825,N_5717);
and U5881 (N_5881,N_5761,N_5788);
xnor U5882 (N_5882,N_5799,N_5748);
nand U5883 (N_5883,N_5720,N_5810);
nor U5884 (N_5884,N_5739,N_5791);
nor U5885 (N_5885,N_5723,N_5738);
nor U5886 (N_5886,N_5732,N_5743);
and U5887 (N_5887,N_5756,N_5711);
xnor U5888 (N_5888,N_5770,N_5769);
nand U5889 (N_5889,N_5725,N_5744);
or U5890 (N_5890,N_5811,N_5747);
and U5891 (N_5891,N_5741,N_5824);
or U5892 (N_5892,N_5814,N_5758);
nand U5893 (N_5893,N_5821,N_5780);
or U5894 (N_5894,N_5707,N_5760);
or U5895 (N_5895,N_5835,N_5802);
xnor U5896 (N_5896,N_5797,N_5839);
nor U5897 (N_5897,N_5806,N_5778);
xor U5898 (N_5898,N_5708,N_5736);
and U5899 (N_5899,N_5710,N_5703);
nor U5900 (N_5900,N_5803,N_5846);
and U5901 (N_5901,N_5765,N_5749);
nand U5902 (N_5902,N_5819,N_5820);
nand U5903 (N_5903,N_5757,N_5795);
or U5904 (N_5904,N_5826,N_5830);
and U5905 (N_5905,N_5709,N_5742);
nor U5906 (N_5906,N_5848,N_5836);
and U5907 (N_5907,N_5849,N_5840);
nand U5908 (N_5908,N_5740,N_5763);
and U5909 (N_5909,N_5729,N_5722);
nor U5910 (N_5910,N_5755,N_5828);
nor U5911 (N_5911,N_5777,N_5789);
and U5912 (N_5912,N_5817,N_5798);
nand U5913 (N_5913,N_5827,N_5831);
nor U5914 (N_5914,N_5845,N_5734);
and U5915 (N_5915,N_5823,N_5807);
nand U5916 (N_5916,N_5753,N_5714);
nand U5917 (N_5917,N_5726,N_5750);
nand U5918 (N_5918,N_5815,N_5737);
or U5919 (N_5919,N_5751,N_5700);
or U5920 (N_5920,N_5782,N_5754);
xnor U5921 (N_5921,N_5784,N_5762);
nand U5922 (N_5922,N_5735,N_5713);
and U5923 (N_5923,N_5786,N_5719);
and U5924 (N_5924,N_5768,N_5721);
nor U5925 (N_5925,N_5840,N_5764);
and U5926 (N_5926,N_5779,N_5710);
nand U5927 (N_5927,N_5830,N_5796);
nand U5928 (N_5928,N_5849,N_5846);
xor U5929 (N_5929,N_5747,N_5725);
nor U5930 (N_5930,N_5795,N_5711);
nor U5931 (N_5931,N_5830,N_5770);
nor U5932 (N_5932,N_5775,N_5761);
and U5933 (N_5933,N_5722,N_5835);
nand U5934 (N_5934,N_5764,N_5722);
and U5935 (N_5935,N_5811,N_5813);
xor U5936 (N_5936,N_5704,N_5794);
or U5937 (N_5937,N_5822,N_5843);
and U5938 (N_5938,N_5730,N_5774);
xnor U5939 (N_5939,N_5818,N_5840);
xor U5940 (N_5940,N_5840,N_5765);
nand U5941 (N_5941,N_5730,N_5765);
or U5942 (N_5942,N_5730,N_5733);
nor U5943 (N_5943,N_5795,N_5827);
or U5944 (N_5944,N_5788,N_5791);
xnor U5945 (N_5945,N_5780,N_5783);
or U5946 (N_5946,N_5833,N_5770);
or U5947 (N_5947,N_5794,N_5727);
nor U5948 (N_5948,N_5783,N_5720);
nor U5949 (N_5949,N_5706,N_5821);
or U5950 (N_5950,N_5780,N_5809);
nand U5951 (N_5951,N_5816,N_5720);
nor U5952 (N_5952,N_5725,N_5844);
xnor U5953 (N_5953,N_5825,N_5758);
nand U5954 (N_5954,N_5778,N_5786);
nand U5955 (N_5955,N_5845,N_5735);
or U5956 (N_5956,N_5757,N_5743);
xnor U5957 (N_5957,N_5841,N_5819);
nor U5958 (N_5958,N_5801,N_5701);
and U5959 (N_5959,N_5759,N_5810);
nand U5960 (N_5960,N_5771,N_5825);
xor U5961 (N_5961,N_5756,N_5770);
xnor U5962 (N_5962,N_5824,N_5787);
and U5963 (N_5963,N_5847,N_5772);
nor U5964 (N_5964,N_5771,N_5795);
nand U5965 (N_5965,N_5808,N_5705);
nor U5966 (N_5966,N_5830,N_5738);
or U5967 (N_5967,N_5751,N_5840);
xnor U5968 (N_5968,N_5708,N_5776);
nand U5969 (N_5969,N_5729,N_5700);
or U5970 (N_5970,N_5793,N_5724);
or U5971 (N_5971,N_5718,N_5830);
or U5972 (N_5972,N_5830,N_5720);
nor U5973 (N_5973,N_5715,N_5736);
and U5974 (N_5974,N_5829,N_5838);
nor U5975 (N_5975,N_5751,N_5750);
or U5976 (N_5976,N_5843,N_5702);
xnor U5977 (N_5977,N_5722,N_5737);
nor U5978 (N_5978,N_5701,N_5815);
nand U5979 (N_5979,N_5811,N_5783);
xor U5980 (N_5980,N_5817,N_5815);
xnor U5981 (N_5981,N_5816,N_5801);
nor U5982 (N_5982,N_5800,N_5741);
xnor U5983 (N_5983,N_5739,N_5732);
and U5984 (N_5984,N_5760,N_5720);
xnor U5985 (N_5985,N_5752,N_5726);
or U5986 (N_5986,N_5823,N_5781);
nand U5987 (N_5987,N_5845,N_5768);
nor U5988 (N_5988,N_5793,N_5790);
xor U5989 (N_5989,N_5714,N_5801);
or U5990 (N_5990,N_5816,N_5744);
and U5991 (N_5991,N_5712,N_5740);
nand U5992 (N_5992,N_5816,N_5811);
and U5993 (N_5993,N_5821,N_5756);
or U5994 (N_5994,N_5784,N_5745);
nand U5995 (N_5995,N_5757,N_5706);
and U5996 (N_5996,N_5706,N_5814);
or U5997 (N_5997,N_5820,N_5766);
nor U5998 (N_5998,N_5732,N_5736);
and U5999 (N_5999,N_5824,N_5712);
or U6000 (N_6000,N_5995,N_5891);
nand U6001 (N_6001,N_5943,N_5866);
nand U6002 (N_6002,N_5966,N_5912);
or U6003 (N_6003,N_5855,N_5944);
nor U6004 (N_6004,N_5996,N_5998);
or U6005 (N_6005,N_5901,N_5962);
nor U6006 (N_6006,N_5868,N_5917);
and U6007 (N_6007,N_5985,N_5940);
nor U6008 (N_6008,N_5880,N_5864);
nand U6009 (N_6009,N_5920,N_5883);
or U6010 (N_6010,N_5911,N_5862);
or U6011 (N_6011,N_5961,N_5914);
xor U6012 (N_6012,N_5982,N_5959);
xor U6013 (N_6013,N_5861,N_5858);
and U6014 (N_6014,N_5930,N_5978);
and U6015 (N_6015,N_5977,N_5976);
or U6016 (N_6016,N_5931,N_5860);
or U6017 (N_6017,N_5980,N_5878);
nor U6018 (N_6018,N_5882,N_5946);
and U6019 (N_6019,N_5863,N_5885);
xor U6020 (N_6020,N_5952,N_5865);
and U6021 (N_6021,N_5884,N_5850);
or U6022 (N_6022,N_5929,N_5945);
xor U6023 (N_6023,N_5898,N_5951);
and U6024 (N_6024,N_5942,N_5876);
nor U6025 (N_6025,N_5986,N_5937);
and U6026 (N_6026,N_5993,N_5974);
or U6027 (N_6027,N_5875,N_5870);
xnor U6028 (N_6028,N_5892,N_5889);
xnor U6029 (N_6029,N_5958,N_5902);
xor U6030 (N_6030,N_5949,N_5894);
nor U6031 (N_6031,N_5893,N_5933);
xnor U6032 (N_6032,N_5923,N_5913);
or U6033 (N_6033,N_5904,N_5886);
xor U6034 (N_6034,N_5910,N_5896);
nand U6035 (N_6035,N_5979,N_5927);
xor U6036 (N_6036,N_5965,N_5992);
nor U6037 (N_6037,N_5888,N_5874);
or U6038 (N_6038,N_5997,N_5887);
xnor U6039 (N_6039,N_5954,N_5922);
xor U6040 (N_6040,N_5881,N_5903);
nor U6041 (N_6041,N_5932,N_5924);
nor U6042 (N_6042,N_5941,N_5999);
nor U6043 (N_6043,N_5950,N_5955);
or U6044 (N_6044,N_5851,N_5934);
or U6045 (N_6045,N_5975,N_5857);
nand U6046 (N_6046,N_5854,N_5908);
nor U6047 (N_6047,N_5915,N_5988);
xor U6048 (N_6048,N_5921,N_5967);
nand U6049 (N_6049,N_5947,N_5928);
nand U6050 (N_6050,N_5968,N_5897);
nor U6051 (N_6051,N_5879,N_5925);
or U6052 (N_6052,N_5948,N_5853);
or U6053 (N_6053,N_5972,N_5926);
xor U6054 (N_6054,N_5873,N_5990);
nand U6055 (N_6055,N_5916,N_5877);
xor U6056 (N_6056,N_5869,N_5935);
or U6057 (N_6057,N_5984,N_5994);
xnor U6058 (N_6058,N_5987,N_5953);
or U6059 (N_6059,N_5960,N_5852);
nand U6060 (N_6060,N_5859,N_5969);
nor U6061 (N_6061,N_5970,N_5964);
and U6062 (N_6062,N_5905,N_5907);
or U6063 (N_6063,N_5971,N_5973);
xor U6064 (N_6064,N_5856,N_5957);
xnor U6065 (N_6065,N_5906,N_5899);
xnor U6066 (N_6066,N_5983,N_5939);
nor U6067 (N_6067,N_5919,N_5963);
nor U6068 (N_6068,N_5991,N_5956);
nor U6069 (N_6069,N_5895,N_5872);
or U6070 (N_6070,N_5890,N_5900);
and U6071 (N_6071,N_5938,N_5981);
or U6072 (N_6072,N_5989,N_5871);
and U6073 (N_6073,N_5918,N_5936);
nor U6074 (N_6074,N_5867,N_5909);
xnor U6075 (N_6075,N_5868,N_5990);
or U6076 (N_6076,N_5858,N_5975);
or U6077 (N_6077,N_5975,N_5996);
xor U6078 (N_6078,N_5989,N_5908);
nor U6079 (N_6079,N_5912,N_5952);
nand U6080 (N_6080,N_5987,N_5948);
xor U6081 (N_6081,N_5998,N_5897);
nand U6082 (N_6082,N_5880,N_5870);
nand U6083 (N_6083,N_5857,N_5950);
nand U6084 (N_6084,N_5858,N_5916);
and U6085 (N_6085,N_5951,N_5964);
nor U6086 (N_6086,N_5939,N_5899);
xor U6087 (N_6087,N_5880,N_5855);
nand U6088 (N_6088,N_5994,N_5961);
and U6089 (N_6089,N_5855,N_5898);
or U6090 (N_6090,N_5894,N_5943);
nand U6091 (N_6091,N_5855,N_5867);
nor U6092 (N_6092,N_5952,N_5979);
nand U6093 (N_6093,N_5983,N_5957);
xor U6094 (N_6094,N_5884,N_5881);
and U6095 (N_6095,N_5895,N_5933);
and U6096 (N_6096,N_5889,N_5859);
xor U6097 (N_6097,N_5982,N_5921);
or U6098 (N_6098,N_5992,N_5967);
and U6099 (N_6099,N_5973,N_5863);
xnor U6100 (N_6100,N_5904,N_5911);
and U6101 (N_6101,N_5931,N_5872);
or U6102 (N_6102,N_5980,N_5950);
xnor U6103 (N_6103,N_5912,N_5855);
or U6104 (N_6104,N_5954,N_5987);
or U6105 (N_6105,N_5881,N_5919);
nor U6106 (N_6106,N_5890,N_5898);
xor U6107 (N_6107,N_5886,N_5905);
nor U6108 (N_6108,N_5918,N_5952);
xnor U6109 (N_6109,N_5876,N_5895);
and U6110 (N_6110,N_5857,N_5997);
xor U6111 (N_6111,N_5852,N_5890);
or U6112 (N_6112,N_5987,N_5883);
or U6113 (N_6113,N_5910,N_5898);
xor U6114 (N_6114,N_5957,N_5893);
nand U6115 (N_6115,N_5953,N_5873);
or U6116 (N_6116,N_5904,N_5853);
and U6117 (N_6117,N_5903,N_5852);
xnor U6118 (N_6118,N_5944,N_5921);
xnor U6119 (N_6119,N_5891,N_5859);
xor U6120 (N_6120,N_5879,N_5953);
or U6121 (N_6121,N_5934,N_5891);
nand U6122 (N_6122,N_5873,N_5954);
xnor U6123 (N_6123,N_5885,N_5901);
or U6124 (N_6124,N_5949,N_5966);
or U6125 (N_6125,N_5880,N_5872);
nand U6126 (N_6126,N_5948,N_5980);
and U6127 (N_6127,N_5865,N_5904);
and U6128 (N_6128,N_5911,N_5924);
and U6129 (N_6129,N_5901,N_5922);
nor U6130 (N_6130,N_5905,N_5879);
and U6131 (N_6131,N_5912,N_5968);
nor U6132 (N_6132,N_5987,N_5867);
and U6133 (N_6133,N_5995,N_5897);
nor U6134 (N_6134,N_5926,N_5870);
xor U6135 (N_6135,N_5927,N_5911);
and U6136 (N_6136,N_5955,N_5915);
xnor U6137 (N_6137,N_5929,N_5944);
xor U6138 (N_6138,N_5998,N_5971);
nand U6139 (N_6139,N_5980,N_5874);
nand U6140 (N_6140,N_5980,N_5934);
nor U6141 (N_6141,N_5949,N_5908);
xor U6142 (N_6142,N_5871,N_5860);
nand U6143 (N_6143,N_5961,N_5949);
and U6144 (N_6144,N_5963,N_5854);
nor U6145 (N_6145,N_5887,N_5953);
nand U6146 (N_6146,N_5975,N_5913);
nand U6147 (N_6147,N_5979,N_5989);
nand U6148 (N_6148,N_5871,N_5893);
nand U6149 (N_6149,N_5871,N_5921);
or U6150 (N_6150,N_6055,N_6087);
and U6151 (N_6151,N_6064,N_6081);
or U6152 (N_6152,N_6024,N_6060);
xnor U6153 (N_6153,N_6083,N_6010);
or U6154 (N_6154,N_6053,N_6144);
nor U6155 (N_6155,N_6124,N_6148);
and U6156 (N_6156,N_6136,N_6098);
nor U6157 (N_6157,N_6044,N_6086);
and U6158 (N_6158,N_6135,N_6054);
or U6159 (N_6159,N_6074,N_6108);
and U6160 (N_6160,N_6132,N_6000);
and U6161 (N_6161,N_6121,N_6014);
or U6162 (N_6162,N_6107,N_6017);
or U6163 (N_6163,N_6113,N_6034);
xor U6164 (N_6164,N_6122,N_6067);
or U6165 (N_6165,N_6048,N_6037);
xnor U6166 (N_6166,N_6123,N_6011);
xnor U6167 (N_6167,N_6103,N_6105);
and U6168 (N_6168,N_6147,N_6004);
or U6169 (N_6169,N_6027,N_6025);
or U6170 (N_6170,N_6005,N_6120);
nor U6171 (N_6171,N_6049,N_6063);
and U6172 (N_6172,N_6021,N_6131);
or U6173 (N_6173,N_6106,N_6045);
or U6174 (N_6174,N_6149,N_6006);
xnor U6175 (N_6175,N_6030,N_6142);
xor U6176 (N_6176,N_6146,N_6042);
nand U6177 (N_6177,N_6057,N_6051);
xor U6178 (N_6178,N_6101,N_6127);
nand U6179 (N_6179,N_6039,N_6077);
nand U6180 (N_6180,N_6009,N_6016);
xnor U6181 (N_6181,N_6084,N_6038);
and U6182 (N_6182,N_6088,N_6036);
and U6183 (N_6183,N_6085,N_6073);
and U6184 (N_6184,N_6007,N_6001);
nor U6185 (N_6185,N_6035,N_6075);
xnor U6186 (N_6186,N_6046,N_6032);
xor U6187 (N_6187,N_6133,N_6110);
and U6188 (N_6188,N_6056,N_6080);
nor U6189 (N_6189,N_6043,N_6118);
nand U6190 (N_6190,N_6140,N_6109);
nand U6191 (N_6191,N_6052,N_6097);
and U6192 (N_6192,N_6090,N_6058);
xnor U6193 (N_6193,N_6066,N_6134);
xnor U6194 (N_6194,N_6031,N_6089);
xnor U6195 (N_6195,N_6041,N_6141);
or U6196 (N_6196,N_6099,N_6104);
xor U6197 (N_6197,N_6139,N_6119);
nand U6198 (N_6198,N_6019,N_6069);
or U6199 (N_6199,N_6128,N_6026);
and U6200 (N_6200,N_6023,N_6003);
xnor U6201 (N_6201,N_6143,N_6070);
xor U6202 (N_6202,N_6130,N_6145);
nor U6203 (N_6203,N_6062,N_6137);
or U6204 (N_6204,N_6008,N_6076);
xor U6205 (N_6205,N_6112,N_6068);
nand U6206 (N_6206,N_6072,N_6013);
nor U6207 (N_6207,N_6092,N_6115);
and U6208 (N_6208,N_6078,N_6071);
or U6209 (N_6209,N_6022,N_6015);
or U6210 (N_6210,N_6020,N_6061);
xor U6211 (N_6211,N_6033,N_6029);
nand U6212 (N_6212,N_6129,N_6093);
nor U6213 (N_6213,N_6138,N_6111);
or U6214 (N_6214,N_6126,N_6018);
and U6215 (N_6215,N_6040,N_6117);
nand U6216 (N_6216,N_6047,N_6102);
nand U6217 (N_6217,N_6065,N_6116);
and U6218 (N_6218,N_6125,N_6002);
or U6219 (N_6219,N_6091,N_6012);
or U6220 (N_6220,N_6059,N_6028);
xnor U6221 (N_6221,N_6050,N_6082);
nand U6222 (N_6222,N_6095,N_6094);
nor U6223 (N_6223,N_6079,N_6114);
nand U6224 (N_6224,N_6100,N_6096);
or U6225 (N_6225,N_6054,N_6104);
xor U6226 (N_6226,N_6088,N_6143);
or U6227 (N_6227,N_6131,N_6136);
nand U6228 (N_6228,N_6089,N_6084);
nand U6229 (N_6229,N_6079,N_6017);
xor U6230 (N_6230,N_6102,N_6146);
xnor U6231 (N_6231,N_6040,N_6123);
nand U6232 (N_6232,N_6033,N_6094);
or U6233 (N_6233,N_6128,N_6002);
nand U6234 (N_6234,N_6042,N_6078);
nand U6235 (N_6235,N_6082,N_6032);
xnor U6236 (N_6236,N_6058,N_6008);
or U6237 (N_6237,N_6076,N_6025);
and U6238 (N_6238,N_6038,N_6148);
or U6239 (N_6239,N_6107,N_6038);
and U6240 (N_6240,N_6086,N_6054);
xnor U6241 (N_6241,N_6047,N_6058);
or U6242 (N_6242,N_6007,N_6106);
nor U6243 (N_6243,N_6105,N_6022);
nor U6244 (N_6244,N_6087,N_6032);
or U6245 (N_6245,N_6095,N_6007);
nand U6246 (N_6246,N_6109,N_6120);
nand U6247 (N_6247,N_6129,N_6090);
or U6248 (N_6248,N_6031,N_6133);
nand U6249 (N_6249,N_6050,N_6016);
and U6250 (N_6250,N_6141,N_6039);
nand U6251 (N_6251,N_6134,N_6042);
xor U6252 (N_6252,N_6043,N_6132);
xnor U6253 (N_6253,N_6007,N_6033);
and U6254 (N_6254,N_6100,N_6099);
or U6255 (N_6255,N_6007,N_6056);
or U6256 (N_6256,N_6101,N_6116);
nand U6257 (N_6257,N_6116,N_6017);
and U6258 (N_6258,N_6022,N_6122);
or U6259 (N_6259,N_6149,N_6091);
or U6260 (N_6260,N_6004,N_6106);
and U6261 (N_6261,N_6102,N_6034);
and U6262 (N_6262,N_6088,N_6005);
or U6263 (N_6263,N_6024,N_6033);
xor U6264 (N_6264,N_6051,N_6021);
xor U6265 (N_6265,N_6060,N_6093);
nor U6266 (N_6266,N_6083,N_6094);
nor U6267 (N_6267,N_6070,N_6148);
nor U6268 (N_6268,N_6081,N_6069);
xnor U6269 (N_6269,N_6033,N_6043);
nand U6270 (N_6270,N_6051,N_6117);
nand U6271 (N_6271,N_6032,N_6111);
xnor U6272 (N_6272,N_6096,N_6101);
nand U6273 (N_6273,N_6144,N_6057);
or U6274 (N_6274,N_6075,N_6066);
nor U6275 (N_6275,N_6136,N_6046);
xnor U6276 (N_6276,N_6058,N_6060);
nand U6277 (N_6277,N_6101,N_6059);
nand U6278 (N_6278,N_6103,N_6031);
and U6279 (N_6279,N_6012,N_6144);
xnor U6280 (N_6280,N_6019,N_6017);
nand U6281 (N_6281,N_6146,N_6043);
xor U6282 (N_6282,N_6088,N_6123);
xor U6283 (N_6283,N_6117,N_6100);
or U6284 (N_6284,N_6070,N_6117);
and U6285 (N_6285,N_6121,N_6113);
and U6286 (N_6286,N_6137,N_6052);
and U6287 (N_6287,N_6098,N_6107);
xnor U6288 (N_6288,N_6095,N_6060);
nand U6289 (N_6289,N_6062,N_6009);
xnor U6290 (N_6290,N_6031,N_6099);
nand U6291 (N_6291,N_6075,N_6052);
and U6292 (N_6292,N_6013,N_6102);
or U6293 (N_6293,N_6009,N_6082);
and U6294 (N_6294,N_6085,N_6062);
nor U6295 (N_6295,N_6040,N_6074);
nor U6296 (N_6296,N_6003,N_6032);
or U6297 (N_6297,N_6000,N_6063);
or U6298 (N_6298,N_6141,N_6074);
and U6299 (N_6299,N_6121,N_6036);
and U6300 (N_6300,N_6156,N_6241);
and U6301 (N_6301,N_6258,N_6245);
nor U6302 (N_6302,N_6223,N_6247);
nand U6303 (N_6303,N_6184,N_6185);
xor U6304 (N_6304,N_6227,N_6262);
nor U6305 (N_6305,N_6165,N_6292);
xor U6306 (N_6306,N_6238,N_6280);
nor U6307 (N_6307,N_6256,N_6270);
or U6308 (N_6308,N_6186,N_6281);
nand U6309 (N_6309,N_6176,N_6161);
xnor U6310 (N_6310,N_6198,N_6208);
nor U6311 (N_6311,N_6298,N_6170);
or U6312 (N_6312,N_6248,N_6171);
nand U6313 (N_6313,N_6154,N_6213);
or U6314 (N_6314,N_6246,N_6288);
xnor U6315 (N_6315,N_6267,N_6285);
or U6316 (N_6316,N_6221,N_6204);
or U6317 (N_6317,N_6210,N_6231);
and U6318 (N_6318,N_6163,N_6181);
nor U6319 (N_6319,N_6230,N_6274);
nand U6320 (N_6320,N_6155,N_6272);
xor U6321 (N_6321,N_6286,N_6196);
nand U6322 (N_6322,N_6158,N_6266);
nor U6323 (N_6323,N_6242,N_6278);
nand U6324 (N_6324,N_6157,N_6260);
and U6325 (N_6325,N_6239,N_6166);
and U6326 (N_6326,N_6287,N_6192);
xor U6327 (N_6327,N_6202,N_6214);
and U6328 (N_6328,N_6261,N_6273);
nand U6329 (N_6329,N_6180,N_6182);
nand U6330 (N_6330,N_6264,N_6199);
nand U6331 (N_6331,N_6159,N_6265);
nand U6332 (N_6332,N_6240,N_6193);
or U6333 (N_6333,N_6234,N_6206);
and U6334 (N_6334,N_6294,N_6191);
nor U6335 (N_6335,N_6277,N_6216);
nand U6336 (N_6336,N_6252,N_6271);
xor U6337 (N_6337,N_6228,N_6195);
xnor U6338 (N_6338,N_6254,N_6177);
and U6339 (N_6339,N_6224,N_6284);
or U6340 (N_6340,N_6168,N_6189);
xnor U6341 (N_6341,N_6212,N_6297);
xor U6342 (N_6342,N_6253,N_6174);
nor U6343 (N_6343,N_6290,N_6237);
nand U6344 (N_6344,N_6222,N_6211);
xor U6345 (N_6345,N_6226,N_6218);
xnor U6346 (N_6346,N_6244,N_6209);
nand U6347 (N_6347,N_6236,N_6203);
nand U6348 (N_6348,N_6250,N_6200);
or U6349 (N_6349,N_6289,N_6233);
xnor U6350 (N_6350,N_6164,N_6295);
xnor U6351 (N_6351,N_6172,N_6291);
or U6352 (N_6352,N_6251,N_6197);
and U6353 (N_6353,N_6150,N_6268);
xor U6354 (N_6354,N_6178,N_6169);
nor U6355 (N_6355,N_6263,N_6219);
and U6356 (N_6356,N_6215,N_6243);
or U6357 (N_6357,N_6282,N_6160);
and U6358 (N_6358,N_6187,N_6293);
nor U6359 (N_6359,N_6207,N_6279);
nor U6360 (N_6360,N_6188,N_6205);
and U6361 (N_6361,N_6257,N_6151);
nand U6362 (N_6362,N_6173,N_6275);
xnor U6363 (N_6363,N_6194,N_6229);
or U6364 (N_6364,N_6162,N_6179);
xor U6365 (N_6365,N_6235,N_6201);
and U6366 (N_6366,N_6259,N_6183);
nand U6367 (N_6367,N_6153,N_6299);
and U6368 (N_6368,N_6249,N_6217);
nand U6369 (N_6369,N_6255,N_6152);
nor U6370 (N_6370,N_6225,N_6190);
xnor U6371 (N_6371,N_6269,N_6232);
nand U6372 (N_6372,N_6167,N_6276);
xnor U6373 (N_6373,N_6283,N_6220);
or U6374 (N_6374,N_6175,N_6296);
or U6375 (N_6375,N_6198,N_6266);
or U6376 (N_6376,N_6191,N_6261);
and U6377 (N_6377,N_6218,N_6235);
and U6378 (N_6378,N_6244,N_6237);
or U6379 (N_6379,N_6197,N_6291);
and U6380 (N_6380,N_6167,N_6229);
or U6381 (N_6381,N_6215,N_6270);
xor U6382 (N_6382,N_6250,N_6162);
xnor U6383 (N_6383,N_6234,N_6163);
and U6384 (N_6384,N_6203,N_6278);
and U6385 (N_6385,N_6299,N_6263);
and U6386 (N_6386,N_6181,N_6290);
xor U6387 (N_6387,N_6251,N_6254);
and U6388 (N_6388,N_6170,N_6285);
or U6389 (N_6389,N_6201,N_6161);
nor U6390 (N_6390,N_6260,N_6291);
or U6391 (N_6391,N_6206,N_6223);
and U6392 (N_6392,N_6192,N_6249);
or U6393 (N_6393,N_6272,N_6255);
nand U6394 (N_6394,N_6271,N_6181);
and U6395 (N_6395,N_6291,N_6238);
nor U6396 (N_6396,N_6269,N_6154);
and U6397 (N_6397,N_6216,N_6184);
nor U6398 (N_6398,N_6258,N_6166);
and U6399 (N_6399,N_6155,N_6256);
and U6400 (N_6400,N_6217,N_6216);
xor U6401 (N_6401,N_6286,N_6170);
nand U6402 (N_6402,N_6263,N_6213);
and U6403 (N_6403,N_6207,N_6260);
nand U6404 (N_6404,N_6165,N_6202);
or U6405 (N_6405,N_6210,N_6239);
xnor U6406 (N_6406,N_6153,N_6154);
nor U6407 (N_6407,N_6212,N_6184);
xor U6408 (N_6408,N_6295,N_6226);
nor U6409 (N_6409,N_6258,N_6187);
and U6410 (N_6410,N_6151,N_6198);
or U6411 (N_6411,N_6158,N_6209);
or U6412 (N_6412,N_6173,N_6254);
nand U6413 (N_6413,N_6255,N_6168);
and U6414 (N_6414,N_6156,N_6264);
and U6415 (N_6415,N_6287,N_6201);
or U6416 (N_6416,N_6205,N_6290);
and U6417 (N_6417,N_6168,N_6273);
or U6418 (N_6418,N_6157,N_6249);
xnor U6419 (N_6419,N_6178,N_6255);
xnor U6420 (N_6420,N_6294,N_6200);
xnor U6421 (N_6421,N_6181,N_6224);
nor U6422 (N_6422,N_6211,N_6150);
nor U6423 (N_6423,N_6199,N_6293);
and U6424 (N_6424,N_6165,N_6266);
or U6425 (N_6425,N_6273,N_6175);
nand U6426 (N_6426,N_6183,N_6214);
xor U6427 (N_6427,N_6160,N_6297);
xnor U6428 (N_6428,N_6283,N_6266);
xor U6429 (N_6429,N_6269,N_6272);
nand U6430 (N_6430,N_6288,N_6284);
xnor U6431 (N_6431,N_6288,N_6289);
nand U6432 (N_6432,N_6223,N_6245);
nand U6433 (N_6433,N_6159,N_6154);
nand U6434 (N_6434,N_6270,N_6296);
nor U6435 (N_6435,N_6155,N_6170);
xnor U6436 (N_6436,N_6173,N_6280);
nor U6437 (N_6437,N_6187,N_6228);
or U6438 (N_6438,N_6176,N_6286);
and U6439 (N_6439,N_6228,N_6192);
nand U6440 (N_6440,N_6210,N_6233);
or U6441 (N_6441,N_6252,N_6266);
nor U6442 (N_6442,N_6237,N_6166);
nor U6443 (N_6443,N_6240,N_6174);
nand U6444 (N_6444,N_6242,N_6212);
and U6445 (N_6445,N_6231,N_6157);
and U6446 (N_6446,N_6158,N_6286);
nor U6447 (N_6447,N_6293,N_6261);
xnor U6448 (N_6448,N_6150,N_6197);
nand U6449 (N_6449,N_6235,N_6275);
or U6450 (N_6450,N_6393,N_6385);
nor U6451 (N_6451,N_6443,N_6383);
or U6452 (N_6452,N_6389,N_6426);
or U6453 (N_6453,N_6362,N_6449);
nand U6454 (N_6454,N_6441,N_6367);
and U6455 (N_6455,N_6388,N_6430);
and U6456 (N_6456,N_6399,N_6360);
xnor U6457 (N_6457,N_6315,N_6419);
xnor U6458 (N_6458,N_6414,N_6342);
nor U6459 (N_6459,N_6378,N_6312);
or U6460 (N_6460,N_6345,N_6358);
or U6461 (N_6461,N_6346,N_6369);
xor U6462 (N_6462,N_6421,N_6311);
and U6463 (N_6463,N_6347,N_6410);
nor U6464 (N_6464,N_6371,N_6364);
or U6465 (N_6465,N_6349,N_6304);
nand U6466 (N_6466,N_6340,N_6350);
xor U6467 (N_6467,N_6444,N_6357);
nand U6468 (N_6468,N_6394,N_6391);
or U6469 (N_6469,N_6417,N_6445);
and U6470 (N_6470,N_6431,N_6423);
xor U6471 (N_6471,N_6386,N_6302);
nor U6472 (N_6472,N_6435,N_6396);
nor U6473 (N_6473,N_6334,N_6353);
nand U6474 (N_6474,N_6406,N_6361);
nand U6475 (N_6475,N_6306,N_6384);
nor U6476 (N_6476,N_6440,N_6381);
nand U6477 (N_6477,N_6438,N_6398);
nand U6478 (N_6478,N_6442,N_6429);
nand U6479 (N_6479,N_6352,N_6338);
nand U6480 (N_6480,N_6310,N_6425);
nor U6481 (N_6481,N_6328,N_6412);
xor U6482 (N_6482,N_6374,N_6330);
nor U6483 (N_6483,N_6355,N_6376);
or U6484 (N_6484,N_6408,N_6401);
xor U6485 (N_6485,N_6303,N_6335);
or U6486 (N_6486,N_6317,N_6395);
nand U6487 (N_6487,N_6427,N_6411);
xnor U6488 (N_6488,N_6446,N_6326);
nand U6489 (N_6489,N_6404,N_6321);
xor U6490 (N_6490,N_6382,N_6424);
or U6491 (N_6491,N_6403,N_6325);
nor U6492 (N_6492,N_6400,N_6316);
xnor U6493 (N_6493,N_6373,N_6343);
xnor U6494 (N_6494,N_6333,N_6415);
xnor U6495 (N_6495,N_6405,N_6448);
nand U6496 (N_6496,N_6324,N_6307);
or U6497 (N_6497,N_6308,N_6387);
or U6498 (N_6498,N_6344,N_6331);
xor U6499 (N_6499,N_6420,N_6436);
nand U6500 (N_6500,N_6318,N_6377);
nor U6501 (N_6501,N_6301,N_6434);
or U6502 (N_6502,N_6323,N_6329);
and U6503 (N_6503,N_6314,N_6337);
and U6504 (N_6504,N_6397,N_6305);
nand U6505 (N_6505,N_6413,N_6422);
nor U6506 (N_6506,N_6359,N_6375);
nor U6507 (N_6507,N_6416,N_6392);
nor U6508 (N_6508,N_6351,N_6366);
xnor U6509 (N_6509,N_6327,N_6368);
xnor U6510 (N_6510,N_6447,N_6339);
xnor U6511 (N_6511,N_6370,N_6356);
or U6512 (N_6512,N_6428,N_6332);
nand U6513 (N_6513,N_6309,N_6363);
or U6514 (N_6514,N_6319,N_6390);
nor U6515 (N_6515,N_6348,N_6432);
xnor U6516 (N_6516,N_6439,N_6379);
nor U6517 (N_6517,N_6322,N_6372);
xor U6518 (N_6518,N_6320,N_6433);
nand U6519 (N_6519,N_6365,N_6418);
nor U6520 (N_6520,N_6313,N_6336);
nand U6521 (N_6521,N_6402,N_6354);
nand U6522 (N_6522,N_6300,N_6437);
and U6523 (N_6523,N_6380,N_6409);
xnor U6524 (N_6524,N_6341,N_6407);
nor U6525 (N_6525,N_6408,N_6419);
or U6526 (N_6526,N_6407,N_6426);
nand U6527 (N_6527,N_6432,N_6373);
nand U6528 (N_6528,N_6329,N_6419);
nand U6529 (N_6529,N_6429,N_6308);
and U6530 (N_6530,N_6301,N_6395);
nand U6531 (N_6531,N_6410,N_6363);
nand U6532 (N_6532,N_6418,N_6417);
xor U6533 (N_6533,N_6447,N_6436);
nand U6534 (N_6534,N_6362,N_6308);
nor U6535 (N_6535,N_6439,N_6324);
nor U6536 (N_6536,N_6317,N_6441);
xor U6537 (N_6537,N_6387,N_6346);
xor U6538 (N_6538,N_6431,N_6358);
and U6539 (N_6539,N_6332,N_6405);
xnor U6540 (N_6540,N_6387,N_6391);
nand U6541 (N_6541,N_6441,N_6343);
nand U6542 (N_6542,N_6341,N_6412);
and U6543 (N_6543,N_6308,N_6352);
xor U6544 (N_6544,N_6388,N_6413);
and U6545 (N_6545,N_6396,N_6401);
and U6546 (N_6546,N_6418,N_6326);
and U6547 (N_6547,N_6305,N_6388);
nor U6548 (N_6548,N_6362,N_6419);
xnor U6549 (N_6549,N_6329,N_6379);
and U6550 (N_6550,N_6365,N_6321);
xor U6551 (N_6551,N_6317,N_6448);
xnor U6552 (N_6552,N_6442,N_6379);
nand U6553 (N_6553,N_6374,N_6392);
nor U6554 (N_6554,N_6397,N_6423);
nand U6555 (N_6555,N_6327,N_6415);
nor U6556 (N_6556,N_6358,N_6409);
nor U6557 (N_6557,N_6354,N_6405);
nand U6558 (N_6558,N_6349,N_6370);
nand U6559 (N_6559,N_6323,N_6386);
nor U6560 (N_6560,N_6325,N_6360);
nor U6561 (N_6561,N_6349,N_6323);
or U6562 (N_6562,N_6329,N_6338);
nand U6563 (N_6563,N_6309,N_6431);
nor U6564 (N_6564,N_6393,N_6312);
nor U6565 (N_6565,N_6336,N_6448);
xor U6566 (N_6566,N_6405,N_6427);
and U6567 (N_6567,N_6310,N_6380);
nor U6568 (N_6568,N_6322,N_6404);
and U6569 (N_6569,N_6316,N_6367);
and U6570 (N_6570,N_6437,N_6330);
and U6571 (N_6571,N_6395,N_6305);
nor U6572 (N_6572,N_6314,N_6349);
xnor U6573 (N_6573,N_6318,N_6385);
nand U6574 (N_6574,N_6429,N_6407);
or U6575 (N_6575,N_6414,N_6392);
and U6576 (N_6576,N_6349,N_6313);
and U6577 (N_6577,N_6435,N_6366);
nand U6578 (N_6578,N_6350,N_6336);
xnor U6579 (N_6579,N_6402,N_6443);
nor U6580 (N_6580,N_6427,N_6333);
xnor U6581 (N_6581,N_6343,N_6347);
xnor U6582 (N_6582,N_6307,N_6419);
xnor U6583 (N_6583,N_6331,N_6449);
and U6584 (N_6584,N_6420,N_6417);
nor U6585 (N_6585,N_6355,N_6370);
and U6586 (N_6586,N_6383,N_6448);
and U6587 (N_6587,N_6323,N_6369);
and U6588 (N_6588,N_6391,N_6357);
nand U6589 (N_6589,N_6340,N_6335);
xor U6590 (N_6590,N_6352,N_6316);
nor U6591 (N_6591,N_6411,N_6339);
or U6592 (N_6592,N_6318,N_6371);
xnor U6593 (N_6593,N_6306,N_6408);
or U6594 (N_6594,N_6396,N_6407);
or U6595 (N_6595,N_6443,N_6441);
or U6596 (N_6596,N_6431,N_6372);
or U6597 (N_6597,N_6302,N_6384);
xnor U6598 (N_6598,N_6411,N_6367);
and U6599 (N_6599,N_6310,N_6445);
nor U6600 (N_6600,N_6551,N_6550);
nor U6601 (N_6601,N_6546,N_6458);
or U6602 (N_6602,N_6489,N_6598);
or U6603 (N_6603,N_6496,N_6516);
xor U6604 (N_6604,N_6510,N_6528);
and U6605 (N_6605,N_6459,N_6545);
nor U6606 (N_6606,N_6560,N_6532);
nand U6607 (N_6607,N_6566,N_6508);
or U6608 (N_6608,N_6514,N_6487);
nor U6609 (N_6609,N_6500,N_6587);
or U6610 (N_6610,N_6585,N_6472);
or U6611 (N_6611,N_6590,N_6513);
nor U6612 (N_6612,N_6524,N_6460);
xor U6613 (N_6613,N_6572,N_6592);
nand U6614 (N_6614,N_6512,N_6491);
nand U6615 (N_6615,N_6461,N_6543);
nand U6616 (N_6616,N_6466,N_6537);
and U6617 (N_6617,N_6577,N_6594);
nor U6618 (N_6618,N_6511,N_6456);
and U6619 (N_6619,N_6507,N_6561);
xnor U6620 (N_6620,N_6515,N_6565);
nor U6621 (N_6621,N_6475,N_6559);
or U6622 (N_6622,N_6553,N_6596);
and U6623 (N_6623,N_6476,N_6504);
nor U6624 (N_6624,N_6567,N_6536);
xnor U6625 (N_6625,N_6479,N_6563);
nor U6626 (N_6626,N_6588,N_6549);
xor U6627 (N_6627,N_6575,N_6548);
nor U6628 (N_6628,N_6529,N_6505);
nand U6629 (N_6629,N_6518,N_6519);
and U6630 (N_6630,N_6584,N_6499);
xnor U6631 (N_6631,N_6469,N_6474);
or U6632 (N_6632,N_6568,N_6520);
or U6633 (N_6633,N_6582,N_6555);
and U6634 (N_6634,N_6579,N_6576);
nand U6635 (N_6635,N_6451,N_6552);
nand U6636 (N_6636,N_6471,N_6564);
and U6637 (N_6637,N_6502,N_6488);
nor U6638 (N_6638,N_6463,N_6591);
nor U6639 (N_6639,N_6509,N_6583);
or U6640 (N_6640,N_6574,N_6478);
nand U6641 (N_6641,N_6465,N_6538);
xor U6642 (N_6642,N_6503,N_6599);
or U6643 (N_6643,N_6557,N_6486);
nand U6644 (N_6644,N_6464,N_6485);
nand U6645 (N_6645,N_6525,N_6480);
and U6646 (N_6646,N_6527,N_6540);
or U6647 (N_6647,N_6454,N_6521);
xor U6648 (N_6648,N_6494,N_6569);
and U6649 (N_6649,N_6493,N_6506);
and U6650 (N_6650,N_6541,N_6539);
or U6651 (N_6651,N_6450,N_6477);
xnor U6652 (N_6652,N_6533,N_6501);
or U6653 (N_6653,N_6573,N_6457);
nor U6654 (N_6654,N_6586,N_6452);
or U6655 (N_6655,N_6470,N_6473);
xor U6656 (N_6656,N_6482,N_6530);
or U6657 (N_6657,N_6562,N_6593);
nor U6658 (N_6658,N_6558,N_6517);
and U6659 (N_6659,N_6483,N_6570);
and U6660 (N_6660,N_6484,N_6490);
nand U6661 (N_6661,N_6455,N_6492);
and U6662 (N_6662,N_6597,N_6554);
and U6663 (N_6663,N_6595,N_6547);
xor U6664 (N_6664,N_6531,N_6535);
or U6665 (N_6665,N_6571,N_6495);
nor U6666 (N_6666,N_6498,N_6467);
and U6667 (N_6667,N_6581,N_6523);
nor U6668 (N_6668,N_6468,N_6580);
nand U6669 (N_6669,N_6589,N_6522);
and U6670 (N_6670,N_6462,N_6578);
nor U6671 (N_6671,N_6497,N_6556);
and U6672 (N_6672,N_6453,N_6534);
and U6673 (N_6673,N_6481,N_6526);
nor U6674 (N_6674,N_6544,N_6542);
or U6675 (N_6675,N_6508,N_6549);
xor U6676 (N_6676,N_6570,N_6496);
nand U6677 (N_6677,N_6579,N_6535);
nor U6678 (N_6678,N_6487,N_6531);
nand U6679 (N_6679,N_6550,N_6584);
xnor U6680 (N_6680,N_6467,N_6450);
xnor U6681 (N_6681,N_6539,N_6512);
or U6682 (N_6682,N_6564,N_6520);
and U6683 (N_6683,N_6584,N_6477);
xor U6684 (N_6684,N_6561,N_6572);
or U6685 (N_6685,N_6533,N_6541);
nand U6686 (N_6686,N_6473,N_6469);
xnor U6687 (N_6687,N_6485,N_6567);
or U6688 (N_6688,N_6494,N_6558);
xnor U6689 (N_6689,N_6481,N_6486);
and U6690 (N_6690,N_6570,N_6536);
nand U6691 (N_6691,N_6475,N_6463);
nand U6692 (N_6692,N_6560,N_6573);
xnor U6693 (N_6693,N_6556,N_6568);
and U6694 (N_6694,N_6458,N_6561);
nor U6695 (N_6695,N_6574,N_6593);
or U6696 (N_6696,N_6462,N_6464);
nor U6697 (N_6697,N_6588,N_6572);
and U6698 (N_6698,N_6517,N_6467);
nand U6699 (N_6699,N_6583,N_6523);
nor U6700 (N_6700,N_6562,N_6457);
or U6701 (N_6701,N_6487,N_6567);
and U6702 (N_6702,N_6464,N_6565);
and U6703 (N_6703,N_6484,N_6480);
and U6704 (N_6704,N_6539,N_6516);
xnor U6705 (N_6705,N_6531,N_6594);
nand U6706 (N_6706,N_6529,N_6562);
and U6707 (N_6707,N_6524,N_6454);
nand U6708 (N_6708,N_6475,N_6566);
or U6709 (N_6709,N_6474,N_6503);
xnor U6710 (N_6710,N_6525,N_6491);
nor U6711 (N_6711,N_6578,N_6497);
and U6712 (N_6712,N_6483,N_6520);
nand U6713 (N_6713,N_6571,N_6549);
xnor U6714 (N_6714,N_6542,N_6455);
and U6715 (N_6715,N_6563,N_6589);
xor U6716 (N_6716,N_6595,N_6491);
or U6717 (N_6717,N_6526,N_6566);
and U6718 (N_6718,N_6549,N_6535);
nand U6719 (N_6719,N_6451,N_6536);
or U6720 (N_6720,N_6486,N_6508);
or U6721 (N_6721,N_6481,N_6452);
nor U6722 (N_6722,N_6597,N_6450);
or U6723 (N_6723,N_6508,N_6458);
or U6724 (N_6724,N_6456,N_6580);
nand U6725 (N_6725,N_6581,N_6533);
nand U6726 (N_6726,N_6544,N_6598);
nand U6727 (N_6727,N_6566,N_6567);
and U6728 (N_6728,N_6593,N_6501);
nor U6729 (N_6729,N_6488,N_6509);
and U6730 (N_6730,N_6578,N_6575);
nor U6731 (N_6731,N_6476,N_6588);
or U6732 (N_6732,N_6488,N_6589);
xnor U6733 (N_6733,N_6469,N_6513);
nor U6734 (N_6734,N_6479,N_6528);
nand U6735 (N_6735,N_6561,N_6551);
nand U6736 (N_6736,N_6575,N_6460);
nor U6737 (N_6737,N_6540,N_6491);
xor U6738 (N_6738,N_6578,N_6485);
nand U6739 (N_6739,N_6589,N_6559);
xor U6740 (N_6740,N_6568,N_6515);
or U6741 (N_6741,N_6470,N_6531);
nor U6742 (N_6742,N_6450,N_6543);
and U6743 (N_6743,N_6592,N_6450);
nand U6744 (N_6744,N_6573,N_6506);
nand U6745 (N_6745,N_6491,N_6486);
xnor U6746 (N_6746,N_6482,N_6472);
xnor U6747 (N_6747,N_6491,N_6542);
and U6748 (N_6748,N_6568,N_6590);
nor U6749 (N_6749,N_6455,N_6597);
or U6750 (N_6750,N_6623,N_6675);
nand U6751 (N_6751,N_6742,N_6649);
xor U6752 (N_6752,N_6657,N_6695);
and U6753 (N_6753,N_6717,N_6653);
nand U6754 (N_6754,N_6705,N_6724);
nor U6755 (N_6755,N_6665,N_6673);
xnor U6756 (N_6756,N_6604,N_6647);
nor U6757 (N_6757,N_6678,N_6721);
nand U6758 (N_6758,N_6738,N_6739);
nand U6759 (N_6759,N_6715,N_6667);
nand U6760 (N_6760,N_6735,N_6691);
nor U6761 (N_6761,N_6666,N_6684);
nand U6762 (N_6762,N_6732,N_6683);
nor U6763 (N_6763,N_6731,N_6674);
and U6764 (N_6764,N_6687,N_6646);
and U6765 (N_6765,N_6636,N_6628);
and U6766 (N_6766,N_6749,N_6658);
and U6767 (N_6767,N_6697,N_6671);
and U6768 (N_6768,N_6670,N_6626);
nand U6769 (N_6769,N_6660,N_6654);
or U6770 (N_6770,N_6639,N_6614);
nor U6771 (N_6771,N_6696,N_6600);
xor U6772 (N_6772,N_6634,N_6679);
nor U6773 (N_6773,N_6747,N_6743);
nor U6774 (N_6774,N_6744,N_6621);
nor U6775 (N_6775,N_6622,N_6608);
nor U6776 (N_6776,N_6734,N_6659);
xnor U6777 (N_6777,N_6704,N_6736);
nor U6778 (N_6778,N_6677,N_6638);
nor U6779 (N_6779,N_6727,N_6722);
nor U6780 (N_6780,N_6681,N_6617);
or U6781 (N_6781,N_6620,N_6726);
xnor U6782 (N_6782,N_6672,N_6698);
xor U6783 (N_6783,N_6720,N_6656);
nor U6784 (N_6784,N_6689,N_6686);
nor U6785 (N_6785,N_6652,N_6707);
nand U6786 (N_6786,N_6709,N_6613);
or U6787 (N_6787,N_6605,N_6713);
xnor U6788 (N_6788,N_6664,N_6692);
or U6789 (N_6789,N_6625,N_6706);
and U6790 (N_6790,N_6746,N_6663);
or U6791 (N_6791,N_6748,N_6693);
nor U6792 (N_6792,N_6733,N_6711);
or U6793 (N_6793,N_6723,N_6635);
and U6794 (N_6794,N_6716,N_6632);
nor U6795 (N_6795,N_6702,N_6603);
or U6796 (N_6796,N_6615,N_6661);
or U6797 (N_6797,N_6741,N_6690);
nor U6798 (N_6798,N_6616,N_6631);
nor U6799 (N_6799,N_6630,N_6730);
nand U6800 (N_6800,N_6694,N_6607);
nand U6801 (N_6801,N_6640,N_6610);
or U6802 (N_6802,N_6662,N_6719);
or U6803 (N_6803,N_6703,N_6611);
or U6804 (N_6804,N_6601,N_6602);
nand U6805 (N_6805,N_6701,N_6682);
or U6806 (N_6806,N_6710,N_6650);
nor U6807 (N_6807,N_6714,N_6624);
or U6808 (N_6808,N_6629,N_6642);
nor U6809 (N_6809,N_6644,N_6618);
nor U6810 (N_6810,N_6729,N_6619);
xnor U6811 (N_6811,N_6648,N_6685);
or U6812 (N_6812,N_6651,N_6606);
nand U6813 (N_6813,N_6688,N_6633);
nor U6814 (N_6814,N_6645,N_6612);
nand U6815 (N_6815,N_6745,N_6641);
nand U6816 (N_6816,N_6708,N_6655);
or U6817 (N_6817,N_6627,N_6668);
nand U6818 (N_6818,N_6737,N_6643);
and U6819 (N_6819,N_6712,N_6699);
or U6820 (N_6820,N_6637,N_6740);
nand U6821 (N_6821,N_6669,N_6700);
xnor U6822 (N_6822,N_6676,N_6725);
or U6823 (N_6823,N_6680,N_6728);
nand U6824 (N_6824,N_6609,N_6718);
and U6825 (N_6825,N_6733,N_6604);
and U6826 (N_6826,N_6728,N_6733);
or U6827 (N_6827,N_6711,N_6622);
xor U6828 (N_6828,N_6709,N_6629);
xor U6829 (N_6829,N_6656,N_6653);
xnor U6830 (N_6830,N_6622,N_6699);
nand U6831 (N_6831,N_6620,N_6737);
xnor U6832 (N_6832,N_6642,N_6644);
xor U6833 (N_6833,N_6676,N_6618);
nand U6834 (N_6834,N_6713,N_6690);
nand U6835 (N_6835,N_6739,N_6630);
nand U6836 (N_6836,N_6667,N_6721);
nor U6837 (N_6837,N_6742,N_6748);
nand U6838 (N_6838,N_6612,N_6696);
nand U6839 (N_6839,N_6730,N_6695);
nand U6840 (N_6840,N_6626,N_6618);
and U6841 (N_6841,N_6693,N_6606);
nor U6842 (N_6842,N_6668,N_6600);
and U6843 (N_6843,N_6611,N_6684);
nand U6844 (N_6844,N_6702,N_6683);
xnor U6845 (N_6845,N_6717,N_6728);
nor U6846 (N_6846,N_6702,N_6728);
xor U6847 (N_6847,N_6607,N_6612);
or U6848 (N_6848,N_6692,N_6748);
nor U6849 (N_6849,N_6729,N_6614);
nand U6850 (N_6850,N_6707,N_6602);
or U6851 (N_6851,N_6666,N_6693);
xor U6852 (N_6852,N_6631,N_6677);
nor U6853 (N_6853,N_6717,N_6705);
nor U6854 (N_6854,N_6719,N_6735);
xnor U6855 (N_6855,N_6624,N_6676);
nor U6856 (N_6856,N_6660,N_6623);
nand U6857 (N_6857,N_6601,N_6614);
nand U6858 (N_6858,N_6692,N_6729);
or U6859 (N_6859,N_6686,N_6634);
and U6860 (N_6860,N_6719,N_6605);
or U6861 (N_6861,N_6620,N_6643);
xnor U6862 (N_6862,N_6744,N_6645);
nand U6863 (N_6863,N_6691,N_6610);
and U6864 (N_6864,N_6650,N_6640);
or U6865 (N_6865,N_6699,N_6639);
or U6866 (N_6866,N_6684,N_6628);
or U6867 (N_6867,N_6704,N_6680);
and U6868 (N_6868,N_6737,N_6702);
or U6869 (N_6869,N_6703,N_6601);
xor U6870 (N_6870,N_6659,N_6749);
xnor U6871 (N_6871,N_6717,N_6678);
xor U6872 (N_6872,N_6653,N_6642);
nor U6873 (N_6873,N_6627,N_6722);
nand U6874 (N_6874,N_6652,N_6653);
xor U6875 (N_6875,N_6672,N_6690);
nor U6876 (N_6876,N_6607,N_6681);
nand U6877 (N_6877,N_6685,N_6616);
and U6878 (N_6878,N_6725,N_6749);
nor U6879 (N_6879,N_6718,N_6677);
xor U6880 (N_6880,N_6695,N_6680);
and U6881 (N_6881,N_6657,N_6667);
nor U6882 (N_6882,N_6684,N_6702);
nand U6883 (N_6883,N_6614,N_6681);
nand U6884 (N_6884,N_6718,N_6678);
or U6885 (N_6885,N_6740,N_6722);
nor U6886 (N_6886,N_6646,N_6745);
xnor U6887 (N_6887,N_6655,N_6693);
nand U6888 (N_6888,N_6674,N_6676);
or U6889 (N_6889,N_6691,N_6686);
or U6890 (N_6890,N_6668,N_6672);
nor U6891 (N_6891,N_6646,N_6707);
xor U6892 (N_6892,N_6749,N_6671);
nand U6893 (N_6893,N_6706,N_6677);
nand U6894 (N_6894,N_6600,N_6717);
xor U6895 (N_6895,N_6693,N_6627);
nor U6896 (N_6896,N_6748,N_6635);
nor U6897 (N_6897,N_6727,N_6677);
nand U6898 (N_6898,N_6605,N_6675);
xnor U6899 (N_6899,N_6669,N_6604);
nor U6900 (N_6900,N_6854,N_6771);
nand U6901 (N_6901,N_6801,N_6850);
and U6902 (N_6902,N_6772,N_6835);
nand U6903 (N_6903,N_6816,N_6840);
nand U6904 (N_6904,N_6799,N_6764);
nor U6905 (N_6905,N_6853,N_6807);
xor U6906 (N_6906,N_6893,N_6873);
xnor U6907 (N_6907,N_6871,N_6811);
or U6908 (N_6908,N_6759,N_6755);
nand U6909 (N_6909,N_6774,N_6776);
nor U6910 (N_6910,N_6808,N_6882);
and U6911 (N_6911,N_6890,N_6821);
and U6912 (N_6912,N_6852,N_6806);
nor U6913 (N_6913,N_6760,N_6812);
nor U6914 (N_6914,N_6851,N_6753);
or U6915 (N_6915,N_6881,N_6877);
and U6916 (N_6916,N_6857,N_6839);
xnor U6917 (N_6917,N_6785,N_6844);
or U6918 (N_6918,N_6797,N_6884);
and U6919 (N_6919,N_6758,N_6896);
xor U6920 (N_6920,N_6793,N_6766);
nand U6921 (N_6921,N_6894,N_6865);
or U6922 (N_6922,N_6826,N_6860);
nor U6923 (N_6923,N_6856,N_6830);
nand U6924 (N_6924,N_6784,N_6790);
xor U6925 (N_6925,N_6792,N_6800);
and U6926 (N_6926,N_6803,N_6846);
xnor U6927 (N_6927,N_6825,N_6804);
nand U6928 (N_6928,N_6858,N_6750);
and U6929 (N_6929,N_6814,N_6891);
nor U6930 (N_6930,N_6775,N_6849);
or U6931 (N_6931,N_6880,N_6751);
nor U6932 (N_6932,N_6878,N_6779);
nand U6933 (N_6933,N_6829,N_6781);
nand U6934 (N_6934,N_6789,N_6824);
and U6935 (N_6935,N_6864,N_6817);
xnor U6936 (N_6936,N_6885,N_6823);
nand U6937 (N_6937,N_6897,N_6791);
nor U6938 (N_6938,N_6859,N_6842);
and U6939 (N_6939,N_6867,N_6813);
and U6940 (N_6940,N_6822,N_6819);
nand U6941 (N_6941,N_6834,N_6795);
and U6942 (N_6942,N_6870,N_6815);
and U6943 (N_6943,N_6761,N_6802);
nor U6944 (N_6944,N_6888,N_6757);
and U6945 (N_6945,N_6843,N_6756);
and U6946 (N_6946,N_6752,N_6892);
xor U6947 (N_6947,N_6848,N_6818);
and U6948 (N_6948,N_6780,N_6838);
nand U6949 (N_6949,N_6866,N_6855);
nor U6950 (N_6950,N_6769,N_6899);
or U6951 (N_6951,N_6845,N_6832);
nor U6952 (N_6952,N_6794,N_6833);
nand U6953 (N_6953,N_6886,N_6898);
nand U6954 (N_6954,N_6768,N_6786);
or U6955 (N_6955,N_6767,N_6754);
nor U6956 (N_6956,N_6810,N_6778);
nand U6957 (N_6957,N_6782,N_6796);
and U6958 (N_6958,N_6798,N_6763);
and U6959 (N_6959,N_6836,N_6895);
and U6960 (N_6960,N_6883,N_6862);
or U6961 (N_6961,N_6805,N_6762);
xnor U6962 (N_6962,N_6809,N_6889);
nor U6963 (N_6963,N_6872,N_6783);
xnor U6964 (N_6964,N_6770,N_6831);
nor U6965 (N_6965,N_6788,N_6841);
nor U6966 (N_6966,N_6787,N_6765);
or U6967 (N_6967,N_6820,N_6887);
or U6968 (N_6968,N_6863,N_6773);
nor U6969 (N_6969,N_6777,N_6847);
and U6970 (N_6970,N_6828,N_6827);
nand U6971 (N_6971,N_6879,N_6861);
nand U6972 (N_6972,N_6876,N_6875);
xor U6973 (N_6973,N_6837,N_6869);
or U6974 (N_6974,N_6874,N_6868);
nand U6975 (N_6975,N_6786,N_6829);
xnor U6976 (N_6976,N_6855,N_6814);
nor U6977 (N_6977,N_6801,N_6887);
nor U6978 (N_6978,N_6766,N_6873);
nand U6979 (N_6979,N_6796,N_6823);
xnor U6980 (N_6980,N_6846,N_6806);
or U6981 (N_6981,N_6846,N_6762);
nand U6982 (N_6982,N_6883,N_6857);
or U6983 (N_6983,N_6785,N_6816);
or U6984 (N_6984,N_6849,N_6774);
nand U6985 (N_6985,N_6814,N_6884);
xnor U6986 (N_6986,N_6831,N_6757);
and U6987 (N_6987,N_6829,N_6831);
nor U6988 (N_6988,N_6752,N_6774);
nor U6989 (N_6989,N_6816,N_6825);
nor U6990 (N_6990,N_6899,N_6876);
xnor U6991 (N_6991,N_6845,N_6815);
and U6992 (N_6992,N_6844,N_6881);
xor U6993 (N_6993,N_6810,N_6771);
xnor U6994 (N_6994,N_6859,N_6788);
and U6995 (N_6995,N_6761,N_6874);
and U6996 (N_6996,N_6765,N_6811);
xnor U6997 (N_6997,N_6881,N_6774);
nor U6998 (N_6998,N_6863,N_6806);
xnor U6999 (N_6999,N_6854,N_6768);
nand U7000 (N_7000,N_6875,N_6848);
and U7001 (N_7001,N_6777,N_6781);
and U7002 (N_7002,N_6786,N_6862);
and U7003 (N_7003,N_6752,N_6882);
and U7004 (N_7004,N_6769,N_6837);
nand U7005 (N_7005,N_6867,N_6860);
nand U7006 (N_7006,N_6842,N_6834);
and U7007 (N_7007,N_6865,N_6771);
or U7008 (N_7008,N_6776,N_6861);
xor U7009 (N_7009,N_6899,N_6800);
and U7010 (N_7010,N_6811,N_6768);
xnor U7011 (N_7011,N_6770,N_6821);
xor U7012 (N_7012,N_6872,N_6823);
nand U7013 (N_7013,N_6806,N_6802);
nand U7014 (N_7014,N_6751,N_6762);
nand U7015 (N_7015,N_6817,N_6769);
or U7016 (N_7016,N_6804,N_6818);
or U7017 (N_7017,N_6809,N_6858);
nand U7018 (N_7018,N_6767,N_6880);
nor U7019 (N_7019,N_6807,N_6774);
nand U7020 (N_7020,N_6792,N_6825);
and U7021 (N_7021,N_6803,N_6812);
and U7022 (N_7022,N_6815,N_6869);
nand U7023 (N_7023,N_6819,N_6778);
nand U7024 (N_7024,N_6886,N_6771);
nand U7025 (N_7025,N_6794,N_6780);
or U7026 (N_7026,N_6773,N_6843);
nor U7027 (N_7027,N_6870,N_6868);
or U7028 (N_7028,N_6834,N_6794);
xor U7029 (N_7029,N_6771,N_6871);
or U7030 (N_7030,N_6838,N_6817);
nand U7031 (N_7031,N_6803,N_6867);
or U7032 (N_7032,N_6875,N_6803);
or U7033 (N_7033,N_6788,N_6814);
nor U7034 (N_7034,N_6763,N_6886);
nor U7035 (N_7035,N_6898,N_6839);
or U7036 (N_7036,N_6847,N_6897);
and U7037 (N_7037,N_6765,N_6815);
or U7038 (N_7038,N_6750,N_6794);
or U7039 (N_7039,N_6751,N_6823);
nor U7040 (N_7040,N_6771,N_6877);
and U7041 (N_7041,N_6842,N_6878);
and U7042 (N_7042,N_6830,N_6785);
xor U7043 (N_7043,N_6804,N_6843);
nand U7044 (N_7044,N_6864,N_6821);
nor U7045 (N_7045,N_6839,N_6888);
nor U7046 (N_7046,N_6852,N_6825);
nand U7047 (N_7047,N_6894,N_6767);
xnor U7048 (N_7048,N_6758,N_6776);
nand U7049 (N_7049,N_6871,N_6821);
or U7050 (N_7050,N_7005,N_7006);
nor U7051 (N_7051,N_6964,N_6967);
nor U7052 (N_7052,N_7028,N_7021);
or U7053 (N_7053,N_6933,N_7040);
or U7054 (N_7054,N_6900,N_6962);
nand U7055 (N_7055,N_7032,N_6941);
nand U7056 (N_7056,N_6990,N_6965);
nor U7057 (N_7057,N_7010,N_7041);
nor U7058 (N_7058,N_6949,N_7030);
xor U7059 (N_7059,N_6945,N_7036);
nor U7060 (N_7060,N_6903,N_7014);
xor U7061 (N_7061,N_6985,N_6926);
and U7062 (N_7062,N_7012,N_6922);
and U7063 (N_7063,N_6935,N_6953);
and U7064 (N_7064,N_6928,N_6942);
nor U7065 (N_7065,N_6947,N_6995);
or U7066 (N_7066,N_6997,N_6939);
and U7067 (N_7067,N_7049,N_6924);
and U7068 (N_7068,N_6996,N_6932);
and U7069 (N_7069,N_6963,N_6981);
and U7070 (N_7070,N_6927,N_6991);
and U7071 (N_7071,N_7027,N_7043);
or U7072 (N_7072,N_6930,N_7039);
and U7073 (N_7073,N_6999,N_6968);
nor U7074 (N_7074,N_7002,N_6977);
or U7075 (N_7075,N_6934,N_7048);
or U7076 (N_7076,N_7047,N_7044);
xnor U7077 (N_7077,N_6960,N_7037);
nand U7078 (N_7078,N_6908,N_7038);
xor U7079 (N_7079,N_7018,N_6975);
nor U7080 (N_7080,N_6971,N_6943);
and U7081 (N_7081,N_7026,N_6936);
or U7082 (N_7082,N_6958,N_7031);
and U7083 (N_7083,N_7009,N_7011);
xnor U7084 (N_7084,N_6987,N_6919);
xor U7085 (N_7085,N_6920,N_6982);
or U7086 (N_7086,N_6961,N_6915);
nor U7087 (N_7087,N_6992,N_7022);
nand U7088 (N_7088,N_7034,N_6929);
and U7089 (N_7089,N_6911,N_7029);
nor U7090 (N_7090,N_6957,N_7016);
and U7091 (N_7091,N_7000,N_6914);
or U7092 (N_7092,N_6970,N_6909);
nand U7093 (N_7093,N_7024,N_7023);
or U7094 (N_7094,N_6921,N_7020);
nor U7095 (N_7095,N_7046,N_6974);
or U7096 (N_7096,N_6986,N_6940);
nor U7097 (N_7097,N_6998,N_7013);
or U7098 (N_7098,N_6980,N_7035);
and U7099 (N_7099,N_6913,N_6969);
xor U7100 (N_7100,N_7017,N_6994);
nand U7101 (N_7101,N_6902,N_6938);
xor U7102 (N_7102,N_6910,N_6955);
xor U7103 (N_7103,N_6976,N_6959);
and U7104 (N_7104,N_6944,N_6950);
nand U7105 (N_7105,N_6972,N_7019);
xor U7106 (N_7106,N_6979,N_6917);
nor U7107 (N_7107,N_6906,N_6983);
or U7108 (N_7108,N_6916,N_6984);
and U7109 (N_7109,N_7042,N_7003);
nor U7110 (N_7110,N_6988,N_6907);
and U7111 (N_7111,N_6954,N_6912);
or U7112 (N_7112,N_6925,N_6923);
or U7113 (N_7113,N_6973,N_7033);
and U7114 (N_7114,N_6989,N_6918);
and U7115 (N_7115,N_6951,N_6966);
and U7116 (N_7116,N_6905,N_6952);
nand U7117 (N_7117,N_7004,N_7045);
xnor U7118 (N_7118,N_7007,N_6937);
or U7119 (N_7119,N_6948,N_6904);
xnor U7120 (N_7120,N_6993,N_7008);
or U7121 (N_7121,N_7015,N_6946);
nand U7122 (N_7122,N_7001,N_7025);
or U7123 (N_7123,N_6978,N_6956);
or U7124 (N_7124,N_6901,N_6931);
nand U7125 (N_7125,N_7034,N_7011);
nand U7126 (N_7126,N_6918,N_6950);
or U7127 (N_7127,N_6970,N_6992);
or U7128 (N_7128,N_6939,N_6921);
xor U7129 (N_7129,N_6942,N_6932);
xor U7130 (N_7130,N_7018,N_6944);
and U7131 (N_7131,N_6983,N_6930);
nor U7132 (N_7132,N_7001,N_7016);
nor U7133 (N_7133,N_7029,N_6948);
or U7134 (N_7134,N_6961,N_6990);
nor U7135 (N_7135,N_7032,N_6947);
nor U7136 (N_7136,N_6966,N_6928);
and U7137 (N_7137,N_6990,N_6944);
and U7138 (N_7138,N_6972,N_6954);
xor U7139 (N_7139,N_7028,N_7007);
or U7140 (N_7140,N_7001,N_6941);
xor U7141 (N_7141,N_6986,N_7034);
or U7142 (N_7142,N_6915,N_6912);
nor U7143 (N_7143,N_7044,N_7048);
or U7144 (N_7144,N_6911,N_7034);
nand U7145 (N_7145,N_6971,N_6960);
nor U7146 (N_7146,N_6972,N_6922);
nor U7147 (N_7147,N_6926,N_7032);
nor U7148 (N_7148,N_6944,N_7003);
nor U7149 (N_7149,N_6976,N_6987);
xnor U7150 (N_7150,N_7002,N_7010);
xnor U7151 (N_7151,N_6935,N_6984);
nand U7152 (N_7152,N_6926,N_7025);
and U7153 (N_7153,N_7013,N_7033);
xor U7154 (N_7154,N_7011,N_6982);
and U7155 (N_7155,N_7008,N_6992);
xor U7156 (N_7156,N_6923,N_6916);
xor U7157 (N_7157,N_7032,N_6919);
xnor U7158 (N_7158,N_6991,N_7000);
and U7159 (N_7159,N_6988,N_6912);
and U7160 (N_7160,N_6998,N_6978);
nand U7161 (N_7161,N_7032,N_6951);
nor U7162 (N_7162,N_7047,N_6996);
or U7163 (N_7163,N_6957,N_7013);
xor U7164 (N_7164,N_6991,N_6978);
and U7165 (N_7165,N_6918,N_7003);
or U7166 (N_7166,N_6937,N_7037);
xnor U7167 (N_7167,N_6992,N_6999);
or U7168 (N_7168,N_6996,N_7013);
and U7169 (N_7169,N_7003,N_7021);
and U7170 (N_7170,N_6925,N_7008);
nor U7171 (N_7171,N_7001,N_7042);
or U7172 (N_7172,N_7035,N_7043);
and U7173 (N_7173,N_7010,N_7005);
nor U7174 (N_7174,N_6959,N_6902);
nor U7175 (N_7175,N_7004,N_7027);
and U7176 (N_7176,N_7019,N_6960);
xnor U7177 (N_7177,N_7020,N_6940);
nor U7178 (N_7178,N_6940,N_6987);
xor U7179 (N_7179,N_6983,N_7003);
or U7180 (N_7180,N_6988,N_6977);
xnor U7181 (N_7181,N_7031,N_7015);
xnor U7182 (N_7182,N_6937,N_6906);
and U7183 (N_7183,N_6936,N_6989);
nand U7184 (N_7184,N_6956,N_7049);
or U7185 (N_7185,N_6902,N_6977);
nand U7186 (N_7186,N_6921,N_6955);
and U7187 (N_7187,N_6905,N_6970);
nand U7188 (N_7188,N_6979,N_7047);
or U7189 (N_7189,N_6940,N_6968);
nor U7190 (N_7190,N_6961,N_6908);
nor U7191 (N_7191,N_6918,N_6969);
xor U7192 (N_7192,N_7038,N_7002);
and U7193 (N_7193,N_6926,N_6979);
nor U7194 (N_7194,N_6964,N_6984);
and U7195 (N_7195,N_6956,N_7010);
nor U7196 (N_7196,N_7008,N_6976);
xnor U7197 (N_7197,N_6964,N_6959);
nand U7198 (N_7198,N_6908,N_6987);
nand U7199 (N_7199,N_6996,N_6995);
nand U7200 (N_7200,N_7129,N_7058);
nor U7201 (N_7201,N_7186,N_7081);
nand U7202 (N_7202,N_7092,N_7175);
nor U7203 (N_7203,N_7144,N_7184);
nand U7204 (N_7204,N_7090,N_7194);
nor U7205 (N_7205,N_7191,N_7059);
or U7206 (N_7206,N_7082,N_7098);
or U7207 (N_7207,N_7104,N_7190);
nor U7208 (N_7208,N_7132,N_7050);
xor U7209 (N_7209,N_7091,N_7139);
nand U7210 (N_7210,N_7130,N_7170);
nor U7211 (N_7211,N_7061,N_7117);
nand U7212 (N_7212,N_7056,N_7096);
nor U7213 (N_7213,N_7079,N_7133);
nand U7214 (N_7214,N_7118,N_7148);
nand U7215 (N_7215,N_7161,N_7097);
nor U7216 (N_7216,N_7125,N_7093);
nand U7217 (N_7217,N_7145,N_7149);
or U7218 (N_7218,N_7135,N_7116);
or U7219 (N_7219,N_7089,N_7155);
nor U7220 (N_7220,N_7126,N_7078);
and U7221 (N_7221,N_7143,N_7177);
xnor U7222 (N_7222,N_7053,N_7094);
xor U7223 (N_7223,N_7159,N_7165);
and U7224 (N_7224,N_7127,N_7121);
nand U7225 (N_7225,N_7084,N_7150);
and U7226 (N_7226,N_7198,N_7110);
and U7227 (N_7227,N_7069,N_7152);
nor U7228 (N_7228,N_7070,N_7123);
and U7229 (N_7229,N_7119,N_7085);
xnor U7230 (N_7230,N_7166,N_7095);
and U7231 (N_7231,N_7106,N_7105);
or U7232 (N_7232,N_7064,N_7108);
nand U7233 (N_7233,N_7124,N_7109);
nor U7234 (N_7234,N_7052,N_7101);
xnor U7235 (N_7235,N_7160,N_7142);
nor U7236 (N_7236,N_7100,N_7107);
nand U7237 (N_7237,N_7122,N_7173);
nor U7238 (N_7238,N_7134,N_7072);
nand U7239 (N_7239,N_7141,N_7163);
or U7240 (N_7240,N_7088,N_7114);
and U7241 (N_7241,N_7181,N_7137);
nor U7242 (N_7242,N_7128,N_7131);
or U7243 (N_7243,N_7169,N_7168);
nand U7244 (N_7244,N_7111,N_7077);
xor U7245 (N_7245,N_7051,N_7156);
and U7246 (N_7246,N_7103,N_7180);
nand U7247 (N_7247,N_7138,N_7120);
or U7248 (N_7248,N_7179,N_7172);
nor U7249 (N_7249,N_7099,N_7063);
nor U7250 (N_7250,N_7071,N_7136);
xnor U7251 (N_7251,N_7167,N_7086);
nor U7252 (N_7252,N_7187,N_7157);
xnor U7253 (N_7253,N_7164,N_7074);
and U7254 (N_7254,N_7151,N_7076);
nor U7255 (N_7255,N_7112,N_7196);
and U7256 (N_7256,N_7113,N_7057);
nand U7257 (N_7257,N_7067,N_7158);
nand U7258 (N_7258,N_7065,N_7062);
and U7259 (N_7259,N_7087,N_7195);
and U7260 (N_7260,N_7176,N_7075);
nor U7261 (N_7261,N_7182,N_7183);
nand U7262 (N_7262,N_7189,N_7055);
or U7263 (N_7263,N_7185,N_7188);
nand U7264 (N_7264,N_7083,N_7193);
and U7265 (N_7265,N_7162,N_7174);
xnor U7266 (N_7266,N_7147,N_7054);
and U7267 (N_7267,N_7192,N_7068);
xnor U7268 (N_7268,N_7178,N_7115);
and U7269 (N_7269,N_7060,N_7146);
nand U7270 (N_7270,N_7102,N_7154);
nor U7271 (N_7271,N_7066,N_7140);
xnor U7272 (N_7272,N_7080,N_7153);
nand U7273 (N_7273,N_7199,N_7197);
xor U7274 (N_7274,N_7073,N_7171);
nor U7275 (N_7275,N_7198,N_7149);
and U7276 (N_7276,N_7138,N_7081);
and U7277 (N_7277,N_7159,N_7172);
or U7278 (N_7278,N_7069,N_7142);
or U7279 (N_7279,N_7142,N_7162);
nor U7280 (N_7280,N_7072,N_7132);
nor U7281 (N_7281,N_7058,N_7104);
and U7282 (N_7282,N_7162,N_7061);
and U7283 (N_7283,N_7107,N_7185);
nand U7284 (N_7284,N_7127,N_7183);
xor U7285 (N_7285,N_7098,N_7114);
nor U7286 (N_7286,N_7176,N_7106);
nor U7287 (N_7287,N_7171,N_7097);
or U7288 (N_7288,N_7126,N_7095);
xor U7289 (N_7289,N_7064,N_7171);
and U7290 (N_7290,N_7070,N_7054);
nor U7291 (N_7291,N_7079,N_7157);
nor U7292 (N_7292,N_7141,N_7110);
and U7293 (N_7293,N_7123,N_7126);
nor U7294 (N_7294,N_7053,N_7170);
nand U7295 (N_7295,N_7075,N_7174);
nand U7296 (N_7296,N_7181,N_7117);
and U7297 (N_7297,N_7123,N_7191);
or U7298 (N_7298,N_7195,N_7110);
nor U7299 (N_7299,N_7124,N_7194);
or U7300 (N_7300,N_7090,N_7073);
and U7301 (N_7301,N_7154,N_7114);
nand U7302 (N_7302,N_7165,N_7130);
or U7303 (N_7303,N_7132,N_7157);
nor U7304 (N_7304,N_7154,N_7095);
nor U7305 (N_7305,N_7074,N_7096);
or U7306 (N_7306,N_7190,N_7154);
nand U7307 (N_7307,N_7061,N_7075);
nand U7308 (N_7308,N_7164,N_7096);
or U7309 (N_7309,N_7186,N_7151);
and U7310 (N_7310,N_7175,N_7166);
nand U7311 (N_7311,N_7184,N_7052);
or U7312 (N_7312,N_7095,N_7122);
nand U7313 (N_7313,N_7153,N_7173);
or U7314 (N_7314,N_7080,N_7096);
nor U7315 (N_7315,N_7138,N_7198);
or U7316 (N_7316,N_7069,N_7138);
xor U7317 (N_7317,N_7094,N_7171);
nor U7318 (N_7318,N_7059,N_7139);
nand U7319 (N_7319,N_7157,N_7156);
xnor U7320 (N_7320,N_7178,N_7159);
and U7321 (N_7321,N_7058,N_7083);
xnor U7322 (N_7322,N_7156,N_7093);
nand U7323 (N_7323,N_7159,N_7120);
nand U7324 (N_7324,N_7172,N_7062);
nand U7325 (N_7325,N_7109,N_7193);
nor U7326 (N_7326,N_7169,N_7160);
or U7327 (N_7327,N_7177,N_7157);
nor U7328 (N_7328,N_7144,N_7123);
and U7329 (N_7329,N_7175,N_7112);
xnor U7330 (N_7330,N_7134,N_7124);
and U7331 (N_7331,N_7150,N_7088);
nand U7332 (N_7332,N_7168,N_7134);
nand U7333 (N_7333,N_7055,N_7185);
and U7334 (N_7334,N_7078,N_7051);
and U7335 (N_7335,N_7101,N_7195);
and U7336 (N_7336,N_7055,N_7079);
or U7337 (N_7337,N_7185,N_7097);
nor U7338 (N_7338,N_7162,N_7066);
or U7339 (N_7339,N_7104,N_7094);
and U7340 (N_7340,N_7131,N_7185);
and U7341 (N_7341,N_7143,N_7160);
xnor U7342 (N_7342,N_7060,N_7176);
and U7343 (N_7343,N_7149,N_7144);
or U7344 (N_7344,N_7175,N_7148);
nor U7345 (N_7345,N_7094,N_7082);
or U7346 (N_7346,N_7197,N_7101);
and U7347 (N_7347,N_7145,N_7185);
xnor U7348 (N_7348,N_7058,N_7146);
nor U7349 (N_7349,N_7151,N_7068);
nor U7350 (N_7350,N_7338,N_7214);
nand U7351 (N_7351,N_7331,N_7291);
xor U7352 (N_7352,N_7298,N_7303);
and U7353 (N_7353,N_7232,N_7229);
and U7354 (N_7354,N_7330,N_7202);
and U7355 (N_7355,N_7341,N_7222);
or U7356 (N_7356,N_7277,N_7239);
or U7357 (N_7357,N_7246,N_7211);
nor U7358 (N_7358,N_7310,N_7299);
nand U7359 (N_7359,N_7294,N_7334);
nand U7360 (N_7360,N_7333,N_7329);
nand U7361 (N_7361,N_7312,N_7348);
nand U7362 (N_7362,N_7268,N_7241);
or U7363 (N_7363,N_7243,N_7321);
and U7364 (N_7364,N_7319,N_7208);
xnor U7365 (N_7365,N_7322,N_7271);
nand U7366 (N_7366,N_7281,N_7335);
and U7367 (N_7367,N_7342,N_7215);
and U7368 (N_7368,N_7219,N_7315);
nand U7369 (N_7369,N_7217,N_7212);
nor U7370 (N_7370,N_7260,N_7289);
xnor U7371 (N_7371,N_7336,N_7225);
or U7372 (N_7372,N_7228,N_7261);
and U7373 (N_7373,N_7248,N_7288);
nor U7374 (N_7374,N_7286,N_7201);
nand U7375 (N_7375,N_7234,N_7269);
and U7376 (N_7376,N_7205,N_7206);
xor U7377 (N_7377,N_7275,N_7272);
and U7378 (N_7378,N_7302,N_7287);
and U7379 (N_7379,N_7324,N_7344);
and U7380 (N_7380,N_7257,N_7307);
nor U7381 (N_7381,N_7332,N_7210);
nand U7382 (N_7382,N_7317,N_7327);
xnor U7383 (N_7383,N_7323,N_7259);
xnor U7384 (N_7384,N_7345,N_7237);
xnor U7385 (N_7385,N_7326,N_7244);
xor U7386 (N_7386,N_7203,N_7224);
or U7387 (N_7387,N_7296,N_7213);
or U7388 (N_7388,N_7264,N_7340);
nand U7389 (N_7389,N_7316,N_7306);
nor U7390 (N_7390,N_7305,N_7295);
nand U7391 (N_7391,N_7270,N_7284);
and U7392 (N_7392,N_7311,N_7318);
and U7393 (N_7393,N_7308,N_7216);
nor U7394 (N_7394,N_7255,N_7245);
nand U7395 (N_7395,N_7263,N_7226);
nand U7396 (N_7396,N_7218,N_7256);
and U7397 (N_7397,N_7320,N_7313);
nor U7398 (N_7398,N_7300,N_7347);
nand U7399 (N_7399,N_7240,N_7273);
and U7400 (N_7400,N_7349,N_7266);
and U7401 (N_7401,N_7301,N_7267);
xor U7402 (N_7402,N_7339,N_7221);
nor U7403 (N_7403,N_7279,N_7247);
xor U7404 (N_7404,N_7290,N_7283);
or U7405 (N_7405,N_7253,N_7265);
and U7406 (N_7406,N_7282,N_7346);
or U7407 (N_7407,N_7278,N_7227);
and U7408 (N_7408,N_7250,N_7235);
xor U7409 (N_7409,N_7200,N_7249);
nor U7410 (N_7410,N_7297,N_7204);
nand U7411 (N_7411,N_7233,N_7285);
nor U7412 (N_7412,N_7337,N_7252);
and U7413 (N_7413,N_7231,N_7343);
nor U7414 (N_7414,N_7238,N_7230);
or U7415 (N_7415,N_7309,N_7242);
or U7416 (N_7416,N_7325,N_7223);
nor U7417 (N_7417,N_7254,N_7262);
nor U7418 (N_7418,N_7251,N_7276);
nor U7419 (N_7419,N_7274,N_7258);
nand U7420 (N_7420,N_7236,N_7207);
nand U7421 (N_7421,N_7293,N_7314);
or U7422 (N_7422,N_7328,N_7209);
nand U7423 (N_7423,N_7280,N_7304);
and U7424 (N_7424,N_7220,N_7292);
xnor U7425 (N_7425,N_7227,N_7333);
nand U7426 (N_7426,N_7214,N_7324);
or U7427 (N_7427,N_7284,N_7336);
nand U7428 (N_7428,N_7261,N_7295);
or U7429 (N_7429,N_7336,N_7218);
nand U7430 (N_7430,N_7225,N_7303);
and U7431 (N_7431,N_7279,N_7313);
or U7432 (N_7432,N_7209,N_7238);
xor U7433 (N_7433,N_7268,N_7237);
xnor U7434 (N_7434,N_7299,N_7220);
xor U7435 (N_7435,N_7235,N_7283);
and U7436 (N_7436,N_7247,N_7246);
xnor U7437 (N_7437,N_7347,N_7330);
nand U7438 (N_7438,N_7336,N_7281);
nor U7439 (N_7439,N_7284,N_7259);
nor U7440 (N_7440,N_7293,N_7321);
nor U7441 (N_7441,N_7284,N_7214);
nor U7442 (N_7442,N_7280,N_7261);
and U7443 (N_7443,N_7294,N_7291);
xnor U7444 (N_7444,N_7311,N_7292);
or U7445 (N_7445,N_7339,N_7313);
and U7446 (N_7446,N_7286,N_7257);
and U7447 (N_7447,N_7282,N_7301);
xnor U7448 (N_7448,N_7217,N_7338);
nand U7449 (N_7449,N_7230,N_7252);
and U7450 (N_7450,N_7347,N_7235);
nand U7451 (N_7451,N_7339,N_7273);
and U7452 (N_7452,N_7293,N_7290);
nor U7453 (N_7453,N_7257,N_7311);
or U7454 (N_7454,N_7344,N_7348);
xor U7455 (N_7455,N_7345,N_7319);
xor U7456 (N_7456,N_7297,N_7216);
nor U7457 (N_7457,N_7278,N_7202);
or U7458 (N_7458,N_7346,N_7223);
or U7459 (N_7459,N_7203,N_7264);
xnor U7460 (N_7460,N_7275,N_7346);
nand U7461 (N_7461,N_7238,N_7285);
or U7462 (N_7462,N_7306,N_7332);
xor U7463 (N_7463,N_7289,N_7330);
and U7464 (N_7464,N_7254,N_7207);
xnor U7465 (N_7465,N_7293,N_7215);
or U7466 (N_7466,N_7299,N_7345);
or U7467 (N_7467,N_7346,N_7233);
and U7468 (N_7468,N_7289,N_7282);
and U7469 (N_7469,N_7292,N_7285);
nand U7470 (N_7470,N_7251,N_7223);
xnor U7471 (N_7471,N_7271,N_7316);
nor U7472 (N_7472,N_7330,N_7291);
or U7473 (N_7473,N_7208,N_7229);
or U7474 (N_7474,N_7258,N_7273);
or U7475 (N_7475,N_7326,N_7223);
nand U7476 (N_7476,N_7283,N_7254);
xnor U7477 (N_7477,N_7279,N_7312);
nand U7478 (N_7478,N_7228,N_7284);
nand U7479 (N_7479,N_7269,N_7248);
nand U7480 (N_7480,N_7341,N_7304);
or U7481 (N_7481,N_7295,N_7328);
or U7482 (N_7482,N_7288,N_7330);
and U7483 (N_7483,N_7221,N_7225);
nor U7484 (N_7484,N_7266,N_7239);
nor U7485 (N_7485,N_7236,N_7315);
xnor U7486 (N_7486,N_7330,N_7205);
xnor U7487 (N_7487,N_7215,N_7345);
xnor U7488 (N_7488,N_7328,N_7348);
or U7489 (N_7489,N_7223,N_7252);
and U7490 (N_7490,N_7285,N_7284);
nand U7491 (N_7491,N_7227,N_7326);
and U7492 (N_7492,N_7207,N_7214);
xor U7493 (N_7493,N_7277,N_7340);
or U7494 (N_7494,N_7241,N_7345);
nand U7495 (N_7495,N_7267,N_7305);
nor U7496 (N_7496,N_7287,N_7339);
xor U7497 (N_7497,N_7267,N_7337);
or U7498 (N_7498,N_7203,N_7291);
and U7499 (N_7499,N_7312,N_7346);
nor U7500 (N_7500,N_7357,N_7453);
or U7501 (N_7501,N_7471,N_7465);
nor U7502 (N_7502,N_7435,N_7414);
and U7503 (N_7503,N_7474,N_7375);
nor U7504 (N_7504,N_7391,N_7410);
and U7505 (N_7505,N_7356,N_7472);
nand U7506 (N_7506,N_7390,N_7402);
xor U7507 (N_7507,N_7439,N_7499);
nor U7508 (N_7508,N_7361,N_7434);
nor U7509 (N_7509,N_7398,N_7416);
nor U7510 (N_7510,N_7492,N_7422);
nand U7511 (N_7511,N_7359,N_7485);
xor U7512 (N_7512,N_7403,N_7476);
nand U7513 (N_7513,N_7473,N_7493);
nor U7514 (N_7514,N_7436,N_7432);
nand U7515 (N_7515,N_7451,N_7480);
xor U7516 (N_7516,N_7353,N_7389);
nor U7517 (N_7517,N_7482,N_7364);
nand U7518 (N_7518,N_7487,N_7415);
nor U7519 (N_7519,N_7406,N_7495);
nand U7520 (N_7520,N_7475,N_7385);
nand U7521 (N_7521,N_7399,N_7396);
nand U7522 (N_7522,N_7351,N_7460);
nor U7523 (N_7523,N_7387,N_7409);
nand U7524 (N_7524,N_7386,N_7426);
xnor U7525 (N_7525,N_7367,N_7405);
and U7526 (N_7526,N_7404,N_7427);
or U7527 (N_7527,N_7382,N_7445);
xor U7528 (N_7528,N_7454,N_7452);
and U7529 (N_7529,N_7464,N_7498);
nor U7530 (N_7530,N_7468,N_7419);
xor U7531 (N_7531,N_7413,N_7370);
nand U7532 (N_7532,N_7490,N_7449);
nor U7533 (N_7533,N_7378,N_7352);
xnor U7534 (N_7534,N_7350,N_7381);
nand U7535 (N_7535,N_7496,N_7440);
or U7536 (N_7536,N_7428,N_7423);
xnor U7537 (N_7537,N_7438,N_7394);
nand U7538 (N_7538,N_7444,N_7355);
and U7539 (N_7539,N_7380,N_7469);
nor U7540 (N_7540,N_7483,N_7358);
or U7541 (N_7541,N_7383,N_7491);
or U7542 (N_7542,N_7411,N_7459);
or U7543 (N_7543,N_7489,N_7488);
xor U7544 (N_7544,N_7368,N_7354);
nor U7545 (N_7545,N_7360,N_7412);
xnor U7546 (N_7546,N_7366,N_7384);
or U7547 (N_7547,N_7446,N_7379);
and U7548 (N_7548,N_7363,N_7433);
or U7549 (N_7549,N_7420,N_7497);
xor U7550 (N_7550,N_7462,N_7429);
xnor U7551 (N_7551,N_7397,N_7421);
xor U7552 (N_7552,N_7457,N_7400);
or U7553 (N_7553,N_7424,N_7417);
and U7554 (N_7554,N_7441,N_7481);
nor U7555 (N_7555,N_7466,N_7407);
and U7556 (N_7556,N_7401,N_7430);
nand U7557 (N_7557,N_7470,N_7362);
xnor U7558 (N_7558,N_7393,N_7437);
nor U7559 (N_7559,N_7467,N_7477);
xor U7560 (N_7560,N_7408,N_7369);
and U7561 (N_7561,N_7478,N_7443);
nand U7562 (N_7562,N_7431,N_7377);
nor U7563 (N_7563,N_7373,N_7374);
xnor U7564 (N_7564,N_7455,N_7418);
xnor U7565 (N_7565,N_7484,N_7486);
nor U7566 (N_7566,N_7395,N_7371);
nand U7567 (N_7567,N_7479,N_7463);
or U7568 (N_7568,N_7461,N_7425);
or U7569 (N_7569,N_7458,N_7448);
or U7570 (N_7570,N_7388,N_7447);
and U7571 (N_7571,N_7494,N_7442);
nor U7572 (N_7572,N_7372,N_7365);
xor U7573 (N_7573,N_7376,N_7450);
nand U7574 (N_7574,N_7456,N_7392);
xor U7575 (N_7575,N_7358,N_7425);
nor U7576 (N_7576,N_7357,N_7374);
nor U7577 (N_7577,N_7427,N_7469);
and U7578 (N_7578,N_7492,N_7465);
xor U7579 (N_7579,N_7383,N_7420);
xor U7580 (N_7580,N_7472,N_7468);
nor U7581 (N_7581,N_7427,N_7498);
and U7582 (N_7582,N_7450,N_7476);
and U7583 (N_7583,N_7380,N_7436);
and U7584 (N_7584,N_7393,N_7366);
or U7585 (N_7585,N_7408,N_7484);
and U7586 (N_7586,N_7436,N_7418);
xor U7587 (N_7587,N_7495,N_7499);
nand U7588 (N_7588,N_7438,N_7435);
nor U7589 (N_7589,N_7423,N_7369);
nand U7590 (N_7590,N_7425,N_7440);
and U7591 (N_7591,N_7398,N_7426);
or U7592 (N_7592,N_7387,N_7361);
nand U7593 (N_7593,N_7354,N_7460);
nor U7594 (N_7594,N_7395,N_7454);
or U7595 (N_7595,N_7453,N_7391);
and U7596 (N_7596,N_7360,N_7497);
xor U7597 (N_7597,N_7376,N_7474);
or U7598 (N_7598,N_7409,N_7485);
xnor U7599 (N_7599,N_7472,N_7454);
nor U7600 (N_7600,N_7432,N_7361);
nor U7601 (N_7601,N_7493,N_7367);
and U7602 (N_7602,N_7482,N_7398);
nor U7603 (N_7603,N_7476,N_7463);
or U7604 (N_7604,N_7386,N_7481);
xor U7605 (N_7605,N_7463,N_7442);
or U7606 (N_7606,N_7443,N_7380);
nand U7607 (N_7607,N_7397,N_7377);
or U7608 (N_7608,N_7358,N_7494);
nor U7609 (N_7609,N_7417,N_7460);
or U7610 (N_7610,N_7380,N_7390);
or U7611 (N_7611,N_7382,N_7424);
nand U7612 (N_7612,N_7477,N_7437);
nand U7613 (N_7613,N_7488,N_7392);
nor U7614 (N_7614,N_7353,N_7425);
and U7615 (N_7615,N_7437,N_7366);
nor U7616 (N_7616,N_7458,N_7492);
and U7617 (N_7617,N_7455,N_7446);
or U7618 (N_7618,N_7399,N_7379);
nand U7619 (N_7619,N_7464,N_7361);
xor U7620 (N_7620,N_7405,N_7474);
xnor U7621 (N_7621,N_7363,N_7498);
and U7622 (N_7622,N_7379,N_7463);
nor U7623 (N_7623,N_7454,N_7392);
nand U7624 (N_7624,N_7464,N_7460);
or U7625 (N_7625,N_7377,N_7399);
nor U7626 (N_7626,N_7368,N_7406);
nand U7627 (N_7627,N_7437,N_7459);
xnor U7628 (N_7628,N_7399,N_7410);
or U7629 (N_7629,N_7431,N_7415);
or U7630 (N_7630,N_7467,N_7384);
nor U7631 (N_7631,N_7454,N_7489);
nand U7632 (N_7632,N_7362,N_7459);
xor U7633 (N_7633,N_7415,N_7389);
nor U7634 (N_7634,N_7461,N_7384);
or U7635 (N_7635,N_7460,N_7388);
nor U7636 (N_7636,N_7404,N_7359);
nand U7637 (N_7637,N_7471,N_7373);
and U7638 (N_7638,N_7476,N_7462);
and U7639 (N_7639,N_7396,N_7496);
and U7640 (N_7640,N_7363,N_7408);
and U7641 (N_7641,N_7409,N_7463);
nand U7642 (N_7642,N_7368,N_7404);
nand U7643 (N_7643,N_7417,N_7467);
or U7644 (N_7644,N_7446,N_7424);
nor U7645 (N_7645,N_7360,N_7470);
xor U7646 (N_7646,N_7370,N_7380);
nor U7647 (N_7647,N_7383,N_7387);
xnor U7648 (N_7648,N_7367,N_7465);
and U7649 (N_7649,N_7427,N_7425);
or U7650 (N_7650,N_7597,N_7534);
nor U7651 (N_7651,N_7639,N_7635);
or U7652 (N_7652,N_7512,N_7541);
or U7653 (N_7653,N_7590,N_7624);
xnor U7654 (N_7654,N_7616,N_7647);
nor U7655 (N_7655,N_7544,N_7609);
and U7656 (N_7656,N_7613,N_7644);
nand U7657 (N_7657,N_7632,N_7628);
nand U7658 (N_7658,N_7587,N_7547);
and U7659 (N_7659,N_7535,N_7551);
xor U7660 (N_7660,N_7640,N_7615);
xor U7661 (N_7661,N_7565,N_7500);
nand U7662 (N_7662,N_7592,N_7508);
or U7663 (N_7663,N_7595,N_7564);
and U7664 (N_7664,N_7543,N_7603);
or U7665 (N_7665,N_7503,N_7571);
nand U7666 (N_7666,N_7510,N_7629);
or U7667 (N_7667,N_7588,N_7516);
and U7668 (N_7668,N_7630,N_7521);
nand U7669 (N_7669,N_7602,N_7507);
nand U7670 (N_7670,N_7612,N_7638);
nand U7671 (N_7671,N_7561,N_7617);
xnor U7672 (N_7672,N_7505,N_7594);
and U7673 (N_7673,N_7637,N_7600);
nand U7674 (N_7674,N_7502,N_7526);
and U7675 (N_7675,N_7531,N_7619);
nand U7676 (N_7676,N_7575,N_7589);
nor U7677 (N_7677,N_7542,N_7566);
or U7678 (N_7678,N_7536,N_7570);
nor U7679 (N_7679,N_7527,N_7643);
nor U7680 (N_7680,N_7524,N_7553);
nor U7681 (N_7681,N_7555,N_7529);
xnor U7682 (N_7682,N_7582,N_7598);
and U7683 (N_7683,N_7549,N_7533);
nand U7684 (N_7684,N_7601,N_7618);
and U7685 (N_7685,N_7614,N_7552);
xnor U7686 (N_7686,N_7559,N_7557);
and U7687 (N_7687,N_7579,N_7611);
or U7688 (N_7688,N_7623,N_7548);
or U7689 (N_7689,N_7581,N_7539);
or U7690 (N_7690,N_7525,N_7519);
nor U7691 (N_7691,N_7620,N_7591);
and U7692 (N_7692,N_7627,N_7608);
and U7693 (N_7693,N_7545,N_7626);
nor U7694 (N_7694,N_7578,N_7554);
nor U7695 (N_7695,N_7522,N_7514);
nand U7696 (N_7696,N_7648,N_7509);
and U7697 (N_7697,N_7631,N_7550);
nand U7698 (N_7698,N_7574,N_7537);
xnor U7699 (N_7699,N_7532,N_7605);
xor U7700 (N_7700,N_7584,N_7599);
nor U7701 (N_7701,N_7560,N_7538);
xor U7702 (N_7702,N_7585,N_7513);
xnor U7703 (N_7703,N_7523,N_7596);
nor U7704 (N_7704,N_7645,N_7556);
and U7705 (N_7705,N_7649,N_7593);
xor U7706 (N_7706,N_7518,N_7607);
nor U7707 (N_7707,N_7572,N_7576);
or U7708 (N_7708,N_7506,N_7563);
nor U7709 (N_7709,N_7562,N_7504);
nor U7710 (N_7710,N_7530,N_7568);
nor U7711 (N_7711,N_7642,N_7558);
or U7712 (N_7712,N_7636,N_7569);
nand U7713 (N_7713,N_7577,N_7646);
or U7714 (N_7714,N_7517,N_7610);
nor U7715 (N_7715,N_7604,N_7606);
or U7716 (N_7716,N_7501,N_7528);
xnor U7717 (N_7717,N_7511,N_7634);
and U7718 (N_7718,N_7546,N_7573);
nor U7719 (N_7719,N_7580,N_7586);
nand U7720 (N_7720,N_7641,N_7621);
nand U7721 (N_7721,N_7540,N_7622);
nand U7722 (N_7722,N_7633,N_7515);
or U7723 (N_7723,N_7567,N_7583);
nor U7724 (N_7724,N_7625,N_7520);
xnor U7725 (N_7725,N_7552,N_7587);
nor U7726 (N_7726,N_7524,N_7559);
and U7727 (N_7727,N_7581,N_7520);
nand U7728 (N_7728,N_7585,N_7620);
or U7729 (N_7729,N_7505,N_7549);
nor U7730 (N_7730,N_7638,N_7602);
xor U7731 (N_7731,N_7616,N_7635);
xor U7732 (N_7732,N_7631,N_7629);
or U7733 (N_7733,N_7609,N_7621);
nor U7734 (N_7734,N_7557,N_7614);
xor U7735 (N_7735,N_7619,N_7631);
nand U7736 (N_7736,N_7506,N_7510);
nand U7737 (N_7737,N_7640,N_7565);
nor U7738 (N_7738,N_7591,N_7563);
nor U7739 (N_7739,N_7619,N_7584);
nor U7740 (N_7740,N_7573,N_7620);
or U7741 (N_7741,N_7516,N_7565);
and U7742 (N_7742,N_7647,N_7641);
nand U7743 (N_7743,N_7614,N_7581);
nor U7744 (N_7744,N_7610,N_7530);
and U7745 (N_7745,N_7569,N_7502);
and U7746 (N_7746,N_7555,N_7516);
xnor U7747 (N_7747,N_7500,N_7570);
or U7748 (N_7748,N_7523,N_7560);
nand U7749 (N_7749,N_7594,N_7577);
and U7750 (N_7750,N_7620,N_7600);
xor U7751 (N_7751,N_7508,N_7566);
and U7752 (N_7752,N_7546,N_7532);
or U7753 (N_7753,N_7505,N_7512);
nand U7754 (N_7754,N_7611,N_7532);
nor U7755 (N_7755,N_7556,N_7567);
xor U7756 (N_7756,N_7557,N_7638);
xor U7757 (N_7757,N_7633,N_7642);
nor U7758 (N_7758,N_7587,N_7648);
or U7759 (N_7759,N_7521,N_7645);
and U7760 (N_7760,N_7541,N_7621);
nor U7761 (N_7761,N_7507,N_7561);
nand U7762 (N_7762,N_7587,N_7543);
nand U7763 (N_7763,N_7640,N_7502);
or U7764 (N_7764,N_7555,N_7605);
nand U7765 (N_7765,N_7518,N_7568);
xor U7766 (N_7766,N_7623,N_7568);
nor U7767 (N_7767,N_7536,N_7584);
nand U7768 (N_7768,N_7512,N_7557);
nand U7769 (N_7769,N_7595,N_7502);
nand U7770 (N_7770,N_7537,N_7629);
and U7771 (N_7771,N_7634,N_7566);
nor U7772 (N_7772,N_7605,N_7526);
xnor U7773 (N_7773,N_7639,N_7582);
nand U7774 (N_7774,N_7501,N_7511);
xnor U7775 (N_7775,N_7579,N_7519);
xnor U7776 (N_7776,N_7612,N_7572);
nor U7777 (N_7777,N_7583,N_7600);
nor U7778 (N_7778,N_7628,N_7592);
or U7779 (N_7779,N_7520,N_7573);
nand U7780 (N_7780,N_7502,N_7530);
nor U7781 (N_7781,N_7612,N_7586);
nor U7782 (N_7782,N_7549,N_7577);
and U7783 (N_7783,N_7504,N_7589);
xor U7784 (N_7784,N_7611,N_7625);
nor U7785 (N_7785,N_7583,N_7525);
or U7786 (N_7786,N_7646,N_7553);
xnor U7787 (N_7787,N_7545,N_7533);
xnor U7788 (N_7788,N_7538,N_7620);
xor U7789 (N_7789,N_7579,N_7642);
or U7790 (N_7790,N_7563,N_7642);
nor U7791 (N_7791,N_7551,N_7554);
and U7792 (N_7792,N_7548,N_7644);
or U7793 (N_7793,N_7598,N_7589);
or U7794 (N_7794,N_7638,N_7620);
or U7795 (N_7795,N_7630,N_7590);
and U7796 (N_7796,N_7548,N_7550);
xor U7797 (N_7797,N_7618,N_7505);
nand U7798 (N_7798,N_7622,N_7541);
xnor U7799 (N_7799,N_7536,N_7550);
or U7800 (N_7800,N_7756,N_7765);
nand U7801 (N_7801,N_7718,N_7726);
xor U7802 (N_7802,N_7670,N_7794);
nor U7803 (N_7803,N_7665,N_7752);
and U7804 (N_7804,N_7706,N_7710);
and U7805 (N_7805,N_7686,N_7714);
xnor U7806 (N_7806,N_7791,N_7763);
or U7807 (N_7807,N_7773,N_7667);
xor U7808 (N_7808,N_7780,N_7783);
and U7809 (N_7809,N_7777,N_7716);
or U7810 (N_7810,N_7717,N_7715);
or U7811 (N_7811,N_7700,N_7661);
and U7812 (N_7812,N_7733,N_7789);
xor U7813 (N_7813,N_7691,N_7734);
or U7814 (N_7814,N_7747,N_7785);
nand U7815 (N_7815,N_7720,N_7799);
nor U7816 (N_7816,N_7663,N_7725);
nor U7817 (N_7817,N_7739,N_7738);
and U7818 (N_7818,N_7659,N_7671);
and U7819 (N_7819,N_7724,N_7702);
nand U7820 (N_7820,N_7759,N_7682);
or U7821 (N_7821,N_7767,N_7786);
nand U7822 (N_7822,N_7798,N_7778);
and U7823 (N_7823,N_7771,N_7737);
nand U7824 (N_7824,N_7711,N_7776);
nand U7825 (N_7825,N_7770,N_7781);
or U7826 (N_7826,N_7701,N_7735);
and U7827 (N_7827,N_7736,N_7692);
and U7828 (N_7828,N_7787,N_7705);
nand U7829 (N_7829,N_7651,N_7774);
and U7830 (N_7830,N_7679,N_7695);
nor U7831 (N_7831,N_7760,N_7779);
xnor U7832 (N_7832,N_7660,N_7782);
or U7833 (N_7833,N_7723,N_7655);
xor U7834 (N_7834,N_7758,N_7708);
or U7835 (N_7835,N_7761,N_7664);
or U7836 (N_7836,N_7675,N_7790);
and U7837 (N_7837,N_7687,N_7743);
nand U7838 (N_7838,N_7668,N_7772);
and U7839 (N_7839,N_7719,N_7754);
nand U7840 (N_7840,N_7666,N_7797);
nand U7841 (N_7841,N_7680,N_7784);
or U7842 (N_7842,N_7697,N_7657);
and U7843 (N_7843,N_7730,N_7768);
xor U7844 (N_7844,N_7650,N_7757);
xnor U7845 (N_7845,N_7683,N_7678);
nor U7846 (N_7846,N_7685,N_7676);
nor U7847 (N_7847,N_7707,N_7775);
nor U7848 (N_7848,N_7689,N_7788);
and U7849 (N_7849,N_7658,N_7745);
nand U7850 (N_7850,N_7662,N_7793);
nand U7851 (N_7851,N_7755,N_7732);
nor U7852 (N_7852,N_7722,N_7690);
or U7853 (N_7853,N_7652,N_7713);
xnor U7854 (N_7854,N_7656,N_7728);
or U7855 (N_7855,N_7703,N_7704);
nand U7856 (N_7856,N_7672,N_7766);
and U7857 (N_7857,N_7693,N_7762);
xnor U7858 (N_7858,N_7696,N_7673);
and U7859 (N_7859,N_7694,N_7669);
xor U7860 (N_7860,N_7746,N_7674);
xor U7861 (N_7861,N_7740,N_7748);
or U7862 (N_7862,N_7653,N_7744);
nor U7863 (N_7863,N_7677,N_7769);
or U7864 (N_7864,N_7721,N_7742);
nor U7865 (N_7865,N_7751,N_7688);
xnor U7866 (N_7866,N_7731,N_7654);
and U7867 (N_7867,N_7698,N_7699);
xnor U7868 (N_7868,N_7795,N_7764);
or U7869 (N_7869,N_7727,N_7712);
or U7870 (N_7870,N_7753,N_7729);
nand U7871 (N_7871,N_7792,N_7749);
or U7872 (N_7872,N_7709,N_7741);
nand U7873 (N_7873,N_7796,N_7681);
and U7874 (N_7874,N_7750,N_7684);
nand U7875 (N_7875,N_7755,N_7691);
nand U7876 (N_7876,N_7727,N_7680);
xor U7877 (N_7877,N_7666,N_7717);
or U7878 (N_7878,N_7674,N_7652);
and U7879 (N_7879,N_7666,N_7740);
nor U7880 (N_7880,N_7792,N_7777);
nand U7881 (N_7881,N_7728,N_7719);
nand U7882 (N_7882,N_7695,N_7658);
nor U7883 (N_7883,N_7650,N_7732);
nor U7884 (N_7884,N_7758,N_7777);
xnor U7885 (N_7885,N_7654,N_7751);
nand U7886 (N_7886,N_7678,N_7654);
nor U7887 (N_7887,N_7657,N_7737);
xor U7888 (N_7888,N_7651,N_7725);
nand U7889 (N_7889,N_7742,N_7683);
nor U7890 (N_7890,N_7743,N_7777);
and U7891 (N_7891,N_7774,N_7680);
or U7892 (N_7892,N_7699,N_7744);
nor U7893 (N_7893,N_7717,N_7676);
nor U7894 (N_7894,N_7762,N_7663);
xor U7895 (N_7895,N_7693,N_7750);
xnor U7896 (N_7896,N_7719,N_7788);
nor U7897 (N_7897,N_7748,N_7744);
and U7898 (N_7898,N_7677,N_7717);
xor U7899 (N_7899,N_7742,N_7677);
and U7900 (N_7900,N_7651,N_7795);
and U7901 (N_7901,N_7783,N_7730);
nand U7902 (N_7902,N_7718,N_7700);
and U7903 (N_7903,N_7764,N_7726);
nand U7904 (N_7904,N_7793,N_7713);
xnor U7905 (N_7905,N_7750,N_7791);
or U7906 (N_7906,N_7659,N_7765);
and U7907 (N_7907,N_7741,N_7653);
nand U7908 (N_7908,N_7711,N_7725);
nand U7909 (N_7909,N_7745,N_7730);
or U7910 (N_7910,N_7700,N_7662);
xor U7911 (N_7911,N_7695,N_7718);
and U7912 (N_7912,N_7676,N_7793);
nor U7913 (N_7913,N_7674,N_7776);
and U7914 (N_7914,N_7712,N_7760);
nand U7915 (N_7915,N_7786,N_7768);
xnor U7916 (N_7916,N_7782,N_7795);
and U7917 (N_7917,N_7753,N_7769);
or U7918 (N_7918,N_7716,N_7798);
xor U7919 (N_7919,N_7664,N_7744);
nand U7920 (N_7920,N_7672,N_7689);
nor U7921 (N_7921,N_7686,N_7699);
or U7922 (N_7922,N_7774,N_7736);
nand U7923 (N_7923,N_7721,N_7668);
and U7924 (N_7924,N_7668,N_7780);
nor U7925 (N_7925,N_7670,N_7776);
xor U7926 (N_7926,N_7762,N_7669);
and U7927 (N_7927,N_7663,N_7688);
xnor U7928 (N_7928,N_7725,N_7664);
nor U7929 (N_7929,N_7696,N_7743);
and U7930 (N_7930,N_7757,N_7687);
or U7931 (N_7931,N_7735,N_7777);
nor U7932 (N_7932,N_7729,N_7663);
and U7933 (N_7933,N_7730,N_7702);
nor U7934 (N_7934,N_7674,N_7781);
or U7935 (N_7935,N_7712,N_7729);
nand U7936 (N_7936,N_7766,N_7753);
and U7937 (N_7937,N_7650,N_7659);
and U7938 (N_7938,N_7692,N_7680);
xor U7939 (N_7939,N_7766,N_7663);
and U7940 (N_7940,N_7789,N_7653);
or U7941 (N_7941,N_7792,N_7769);
and U7942 (N_7942,N_7777,N_7665);
nand U7943 (N_7943,N_7731,N_7660);
nor U7944 (N_7944,N_7695,N_7671);
nor U7945 (N_7945,N_7709,N_7712);
and U7946 (N_7946,N_7728,N_7702);
and U7947 (N_7947,N_7719,N_7699);
nor U7948 (N_7948,N_7745,N_7765);
xnor U7949 (N_7949,N_7681,N_7694);
and U7950 (N_7950,N_7831,N_7918);
and U7951 (N_7951,N_7822,N_7898);
or U7952 (N_7952,N_7938,N_7901);
nor U7953 (N_7953,N_7874,N_7817);
nand U7954 (N_7954,N_7800,N_7812);
nor U7955 (N_7955,N_7868,N_7891);
xor U7956 (N_7956,N_7866,N_7862);
nand U7957 (N_7957,N_7872,N_7844);
nor U7958 (N_7958,N_7813,N_7854);
and U7959 (N_7959,N_7913,N_7924);
xnor U7960 (N_7960,N_7807,N_7881);
xor U7961 (N_7961,N_7909,N_7832);
nand U7962 (N_7962,N_7803,N_7809);
nand U7963 (N_7963,N_7839,N_7821);
or U7964 (N_7964,N_7873,N_7816);
and U7965 (N_7965,N_7916,N_7882);
nor U7966 (N_7966,N_7945,N_7889);
or U7967 (N_7967,N_7936,N_7931);
and U7968 (N_7968,N_7858,N_7826);
and U7969 (N_7969,N_7937,N_7885);
or U7970 (N_7970,N_7919,N_7801);
xnor U7971 (N_7971,N_7879,N_7871);
nand U7972 (N_7972,N_7846,N_7927);
or U7973 (N_7973,N_7928,N_7864);
and U7974 (N_7974,N_7875,N_7946);
or U7975 (N_7975,N_7920,N_7930);
or U7976 (N_7976,N_7895,N_7841);
or U7977 (N_7977,N_7845,N_7933);
xor U7978 (N_7978,N_7894,N_7903);
and U7979 (N_7979,N_7949,N_7827);
and U7980 (N_7980,N_7917,N_7914);
xor U7981 (N_7981,N_7942,N_7867);
or U7982 (N_7982,N_7848,N_7834);
nand U7983 (N_7983,N_7940,N_7907);
nor U7984 (N_7984,N_7947,N_7838);
or U7985 (N_7985,N_7908,N_7906);
nor U7986 (N_7986,N_7855,N_7912);
nand U7987 (N_7987,N_7939,N_7880);
nor U7988 (N_7988,N_7828,N_7934);
xor U7989 (N_7989,N_7897,N_7863);
xor U7990 (N_7990,N_7837,N_7825);
nand U7991 (N_7991,N_7925,N_7853);
nor U7992 (N_7992,N_7888,N_7835);
and U7993 (N_7993,N_7829,N_7840);
and U7994 (N_7994,N_7824,N_7926);
and U7995 (N_7995,N_7887,N_7843);
and U7996 (N_7996,N_7860,N_7886);
nand U7997 (N_7997,N_7904,N_7850);
xor U7998 (N_7998,N_7856,N_7819);
or U7999 (N_7999,N_7842,N_7911);
or U8000 (N_8000,N_7847,N_7818);
and U8001 (N_8001,N_7833,N_7948);
and U8002 (N_8002,N_7857,N_7805);
or U8003 (N_8003,N_7902,N_7941);
nor U8004 (N_8004,N_7890,N_7899);
nand U8005 (N_8005,N_7814,N_7923);
nand U8006 (N_8006,N_7883,N_7922);
nand U8007 (N_8007,N_7877,N_7892);
or U8008 (N_8008,N_7878,N_7820);
nor U8009 (N_8009,N_7929,N_7852);
xor U8010 (N_8010,N_7804,N_7810);
and U8011 (N_8011,N_7932,N_7806);
or U8012 (N_8012,N_7944,N_7921);
or U8013 (N_8013,N_7808,N_7870);
and U8014 (N_8014,N_7861,N_7935);
nor U8015 (N_8015,N_7859,N_7836);
or U8016 (N_8016,N_7830,N_7884);
and U8017 (N_8017,N_7815,N_7943);
xor U8018 (N_8018,N_7849,N_7802);
xor U8019 (N_8019,N_7915,N_7893);
nor U8020 (N_8020,N_7910,N_7823);
and U8021 (N_8021,N_7851,N_7876);
or U8022 (N_8022,N_7811,N_7869);
nand U8023 (N_8023,N_7900,N_7905);
nand U8024 (N_8024,N_7865,N_7896);
or U8025 (N_8025,N_7821,N_7825);
nand U8026 (N_8026,N_7910,N_7913);
nor U8027 (N_8027,N_7839,N_7923);
or U8028 (N_8028,N_7875,N_7823);
nand U8029 (N_8029,N_7863,N_7914);
or U8030 (N_8030,N_7832,N_7863);
or U8031 (N_8031,N_7894,N_7802);
nand U8032 (N_8032,N_7916,N_7819);
or U8033 (N_8033,N_7884,N_7900);
nor U8034 (N_8034,N_7905,N_7812);
nor U8035 (N_8035,N_7815,N_7866);
nor U8036 (N_8036,N_7838,N_7813);
nor U8037 (N_8037,N_7867,N_7907);
nor U8038 (N_8038,N_7882,N_7935);
or U8039 (N_8039,N_7864,N_7868);
nand U8040 (N_8040,N_7838,N_7857);
xnor U8041 (N_8041,N_7855,N_7821);
or U8042 (N_8042,N_7900,N_7848);
or U8043 (N_8043,N_7916,N_7900);
or U8044 (N_8044,N_7912,N_7846);
nor U8045 (N_8045,N_7884,N_7848);
nor U8046 (N_8046,N_7944,N_7817);
nor U8047 (N_8047,N_7896,N_7833);
nand U8048 (N_8048,N_7833,N_7814);
xnor U8049 (N_8049,N_7897,N_7898);
nand U8050 (N_8050,N_7930,N_7912);
xnor U8051 (N_8051,N_7833,N_7863);
nand U8052 (N_8052,N_7856,N_7916);
or U8053 (N_8053,N_7892,N_7875);
nand U8054 (N_8054,N_7846,N_7865);
nor U8055 (N_8055,N_7883,N_7949);
xnor U8056 (N_8056,N_7897,N_7822);
and U8057 (N_8057,N_7937,N_7912);
xor U8058 (N_8058,N_7874,N_7883);
nand U8059 (N_8059,N_7935,N_7944);
nor U8060 (N_8060,N_7896,N_7868);
nand U8061 (N_8061,N_7862,N_7900);
nand U8062 (N_8062,N_7809,N_7862);
or U8063 (N_8063,N_7839,N_7888);
xnor U8064 (N_8064,N_7907,N_7816);
nand U8065 (N_8065,N_7930,N_7804);
or U8066 (N_8066,N_7915,N_7823);
nor U8067 (N_8067,N_7880,N_7887);
or U8068 (N_8068,N_7826,N_7906);
and U8069 (N_8069,N_7929,N_7877);
and U8070 (N_8070,N_7937,N_7893);
and U8071 (N_8071,N_7858,N_7841);
xor U8072 (N_8072,N_7929,N_7890);
xor U8073 (N_8073,N_7849,N_7819);
or U8074 (N_8074,N_7886,N_7872);
nand U8075 (N_8075,N_7943,N_7877);
and U8076 (N_8076,N_7835,N_7848);
nand U8077 (N_8077,N_7817,N_7949);
nand U8078 (N_8078,N_7867,N_7825);
or U8079 (N_8079,N_7868,N_7847);
and U8080 (N_8080,N_7858,N_7863);
nand U8081 (N_8081,N_7857,N_7908);
and U8082 (N_8082,N_7947,N_7863);
nor U8083 (N_8083,N_7854,N_7928);
xor U8084 (N_8084,N_7919,N_7888);
or U8085 (N_8085,N_7823,N_7830);
or U8086 (N_8086,N_7888,N_7930);
and U8087 (N_8087,N_7897,N_7868);
or U8088 (N_8088,N_7901,N_7845);
xnor U8089 (N_8089,N_7888,N_7866);
nand U8090 (N_8090,N_7899,N_7827);
xor U8091 (N_8091,N_7876,N_7906);
xor U8092 (N_8092,N_7902,N_7898);
nand U8093 (N_8093,N_7821,N_7833);
nand U8094 (N_8094,N_7875,N_7905);
or U8095 (N_8095,N_7858,N_7888);
or U8096 (N_8096,N_7938,N_7832);
and U8097 (N_8097,N_7825,N_7919);
nand U8098 (N_8098,N_7844,N_7902);
nor U8099 (N_8099,N_7832,N_7883);
or U8100 (N_8100,N_8087,N_7954);
or U8101 (N_8101,N_8033,N_7982);
or U8102 (N_8102,N_8001,N_8036);
xnor U8103 (N_8103,N_8012,N_8042);
nor U8104 (N_8104,N_8083,N_8008);
xnor U8105 (N_8105,N_8048,N_7964);
and U8106 (N_8106,N_8027,N_8068);
and U8107 (N_8107,N_7963,N_7961);
or U8108 (N_8108,N_7960,N_7950);
nand U8109 (N_8109,N_7997,N_7966);
nand U8110 (N_8110,N_8032,N_7969);
nand U8111 (N_8111,N_8056,N_8054);
or U8112 (N_8112,N_7955,N_8065);
xnor U8113 (N_8113,N_8069,N_8017);
nand U8114 (N_8114,N_8019,N_8058);
xnor U8115 (N_8115,N_7993,N_8067);
nor U8116 (N_8116,N_7986,N_8046);
xor U8117 (N_8117,N_8084,N_8039);
xnor U8118 (N_8118,N_8085,N_8002);
xor U8119 (N_8119,N_7971,N_8013);
or U8120 (N_8120,N_8057,N_8071);
and U8121 (N_8121,N_8040,N_7953);
nor U8122 (N_8122,N_8023,N_7985);
xnor U8123 (N_8123,N_8079,N_7977);
and U8124 (N_8124,N_8059,N_8096);
and U8125 (N_8125,N_8031,N_8082);
nand U8126 (N_8126,N_8037,N_7983);
or U8127 (N_8127,N_8041,N_8081);
xor U8128 (N_8128,N_7989,N_7958);
or U8129 (N_8129,N_7970,N_8094);
xor U8130 (N_8130,N_8070,N_7990);
xnor U8131 (N_8131,N_7972,N_7956);
and U8132 (N_8132,N_8074,N_8011);
and U8133 (N_8133,N_8007,N_8003);
nand U8134 (N_8134,N_8015,N_7978);
or U8135 (N_8135,N_7968,N_8075);
xor U8136 (N_8136,N_8016,N_8086);
nor U8137 (N_8137,N_8073,N_8098);
nor U8138 (N_8138,N_8030,N_7974);
and U8139 (N_8139,N_7952,N_8095);
and U8140 (N_8140,N_7981,N_8022);
nand U8141 (N_8141,N_8091,N_7962);
and U8142 (N_8142,N_8009,N_7979);
nor U8143 (N_8143,N_7976,N_8004);
nand U8144 (N_8144,N_8029,N_8062);
nor U8145 (N_8145,N_7999,N_7965);
nand U8146 (N_8146,N_8034,N_8099);
and U8147 (N_8147,N_8090,N_7973);
nand U8148 (N_8148,N_8018,N_7957);
nand U8149 (N_8149,N_8053,N_8035);
or U8150 (N_8150,N_8006,N_8049);
and U8151 (N_8151,N_8066,N_8072);
and U8152 (N_8152,N_7959,N_8088);
and U8153 (N_8153,N_7975,N_8092);
nor U8154 (N_8154,N_7991,N_8064);
xor U8155 (N_8155,N_8077,N_7998);
xnor U8156 (N_8156,N_8021,N_8050);
and U8157 (N_8157,N_8028,N_8014);
and U8158 (N_8158,N_7988,N_8044);
or U8159 (N_8159,N_8051,N_7995);
nand U8160 (N_8160,N_7980,N_8043);
nor U8161 (N_8161,N_8010,N_7987);
xor U8162 (N_8162,N_8061,N_8060);
xnor U8163 (N_8163,N_8045,N_7994);
xor U8164 (N_8164,N_8080,N_8000);
xor U8165 (N_8165,N_8026,N_8055);
xnor U8166 (N_8166,N_8005,N_7992);
or U8167 (N_8167,N_8024,N_8052);
or U8168 (N_8168,N_7967,N_8097);
or U8169 (N_8169,N_7984,N_7951);
nand U8170 (N_8170,N_8076,N_8093);
xnor U8171 (N_8171,N_7996,N_8063);
or U8172 (N_8172,N_8089,N_8078);
nand U8173 (N_8173,N_8020,N_8047);
xor U8174 (N_8174,N_8038,N_8025);
and U8175 (N_8175,N_7970,N_7988);
nor U8176 (N_8176,N_8052,N_7989);
xnor U8177 (N_8177,N_7976,N_7967);
xnor U8178 (N_8178,N_8048,N_7982);
and U8179 (N_8179,N_7974,N_7980);
and U8180 (N_8180,N_7958,N_8016);
nand U8181 (N_8181,N_8025,N_7972);
nor U8182 (N_8182,N_7991,N_7981);
xor U8183 (N_8183,N_8031,N_8057);
or U8184 (N_8184,N_7970,N_8067);
xor U8185 (N_8185,N_8029,N_7993);
nor U8186 (N_8186,N_8003,N_8094);
and U8187 (N_8187,N_7962,N_7974);
and U8188 (N_8188,N_7973,N_8095);
xnor U8189 (N_8189,N_7959,N_8034);
and U8190 (N_8190,N_7985,N_8071);
xnor U8191 (N_8191,N_8084,N_7961);
or U8192 (N_8192,N_8067,N_8022);
nand U8193 (N_8193,N_8064,N_7980);
nor U8194 (N_8194,N_8078,N_7973);
or U8195 (N_8195,N_7968,N_8069);
nor U8196 (N_8196,N_8078,N_7983);
or U8197 (N_8197,N_7995,N_7992);
xnor U8198 (N_8198,N_7979,N_8085);
nand U8199 (N_8199,N_8018,N_7995);
and U8200 (N_8200,N_8058,N_8077);
or U8201 (N_8201,N_7989,N_8004);
or U8202 (N_8202,N_8047,N_8092);
or U8203 (N_8203,N_8064,N_8027);
xnor U8204 (N_8204,N_7993,N_8025);
nor U8205 (N_8205,N_7966,N_8011);
and U8206 (N_8206,N_7985,N_8025);
nor U8207 (N_8207,N_7996,N_7951);
and U8208 (N_8208,N_8064,N_7995);
xor U8209 (N_8209,N_8091,N_8045);
nor U8210 (N_8210,N_7955,N_8069);
or U8211 (N_8211,N_7963,N_7959);
or U8212 (N_8212,N_8041,N_8033);
xor U8213 (N_8213,N_7998,N_8056);
nor U8214 (N_8214,N_8021,N_7973);
nand U8215 (N_8215,N_8061,N_8063);
and U8216 (N_8216,N_8096,N_8056);
or U8217 (N_8217,N_8071,N_8099);
and U8218 (N_8218,N_8070,N_8088);
and U8219 (N_8219,N_7978,N_8041);
and U8220 (N_8220,N_8065,N_7950);
nor U8221 (N_8221,N_7960,N_8053);
and U8222 (N_8222,N_8000,N_8042);
nand U8223 (N_8223,N_8099,N_8042);
xnor U8224 (N_8224,N_8096,N_7961);
xnor U8225 (N_8225,N_7983,N_8097);
nand U8226 (N_8226,N_7959,N_8049);
xnor U8227 (N_8227,N_8011,N_8041);
or U8228 (N_8228,N_8015,N_8032);
xor U8229 (N_8229,N_8047,N_8005);
xnor U8230 (N_8230,N_8049,N_7999);
and U8231 (N_8231,N_8019,N_7995);
xnor U8232 (N_8232,N_8055,N_8088);
or U8233 (N_8233,N_7959,N_8089);
nor U8234 (N_8234,N_8035,N_8048);
nor U8235 (N_8235,N_8077,N_8019);
or U8236 (N_8236,N_7951,N_8086);
or U8237 (N_8237,N_7955,N_8001);
xnor U8238 (N_8238,N_8033,N_8011);
nand U8239 (N_8239,N_7955,N_8072);
nor U8240 (N_8240,N_8059,N_7995);
nor U8241 (N_8241,N_8074,N_8092);
nand U8242 (N_8242,N_7971,N_8034);
xor U8243 (N_8243,N_7994,N_8009);
or U8244 (N_8244,N_8034,N_8003);
xnor U8245 (N_8245,N_8000,N_7999);
nor U8246 (N_8246,N_8029,N_8060);
xor U8247 (N_8247,N_8096,N_8019);
nand U8248 (N_8248,N_8084,N_7990);
and U8249 (N_8249,N_7999,N_7988);
xnor U8250 (N_8250,N_8115,N_8125);
or U8251 (N_8251,N_8229,N_8116);
nor U8252 (N_8252,N_8205,N_8148);
nand U8253 (N_8253,N_8104,N_8233);
xor U8254 (N_8254,N_8149,N_8172);
nand U8255 (N_8255,N_8230,N_8166);
or U8256 (N_8256,N_8112,N_8177);
xor U8257 (N_8257,N_8106,N_8170);
xor U8258 (N_8258,N_8173,N_8196);
and U8259 (N_8259,N_8247,N_8193);
nand U8260 (N_8260,N_8227,N_8128);
nand U8261 (N_8261,N_8130,N_8198);
and U8262 (N_8262,N_8140,N_8246);
and U8263 (N_8263,N_8175,N_8113);
and U8264 (N_8264,N_8179,N_8162);
xnor U8265 (N_8265,N_8176,N_8123);
and U8266 (N_8266,N_8185,N_8117);
and U8267 (N_8267,N_8114,N_8225);
nor U8268 (N_8268,N_8232,N_8110);
and U8269 (N_8269,N_8142,N_8226);
nand U8270 (N_8270,N_8224,N_8127);
and U8271 (N_8271,N_8222,N_8152);
xor U8272 (N_8272,N_8167,N_8191);
and U8273 (N_8273,N_8192,N_8101);
xor U8274 (N_8274,N_8122,N_8118);
or U8275 (N_8275,N_8241,N_8200);
nor U8276 (N_8276,N_8219,N_8223);
nor U8277 (N_8277,N_8242,N_8245);
and U8278 (N_8278,N_8195,N_8214);
nand U8279 (N_8279,N_8157,N_8206);
xnor U8280 (N_8280,N_8169,N_8138);
nand U8281 (N_8281,N_8102,N_8188);
and U8282 (N_8282,N_8126,N_8178);
xor U8283 (N_8283,N_8215,N_8109);
nor U8284 (N_8284,N_8124,N_8105);
nor U8285 (N_8285,N_8100,N_8136);
or U8286 (N_8286,N_8171,N_8147);
or U8287 (N_8287,N_8207,N_8133);
xor U8288 (N_8288,N_8190,N_8180);
xnor U8289 (N_8289,N_8160,N_8135);
or U8290 (N_8290,N_8197,N_8249);
xnor U8291 (N_8291,N_8211,N_8201);
nor U8292 (N_8292,N_8209,N_8202);
nor U8293 (N_8293,N_8213,N_8164);
nand U8294 (N_8294,N_8131,N_8199);
and U8295 (N_8295,N_8186,N_8120);
and U8296 (N_8296,N_8174,N_8103);
nor U8297 (N_8297,N_8203,N_8163);
nand U8298 (N_8298,N_8240,N_8220);
nor U8299 (N_8299,N_8243,N_8137);
or U8300 (N_8300,N_8151,N_8239);
and U8301 (N_8301,N_8187,N_8237);
nand U8302 (N_8302,N_8119,N_8221);
xnor U8303 (N_8303,N_8235,N_8168);
nand U8304 (N_8304,N_8210,N_8181);
or U8305 (N_8305,N_8111,N_8212);
nor U8306 (N_8306,N_8165,N_8143);
and U8307 (N_8307,N_8217,N_8139);
nand U8308 (N_8308,N_8236,N_8108);
or U8309 (N_8309,N_8150,N_8154);
or U8310 (N_8310,N_8182,N_8216);
and U8311 (N_8311,N_8158,N_8129);
and U8312 (N_8312,N_8144,N_8189);
xor U8313 (N_8313,N_8132,N_8153);
nor U8314 (N_8314,N_8146,N_8121);
xnor U8315 (N_8315,N_8107,N_8183);
nor U8316 (N_8316,N_8155,N_8134);
or U8317 (N_8317,N_8194,N_8141);
and U8318 (N_8318,N_8218,N_8156);
xor U8319 (N_8319,N_8238,N_8145);
nor U8320 (N_8320,N_8234,N_8208);
or U8321 (N_8321,N_8244,N_8231);
nor U8322 (N_8322,N_8228,N_8184);
nand U8323 (N_8323,N_8248,N_8161);
nand U8324 (N_8324,N_8159,N_8204);
or U8325 (N_8325,N_8225,N_8153);
and U8326 (N_8326,N_8201,N_8163);
and U8327 (N_8327,N_8201,N_8204);
nand U8328 (N_8328,N_8150,N_8185);
nor U8329 (N_8329,N_8128,N_8197);
xnor U8330 (N_8330,N_8151,N_8211);
and U8331 (N_8331,N_8249,N_8240);
and U8332 (N_8332,N_8227,N_8219);
nor U8333 (N_8333,N_8224,N_8216);
or U8334 (N_8334,N_8100,N_8245);
nor U8335 (N_8335,N_8170,N_8203);
xor U8336 (N_8336,N_8216,N_8223);
nand U8337 (N_8337,N_8246,N_8208);
nor U8338 (N_8338,N_8199,N_8102);
nand U8339 (N_8339,N_8137,N_8192);
nand U8340 (N_8340,N_8118,N_8191);
or U8341 (N_8341,N_8139,N_8107);
xor U8342 (N_8342,N_8180,N_8101);
nand U8343 (N_8343,N_8184,N_8163);
nor U8344 (N_8344,N_8192,N_8225);
xnor U8345 (N_8345,N_8121,N_8201);
and U8346 (N_8346,N_8236,N_8222);
xor U8347 (N_8347,N_8143,N_8146);
nand U8348 (N_8348,N_8151,N_8142);
or U8349 (N_8349,N_8141,N_8189);
or U8350 (N_8350,N_8146,N_8205);
nand U8351 (N_8351,N_8239,N_8177);
and U8352 (N_8352,N_8217,N_8165);
nor U8353 (N_8353,N_8149,N_8153);
xnor U8354 (N_8354,N_8100,N_8175);
nor U8355 (N_8355,N_8138,N_8104);
xnor U8356 (N_8356,N_8236,N_8195);
and U8357 (N_8357,N_8188,N_8146);
nand U8358 (N_8358,N_8104,N_8134);
or U8359 (N_8359,N_8165,N_8245);
and U8360 (N_8360,N_8244,N_8104);
nand U8361 (N_8361,N_8236,N_8243);
nor U8362 (N_8362,N_8215,N_8186);
or U8363 (N_8363,N_8127,N_8200);
xnor U8364 (N_8364,N_8200,N_8186);
nor U8365 (N_8365,N_8122,N_8107);
xnor U8366 (N_8366,N_8136,N_8144);
nand U8367 (N_8367,N_8213,N_8122);
or U8368 (N_8368,N_8126,N_8195);
or U8369 (N_8369,N_8164,N_8193);
or U8370 (N_8370,N_8203,N_8200);
or U8371 (N_8371,N_8110,N_8219);
and U8372 (N_8372,N_8208,N_8188);
nand U8373 (N_8373,N_8112,N_8239);
nor U8374 (N_8374,N_8127,N_8142);
xor U8375 (N_8375,N_8243,N_8249);
and U8376 (N_8376,N_8175,N_8210);
or U8377 (N_8377,N_8158,N_8214);
or U8378 (N_8378,N_8129,N_8204);
xor U8379 (N_8379,N_8123,N_8248);
nor U8380 (N_8380,N_8104,N_8198);
and U8381 (N_8381,N_8183,N_8202);
and U8382 (N_8382,N_8242,N_8115);
xor U8383 (N_8383,N_8166,N_8165);
xnor U8384 (N_8384,N_8125,N_8187);
or U8385 (N_8385,N_8106,N_8113);
nor U8386 (N_8386,N_8140,N_8133);
nor U8387 (N_8387,N_8104,N_8179);
or U8388 (N_8388,N_8127,N_8249);
nand U8389 (N_8389,N_8244,N_8236);
or U8390 (N_8390,N_8127,N_8188);
nor U8391 (N_8391,N_8189,N_8148);
and U8392 (N_8392,N_8105,N_8205);
or U8393 (N_8393,N_8114,N_8244);
nand U8394 (N_8394,N_8169,N_8191);
xor U8395 (N_8395,N_8178,N_8174);
or U8396 (N_8396,N_8229,N_8196);
or U8397 (N_8397,N_8116,N_8134);
nand U8398 (N_8398,N_8156,N_8209);
and U8399 (N_8399,N_8123,N_8191);
nand U8400 (N_8400,N_8371,N_8336);
nand U8401 (N_8401,N_8323,N_8311);
nand U8402 (N_8402,N_8340,N_8356);
nor U8403 (N_8403,N_8398,N_8316);
and U8404 (N_8404,N_8285,N_8363);
and U8405 (N_8405,N_8362,N_8360);
and U8406 (N_8406,N_8333,N_8388);
or U8407 (N_8407,N_8276,N_8332);
nand U8408 (N_8408,N_8295,N_8394);
or U8409 (N_8409,N_8357,N_8320);
nor U8410 (N_8410,N_8325,N_8393);
xor U8411 (N_8411,N_8344,N_8261);
or U8412 (N_8412,N_8339,N_8262);
and U8413 (N_8413,N_8345,N_8352);
nor U8414 (N_8414,N_8373,N_8370);
or U8415 (N_8415,N_8268,N_8353);
or U8416 (N_8416,N_8264,N_8267);
nor U8417 (N_8417,N_8305,N_8342);
and U8418 (N_8418,N_8379,N_8318);
and U8419 (N_8419,N_8386,N_8365);
xor U8420 (N_8420,N_8251,N_8266);
nor U8421 (N_8421,N_8296,N_8389);
xor U8422 (N_8422,N_8322,N_8275);
nor U8423 (N_8423,N_8335,N_8255);
nand U8424 (N_8424,N_8330,N_8263);
or U8425 (N_8425,N_8271,N_8286);
nand U8426 (N_8426,N_8265,N_8297);
nor U8427 (N_8427,N_8390,N_8272);
xnor U8428 (N_8428,N_8299,N_8348);
nand U8429 (N_8429,N_8376,N_8387);
nor U8430 (N_8430,N_8378,N_8312);
or U8431 (N_8431,N_8396,N_8327);
nor U8432 (N_8432,N_8274,N_8382);
xor U8433 (N_8433,N_8321,N_8253);
xor U8434 (N_8434,N_8331,N_8392);
or U8435 (N_8435,N_8367,N_8315);
xnor U8436 (N_8436,N_8338,N_8347);
xor U8437 (N_8437,N_8313,N_8281);
xor U8438 (N_8438,N_8397,N_8283);
and U8439 (N_8439,N_8391,N_8328);
xor U8440 (N_8440,N_8346,N_8309);
xor U8441 (N_8441,N_8364,N_8301);
nor U8442 (N_8442,N_8257,N_8359);
or U8443 (N_8443,N_8399,N_8302);
nor U8444 (N_8444,N_8288,N_8258);
xnor U8445 (N_8445,N_8350,N_8290);
nand U8446 (N_8446,N_8254,N_8374);
nor U8447 (N_8447,N_8384,N_8292);
nand U8448 (N_8448,N_8372,N_8343);
xnor U8449 (N_8449,N_8307,N_8334);
nand U8450 (N_8450,N_8280,N_8260);
or U8451 (N_8451,N_8369,N_8358);
xnor U8452 (N_8452,N_8279,N_8270);
or U8453 (N_8453,N_8304,N_8375);
and U8454 (N_8454,N_8250,N_8273);
and U8455 (N_8455,N_8368,N_8317);
or U8456 (N_8456,N_8308,N_8351);
nand U8457 (N_8457,N_8341,N_8366);
or U8458 (N_8458,N_8329,N_8355);
xnor U8459 (N_8459,N_8337,N_8269);
or U8460 (N_8460,N_8293,N_8303);
or U8461 (N_8461,N_8294,N_8282);
nor U8462 (N_8462,N_8380,N_8319);
xnor U8463 (N_8463,N_8300,N_8349);
or U8464 (N_8464,N_8395,N_8287);
nand U8465 (N_8465,N_8289,N_8291);
xor U8466 (N_8466,N_8381,N_8361);
nand U8467 (N_8467,N_8306,N_8324);
or U8468 (N_8468,N_8298,N_8314);
xnor U8469 (N_8469,N_8354,N_8377);
xnor U8470 (N_8470,N_8256,N_8278);
nand U8471 (N_8471,N_8277,N_8383);
nor U8472 (N_8472,N_8252,N_8326);
nor U8473 (N_8473,N_8385,N_8310);
nand U8474 (N_8474,N_8259,N_8284);
and U8475 (N_8475,N_8283,N_8292);
nand U8476 (N_8476,N_8399,N_8307);
xor U8477 (N_8477,N_8329,N_8396);
xor U8478 (N_8478,N_8309,N_8349);
or U8479 (N_8479,N_8397,N_8325);
xnor U8480 (N_8480,N_8317,N_8301);
nor U8481 (N_8481,N_8329,N_8293);
xnor U8482 (N_8482,N_8344,N_8363);
or U8483 (N_8483,N_8324,N_8337);
or U8484 (N_8484,N_8356,N_8344);
nor U8485 (N_8485,N_8329,N_8269);
nand U8486 (N_8486,N_8251,N_8334);
xor U8487 (N_8487,N_8391,N_8397);
and U8488 (N_8488,N_8257,N_8270);
or U8489 (N_8489,N_8391,N_8258);
nor U8490 (N_8490,N_8357,N_8256);
nor U8491 (N_8491,N_8334,N_8293);
and U8492 (N_8492,N_8269,N_8303);
nor U8493 (N_8493,N_8255,N_8270);
or U8494 (N_8494,N_8268,N_8377);
nor U8495 (N_8495,N_8258,N_8327);
or U8496 (N_8496,N_8318,N_8327);
nor U8497 (N_8497,N_8396,N_8278);
and U8498 (N_8498,N_8278,N_8261);
nand U8499 (N_8499,N_8263,N_8375);
xnor U8500 (N_8500,N_8350,N_8330);
nand U8501 (N_8501,N_8328,N_8289);
xnor U8502 (N_8502,N_8372,N_8352);
xnor U8503 (N_8503,N_8269,N_8352);
nor U8504 (N_8504,N_8283,N_8325);
and U8505 (N_8505,N_8370,N_8312);
xor U8506 (N_8506,N_8288,N_8309);
or U8507 (N_8507,N_8312,N_8366);
nand U8508 (N_8508,N_8281,N_8332);
and U8509 (N_8509,N_8399,N_8377);
or U8510 (N_8510,N_8334,N_8263);
nand U8511 (N_8511,N_8345,N_8371);
or U8512 (N_8512,N_8328,N_8306);
xor U8513 (N_8513,N_8341,N_8312);
nand U8514 (N_8514,N_8307,N_8274);
nand U8515 (N_8515,N_8344,N_8278);
nor U8516 (N_8516,N_8256,N_8398);
nand U8517 (N_8517,N_8311,N_8305);
nor U8518 (N_8518,N_8274,N_8335);
and U8519 (N_8519,N_8333,N_8296);
and U8520 (N_8520,N_8350,N_8316);
nand U8521 (N_8521,N_8379,N_8390);
or U8522 (N_8522,N_8277,N_8363);
nor U8523 (N_8523,N_8289,N_8338);
nand U8524 (N_8524,N_8361,N_8360);
and U8525 (N_8525,N_8379,N_8255);
xor U8526 (N_8526,N_8382,N_8371);
nand U8527 (N_8527,N_8354,N_8313);
xor U8528 (N_8528,N_8327,N_8357);
and U8529 (N_8529,N_8327,N_8365);
nand U8530 (N_8530,N_8398,N_8326);
nor U8531 (N_8531,N_8296,N_8323);
nand U8532 (N_8532,N_8387,N_8357);
nor U8533 (N_8533,N_8314,N_8293);
and U8534 (N_8534,N_8257,N_8338);
and U8535 (N_8535,N_8371,N_8352);
or U8536 (N_8536,N_8378,N_8344);
or U8537 (N_8537,N_8273,N_8310);
nor U8538 (N_8538,N_8296,N_8346);
and U8539 (N_8539,N_8304,N_8331);
and U8540 (N_8540,N_8310,N_8378);
xnor U8541 (N_8541,N_8369,N_8260);
and U8542 (N_8542,N_8348,N_8262);
and U8543 (N_8543,N_8374,N_8302);
nor U8544 (N_8544,N_8385,N_8303);
xnor U8545 (N_8545,N_8271,N_8305);
and U8546 (N_8546,N_8379,N_8320);
xnor U8547 (N_8547,N_8338,N_8263);
nor U8548 (N_8548,N_8320,N_8350);
or U8549 (N_8549,N_8382,N_8303);
xnor U8550 (N_8550,N_8441,N_8503);
nor U8551 (N_8551,N_8417,N_8421);
nor U8552 (N_8552,N_8459,N_8416);
nand U8553 (N_8553,N_8487,N_8483);
or U8554 (N_8554,N_8400,N_8440);
or U8555 (N_8555,N_8431,N_8497);
xor U8556 (N_8556,N_8485,N_8525);
xor U8557 (N_8557,N_8473,N_8438);
nand U8558 (N_8558,N_8546,N_8463);
nand U8559 (N_8559,N_8527,N_8450);
or U8560 (N_8560,N_8436,N_8469);
or U8561 (N_8561,N_8401,N_8434);
and U8562 (N_8562,N_8449,N_8447);
or U8563 (N_8563,N_8460,N_8515);
or U8564 (N_8564,N_8536,N_8549);
nand U8565 (N_8565,N_8462,N_8425);
nor U8566 (N_8566,N_8540,N_8454);
nor U8567 (N_8567,N_8418,N_8465);
xnor U8568 (N_8568,N_8533,N_8486);
xor U8569 (N_8569,N_8482,N_8535);
and U8570 (N_8570,N_8439,N_8492);
and U8571 (N_8571,N_8461,N_8548);
nand U8572 (N_8572,N_8408,N_8423);
xor U8573 (N_8573,N_8537,N_8442);
and U8574 (N_8574,N_8522,N_8452);
or U8575 (N_8575,N_8538,N_8526);
nand U8576 (N_8576,N_8455,N_8518);
nand U8577 (N_8577,N_8498,N_8470);
nand U8578 (N_8578,N_8477,N_8491);
xor U8579 (N_8579,N_8542,N_8507);
nand U8580 (N_8580,N_8410,N_8456);
nand U8581 (N_8581,N_8453,N_8409);
xor U8582 (N_8582,N_8475,N_8407);
nor U8583 (N_8583,N_8494,N_8468);
and U8584 (N_8584,N_8541,N_8504);
nor U8585 (N_8585,N_8406,N_8457);
or U8586 (N_8586,N_8509,N_8432);
nand U8587 (N_8587,N_8495,N_8530);
nor U8588 (N_8588,N_8404,N_8435);
or U8589 (N_8589,N_8443,N_8430);
and U8590 (N_8590,N_8528,N_8414);
and U8591 (N_8591,N_8471,N_8499);
or U8592 (N_8592,N_8479,N_8405);
nand U8593 (N_8593,N_8481,N_8412);
or U8594 (N_8594,N_8484,N_8508);
nand U8595 (N_8595,N_8428,N_8458);
and U8596 (N_8596,N_8480,N_8501);
xor U8597 (N_8597,N_8516,N_8513);
xnor U8598 (N_8598,N_8532,N_8433);
and U8599 (N_8599,N_8427,N_8420);
and U8600 (N_8600,N_8493,N_8545);
nor U8601 (N_8601,N_8444,N_8539);
and U8602 (N_8602,N_8520,N_8500);
and U8603 (N_8603,N_8415,N_8472);
or U8604 (N_8604,N_8413,N_8402);
and U8605 (N_8605,N_8411,N_8517);
and U8606 (N_8606,N_8464,N_8512);
nand U8607 (N_8607,N_8524,N_8424);
or U8608 (N_8608,N_8451,N_8490);
and U8609 (N_8609,N_8489,N_8437);
xnor U8610 (N_8610,N_8502,N_8478);
xnor U8611 (N_8611,N_8544,N_8534);
nor U8612 (N_8612,N_8426,N_8506);
xor U8613 (N_8613,N_8505,N_8543);
xnor U8614 (N_8614,N_8474,N_8547);
and U8615 (N_8615,N_8403,N_8476);
or U8616 (N_8616,N_8511,N_8488);
nor U8617 (N_8617,N_8445,N_8529);
or U8618 (N_8618,N_8448,N_8496);
or U8619 (N_8619,N_8519,N_8422);
and U8620 (N_8620,N_8429,N_8467);
or U8621 (N_8621,N_8419,N_8521);
or U8622 (N_8622,N_8466,N_8510);
xor U8623 (N_8623,N_8446,N_8514);
xnor U8624 (N_8624,N_8523,N_8531);
nor U8625 (N_8625,N_8549,N_8476);
nor U8626 (N_8626,N_8505,N_8539);
nand U8627 (N_8627,N_8536,N_8441);
nor U8628 (N_8628,N_8450,N_8514);
and U8629 (N_8629,N_8508,N_8431);
and U8630 (N_8630,N_8491,N_8535);
or U8631 (N_8631,N_8407,N_8531);
nand U8632 (N_8632,N_8525,N_8518);
nor U8633 (N_8633,N_8445,N_8495);
xor U8634 (N_8634,N_8465,N_8478);
or U8635 (N_8635,N_8473,N_8436);
nor U8636 (N_8636,N_8517,N_8524);
nand U8637 (N_8637,N_8442,N_8502);
nand U8638 (N_8638,N_8433,N_8421);
nand U8639 (N_8639,N_8522,N_8400);
nor U8640 (N_8640,N_8524,N_8527);
and U8641 (N_8641,N_8402,N_8461);
nand U8642 (N_8642,N_8506,N_8464);
and U8643 (N_8643,N_8511,N_8501);
and U8644 (N_8644,N_8523,N_8434);
and U8645 (N_8645,N_8419,N_8462);
and U8646 (N_8646,N_8543,N_8420);
nand U8647 (N_8647,N_8421,N_8530);
and U8648 (N_8648,N_8415,N_8478);
or U8649 (N_8649,N_8411,N_8464);
xor U8650 (N_8650,N_8444,N_8500);
or U8651 (N_8651,N_8406,N_8489);
or U8652 (N_8652,N_8452,N_8407);
nor U8653 (N_8653,N_8498,N_8416);
and U8654 (N_8654,N_8452,N_8520);
xnor U8655 (N_8655,N_8532,N_8458);
xor U8656 (N_8656,N_8432,N_8464);
xor U8657 (N_8657,N_8527,N_8539);
nand U8658 (N_8658,N_8415,N_8524);
nor U8659 (N_8659,N_8426,N_8418);
and U8660 (N_8660,N_8518,N_8504);
nor U8661 (N_8661,N_8490,N_8492);
nor U8662 (N_8662,N_8437,N_8472);
xnor U8663 (N_8663,N_8402,N_8405);
nand U8664 (N_8664,N_8407,N_8496);
and U8665 (N_8665,N_8506,N_8548);
or U8666 (N_8666,N_8535,N_8496);
nand U8667 (N_8667,N_8446,N_8525);
or U8668 (N_8668,N_8402,N_8487);
and U8669 (N_8669,N_8508,N_8429);
or U8670 (N_8670,N_8539,N_8508);
and U8671 (N_8671,N_8527,N_8523);
nor U8672 (N_8672,N_8447,N_8484);
nand U8673 (N_8673,N_8518,N_8522);
and U8674 (N_8674,N_8544,N_8514);
nand U8675 (N_8675,N_8416,N_8427);
nand U8676 (N_8676,N_8521,N_8458);
xnor U8677 (N_8677,N_8534,N_8434);
or U8678 (N_8678,N_8524,N_8461);
or U8679 (N_8679,N_8505,N_8439);
and U8680 (N_8680,N_8483,N_8427);
and U8681 (N_8681,N_8523,N_8437);
xor U8682 (N_8682,N_8455,N_8419);
or U8683 (N_8683,N_8539,N_8523);
or U8684 (N_8684,N_8488,N_8479);
xor U8685 (N_8685,N_8445,N_8428);
and U8686 (N_8686,N_8465,N_8488);
xnor U8687 (N_8687,N_8547,N_8511);
nand U8688 (N_8688,N_8489,N_8472);
and U8689 (N_8689,N_8412,N_8430);
xnor U8690 (N_8690,N_8513,N_8458);
nand U8691 (N_8691,N_8461,N_8438);
xnor U8692 (N_8692,N_8471,N_8411);
nor U8693 (N_8693,N_8517,N_8508);
nor U8694 (N_8694,N_8411,N_8515);
and U8695 (N_8695,N_8532,N_8482);
nand U8696 (N_8696,N_8517,N_8487);
nor U8697 (N_8697,N_8517,N_8455);
or U8698 (N_8698,N_8414,N_8504);
nor U8699 (N_8699,N_8415,N_8436);
and U8700 (N_8700,N_8618,N_8593);
and U8701 (N_8701,N_8594,N_8597);
xor U8702 (N_8702,N_8664,N_8604);
or U8703 (N_8703,N_8611,N_8631);
or U8704 (N_8704,N_8655,N_8670);
nor U8705 (N_8705,N_8698,N_8586);
and U8706 (N_8706,N_8651,N_8676);
nor U8707 (N_8707,N_8588,N_8689);
xor U8708 (N_8708,N_8691,N_8687);
xnor U8709 (N_8709,N_8603,N_8641);
xnor U8710 (N_8710,N_8553,N_8650);
nand U8711 (N_8711,N_8566,N_8645);
xnor U8712 (N_8712,N_8632,N_8551);
nand U8713 (N_8713,N_8666,N_8598);
and U8714 (N_8714,N_8591,N_8682);
and U8715 (N_8715,N_8679,N_8585);
or U8716 (N_8716,N_8596,N_8663);
nand U8717 (N_8717,N_8644,N_8690);
or U8718 (N_8718,N_8681,N_8621);
and U8719 (N_8719,N_8610,N_8667);
xor U8720 (N_8720,N_8619,N_8550);
nand U8721 (N_8721,N_8606,N_8646);
nor U8722 (N_8722,N_8638,N_8626);
and U8723 (N_8723,N_8614,N_8648);
nor U8724 (N_8724,N_8672,N_8570);
nand U8725 (N_8725,N_8674,N_8683);
nand U8726 (N_8726,N_8686,N_8581);
and U8727 (N_8727,N_8656,N_8624);
nand U8728 (N_8728,N_8565,N_8560);
xor U8729 (N_8729,N_8562,N_8564);
xnor U8730 (N_8730,N_8633,N_8639);
and U8731 (N_8731,N_8622,N_8643);
or U8732 (N_8732,N_8654,N_8612);
nand U8733 (N_8733,N_8625,N_8629);
or U8734 (N_8734,N_8579,N_8617);
nor U8735 (N_8735,N_8589,N_8595);
or U8736 (N_8736,N_8605,N_8561);
or U8737 (N_8737,N_8615,N_8573);
nor U8738 (N_8738,N_8559,N_8671);
xor U8739 (N_8739,N_8678,N_8652);
nor U8740 (N_8740,N_8574,N_8607);
and U8741 (N_8741,N_8693,N_8695);
nor U8742 (N_8742,N_8653,N_8554);
and U8743 (N_8743,N_8576,N_8568);
and U8744 (N_8744,N_8601,N_8657);
xor U8745 (N_8745,N_8685,N_8613);
or U8746 (N_8746,N_8584,N_8692);
and U8747 (N_8747,N_8602,N_8630);
and U8748 (N_8748,N_8600,N_8649);
or U8749 (N_8749,N_8571,N_8659);
xnor U8750 (N_8750,N_8577,N_8642);
and U8751 (N_8751,N_8694,N_8640);
nor U8752 (N_8752,N_8677,N_8662);
nor U8753 (N_8753,N_8658,N_8635);
or U8754 (N_8754,N_8699,N_8620);
nand U8755 (N_8755,N_8675,N_8563);
nor U8756 (N_8756,N_8575,N_8697);
or U8757 (N_8757,N_8647,N_8590);
xnor U8758 (N_8758,N_8616,N_8634);
and U8759 (N_8759,N_8578,N_8599);
nand U8760 (N_8760,N_8583,N_8661);
nor U8761 (N_8761,N_8609,N_8680);
nand U8762 (N_8762,N_8627,N_8592);
nor U8763 (N_8763,N_8557,N_8558);
nand U8764 (N_8764,N_8587,N_8623);
nor U8765 (N_8765,N_8665,N_8673);
and U8766 (N_8766,N_8660,N_8637);
xnor U8767 (N_8767,N_8556,N_8552);
and U8768 (N_8768,N_8608,N_8555);
and U8769 (N_8769,N_8668,N_8580);
and U8770 (N_8770,N_8572,N_8636);
or U8771 (N_8771,N_8569,N_8582);
nor U8772 (N_8772,N_8567,N_8688);
xor U8773 (N_8773,N_8696,N_8669);
nand U8774 (N_8774,N_8628,N_8684);
and U8775 (N_8775,N_8594,N_8591);
and U8776 (N_8776,N_8654,N_8599);
nor U8777 (N_8777,N_8666,N_8665);
or U8778 (N_8778,N_8591,N_8593);
and U8779 (N_8779,N_8573,N_8634);
or U8780 (N_8780,N_8608,N_8697);
xor U8781 (N_8781,N_8600,N_8570);
nand U8782 (N_8782,N_8659,N_8561);
nand U8783 (N_8783,N_8600,N_8698);
xnor U8784 (N_8784,N_8698,N_8589);
xor U8785 (N_8785,N_8583,N_8656);
nand U8786 (N_8786,N_8597,N_8553);
xnor U8787 (N_8787,N_8564,N_8673);
nor U8788 (N_8788,N_8634,N_8598);
nor U8789 (N_8789,N_8644,N_8675);
nand U8790 (N_8790,N_8643,N_8645);
nor U8791 (N_8791,N_8569,N_8597);
nand U8792 (N_8792,N_8564,N_8666);
xnor U8793 (N_8793,N_8605,N_8691);
nor U8794 (N_8794,N_8672,N_8580);
and U8795 (N_8795,N_8617,N_8662);
xnor U8796 (N_8796,N_8560,N_8695);
nand U8797 (N_8797,N_8566,N_8629);
and U8798 (N_8798,N_8676,N_8678);
xor U8799 (N_8799,N_8694,N_8664);
xnor U8800 (N_8800,N_8672,N_8640);
nand U8801 (N_8801,N_8664,N_8591);
nor U8802 (N_8802,N_8698,N_8654);
and U8803 (N_8803,N_8557,N_8669);
nand U8804 (N_8804,N_8653,N_8652);
xnor U8805 (N_8805,N_8627,N_8552);
or U8806 (N_8806,N_8597,N_8618);
nand U8807 (N_8807,N_8656,N_8648);
nor U8808 (N_8808,N_8663,N_8680);
nand U8809 (N_8809,N_8592,N_8589);
nor U8810 (N_8810,N_8657,N_8554);
nor U8811 (N_8811,N_8650,N_8638);
nor U8812 (N_8812,N_8624,N_8579);
xnor U8813 (N_8813,N_8559,N_8697);
or U8814 (N_8814,N_8641,N_8555);
or U8815 (N_8815,N_8595,N_8558);
or U8816 (N_8816,N_8576,N_8614);
and U8817 (N_8817,N_8554,N_8678);
nor U8818 (N_8818,N_8562,N_8637);
nor U8819 (N_8819,N_8553,N_8667);
or U8820 (N_8820,N_8559,N_8614);
xor U8821 (N_8821,N_8598,N_8695);
xnor U8822 (N_8822,N_8631,N_8641);
and U8823 (N_8823,N_8599,N_8684);
nand U8824 (N_8824,N_8681,N_8645);
nor U8825 (N_8825,N_8670,N_8628);
nand U8826 (N_8826,N_8605,N_8593);
or U8827 (N_8827,N_8571,N_8698);
nor U8828 (N_8828,N_8690,N_8638);
nand U8829 (N_8829,N_8688,N_8649);
or U8830 (N_8830,N_8695,N_8573);
xnor U8831 (N_8831,N_8555,N_8582);
or U8832 (N_8832,N_8589,N_8682);
xnor U8833 (N_8833,N_8635,N_8683);
nor U8834 (N_8834,N_8676,N_8566);
and U8835 (N_8835,N_8650,N_8577);
nand U8836 (N_8836,N_8579,N_8557);
and U8837 (N_8837,N_8626,N_8631);
or U8838 (N_8838,N_8646,N_8567);
nor U8839 (N_8839,N_8562,N_8596);
xnor U8840 (N_8840,N_8682,N_8592);
nor U8841 (N_8841,N_8609,N_8574);
xor U8842 (N_8842,N_8597,N_8599);
nor U8843 (N_8843,N_8636,N_8623);
and U8844 (N_8844,N_8652,N_8613);
or U8845 (N_8845,N_8698,N_8603);
or U8846 (N_8846,N_8684,N_8568);
and U8847 (N_8847,N_8674,N_8668);
xnor U8848 (N_8848,N_8654,N_8601);
or U8849 (N_8849,N_8650,N_8580);
and U8850 (N_8850,N_8723,N_8747);
or U8851 (N_8851,N_8818,N_8835);
xnor U8852 (N_8852,N_8791,N_8736);
nand U8853 (N_8853,N_8762,N_8756);
and U8854 (N_8854,N_8705,N_8729);
xnor U8855 (N_8855,N_8721,N_8734);
xnor U8856 (N_8856,N_8772,N_8733);
and U8857 (N_8857,N_8821,N_8775);
nand U8858 (N_8858,N_8797,N_8789);
nand U8859 (N_8859,N_8710,N_8776);
nand U8860 (N_8860,N_8842,N_8809);
xnor U8861 (N_8861,N_8819,N_8716);
or U8862 (N_8862,N_8711,N_8726);
or U8863 (N_8863,N_8731,N_8754);
nand U8864 (N_8864,N_8714,N_8781);
and U8865 (N_8865,N_8829,N_8800);
or U8866 (N_8866,N_8758,N_8771);
or U8867 (N_8867,N_8783,N_8832);
nand U8868 (N_8868,N_8828,N_8815);
and U8869 (N_8869,N_8796,N_8798);
or U8870 (N_8870,N_8814,N_8816);
and U8871 (N_8871,N_8724,N_8746);
nand U8872 (N_8872,N_8703,N_8712);
nor U8873 (N_8873,N_8786,N_8744);
xnor U8874 (N_8874,N_8806,N_8836);
xor U8875 (N_8875,N_8763,N_8840);
nor U8876 (N_8876,N_8745,N_8825);
nor U8877 (N_8877,N_8849,N_8838);
nand U8878 (N_8878,N_8777,N_8755);
nor U8879 (N_8879,N_8837,N_8715);
nor U8880 (N_8880,N_8782,N_8811);
xnor U8881 (N_8881,N_8707,N_8769);
nor U8882 (N_8882,N_8741,N_8831);
nor U8883 (N_8883,N_8847,N_8784);
and U8884 (N_8884,N_8764,N_8752);
xnor U8885 (N_8885,N_8846,N_8848);
and U8886 (N_8886,N_8702,N_8804);
nor U8887 (N_8887,N_8767,N_8761);
or U8888 (N_8888,N_8802,N_8748);
nor U8889 (N_8889,N_8719,N_8817);
nand U8890 (N_8890,N_8704,N_8795);
or U8891 (N_8891,N_8737,N_8740);
xnor U8892 (N_8892,N_8725,N_8830);
and U8893 (N_8893,N_8822,N_8751);
xor U8894 (N_8894,N_8768,N_8774);
nor U8895 (N_8895,N_8827,N_8738);
xor U8896 (N_8896,N_8728,N_8735);
or U8897 (N_8897,N_8765,N_8720);
nor U8898 (N_8898,N_8730,N_8760);
xnor U8899 (N_8899,N_8808,N_8779);
nor U8900 (N_8900,N_8845,N_8844);
or U8901 (N_8901,N_8732,N_8757);
and U8902 (N_8902,N_8801,N_8820);
xor U8903 (N_8903,N_8807,N_8833);
nor U8904 (N_8904,N_8722,N_8803);
or U8905 (N_8905,N_8799,N_8790);
nand U8906 (N_8906,N_8787,N_8701);
xnor U8907 (N_8907,N_8700,N_8713);
and U8908 (N_8908,N_8834,N_8823);
nand U8909 (N_8909,N_8785,N_8709);
nor U8910 (N_8910,N_8718,N_8826);
nor U8911 (N_8911,N_8742,N_8843);
or U8912 (N_8912,N_8727,N_8739);
or U8913 (N_8913,N_8766,N_8749);
and U8914 (N_8914,N_8810,N_8717);
or U8915 (N_8915,N_8773,N_8794);
nor U8916 (N_8916,N_8759,N_8706);
xor U8917 (N_8917,N_8805,N_8770);
xor U8918 (N_8918,N_8743,N_8788);
nor U8919 (N_8919,N_8812,N_8708);
nor U8920 (N_8920,N_8839,N_8753);
and U8921 (N_8921,N_8793,N_8824);
xnor U8922 (N_8922,N_8841,N_8780);
nand U8923 (N_8923,N_8778,N_8792);
xnor U8924 (N_8924,N_8813,N_8750);
nand U8925 (N_8925,N_8734,N_8742);
nand U8926 (N_8926,N_8791,N_8772);
nor U8927 (N_8927,N_8751,N_8702);
nor U8928 (N_8928,N_8733,N_8845);
nor U8929 (N_8929,N_8768,N_8754);
nor U8930 (N_8930,N_8795,N_8833);
or U8931 (N_8931,N_8729,N_8780);
or U8932 (N_8932,N_8746,N_8714);
xnor U8933 (N_8933,N_8761,N_8705);
or U8934 (N_8934,N_8704,N_8703);
or U8935 (N_8935,N_8767,N_8720);
and U8936 (N_8936,N_8776,N_8844);
nor U8937 (N_8937,N_8719,N_8815);
nand U8938 (N_8938,N_8841,N_8712);
nand U8939 (N_8939,N_8824,N_8750);
or U8940 (N_8940,N_8759,N_8790);
xor U8941 (N_8941,N_8773,N_8822);
nand U8942 (N_8942,N_8751,N_8739);
nand U8943 (N_8943,N_8728,N_8736);
and U8944 (N_8944,N_8809,N_8794);
xnor U8945 (N_8945,N_8828,N_8789);
nor U8946 (N_8946,N_8702,N_8781);
nand U8947 (N_8947,N_8724,N_8785);
nand U8948 (N_8948,N_8703,N_8846);
and U8949 (N_8949,N_8729,N_8700);
nor U8950 (N_8950,N_8768,N_8837);
nand U8951 (N_8951,N_8720,N_8756);
nand U8952 (N_8952,N_8815,N_8809);
xnor U8953 (N_8953,N_8835,N_8720);
nand U8954 (N_8954,N_8814,N_8818);
nand U8955 (N_8955,N_8709,N_8727);
nor U8956 (N_8956,N_8774,N_8716);
and U8957 (N_8957,N_8723,N_8704);
and U8958 (N_8958,N_8788,N_8717);
nand U8959 (N_8959,N_8762,N_8836);
and U8960 (N_8960,N_8708,N_8821);
or U8961 (N_8961,N_8824,N_8762);
xor U8962 (N_8962,N_8749,N_8821);
xor U8963 (N_8963,N_8755,N_8742);
xor U8964 (N_8964,N_8760,N_8741);
nand U8965 (N_8965,N_8813,N_8752);
nand U8966 (N_8966,N_8808,N_8743);
nor U8967 (N_8967,N_8715,N_8732);
nand U8968 (N_8968,N_8718,N_8709);
nand U8969 (N_8969,N_8788,N_8752);
xor U8970 (N_8970,N_8840,N_8847);
or U8971 (N_8971,N_8704,N_8823);
nor U8972 (N_8972,N_8835,N_8797);
xor U8973 (N_8973,N_8775,N_8782);
and U8974 (N_8974,N_8739,N_8769);
nor U8975 (N_8975,N_8812,N_8803);
or U8976 (N_8976,N_8829,N_8823);
and U8977 (N_8977,N_8825,N_8801);
xnor U8978 (N_8978,N_8761,N_8759);
nand U8979 (N_8979,N_8704,N_8759);
or U8980 (N_8980,N_8787,N_8774);
and U8981 (N_8981,N_8761,N_8824);
or U8982 (N_8982,N_8762,N_8734);
nor U8983 (N_8983,N_8739,N_8741);
xor U8984 (N_8984,N_8740,N_8799);
nand U8985 (N_8985,N_8731,N_8730);
nor U8986 (N_8986,N_8738,N_8739);
or U8987 (N_8987,N_8826,N_8723);
xor U8988 (N_8988,N_8707,N_8761);
or U8989 (N_8989,N_8734,N_8727);
xor U8990 (N_8990,N_8774,N_8756);
and U8991 (N_8991,N_8752,N_8767);
or U8992 (N_8992,N_8782,N_8746);
and U8993 (N_8993,N_8736,N_8780);
nand U8994 (N_8994,N_8799,N_8834);
and U8995 (N_8995,N_8736,N_8726);
nand U8996 (N_8996,N_8747,N_8833);
nand U8997 (N_8997,N_8757,N_8767);
or U8998 (N_8998,N_8761,N_8828);
nand U8999 (N_8999,N_8829,N_8848);
nor U9000 (N_9000,N_8995,N_8896);
nor U9001 (N_9001,N_8994,N_8874);
or U9002 (N_9002,N_8993,N_8938);
nor U9003 (N_9003,N_8922,N_8986);
xor U9004 (N_9004,N_8870,N_8886);
nand U9005 (N_9005,N_8982,N_8970);
nor U9006 (N_9006,N_8991,N_8876);
and U9007 (N_9007,N_8914,N_8998);
or U9008 (N_9008,N_8887,N_8900);
or U9009 (N_9009,N_8908,N_8983);
or U9010 (N_9010,N_8906,N_8942);
and U9011 (N_9011,N_8909,N_8917);
or U9012 (N_9012,N_8944,N_8890);
xor U9013 (N_9013,N_8984,N_8954);
nor U9014 (N_9014,N_8903,N_8877);
or U9015 (N_9015,N_8901,N_8902);
and U9016 (N_9016,N_8962,N_8948);
nand U9017 (N_9017,N_8885,N_8958);
xor U9018 (N_9018,N_8881,N_8920);
nor U9019 (N_9019,N_8976,N_8980);
nor U9020 (N_9020,N_8977,N_8872);
nand U9021 (N_9021,N_8892,N_8963);
and U9022 (N_9022,N_8936,N_8852);
nand U9023 (N_9023,N_8947,N_8974);
or U9024 (N_9024,N_8987,N_8926);
nor U9025 (N_9025,N_8981,N_8882);
and U9026 (N_9026,N_8919,N_8918);
and U9027 (N_9027,N_8952,N_8941);
xor U9028 (N_9028,N_8992,N_8990);
and U9029 (N_9029,N_8973,N_8854);
or U9030 (N_9030,N_8862,N_8940);
xnor U9031 (N_9031,N_8939,N_8866);
nand U9032 (N_9032,N_8873,N_8979);
xnor U9033 (N_9033,N_8921,N_8907);
nor U9034 (N_9034,N_8949,N_8931);
nor U9035 (N_9035,N_8916,N_8988);
nor U9036 (N_9036,N_8965,N_8996);
and U9037 (N_9037,N_8894,N_8899);
or U9038 (N_9038,N_8878,N_8972);
and U9039 (N_9039,N_8868,N_8880);
nand U9040 (N_9040,N_8967,N_8932);
or U9041 (N_9041,N_8997,N_8957);
nand U9042 (N_9042,N_8863,N_8966);
or U9043 (N_9043,N_8859,N_8905);
xor U9044 (N_9044,N_8884,N_8961);
nor U9045 (N_9045,N_8937,N_8860);
or U9046 (N_9046,N_8985,N_8891);
nor U9047 (N_9047,N_8889,N_8867);
and U9048 (N_9048,N_8865,N_8913);
nand U9049 (N_9049,N_8915,N_8893);
or U9050 (N_9050,N_8910,N_8950);
or U9051 (N_9051,N_8969,N_8898);
nor U9052 (N_9052,N_8929,N_8968);
nor U9053 (N_9053,N_8856,N_8895);
xor U9054 (N_9054,N_8951,N_8904);
xnor U9055 (N_9055,N_8924,N_8959);
or U9056 (N_9056,N_8999,N_8912);
xnor U9057 (N_9057,N_8897,N_8955);
nor U9058 (N_9058,N_8911,N_8869);
and U9059 (N_9059,N_8875,N_8851);
nor U9060 (N_9060,N_8857,N_8888);
xor U9061 (N_9061,N_8975,N_8883);
nor U9062 (N_9062,N_8850,N_8933);
xor U9063 (N_9063,N_8923,N_8989);
nor U9064 (N_9064,N_8855,N_8858);
nand U9065 (N_9065,N_8946,N_8953);
and U9066 (N_9066,N_8928,N_8964);
nor U9067 (N_9067,N_8861,N_8927);
nor U9068 (N_9068,N_8978,N_8943);
nor U9069 (N_9069,N_8853,N_8960);
nor U9070 (N_9070,N_8930,N_8934);
and U9071 (N_9071,N_8935,N_8925);
or U9072 (N_9072,N_8945,N_8864);
and U9073 (N_9073,N_8871,N_8956);
nand U9074 (N_9074,N_8971,N_8879);
nor U9075 (N_9075,N_8867,N_8862);
or U9076 (N_9076,N_8868,N_8917);
and U9077 (N_9077,N_8864,N_8870);
nand U9078 (N_9078,N_8895,N_8986);
nand U9079 (N_9079,N_8863,N_8876);
xor U9080 (N_9080,N_8874,N_8993);
nor U9081 (N_9081,N_8958,N_8859);
nor U9082 (N_9082,N_8967,N_8991);
nor U9083 (N_9083,N_8875,N_8951);
or U9084 (N_9084,N_8963,N_8855);
and U9085 (N_9085,N_8930,N_8971);
nand U9086 (N_9086,N_8959,N_8994);
and U9087 (N_9087,N_8913,N_8946);
nand U9088 (N_9088,N_8951,N_8978);
and U9089 (N_9089,N_8902,N_8893);
nand U9090 (N_9090,N_8887,N_8894);
nor U9091 (N_9091,N_8960,N_8868);
nor U9092 (N_9092,N_8890,N_8873);
nand U9093 (N_9093,N_8954,N_8993);
nand U9094 (N_9094,N_8897,N_8937);
or U9095 (N_9095,N_8925,N_8977);
xnor U9096 (N_9096,N_8866,N_8888);
and U9097 (N_9097,N_8853,N_8980);
xor U9098 (N_9098,N_8907,N_8893);
nand U9099 (N_9099,N_8929,N_8976);
xnor U9100 (N_9100,N_8939,N_8990);
xnor U9101 (N_9101,N_8989,N_8913);
and U9102 (N_9102,N_8949,N_8963);
nand U9103 (N_9103,N_8873,N_8961);
or U9104 (N_9104,N_8862,N_8864);
nor U9105 (N_9105,N_8854,N_8992);
xor U9106 (N_9106,N_8959,N_8867);
and U9107 (N_9107,N_8889,N_8969);
and U9108 (N_9108,N_8879,N_8947);
xnor U9109 (N_9109,N_8863,N_8888);
nand U9110 (N_9110,N_8983,N_8947);
xor U9111 (N_9111,N_8927,N_8857);
nor U9112 (N_9112,N_8870,N_8975);
nor U9113 (N_9113,N_8965,N_8927);
and U9114 (N_9114,N_8945,N_8858);
nor U9115 (N_9115,N_8941,N_8994);
or U9116 (N_9116,N_8850,N_8944);
or U9117 (N_9117,N_8941,N_8871);
nor U9118 (N_9118,N_8930,N_8998);
and U9119 (N_9119,N_8889,N_8927);
nand U9120 (N_9120,N_8923,N_8931);
nor U9121 (N_9121,N_8885,N_8902);
xnor U9122 (N_9122,N_8850,N_8967);
or U9123 (N_9123,N_8851,N_8932);
and U9124 (N_9124,N_8865,N_8877);
nand U9125 (N_9125,N_8962,N_8998);
or U9126 (N_9126,N_8973,N_8865);
nand U9127 (N_9127,N_8910,N_8907);
or U9128 (N_9128,N_8887,N_8972);
xor U9129 (N_9129,N_8856,N_8987);
nand U9130 (N_9130,N_8898,N_8880);
xnor U9131 (N_9131,N_8977,N_8986);
nand U9132 (N_9132,N_8922,N_8992);
nand U9133 (N_9133,N_8955,N_8970);
nand U9134 (N_9134,N_8959,N_8904);
nand U9135 (N_9135,N_8860,N_8904);
nand U9136 (N_9136,N_8925,N_8862);
or U9137 (N_9137,N_8948,N_8865);
or U9138 (N_9138,N_8949,N_8899);
or U9139 (N_9139,N_8875,N_8960);
or U9140 (N_9140,N_8907,N_8996);
nor U9141 (N_9141,N_8928,N_8950);
xor U9142 (N_9142,N_8949,N_8862);
and U9143 (N_9143,N_8903,N_8991);
or U9144 (N_9144,N_8939,N_8931);
xnor U9145 (N_9145,N_8869,N_8915);
xor U9146 (N_9146,N_8964,N_8969);
and U9147 (N_9147,N_8852,N_8911);
or U9148 (N_9148,N_8857,N_8859);
and U9149 (N_9149,N_8871,N_8915);
and U9150 (N_9150,N_9136,N_9138);
nor U9151 (N_9151,N_9139,N_9149);
or U9152 (N_9152,N_9009,N_9028);
nor U9153 (N_9153,N_9104,N_9075);
nor U9154 (N_9154,N_9089,N_9120);
or U9155 (N_9155,N_9010,N_9035);
or U9156 (N_9156,N_9116,N_9088);
nand U9157 (N_9157,N_9025,N_9077);
xor U9158 (N_9158,N_9023,N_9118);
nor U9159 (N_9159,N_9141,N_9100);
nand U9160 (N_9160,N_9004,N_9061);
nand U9161 (N_9161,N_9115,N_9081);
or U9162 (N_9162,N_9091,N_9132);
nor U9163 (N_9163,N_9016,N_9073);
xnor U9164 (N_9164,N_9027,N_9003);
nand U9165 (N_9165,N_9031,N_9064);
nor U9166 (N_9166,N_9033,N_9040);
xnor U9167 (N_9167,N_9058,N_9057);
and U9168 (N_9168,N_9026,N_9076);
nand U9169 (N_9169,N_9008,N_9092);
or U9170 (N_9170,N_9067,N_9130);
and U9171 (N_9171,N_9012,N_9127);
nor U9172 (N_9172,N_9110,N_9085);
or U9173 (N_9173,N_9071,N_9046);
nor U9174 (N_9174,N_9122,N_9093);
or U9175 (N_9175,N_9063,N_9123);
and U9176 (N_9176,N_9108,N_9137);
nor U9177 (N_9177,N_9011,N_9021);
nor U9178 (N_9178,N_9129,N_9090);
or U9179 (N_9179,N_9074,N_9142);
nor U9180 (N_9180,N_9128,N_9000);
nor U9181 (N_9181,N_9102,N_9119);
nand U9182 (N_9182,N_9062,N_9133);
and U9183 (N_9183,N_9015,N_9148);
nand U9184 (N_9184,N_9017,N_9041);
xnor U9185 (N_9185,N_9019,N_9106);
or U9186 (N_9186,N_9047,N_9079);
or U9187 (N_9187,N_9042,N_9134);
nand U9188 (N_9188,N_9098,N_9094);
nor U9189 (N_9189,N_9069,N_9014);
nor U9190 (N_9190,N_9029,N_9053);
or U9191 (N_9191,N_9070,N_9007);
nor U9192 (N_9192,N_9036,N_9051);
or U9193 (N_9193,N_9101,N_9131);
nand U9194 (N_9194,N_9140,N_9005);
xnor U9195 (N_9195,N_9066,N_9013);
nor U9196 (N_9196,N_9114,N_9099);
and U9197 (N_9197,N_9049,N_9111);
xor U9198 (N_9198,N_9048,N_9146);
and U9199 (N_9199,N_9113,N_9045);
xnor U9200 (N_9200,N_9037,N_9126);
or U9201 (N_9201,N_9044,N_9050);
and U9202 (N_9202,N_9022,N_9043);
or U9203 (N_9203,N_9034,N_9068);
or U9204 (N_9204,N_9087,N_9065);
nor U9205 (N_9205,N_9147,N_9055);
or U9206 (N_9206,N_9084,N_9060);
and U9207 (N_9207,N_9002,N_9145);
nand U9208 (N_9208,N_9006,N_9054);
xor U9209 (N_9209,N_9082,N_9018);
nor U9210 (N_9210,N_9096,N_9038);
and U9211 (N_9211,N_9086,N_9143);
nand U9212 (N_9212,N_9105,N_9135);
nor U9213 (N_9213,N_9097,N_9109);
nor U9214 (N_9214,N_9107,N_9052);
and U9215 (N_9215,N_9103,N_9112);
and U9216 (N_9216,N_9032,N_9039);
nor U9217 (N_9217,N_9072,N_9024);
nor U9218 (N_9218,N_9020,N_9078);
and U9219 (N_9219,N_9124,N_9030);
nor U9220 (N_9220,N_9095,N_9125);
and U9221 (N_9221,N_9001,N_9117);
nor U9222 (N_9222,N_9144,N_9080);
nand U9223 (N_9223,N_9059,N_9083);
nand U9224 (N_9224,N_9056,N_9121);
xor U9225 (N_9225,N_9000,N_9025);
or U9226 (N_9226,N_9100,N_9136);
nor U9227 (N_9227,N_9146,N_9036);
nor U9228 (N_9228,N_9019,N_9057);
nor U9229 (N_9229,N_9103,N_9119);
nand U9230 (N_9230,N_9073,N_9144);
or U9231 (N_9231,N_9045,N_9103);
nor U9232 (N_9232,N_9001,N_9092);
nand U9233 (N_9233,N_9027,N_9024);
xor U9234 (N_9234,N_9026,N_9075);
xnor U9235 (N_9235,N_9145,N_9012);
nor U9236 (N_9236,N_9014,N_9056);
and U9237 (N_9237,N_9112,N_9077);
nand U9238 (N_9238,N_9072,N_9096);
xor U9239 (N_9239,N_9128,N_9013);
xor U9240 (N_9240,N_9066,N_9109);
and U9241 (N_9241,N_9019,N_9028);
nor U9242 (N_9242,N_9138,N_9094);
xor U9243 (N_9243,N_9087,N_9081);
or U9244 (N_9244,N_9129,N_9084);
xor U9245 (N_9245,N_9125,N_9136);
or U9246 (N_9246,N_9066,N_9009);
nor U9247 (N_9247,N_9057,N_9121);
nand U9248 (N_9248,N_9015,N_9033);
xnor U9249 (N_9249,N_9021,N_9084);
nor U9250 (N_9250,N_9048,N_9035);
xnor U9251 (N_9251,N_9089,N_9041);
nand U9252 (N_9252,N_9070,N_9140);
xor U9253 (N_9253,N_9115,N_9076);
nor U9254 (N_9254,N_9141,N_9098);
nor U9255 (N_9255,N_9117,N_9109);
nor U9256 (N_9256,N_9030,N_9135);
nor U9257 (N_9257,N_9139,N_9102);
xor U9258 (N_9258,N_9147,N_9037);
nand U9259 (N_9259,N_9063,N_9145);
xnor U9260 (N_9260,N_9004,N_9047);
xnor U9261 (N_9261,N_9132,N_9137);
or U9262 (N_9262,N_9016,N_9007);
or U9263 (N_9263,N_9040,N_9129);
nand U9264 (N_9264,N_9022,N_9054);
xnor U9265 (N_9265,N_9127,N_9033);
xor U9266 (N_9266,N_9123,N_9079);
xor U9267 (N_9267,N_9018,N_9144);
and U9268 (N_9268,N_9036,N_9099);
or U9269 (N_9269,N_9003,N_9026);
nor U9270 (N_9270,N_9125,N_9003);
nor U9271 (N_9271,N_9113,N_9035);
or U9272 (N_9272,N_9086,N_9041);
nor U9273 (N_9273,N_9135,N_9100);
xor U9274 (N_9274,N_9055,N_9142);
xnor U9275 (N_9275,N_9102,N_9096);
or U9276 (N_9276,N_9025,N_9103);
nand U9277 (N_9277,N_9036,N_9147);
xor U9278 (N_9278,N_9105,N_9094);
nand U9279 (N_9279,N_9147,N_9045);
nand U9280 (N_9280,N_9044,N_9032);
nor U9281 (N_9281,N_9099,N_9041);
nand U9282 (N_9282,N_9079,N_9119);
nand U9283 (N_9283,N_9033,N_9004);
nand U9284 (N_9284,N_9039,N_9111);
xor U9285 (N_9285,N_9132,N_9001);
nand U9286 (N_9286,N_9002,N_9103);
nor U9287 (N_9287,N_9103,N_9048);
and U9288 (N_9288,N_9002,N_9117);
xor U9289 (N_9289,N_9022,N_9012);
xnor U9290 (N_9290,N_9039,N_9036);
and U9291 (N_9291,N_9077,N_9114);
and U9292 (N_9292,N_9135,N_9122);
nand U9293 (N_9293,N_9117,N_9032);
or U9294 (N_9294,N_9119,N_9061);
xnor U9295 (N_9295,N_9064,N_9005);
xnor U9296 (N_9296,N_9089,N_9135);
or U9297 (N_9297,N_9097,N_9075);
nor U9298 (N_9298,N_9060,N_9091);
nand U9299 (N_9299,N_9036,N_9101);
nand U9300 (N_9300,N_9152,N_9247);
or U9301 (N_9301,N_9157,N_9256);
nor U9302 (N_9302,N_9243,N_9246);
and U9303 (N_9303,N_9264,N_9262);
nand U9304 (N_9304,N_9297,N_9227);
xnor U9305 (N_9305,N_9188,N_9191);
or U9306 (N_9306,N_9223,N_9274);
and U9307 (N_9307,N_9289,N_9212);
and U9308 (N_9308,N_9280,N_9174);
nand U9309 (N_9309,N_9200,N_9202);
and U9310 (N_9310,N_9275,N_9203);
or U9311 (N_9311,N_9167,N_9238);
and U9312 (N_9312,N_9261,N_9279);
nor U9313 (N_9313,N_9184,N_9164);
and U9314 (N_9314,N_9160,N_9150);
nand U9315 (N_9315,N_9194,N_9286);
or U9316 (N_9316,N_9296,N_9232);
and U9317 (N_9317,N_9187,N_9178);
nor U9318 (N_9318,N_9193,N_9166);
and U9319 (N_9319,N_9176,N_9198);
and U9320 (N_9320,N_9171,N_9213);
or U9321 (N_9321,N_9165,N_9293);
nor U9322 (N_9322,N_9158,N_9295);
nor U9323 (N_9323,N_9237,N_9162);
nor U9324 (N_9324,N_9268,N_9151);
nand U9325 (N_9325,N_9281,N_9250);
xnor U9326 (N_9326,N_9248,N_9195);
nand U9327 (N_9327,N_9266,N_9251);
and U9328 (N_9328,N_9168,N_9244);
nand U9329 (N_9329,N_9245,N_9271);
nand U9330 (N_9330,N_9172,N_9221);
and U9331 (N_9331,N_9199,N_9185);
and U9332 (N_9332,N_9282,N_9263);
nor U9333 (N_9333,N_9241,N_9216);
xor U9334 (N_9334,N_9215,N_9240);
nand U9335 (N_9335,N_9291,N_9255);
or U9336 (N_9336,N_9299,N_9177);
and U9337 (N_9337,N_9163,N_9156);
and U9338 (N_9338,N_9235,N_9269);
xor U9339 (N_9339,N_9214,N_9205);
or U9340 (N_9340,N_9276,N_9153);
and U9341 (N_9341,N_9182,N_9225);
and U9342 (N_9342,N_9207,N_9239);
nand U9343 (N_9343,N_9169,N_9196);
xor U9344 (N_9344,N_9186,N_9224);
nor U9345 (N_9345,N_9277,N_9298);
xor U9346 (N_9346,N_9283,N_9220);
or U9347 (N_9347,N_9218,N_9222);
xor U9348 (N_9348,N_9287,N_9285);
xnor U9349 (N_9349,N_9267,N_9155);
xnor U9350 (N_9350,N_9272,N_9290);
and U9351 (N_9351,N_9292,N_9179);
or U9352 (N_9352,N_9159,N_9294);
and U9353 (N_9353,N_9217,N_9208);
nand U9354 (N_9354,N_9252,N_9228);
nand U9355 (N_9355,N_9180,N_9206);
xnor U9356 (N_9356,N_9183,N_9229);
xnor U9357 (N_9357,N_9209,N_9197);
xnor U9358 (N_9358,N_9249,N_9161);
xnor U9359 (N_9359,N_9259,N_9226);
xor U9360 (N_9360,N_9284,N_9242);
xor U9361 (N_9361,N_9204,N_9270);
nand U9362 (N_9362,N_9265,N_9170);
xor U9363 (N_9363,N_9233,N_9230);
nand U9364 (N_9364,N_9288,N_9254);
and U9365 (N_9365,N_9219,N_9192);
nor U9366 (N_9366,N_9201,N_9210);
or U9367 (N_9367,N_9211,N_9273);
and U9368 (N_9368,N_9190,N_9253);
and U9369 (N_9369,N_9175,N_9231);
or U9370 (N_9370,N_9236,N_9278);
and U9371 (N_9371,N_9260,N_9181);
xnor U9372 (N_9372,N_9234,N_9173);
or U9373 (N_9373,N_9154,N_9189);
xnor U9374 (N_9374,N_9258,N_9257);
and U9375 (N_9375,N_9255,N_9225);
nor U9376 (N_9376,N_9284,N_9173);
and U9377 (N_9377,N_9203,N_9174);
or U9378 (N_9378,N_9273,N_9252);
nand U9379 (N_9379,N_9163,N_9273);
nor U9380 (N_9380,N_9299,N_9272);
xnor U9381 (N_9381,N_9291,N_9285);
or U9382 (N_9382,N_9263,N_9156);
xnor U9383 (N_9383,N_9210,N_9156);
nand U9384 (N_9384,N_9233,N_9221);
or U9385 (N_9385,N_9288,N_9258);
nor U9386 (N_9386,N_9157,N_9229);
nand U9387 (N_9387,N_9160,N_9193);
and U9388 (N_9388,N_9216,N_9212);
nand U9389 (N_9389,N_9163,N_9255);
or U9390 (N_9390,N_9275,N_9201);
xnor U9391 (N_9391,N_9215,N_9288);
nor U9392 (N_9392,N_9160,N_9298);
and U9393 (N_9393,N_9297,N_9282);
xnor U9394 (N_9394,N_9188,N_9234);
and U9395 (N_9395,N_9193,N_9154);
and U9396 (N_9396,N_9193,N_9164);
xor U9397 (N_9397,N_9293,N_9262);
xor U9398 (N_9398,N_9230,N_9280);
nand U9399 (N_9399,N_9192,N_9198);
and U9400 (N_9400,N_9199,N_9245);
xor U9401 (N_9401,N_9187,N_9276);
and U9402 (N_9402,N_9220,N_9161);
xor U9403 (N_9403,N_9218,N_9163);
xnor U9404 (N_9404,N_9223,N_9259);
nor U9405 (N_9405,N_9220,N_9238);
xor U9406 (N_9406,N_9249,N_9209);
nand U9407 (N_9407,N_9239,N_9168);
and U9408 (N_9408,N_9237,N_9153);
or U9409 (N_9409,N_9258,N_9166);
xor U9410 (N_9410,N_9270,N_9245);
and U9411 (N_9411,N_9249,N_9247);
or U9412 (N_9412,N_9191,N_9279);
xnor U9413 (N_9413,N_9250,N_9251);
and U9414 (N_9414,N_9267,N_9274);
nor U9415 (N_9415,N_9277,N_9178);
nor U9416 (N_9416,N_9177,N_9211);
and U9417 (N_9417,N_9157,N_9176);
or U9418 (N_9418,N_9291,N_9288);
xnor U9419 (N_9419,N_9288,N_9185);
and U9420 (N_9420,N_9221,N_9150);
nand U9421 (N_9421,N_9291,N_9182);
or U9422 (N_9422,N_9239,N_9281);
and U9423 (N_9423,N_9213,N_9293);
xnor U9424 (N_9424,N_9281,N_9192);
or U9425 (N_9425,N_9171,N_9253);
xor U9426 (N_9426,N_9205,N_9257);
nor U9427 (N_9427,N_9217,N_9265);
and U9428 (N_9428,N_9251,N_9273);
nand U9429 (N_9429,N_9286,N_9281);
nand U9430 (N_9430,N_9159,N_9172);
nand U9431 (N_9431,N_9211,N_9155);
nand U9432 (N_9432,N_9246,N_9264);
nor U9433 (N_9433,N_9286,N_9213);
or U9434 (N_9434,N_9239,N_9278);
and U9435 (N_9435,N_9269,N_9193);
nor U9436 (N_9436,N_9254,N_9161);
nor U9437 (N_9437,N_9209,N_9236);
nand U9438 (N_9438,N_9286,N_9153);
xnor U9439 (N_9439,N_9173,N_9216);
or U9440 (N_9440,N_9196,N_9179);
xnor U9441 (N_9441,N_9200,N_9229);
or U9442 (N_9442,N_9176,N_9277);
or U9443 (N_9443,N_9215,N_9255);
xor U9444 (N_9444,N_9270,N_9165);
nand U9445 (N_9445,N_9238,N_9152);
or U9446 (N_9446,N_9209,N_9298);
nand U9447 (N_9447,N_9195,N_9265);
nor U9448 (N_9448,N_9299,N_9181);
xnor U9449 (N_9449,N_9150,N_9255);
nand U9450 (N_9450,N_9411,N_9385);
nor U9451 (N_9451,N_9422,N_9446);
or U9452 (N_9452,N_9316,N_9426);
nand U9453 (N_9453,N_9383,N_9374);
nand U9454 (N_9454,N_9364,N_9325);
nand U9455 (N_9455,N_9320,N_9376);
nor U9456 (N_9456,N_9363,N_9403);
and U9457 (N_9457,N_9351,N_9307);
and U9458 (N_9458,N_9342,N_9314);
or U9459 (N_9459,N_9408,N_9350);
nor U9460 (N_9460,N_9396,N_9410);
xor U9461 (N_9461,N_9402,N_9330);
xnor U9462 (N_9462,N_9423,N_9415);
xnor U9463 (N_9463,N_9317,N_9355);
and U9464 (N_9464,N_9348,N_9300);
xnor U9465 (N_9465,N_9334,N_9438);
or U9466 (N_9466,N_9302,N_9335);
and U9467 (N_9467,N_9333,N_9336);
nor U9468 (N_9468,N_9379,N_9310);
or U9469 (N_9469,N_9405,N_9323);
xor U9470 (N_9470,N_9417,N_9322);
nor U9471 (N_9471,N_9409,N_9381);
nand U9472 (N_9472,N_9394,N_9388);
nor U9473 (N_9473,N_9341,N_9354);
nand U9474 (N_9474,N_9436,N_9440);
xor U9475 (N_9475,N_9367,N_9435);
or U9476 (N_9476,N_9398,N_9352);
nand U9477 (N_9477,N_9311,N_9413);
or U9478 (N_9478,N_9445,N_9444);
nand U9479 (N_9479,N_9390,N_9395);
xor U9480 (N_9480,N_9419,N_9339);
xnor U9481 (N_9481,N_9368,N_9412);
nand U9482 (N_9482,N_9359,N_9329);
nor U9483 (N_9483,N_9305,N_9340);
xnor U9484 (N_9484,N_9344,N_9439);
and U9485 (N_9485,N_9433,N_9312);
nor U9486 (N_9486,N_9434,N_9373);
nand U9487 (N_9487,N_9369,N_9400);
nor U9488 (N_9488,N_9399,N_9432);
nor U9489 (N_9489,N_9331,N_9437);
nor U9490 (N_9490,N_9441,N_9308);
nor U9491 (N_9491,N_9382,N_9321);
nand U9492 (N_9492,N_9420,N_9380);
or U9493 (N_9493,N_9353,N_9361);
xor U9494 (N_9494,N_9377,N_9304);
or U9495 (N_9495,N_9356,N_9345);
xor U9496 (N_9496,N_9346,N_9332);
or U9497 (N_9497,N_9318,N_9407);
nor U9498 (N_9498,N_9391,N_9429);
nand U9499 (N_9499,N_9349,N_9428);
xor U9500 (N_9500,N_9418,N_9384);
nor U9501 (N_9501,N_9393,N_9371);
nor U9502 (N_9502,N_9313,N_9404);
xor U9503 (N_9503,N_9401,N_9372);
or U9504 (N_9504,N_9414,N_9328);
xor U9505 (N_9505,N_9424,N_9315);
or U9506 (N_9506,N_9324,N_9389);
nor U9507 (N_9507,N_9309,N_9362);
and U9508 (N_9508,N_9447,N_9406);
nand U9509 (N_9509,N_9326,N_9370);
and U9510 (N_9510,N_9449,N_9430);
xnor U9511 (N_9511,N_9425,N_9357);
xor U9512 (N_9512,N_9360,N_9303);
nor U9513 (N_9513,N_9378,N_9306);
or U9514 (N_9514,N_9397,N_9421);
nand U9515 (N_9515,N_9442,N_9319);
and U9516 (N_9516,N_9386,N_9431);
xnor U9517 (N_9517,N_9338,N_9448);
xor U9518 (N_9518,N_9392,N_9327);
and U9519 (N_9519,N_9347,N_9387);
or U9520 (N_9520,N_9343,N_9337);
and U9521 (N_9521,N_9427,N_9301);
or U9522 (N_9522,N_9358,N_9375);
nand U9523 (N_9523,N_9416,N_9443);
and U9524 (N_9524,N_9365,N_9366);
nor U9525 (N_9525,N_9448,N_9446);
and U9526 (N_9526,N_9424,N_9422);
nor U9527 (N_9527,N_9442,N_9374);
or U9528 (N_9528,N_9367,N_9408);
and U9529 (N_9529,N_9301,N_9358);
or U9530 (N_9530,N_9408,N_9418);
nor U9531 (N_9531,N_9342,N_9438);
and U9532 (N_9532,N_9369,N_9442);
and U9533 (N_9533,N_9372,N_9344);
nor U9534 (N_9534,N_9320,N_9421);
nand U9535 (N_9535,N_9318,N_9397);
xnor U9536 (N_9536,N_9389,N_9362);
or U9537 (N_9537,N_9394,N_9321);
nor U9538 (N_9538,N_9400,N_9444);
or U9539 (N_9539,N_9326,N_9338);
and U9540 (N_9540,N_9387,N_9335);
and U9541 (N_9541,N_9402,N_9368);
and U9542 (N_9542,N_9424,N_9381);
xnor U9543 (N_9543,N_9341,N_9417);
and U9544 (N_9544,N_9317,N_9342);
nor U9545 (N_9545,N_9405,N_9431);
and U9546 (N_9546,N_9401,N_9377);
xnor U9547 (N_9547,N_9359,N_9335);
nand U9548 (N_9548,N_9437,N_9371);
nor U9549 (N_9549,N_9343,N_9334);
xor U9550 (N_9550,N_9313,N_9336);
or U9551 (N_9551,N_9369,N_9301);
nand U9552 (N_9552,N_9420,N_9444);
nor U9553 (N_9553,N_9410,N_9397);
or U9554 (N_9554,N_9446,N_9379);
xor U9555 (N_9555,N_9447,N_9398);
or U9556 (N_9556,N_9337,N_9410);
and U9557 (N_9557,N_9363,N_9319);
nand U9558 (N_9558,N_9300,N_9377);
xor U9559 (N_9559,N_9390,N_9352);
or U9560 (N_9560,N_9334,N_9318);
and U9561 (N_9561,N_9399,N_9330);
or U9562 (N_9562,N_9449,N_9312);
or U9563 (N_9563,N_9374,N_9378);
or U9564 (N_9564,N_9348,N_9406);
xor U9565 (N_9565,N_9432,N_9349);
xor U9566 (N_9566,N_9429,N_9384);
xor U9567 (N_9567,N_9339,N_9390);
nor U9568 (N_9568,N_9436,N_9334);
xor U9569 (N_9569,N_9303,N_9331);
nor U9570 (N_9570,N_9398,N_9433);
nor U9571 (N_9571,N_9397,N_9377);
or U9572 (N_9572,N_9376,N_9381);
and U9573 (N_9573,N_9437,N_9319);
or U9574 (N_9574,N_9412,N_9394);
and U9575 (N_9575,N_9387,N_9436);
xor U9576 (N_9576,N_9368,N_9420);
nor U9577 (N_9577,N_9423,N_9361);
or U9578 (N_9578,N_9393,N_9304);
nand U9579 (N_9579,N_9408,N_9375);
xor U9580 (N_9580,N_9387,N_9351);
nor U9581 (N_9581,N_9305,N_9428);
nor U9582 (N_9582,N_9342,N_9413);
nor U9583 (N_9583,N_9389,N_9364);
nor U9584 (N_9584,N_9398,N_9386);
nand U9585 (N_9585,N_9338,N_9344);
xnor U9586 (N_9586,N_9410,N_9372);
xnor U9587 (N_9587,N_9339,N_9319);
or U9588 (N_9588,N_9324,N_9397);
xor U9589 (N_9589,N_9417,N_9345);
nand U9590 (N_9590,N_9337,N_9390);
or U9591 (N_9591,N_9407,N_9409);
or U9592 (N_9592,N_9447,N_9383);
xor U9593 (N_9593,N_9317,N_9387);
nor U9594 (N_9594,N_9404,N_9407);
nand U9595 (N_9595,N_9315,N_9356);
or U9596 (N_9596,N_9381,N_9322);
or U9597 (N_9597,N_9449,N_9406);
nor U9598 (N_9598,N_9342,N_9372);
or U9599 (N_9599,N_9416,N_9389);
nand U9600 (N_9600,N_9505,N_9529);
xnor U9601 (N_9601,N_9546,N_9582);
and U9602 (N_9602,N_9536,N_9491);
and U9603 (N_9603,N_9469,N_9595);
nand U9604 (N_9604,N_9538,N_9470);
or U9605 (N_9605,N_9526,N_9462);
nand U9606 (N_9606,N_9553,N_9527);
nand U9607 (N_9607,N_9555,N_9480);
xnor U9608 (N_9608,N_9569,N_9599);
xnor U9609 (N_9609,N_9572,N_9587);
nand U9610 (N_9610,N_9583,N_9509);
nand U9611 (N_9611,N_9537,N_9507);
nand U9612 (N_9612,N_9559,N_9460);
and U9613 (N_9613,N_9524,N_9567);
xnor U9614 (N_9614,N_9471,N_9459);
nor U9615 (N_9615,N_9482,N_9494);
nor U9616 (N_9616,N_9566,N_9520);
and U9617 (N_9617,N_9478,N_9543);
nand U9618 (N_9618,N_9458,N_9532);
and U9619 (N_9619,N_9535,N_9517);
and U9620 (N_9620,N_9514,N_9579);
nand U9621 (N_9621,N_9588,N_9544);
nor U9622 (N_9622,N_9521,N_9574);
and U9623 (N_9623,N_9522,N_9486);
xor U9624 (N_9624,N_9531,N_9493);
nand U9625 (N_9625,N_9558,N_9593);
and U9626 (N_9626,N_9584,N_9499);
nand U9627 (N_9627,N_9551,N_9561);
nand U9628 (N_9628,N_9475,N_9528);
nor U9629 (N_9629,N_9594,N_9590);
xnor U9630 (N_9630,N_9511,N_9563);
nor U9631 (N_9631,N_9541,N_9534);
nor U9632 (N_9632,N_9504,N_9464);
nor U9633 (N_9633,N_9473,N_9465);
nand U9634 (N_9634,N_9502,N_9503);
nor U9635 (N_9635,N_9508,N_9463);
and U9636 (N_9636,N_9455,N_9516);
nor U9637 (N_9637,N_9576,N_9523);
nor U9638 (N_9638,N_9530,N_9487);
xor U9639 (N_9639,N_9545,N_9560);
nand U9640 (N_9640,N_9498,N_9557);
nand U9641 (N_9641,N_9457,N_9581);
nand U9642 (N_9642,N_9492,N_9506);
and U9643 (N_9643,N_9512,N_9585);
nor U9644 (N_9644,N_9580,N_9454);
nand U9645 (N_9645,N_9515,N_9452);
nand U9646 (N_9646,N_9468,N_9483);
nor U9647 (N_9647,N_9496,N_9539);
xnor U9648 (N_9648,N_9476,N_9562);
xor U9649 (N_9649,N_9533,N_9525);
nand U9650 (N_9650,N_9573,N_9571);
nand U9651 (N_9651,N_9552,N_9461);
nand U9652 (N_9652,N_9518,N_9513);
nor U9653 (N_9653,N_9570,N_9497);
or U9654 (N_9654,N_9565,N_9564);
nor U9655 (N_9655,N_9597,N_9591);
and U9656 (N_9656,N_9501,N_9456);
nand U9657 (N_9657,N_9575,N_9488);
and U9658 (N_9658,N_9467,N_9548);
nand U9659 (N_9659,N_9540,N_9477);
nand U9660 (N_9660,N_9589,N_9484);
or U9661 (N_9661,N_9577,N_9481);
xor U9662 (N_9662,N_9450,N_9453);
and U9663 (N_9663,N_9556,N_9568);
or U9664 (N_9664,N_9479,N_9472);
nand U9665 (N_9665,N_9451,N_9474);
nand U9666 (N_9666,N_9490,N_9554);
nor U9667 (N_9667,N_9592,N_9500);
nand U9668 (N_9668,N_9598,N_9596);
and U9669 (N_9669,N_9578,N_9489);
or U9670 (N_9670,N_9495,N_9550);
or U9671 (N_9671,N_9542,N_9547);
and U9672 (N_9672,N_9510,N_9466);
and U9673 (N_9673,N_9549,N_9519);
or U9674 (N_9674,N_9586,N_9485);
xor U9675 (N_9675,N_9571,N_9585);
and U9676 (N_9676,N_9559,N_9505);
and U9677 (N_9677,N_9538,N_9493);
xnor U9678 (N_9678,N_9501,N_9516);
or U9679 (N_9679,N_9457,N_9560);
or U9680 (N_9680,N_9496,N_9521);
nor U9681 (N_9681,N_9535,N_9559);
xnor U9682 (N_9682,N_9479,N_9552);
and U9683 (N_9683,N_9516,N_9542);
nand U9684 (N_9684,N_9536,N_9518);
or U9685 (N_9685,N_9465,N_9554);
xnor U9686 (N_9686,N_9544,N_9562);
and U9687 (N_9687,N_9537,N_9498);
nor U9688 (N_9688,N_9494,N_9590);
or U9689 (N_9689,N_9509,N_9595);
xnor U9690 (N_9690,N_9496,N_9526);
nor U9691 (N_9691,N_9571,N_9549);
xnor U9692 (N_9692,N_9474,N_9463);
xnor U9693 (N_9693,N_9528,N_9540);
and U9694 (N_9694,N_9489,N_9501);
or U9695 (N_9695,N_9498,N_9542);
nor U9696 (N_9696,N_9461,N_9464);
and U9697 (N_9697,N_9461,N_9518);
xor U9698 (N_9698,N_9514,N_9586);
and U9699 (N_9699,N_9538,N_9500);
xnor U9700 (N_9700,N_9503,N_9572);
or U9701 (N_9701,N_9510,N_9491);
xnor U9702 (N_9702,N_9525,N_9599);
xnor U9703 (N_9703,N_9467,N_9577);
nor U9704 (N_9704,N_9480,N_9597);
or U9705 (N_9705,N_9558,N_9463);
nor U9706 (N_9706,N_9597,N_9574);
xor U9707 (N_9707,N_9512,N_9545);
or U9708 (N_9708,N_9496,N_9477);
xor U9709 (N_9709,N_9502,N_9477);
or U9710 (N_9710,N_9591,N_9484);
nor U9711 (N_9711,N_9498,N_9551);
and U9712 (N_9712,N_9471,N_9506);
xor U9713 (N_9713,N_9525,N_9472);
nor U9714 (N_9714,N_9541,N_9454);
nor U9715 (N_9715,N_9528,N_9465);
xor U9716 (N_9716,N_9466,N_9560);
nand U9717 (N_9717,N_9453,N_9465);
nor U9718 (N_9718,N_9535,N_9456);
xor U9719 (N_9719,N_9534,N_9586);
nand U9720 (N_9720,N_9474,N_9485);
nor U9721 (N_9721,N_9588,N_9463);
or U9722 (N_9722,N_9565,N_9557);
nor U9723 (N_9723,N_9559,N_9562);
or U9724 (N_9724,N_9550,N_9489);
and U9725 (N_9725,N_9567,N_9456);
nor U9726 (N_9726,N_9510,N_9473);
xnor U9727 (N_9727,N_9571,N_9472);
nand U9728 (N_9728,N_9463,N_9509);
nor U9729 (N_9729,N_9537,N_9492);
or U9730 (N_9730,N_9456,N_9474);
or U9731 (N_9731,N_9557,N_9553);
nand U9732 (N_9732,N_9527,N_9570);
nor U9733 (N_9733,N_9451,N_9542);
nand U9734 (N_9734,N_9559,N_9588);
or U9735 (N_9735,N_9552,N_9509);
or U9736 (N_9736,N_9529,N_9589);
xor U9737 (N_9737,N_9553,N_9582);
or U9738 (N_9738,N_9484,N_9531);
nand U9739 (N_9739,N_9566,N_9492);
nor U9740 (N_9740,N_9494,N_9541);
nor U9741 (N_9741,N_9550,N_9570);
nor U9742 (N_9742,N_9581,N_9589);
xor U9743 (N_9743,N_9461,N_9524);
nor U9744 (N_9744,N_9475,N_9533);
nor U9745 (N_9745,N_9594,N_9495);
or U9746 (N_9746,N_9580,N_9483);
and U9747 (N_9747,N_9484,N_9481);
nor U9748 (N_9748,N_9476,N_9521);
xor U9749 (N_9749,N_9510,N_9589);
nand U9750 (N_9750,N_9620,N_9608);
and U9751 (N_9751,N_9680,N_9616);
xnor U9752 (N_9752,N_9646,N_9627);
nand U9753 (N_9753,N_9610,N_9731);
and U9754 (N_9754,N_9701,N_9665);
and U9755 (N_9755,N_9699,N_9602);
or U9756 (N_9756,N_9619,N_9722);
and U9757 (N_9757,N_9723,N_9672);
nand U9758 (N_9758,N_9741,N_9661);
and U9759 (N_9759,N_9637,N_9670);
xnor U9760 (N_9760,N_9635,N_9651);
nor U9761 (N_9761,N_9694,N_9708);
xor U9762 (N_9762,N_9748,N_9682);
nand U9763 (N_9763,N_9609,N_9747);
or U9764 (N_9764,N_9638,N_9712);
xnor U9765 (N_9765,N_9705,N_9629);
nor U9766 (N_9766,N_9632,N_9621);
nor U9767 (N_9767,N_9691,N_9659);
xnor U9768 (N_9768,N_9710,N_9640);
or U9769 (N_9769,N_9744,N_9614);
and U9770 (N_9770,N_9606,N_9657);
nor U9771 (N_9771,N_9678,N_9633);
or U9772 (N_9772,N_9732,N_9667);
nor U9773 (N_9773,N_9643,N_9700);
nor U9774 (N_9774,N_9702,N_9668);
nor U9775 (N_9775,N_9607,N_9707);
or U9776 (N_9776,N_9730,N_9746);
and U9777 (N_9777,N_9656,N_9697);
nor U9778 (N_9778,N_9687,N_9726);
xor U9779 (N_9779,N_9634,N_9688);
xnor U9780 (N_9780,N_9721,N_9692);
nand U9781 (N_9781,N_9704,N_9683);
or U9782 (N_9782,N_9689,N_9745);
nor U9783 (N_9783,N_9729,N_9605);
and U9784 (N_9784,N_9662,N_9649);
and U9785 (N_9785,N_9639,N_9641);
nor U9786 (N_9786,N_9618,N_9671);
or U9787 (N_9787,N_9622,N_9615);
xnor U9788 (N_9788,N_9644,N_9600);
nor U9789 (N_9789,N_9626,N_9737);
xnor U9790 (N_9790,N_9717,N_9736);
xnor U9791 (N_9791,N_9716,N_9738);
nor U9792 (N_9792,N_9695,N_9718);
or U9793 (N_9793,N_9623,N_9735);
nor U9794 (N_9794,N_9673,N_9679);
xor U9795 (N_9795,N_9603,N_9681);
xnor U9796 (N_9796,N_9653,N_9719);
nor U9797 (N_9797,N_9674,N_9685);
or U9798 (N_9798,N_9636,N_9739);
or U9799 (N_9799,N_9728,N_9642);
or U9800 (N_9800,N_9714,N_9611);
nand U9801 (N_9801,N_9676,N_9630);
xor U9802 (N_9802,N_9650,N_9696);
nor U9803 (N_9803,N_9647,N_9742);
nor U9804 (N_9804,N_9743,N_9654);
nand U9805 (N_9805,N_9652,N_9727);
xnor U9806 (N_9806,N_9733,N_9604);
and U9807 (N_9807,N_9709,N_9711);
xor U9808 (N_9808,N_9724,N_9648);
nand U9809 (N_9809,N_9686,N_9690);
xnor U9810 (N_9810,N_9601,N_9658);
nor U9811 (N_9811,N_9706,N_9660);
nor U9812 (N_9812,N_9666,N_9725);
and U9813 (N_9813,N_9749,N_9655);
nand U9814 (N_9814,N_9645,N_9720);
or U9815 (N_9815,N_9612,N_9734);
nor U9816 (N_9816,N_9617,N_9713);
nor U9817 (N_9817,N_9628,N_9624);
nor U9818 (N_9818,N_9675,N_9677);
and U9819 (N_9819,N_9740,N_9703);
and U9820 (N_9820,N_9684,N_9631);
nor U9821 (N_9821,N_9693,N_9663);
and U9822 (N_9822,N_9625,N_9669);
nor U9823 (N_9823,N_9715,N_9698);
and U9824 (N_9824,N_9613,N_9664);
or U9825 (N_9825,N_9623,N_9745);
and U9826 (N_9826,N_9694,N_9727);
nor U9827 (N_9827,N_9706,N_9661);
and U9828 (N_9828,N_9727,N_9610);
xnor U9829 (N_9829,N_9705,N_9687);
nor U9830 (N_9830,N_9694,N_9650);
nor U9831 (N_9831,N_9725,N_9684);
nor U9832 (N_9832,N_9608,N_9606);
and U9833 (N_9833,N_9688,N_9723);
and U9834 (N_9834,N_9636,N_9736);
and U9835 (N_9835,N_9627,N_9658);
and U9836 (N_9836,N_9712,N_9636);
nand U9837 (N_9837,N_9642,N_9680);
and U9838 (N_9838,N_9745,N_9691);
or U9839 (N_9839,N_9680,N_9718);
xnor U9840 (N_9840,N_9696,N_9660);
nor U9841 (N_9841,N_9688,N_9616);
or U9842 (N_9842,N_9696,N_9604);
nand U9843 (N_9843,N_9623,N_9708);
or U9844 (N_9844,N_9679,N_9672);
or U9845 (N_9845,N_9738,N_9605);
or U9846 (N_9846,N_9730,N_9683);
or U9847 (N_9847,N_9621,N_9655);
nor U9848 (N_9848,N_9646,N_9702);
nor U9849 (N_9849,N_9626,N_9647);
or U9850 (N_9850,N_9689,N_9670);
nor U9851 (N_9851,N_9664,N_9655);
nor U9852 (N_9852,N_9606,N_9713);
nand U9853 (N_9853,N_9666,N_9693);
and U9854 (N_9854,N_9613,N_9697);
nand U9855 (N_9855,N_9747,N_9640);
or U9856 (N_9856,N_9608,N_9695);
or U9857 (N_9857,N_9638,N_9628);
nand U9858 (N_9858,N_9642,N_9681);
nor U9859 (N_9859,N_9746,N_9669);
or U9860 (N_9860,N_9678,N_9714);
xnor U9861 (N_9861,N_9703,N_9710);
xnor U9862 (N_9862,N_9624,N_9610);
nor U9863 (N_9863,N_9715,N_9663);
xor U9864 (N_9864,N_9661,N_9715);
and U9865 (N_9865,N_9662,N_9625);
xor U9866 (N_9866,N_9605,N_9611);
nor U9867 (N_9867,N_9611,N_9641);
or U9868 (N_9868,N_9739,N_9669);
nor U9869 (N_9869,N_9728,N_9739);
and U9870 (N_9870,N_9740,N_9712);
nor U9871 (N_9871,N_9614,N_9731);
and U9872 (N_9872,N_9744,N_9746);
xor U9873 (N_9873,N_9624,N_9728);
and U9874 (N_9874,N_9654,N_9644);
nor U9875 (N_9875,N_9743,N_9632);
nor U9876 (N_9876,N_9662,N_9644);
and U9877 (N_9877,N_9657,N_9663);
or U9878 (N_9878,N_9661,N_9659);
or U9879 (N_9879,N_9698,N_9650);
xor U9880 (N_9880,N_9744,N_9699);
nor U9881 (N_9881,N_9638,N_9650);
nand U9882 (N_9882,N_9674,N_9669);
nor U9883 (N_9883,N_9632,N_9684);
xor U9884 (N_9884,N_9624,N_9614);
nor U9885 (N_9885,N_9739,N_9646);
and U9886 (N_9886,N_9665,N_9654);
and U9887 (N_9887,N_9702,N_9658);
nand U9888 (N_9888,N_9650,N_9741);
or U9889 (N_9889,N_9621,N_9730);
and U9890 (N_9890,N_9701,N_9688);
xor U9891 (N_9891,N_9673,N_9680);
xnor U9892 (N_9892,N_9731,N_9734);
xnor U9893 (N_9893,N_9738,N_9626);
nor U9894 (N_9894,N_9619,N_9636);
xor U9895 (N_9895,N_9680,N_9742);
nand U9896 (N_9896,N_9643,N_9667);
xnor U9897 (N_9897,N_9626,N_9744);
or U9898 (N_9898,N_9715,N_9690);
and U9899 (N_9899,N_9613,N_9635);
nor U9900 (N_9900,N_9865,N_9894);
and U9901 (N_9901,N_9887,N_9843);
and U9902 (N_9902,N_9847,N_9837);
and U9903 (N_9903,N_9817,N_9803);
and U9904 (N_9904,N_9793,N_9758);
nand U9905 (N_9905,N_9759,N_9804);
nor U9906 (N_9906,N_9825,N_9845);
xor U9907 (N_9907,N_9770,N_9756);
nand U9908 (N_9908,N_9874,N_9812);
nand U9909 (N_9909,N_9879,N_9839);
xnor U9910 (N_9910,N_9762,N_9842);
nand U9911 (N_9911,N_9757,N_9884);
xor U9912 (N_9912,N_9811,N_9795);
nor U9913 (N_9913,N_9836,N_9790);
or U9914 (N_9914,N_9857,N_9750);
or U9915 (N_9915,N_9821,N_9877);
and U9916 (N_9916,N_9870,N_9818);
and U9917 (N_9917,N_9778,N_9773);
nand U9918 (N_9918,N_9855,N_9810);
nor U9919 (N_9919,N_9827,N_9791);
nor U9920 (N_9920,N_9813,N_9823);
and U9921 (N_9921,N_9890,N_9776);
nand U9922 (N_9922,N_9807,N_9786);
and U9923 (N_9923,N_9799,N_9832);
xnor U9924 (N_9924,N_9753,N_9826);
nand U9925 (N_9925,N_9888,N_9809);
nor U9926 (N_9926,N_9828,N_9882);
xor U9927 (N_9927,N_9858,N_9797);
and U9928 (N_9928,N_9783,N_9895);
nand U9929 (N_9929,N_9849,N_9841);
nand U9930 (N_9930,N_9768,N_9781);
or U9931 (N_9931,N_9796,N_9852);
nand U9932 (N_9932,N_9751,N_9835);
or U9933 (N_9933,N_9863,N_9801);
nor U9934 (N_9934,N_9830,N_9775);
and U9935 (N_9935,N_9856,N_9764);
xor U9936 (N_9936,N_9815,N_9864);
xor U9937 (N_9937,N_9785,N_9765);
or U9938 (N_9938,N_9871,N_9771);
xor U9939 (N_9939,N_9896,N_9754);
and U9940 (N_9940,N_9780,N_9760);
nor U9941 (N_9941,N_9875,N_9850);
xnor U9942 (N_9942,N_9885,N_9862);
nand U9943 (N_9943,N_9808,N_9868);
nor U9944 (N_9944,N_9766,N_9854);
nor U9945 (N_9945,N_9886,N_9769);
and U9946 (N_9946,N_9767,N_9831);
and U9947 (N_9947,N_9784,N_9824);
and U9948 (N_9948,N_9774,N_9800);
xnor U9949 (N_9949,N_9806,N_9789);
nand U9950 (N_9950,N_9820,N_9866);
xnor U9951 (N_9951,N_9840,N_9763);
nor U9952 (N_9952,N_9805,N_9892);
xor U9953 (N_9953,N_9891,N_9819);
and U9954 (N_9954,N_9844,N_9893);
nor U9955 (N_9955,N_9802,N_9873);
nand U9956 (N_9956,N_9867,N_9859);
and U9957 (N_9957,N_9883,N_9829);
xor U9958 (N_9958,N_9772,N_9782);
or U9959 (N_9959,N_9787,N_9869);
and U9960 (N_9960,N_9897,N_9833);
xor U9961 (N_9961,N_9794,N_9853);
nor U9962 (N_9962,N_9814,N_9834);
xor U9963 (N_9963,N_9848,N_9822);
nor U9964 (N_9964,N_9876,N_9777);
xor U9965 (N_9965,N_9846,N_9872);
nand U9966 (N_9966,N_9899,N_9878);
xnor U9967 (N_9967,N_9779,N_9755);
and U9968 (N_9968,N_9816,N_9860);
and U9969 (N_9969,N_9798,N_9838);
or U9970 (N_9970,N_9898,N_9889);
xnor U9971 (N_9971,N_9881,N_9851);
nor U9972 (N_9972,N_9761,N_9752);
or U9973 (N_9973,N_9788,N_9792);
nand U9974 (N_9974,N_9880,N_9861);
nand U9975 (N_9975,N_9884,N_9789);
nand U9976 (N_9976,N_9782,N_9801);
nand U9977 (N_9977,N_9841,N_9889);
or U9978 (N_9978,N_9894,N_9877);
xor U9979 (N_9979,N_9761,N_9759);
nand U9980 (N_9980,N_9789,N_9758);
nand U9981 (N_9981,N_9789,N_9830);
and U9982 (N_9982,N_9776,N_9852);
xor U9983 (N_9983,N_9754,N_9832);
and U9984 (N_9984,N_9876,N_9751);
nor U9985 (N_9985,N_9760,N_9836);
nand U9986 (N_9986,N_9880,N_9847);
nand U9987 (N_9987,N_9847,N_9830);
nand U9988 (N_9988,N_9797,N_9793);
nor U9989 (N_9989,N_9839,N_9787);
and U9990 (N_9990,N_9847,N_9767);
nor U9991 (N_9991,N_9877,N_9751);
nor U9992 (N_9992,N_9766,N_9794);
xor U9993 (N_9993,N_9860,N_9772);
and U9994 (N_9994,N_9887,N_9876);
xnor U9995 (N_9995,N_9782,N_9869);
nand U9996 (N_9996,N_9815,N_9876);
or U9997 (N_9997,N_9807,N_9832);
or U9998 (N_9998,N_9767,N_9753);
xor U9999 (N_9999,N_9862,N_9893);
or U10000 (N_10000,N_9820,N_9767);
nand U10001 (N_10001,N_9851,N_9763);
or U10002 (N_10002,N_9885,N_9830);
xnor U10003 (N_10003,N_9873,N_9786);
nor U10004 (N_10004,N_9796,N_9843);
or U10005 (N_10005,N_9793,N_9824);
or U10006 (N_10006,N_9843,N_9879);
nand U10007 (N_10007,N_9760,N_9797);
and U10008 (N_10008,N_9884,N_9752);
xor U10009 (N_10009,N_9797,N_9877);
and U10010 (N_10010,N_9846,N_9784);
xor U10011 (N_10011,N_9842,N_9790);
xor U10012 (N_10012,N_9882,N_9785);
nand U10013 (N_10013,N_9760,N_9892);
nand U10014 (N_10014,N_9870,N_9851);
xnor U10015 (N_10015,N_9800,N_9898);
nand U10016 (N_10016,N_9769,N_9839);
nor U10017 (N_10017,N_9763,N_9778);
xnor U10018 (N_10018,N_9761,N_9898);
or U10019 (N_10019,N_9838,N_9866);
nand U10020 (N_10020,N_9850,N_9852);
nand U10021 (N_10021,N_9878,N_9778);
nand U10022 (N_10022,N_9799,N_9802);
or U10023 (N_10023,N_9807,N_9869);
and U10024 (N_10024,N_9890,N_9885);
xnor U10025 (N_10025,N_9896,N_9751);
xor U10026 (N_10026,N_9888,N_9858);
xnor U10027 (N_10027,N_9881,N_9815);
nand U10028 (N_10028,N_9766,N_9884);
xor U10029 (N_10029,N_9884,N_9777);
nor U10030 (N_10030,N_9815,N_9845);
nand U10031 (N_10031,N_9870,N_9755);
or U10032 (N_10032,N_9758,N_9861);
xnor U10033 (N_10033,N_9816,N_9785);
xnor U10034 (N_10034,N_9833,N_9842);
nor U10035 (N_10035,N_9865,N_9843);
or U10036 (N_10036,N_9810,N_9825);
and U10037 (N_10037,N_9773,N_9832);
or U10038 (N_10038,N_9784,N_9795);
and U10039 (N_10039,N_9760,N_9796);
and U10040 (N_10040,N_9855,N_9846);
or U10041 (N_10041,N_9820,N_9856);
nor U10042 (N_10042,N_9862,N_9839);
nor U10043 (N_10043,N_9872,N_9756);
or U10044 (N_10044,N_9890,N_9863);
or U10045 (N_10045,N_9793,N_9897);
or U10046 (N_10046,N_9807,N_9751);
or U10047 (N_10047,N_9822,N_9774);
nor U10048 (N_10048,N_9783,N_9866);
nand U10049 (N_10049,N_9844,N_9870);
or U10050 (N_10050,N_10023,N_9921);
xor U10051 (N_10051,N_10036,N_9934);
xor U10052 (N_10052,N_9963,N_10044);
nand U10053 (N_10053,N_9905,N_10015);
xnor U10054 (N_10054,N_10003,N_9944);
nand U10055 (N_10055,N_9901,N_10021);
xnor U10056 (N_10056,N_9939,N_9910);
xor U10057 (N_10057,N_10035,N_9922);
nor U10058 (N_10058,N_10001,N_10048);
and U10059 (N_10059,N_9940,N_9972);
xnor U10060 (N_10060,N_9938,N_9912);
and U10061 (N_10061,N_9937,N_10007);
nor U10062 (N_10062,N_9994,N_10029);
or U10063 (N_10063,N_9943,N_9970);
xnor U10064 (N_10064,N_10042,N_9908);
nand U10065 (N_10065,N_10031,N_9979);
nor U10066 (N_10066,N_10011,N_10025);
xnor U10067 (N_10067,N_9993,N_10024);
nor U10068 (N_10068,N_9911,N_9955);
and U10069 (N_10069,N_9920,N_9960);
nand U10070 (N_10070,N_10010,N_9991);
nor U10071 (N_10071,N_10004,N_9999);
nor U10072 (N_10072,N_10034,N_9957);
or U10073 (N_10073,N_9981,N_9917);
nand U10074 (N_10074,N_9988,N_9968);
nor U10075 (N_10075,N_9973,N_9998);
nand U10076 (N_10076,N_9965,N_9942);
xor U10077 (N_10077,N_9913,N_9907);
and U10078 (N_10078,N_9924,N_9962);
nand U10079 (N_10079,N_9914,N_10005);
and U10080 (N_10080,N_9926,N_9977);
or U10081 (N_10081,N_10019,N_9927);
nor U10082 (N_10082,N_9982,N_9986);
nor U10083 (N_10083,N_9976,N_10039);
and U10084 (N_10084,N_9916,N_9936);
or U10085 (N_10085,N_9956,N_9930);
nor U10086 (N_10086,N_9971,N_9949);
xor U10087 (N_10087,N_10026,N_9947);
xnor U10088 (N_10088,N_9909,N_9990);
and U10089 (N_10089,N_10045,N_9997);
and U10090 (N_10090,N_10041,N_9904);
nand U10091 (N_10091,N_9996,N_10030);
and U10092 (N_10092,N_9900,N_9967);
xnor U10093 (N_10093,N_9902,N_10012);
or U10094 (N_10094,N_9975,N_9923);
nor U10095 (N_10095,N_10018,N_9966);
nor U10096 (N_10096,N_9974,N_9989);
and U10097 (N_10097,N_10002,N_9959);
nor U10098 (N_10098,N_9918,N_10020);
nor U10099 (N_10099,N_10014,N_9961);
or U10100 (N_10100,N_9951,N_9903);
or U10101 (N_10101,N_9958,N_9906);
xnor U10102 (N_10102,N_9929,N_9948);
or U10103 (N_10103,N_9933,N_10037);
nand U10104 (N_10104,N_10043,N_9932);
nand U10105 (N_10105,N_10000,N_9992);
nor U10106 (N_10106,N_10006,N_9915);
nand U10107 (N_10107,N_9978,N_9987);
or U10108 (N_10108,N_9941,N_9995);
xnor U10109 (N_10109,N_10008,N_10016);
nor U10110 (N_10110,N_9919,N_9946);
and U10111 (N_10111,N_10033,N_9985);
xnor U10112 (N_10112,N_9925,N_9980);
or U10113 (N_10113,N_9935,N_9954);
nor U10114 (N_10114,N_10017,N_9983);
xor U10115 (N_10115,N_10049,N_10022);
or U10116 (N_10116,N_9984,N_10047);
nor U10117 (N_10117,N_10009,N_9928);
or U10118 (N_10118,N_9950,N_10040);
nor U10119 (N_10119,N_9931,N_10013);
and U10120 (N_10120,N_10028,N_10038);
xnor U10121 (N_10121,N_9952,N_9964);
nor U10122 (N_10122,N_9953,N_10032);
nand U10123 (N_10123,N_9945,N_9969);
and U10124 (N_10124,N_10027,N_10046);
nand U10125 (N_10125,N_9929,N_9925);
xnor U10126 (N_10126,N_9994,N_9906);
or U10127 (N_10127,N_9955,N_9958);
nor U10128 (N_10128,N_9976,N_9955);
nand U10129 (N_10129,N_9961,N_10037);
or U10130 (N_10130,N_10005,N_10017);
and U10131 (N_10131,N_10047,N_9906);
and U10132 (N_10132,N_9999,N_9988);
and U10133 (N_10133,N_9972,N_9939);
xnor U10134 (N_10134,N_10025,N_10013);
and U10135 (N_10135,N_9945,N_9960);
and U10136 (N_10136,N_9973,N_9935);
nand U10137 (N_10137,N_9903,N_10016);
nor U10138 (N_10138,N_9928,N_10033);
xor U10139 (N_10139,N_9948,N_9955);
and U10140 (N_10140,N_9974,N_9937);
or U10141 (N_10141,N_10040,N_9983);
and U10142 (N_10142,N_9903,N_9935);
or U10143 (N_10143,N_9972,N_10033);
nand U10144 (N_10144,N_9964,N_9921);
xnor U10145 (N_10145,N_9947,N_9941);
and U10146 (N_10146,N_9972,N_9954);
xnor U10147 (N_10147,N_10033,N_9966);
and U10148 (N_10148,N_10037,N_9916);
nand U10149 (N_10149,N_10038,N_9966);
nor U10150 (N_10150,N_9979,N_9982);
nor U10151 (N_10151,N_9964,N_9948);
nor U10152 (N_10152,N_9919,N_9979);
nand U10153 (N_10153,N_9977,N_9987);
nand U10154 (N_10154,N_9924,N_9990);
nor U10155 (N_10155,N_10045,N_9941);
xnor U10156 (N_10156,N_9903,N_9948);
nand U10157 (N_10157,N_9904,N_9943);
and U10158 (N_10158,N_9973,N_9959);
xor U10159 (N_10159,N_9943,N_9925);
nand U10160 (N_10160,N_9928,N_10019);
and U10161 (N_10161,N_9985,N_10018);
nand U10162 (N_10162,N_9947,N_9917);
nand U10163 (N_10163,N_9989,N_10022);
and U10164 (N_10164,N_9905,N_10047);
and U10165 (N_10165,N_10018,N_9962);
nand U10166 (N_10166,N_9996,N_10034);
nand U10167 (N_10167,N_9976,N_10025);
and U10168 (N_10168,N_10010,N_9917);
nand U10169 (N_10169,N_10003,N_9991);
nand U10170 (N_10170,N_9988,N_10046);
and U10171 (N_10171,N_10034,N_9962);
and U10172 (N_10172,N_10010,N_9954);
or U10173 (N_10173,N_9965,N_10022);
xor U10174 (N_10174,N_9940,N_9909);
and U10175 (N_10175,N_10017,N_9978);
nand U10176 (N_10176,N_10019,N_9980);
and U10177 (N_10177,N_9912,N_9941);
and U10178 (N_10178,N_9984,N_10021);
nand U10179 (N_10179,N_9952,N_9973);
or U10180 (N_10180,N_9936,N_9942);
xor U10181 (N_10181,N_10026,N_10010);
nor U10182 (N_10182,N_10046,N_10023);
and U10183 (N_10183,N_10017,N_9945);
and U10184 (N_10184,N_9968,N_9959);
xor U10185 (N_10185,N_10035,N_9989);
and U10186 (N_10186,N_10013,N_10000);
or U10187 (N_10187,N_9986,N_9944);
xnor U10188 (N_10188,N_10034,N_9946);
nor U10189 (N_10189,N_9909,N_10013);
xor U10190 (N_10190,N_9953,N_10014);
xor U10191 (N_10191,N_9981,N_10031);
or U10192 (N_10192,N_9957,N_10039);
nor U10193 (N_10193,N_9924,N_9989);
and U10194 (N_10194,N_9971,N_10010);
and U10195 (N_10195,N_9978,N_9947);
xor U10196 (N_10196,N_9959,N_10044);
or U10197 (N_10197,N_9935,N_10020);
nand U10198 (N_10198,N_9949,N_9924);
and U10199 (N_10199,N_9926,N_10000);
nor U10200 (N_10200,N_10125,N_10124);
xor U10201 (N_10201,N_10131,N_10174);
xnor U10202 (N_10202,N_10107,N_10064);
nand U10203 (N_10203,N_10065,N_10159);
and U10204 (N_10204,N_10140,N_10123);
nor U10205 (N_10205,N_10082,N_10105);
and U10206 (N_10206,N_10068,N_10146);
and U10207 (N_10207,N_10154,N_10167);
nor U10208 (N_10208,N_10108,N_10066);
nand U10209 (N_10209,N_10147,N_10151);
nor U10210 (N_10210,N_10080,N_10199);
xor U10211 (N_10211,N_10136,N_10067);
or U10212 (N_10212,N_10073,N_10087);
xor U10213 (N_10213,N_10061,N_10168);
or U10214 (N_10214,N_10163,N_10176);
or U10215 (N_10215,N_10091,N_10117);
and U10216 (N_10216,N_10113,N_10083);
or U10217 (N_10217,N_10070,N_10056);
nor U10218 (N_10218,N_10075,N_10187);
and U10219 (N_10219,N_10130,N_10170);
xnor U10220 (N_10220,N_10173,N_10138);
nand U10221 (N_10221,N_10057,N_10099);
or U10222 (N_10222,N_10137,N_10181);
and U10223 (N_10223,N_10104,N_10197);
xnor U10224 (N_10224,N_10189,N_10177);
nand U10225 (N_10225,N_10172,N_10102);
or U10226 (N_10226,N_10072,N_10185);
and U10227 (N_10227,N_10152,N_10096);
or U10228 (N_10228,N_10121,N_10122);
and U10229 (N_10229,N_10179,N_10142);
nand U10230 (N_10230,N_10115,N_10149);
nand U10231 (N_10231,N_10180,N_10054);
and U10232 (N_10232,N_10058,N_10133);
and U10233 (N_10233,N_10088,N_10079);
nand U10234 (N_10234,N_10119,N_10114);
xor U10235 (N_10235,N_10053,N_10192);
nor U10236 (N_10236,N_10171,N_10162);
xnor U10237 (N_10237,N_10116,N_10160);
nor U10238 (N_10238,N_10093,N_10059);
or U10239 (N_10239,N_10109,N_10145);
nor U10240 (N_10240,N_10186,N_10164);
and U10241 (N_10241,N_10112,N_10153);
or U10242 (N_10242,N_10090,N_10081);
nand U10243 (N_10243,N_10094,N_10051);
or U10244 (N_10244,N_10084,N_10158);
nand U10245 (N_10245,N_10078,N_10156);
and U10246 (N_10246,N_10120,N_10071);
or U10247 (N_10247,N_10118,N_10062);
and U10248 (N_10248,N_10100,N_10098);
and U10249 (N_10249,N_10148,N_10182);
nand U10250 (N_10250,N_10128,N_10076);
or U10251 (N_10251,N_10103,N_10074);
xor U10252 (N_10252,N_10063,N_10139);
nor U10253 (N_10253,N_10155,N_10069);
xor U10254 (N_10254,N_10183,N_10143);
nand U10255 (N_10255,N_10106,N_10193);
or U10256 (N_10256,N_10127,N_10198);
or U10257 (N_10257,N_10129,N_10191);
nor U10258 (N_10258,N_10052,N_10111);
xnor U10259 (N_10259,N_10161,N_10165);
nor U10260 (N_10260,N_10095,N_10077);
nand U10261 (N_10261,N_10101,N_10150);
and U10262 (N_10262,N_10060,N_10086);
nand U10263 (N_10263,N_10190,N_10184);
and U10264 (N_10264,N_10126,N_10055);
or U10265 (N_10265,N_10141,N_10157);
xor U10266 (N_10266,N_10097,N_10144);
nand U10267 (N_10267,N_10194,N_10196);
nand U10268 (N_10268,N_10050,N_10175);
nand U10269 (N_10269,N_10178,N_10132);
or U10270 (N_10270,N_10166,N_10188);
nand U10271 (N_10271,N_10134,N_10169);
nand U10272 (N_10272,N_10092,N_10089);
nor U10273 (N_10273,N_10135,N_10110);
or U10274 (N_10274,N_10195,N_10085);
nand U10275 (N_10275,N_10176,N_10124);
nor U10276 (N_10276,N_10142,N_10113);
nor U10277 (N_10277,N_10092,N_10126);
nor U10278 (N_10278,N_10074,N_10119);
nor U10279 (N_10279,N_10134,N_10184);
nand U10280 (N_10280,N_10166,N_10067);
nor U10281 (N_10281,N_10064,N_10147);
nand U10282 (N_10282,N_10052,N_10137);
and U10283 (N_10283,N_10090,N_10171);
nand U10284 (N_10284,N_10190,N_10150);
nor U10285 (N_10285,N_10074,N_10066);
or U10286 (N_10286,N_10115,N_10117);
xnor U10287 (N_10287,N_10080,N_10115);
and U10288 (N_10288,N_10106,N_10181);
or U10289 (N_10289,N_10134,N_10179);
nand U10290 (N_10290,N_10059,N_10118);
or U10291 (N_10291,N_10065,N_10068);
xor U10292 (N_10292,N_10140,N_10180);
or U10293 (N_10293,N_10152,N_10093);
nand U10294 (N_10294,N_10125,N_10131);
and U10295 (N_10295,N_10186,N_10057);
nor U10296 (N_10296,N_10160,N_10069);
and U10297 (N_10297,N_10168,N_10102);
xor U10298 (N_10298,N_10122,N_10079);
nand U10299 (N_10299,N_10105,N_10137);
xor U10300 (N_10300,N_10138,N_10157);
or U10301 (N_10301,N_10057,N_10138);
xor U10302 (N_10302,N_10110,N_10112);
nor U10303 (N_10303,N_10116,N_10059);
and U10304 (N_10304,N_10166,N_10092);
nand U10305 (N_10305,N_10125,N_10098);
nand U10306 (N_10306,N_10172,N_10113);
nor U10307 (N_10307,N_10155,N_10178);
or U10308 (N_10308,N_10093,N_10110);
or U10309 (N_10309,N_10154,N_10132);
and U10310 (N_10310,N_10119,N_10105);
nor U10311 (N_10311,N_10051,N_10052);
and U10312 (N_10312,N_10052,N_10102);
and U10313 (N_10313,N_10165,N_10175);
or U10314 (N_10314,N_10061,N_10156);
or U10315 (N_10315,N_10101,N_10124);
and U10316 (N_10316,N_10167,N_10173);
xnor U10317 (N_10317,N_10089,N_10052);
nor U10318 (N_10318,N_10060,N_10056);
xnor U10319 (N_10319,N_10066,N_10184);
and U10320 (N_10320,N_10195,N_10199);
and U10321 (N_10321,N_10197,N_10124);
nand U10322 (N_10322,N_10130,N_10121);
and U10323 (N_10323,N_10079,N_10132);
nor U10324 (N_10324,N_10128,N_10067);
and U10325 (N_10325,N_10184,N_10193);
nand U10326 (N_10326,N_10050,N_10170);
nand U10327 (N_10327,N_10122,N_10110);
nor U10328 (N_10328,N_10178,N_10092);
xor U10329 (N_10329,N_10129,N_10076);
and U10330 (N_10330,N_10078,N_10107);
or U10331 (N_10331,N_10199,N_10118);
nand U10332 (N_10332,N_10078,N_10125);
xnor U10333 (N_10333,N_10149,N_10170);
and U10334 (N_10334,N_10115,N_10155);
nand U10335 (N_10335,N_10161,N_10102);
nor U10336 (N_10336,N_10102,N_10179);
and U10337 (N_10337,N_10077,N_10073);
xor U10338 (N_10338,N_10053,N_10188);
nor U10339 (N_10339,N_10109,N_10124);
xnor U10340 (N_10340,N_10051,N_10108);
xor U10341 (N_10341,N_10098,N_10069);
nor U10342 (N_10342,N_10176,N_10095);
xor U10343 (N_10343,N_10174,N_10126);
xnor U10344 (N_10344,N_10063,N_10087);
xor U10345 (N_10345,N_10160,N_10161);
nand U10346 (N_10346,N_10161,N_10113);
and U10347 (N_10347,N_10163,N_10186);
and U10348 (N_10348,N_10144,N_10110);
nand U10349 (N_10349,N_10107,N_10065);
nand U10350 (N_10350,N_10292,N_10262);
xnor U10351 (N_10351,N_10297,N_10288);
and U10352 (N_10352,N_10268,N_10317);
nor U10353 (N_10353,N_10338,N_10321);
nor U10354 (N_10354,N_10216,N_10291);
xor U10355 (N_10355,N_10306,N_10227);
nor U10356 (N_10356,N_10319,N_10290);
nor U10357 (N_10357,N_10260,N_10264);
xnor U10358 (N_10358,N_10300,N_10265);
and U10359 (N_10359,N_10330,N_10276);
and U10360 (N_10360,N_10269,N_10334);
nand U10361 (N_10361,N_10206,N_10324);
or U10362 (N_10362,N_10201,N_10280);
nand U10363 (N_10363,N_10222,N_10301);
nor U10364 (N_10364,N_10245,N_10247);
nor U10365 (N_10365,N_10256,N_10255);
xnor U10366 (N_10366,N_10348,N_10345);
nor U10367 (N_10367,N_10248,N_10271);
xor U10368 (N_10368,N_10293,N_10230);
nand U10369 (N_10369,N_10274,N_10342);
xor U10370 (N_10370,N_10322,N_10331);
and U10371 (N_10371,N_10327,N_10340);
and U10372 (N_10372,N_10346,N_10349);
and U10373 (N_10373,N_10205,N_10305);
nor U10374 (N_10374,N_10261,N_10323);
or U10375 (N_10375,N_10244,N_10335);
nor U10376 (N_10376,N_10343,N_10217);
xor U10377 (N_10377,N_10235,N_10233);
and U10378 (N_10378,N_10229,N_10209);
or U10379 (N_10379,N_10314,N_10202);
and U10380 (N_10380,N_10226,N_10279);
or U10381 (N_10381,N_10302,N_10219);
and U10382 (N_10382,N_10309,N_10273);
nand U10383 (N_10383,N_10312,N_10303);
or U10384 (N_10384,N_10294,N_10249);
and U10385 (N_10385,N_10231,N_10210);
and U10386 (N_10386,N_10278,N_10281);
nor U10387 (N_10387,N_10267,N_10214);
nand U10388 (N_10388,N_10285,N_10266);
xnor U10389 (N_10389,N_10283,N_10339);
xnor U10390 (N_10390,N_10246,N_10307);
nor U10391 (N_10391,N_10298,N_10251);
nor U10392 (N_10392,N_10259,N_10337);
nor U10393 (N_10393,N_10313,N_10326);
nor U10394 (N_10394,N_10284,N_10289);
xnor U10395 (N_10395,N_10237,N_10253);
and U10396 (N_10396,N_10234,N_10329);
nand U10397 (N_10397,N_10213,N_10287);
and U10398 (N_10398,N_10208,N_10304);
or U10399 (N_10399,N_10221,N_10320);
xnor U10400 (N_10400,N_10203,N_10296);
and U10401 (N_10401,N_10207,N_10270);
nor U10402 (N_10402,N_10275,N_10218);
nand U10403 (N_10403,N_10347,N_10272);
and U10404 (N_10404,N_10240,N_10336);
nor U10405 (N_10405,N_10282,N_10310);
nor U10406 (N_10406,N_10341,N_10241);
nand U10407 (N_10407,N_10220,N_10295);
xor U10408 (N_10408,N_10243,N_10250);
xor U10409 (N_10409,N_10200,N_10311);
and U10410 (N_10410,N_10316,N_10299);
nor U10411 (N_10411,N_10257,N_10318);
and U10412 (N_10412,N_10228,N_10258);
or U10413 (N_10413,N_10254,N_10277);
nor U10414 (N_10414,N_10236,N_10332);
and U10415 (N_10415,N_10215,N_10325);
nor U10416 (N_10416,N_10204,N_10286);
or U10417 (N_10417,N_10239,N_10224);
or U10418 (N_10418,N_10308,N_10232);
nand U10419 (N_10419,N_10223,N_10238);
nor U10420 (N_10420,N_10263,N_10242);
nand U10421 (N_10421,N_10225,N_10211);
nor U10422 (N_10422,N_10315,N_10252);
nand U10423 (N_10423,N_10328,N_10333);
and U10424 (N_10424,N_10344,N_10212);
xnor U10425 (N_10425,N_10321,N_10300);
nand U10426 (N_10426,N_10260,N_10265);
and U10427 (N_10427,N_10342,N_10323);
xor U10428 (N_10428,N_10252,N_10214);
or U10429 (N_10429,N_10264,N_10317);
xor U10430 (N_10430,N_10290,N_10257);
nor U10431 (N_10431,N_10266,N_10267);
nor U10432 (N_10432,N_10298,N_10301);
nand U10433 (N_10433,N_10253,N_10324);
and U10434 (N_10434,N_10253,N_10221);
nor U10435 (N_10435,N_10214,N_10328);
and U10436 (N_10436,N_10321,N_10317);
nand U10437 (N_10437,N_10259,N_10237);
or U10438 (N_10438,N_10237,N_10216);
nand U10439 (N_10439,N_10286,N_10297);
or U10440 (N_10440,N_10299,N_10308);
or U10441 (N_10441,N_10213,N_10203);
or U10442 (N_10442,N_10331,N_10226);
xor U10443 (N_10443,N_10345,N_10246);
or U10444 (N_10444,N_10240,N_10222);
and U10445 (N_10445,N_10301,N_10325);
nand U10446 (N_10446,N_10260,N_10323);
or U10447 (N_10447,N_10287,N_10272);
and U10448 (N_10448,N_10311,N_10288);
and U10449 (N_10449,N_10311,N_10245);
or U10450 (N_10450,N_10282,N_10255);
nand U10451 (N_10451,N_10318,N_10244);
or U10452 (N_10452,N_10254,N_10344);
xor U10453 (N_10453,N_10337,N_10266);
or U10454 (N_10454,N_10336,N_10217);
nand U10455 (N_10455,N_10237,N_10297);
xor U10456 (N_10456,N_10308,N_10259);
nand U10457 (N_10457,N_10308,N_10249);
nand U10458 (N_10458,N_10207,N_10267);
nor U10459 (N_10459,N_10331,N_10309);
nand U10460 (N_10460,N_10202,N_10279);
or U10461 (N_10461,N_10315,N_10283);
and U10462 (N_10462,N_10347,N_10218);
or U10463 (N_10463,N_10245,N_10207);
nand U10464 (N_10464,N_10332,N_10305);
nor U10465 (N_10465,N_10329,N_10220);
xor U10466 (N_10466,N_10291,N_10261);
nor U10467 (N_10467,N_10222,N_10333);
or U10468 (N_10468,N_10308,N_10345);
or U10469 (N_10469,N_10222,N_10287);
nor U10470 (N_10470,N_10289,N_10335);
nor U10471 (N_10471,N_10200,N_10337);
xor U10472 (N_10472,N_10288,N_10229);
nor U10473 (N_10473,N_10217,N_10253);
xor U10474 (N_10474,N_10285,N_10243);
or U10475 (N_10475,N_10234,N_10251);
or U10476 (N_10476,N_10283,N_10306);
nor U10477 (N_10477,N_10278,N_10223);
nand U10478 (N_10478,N_10238,N_10263);
nand U10479 (N_10479,N_10286,N_10279);
nor U10480 (N_10480,N_10349,N_10252);
or U10481 (N_10481,N_10323,N_10320);
or U10482 (N_10482,N_10266,N_10301);
nor U10483 (N_10483,N_10273,N_10231);
or U10484 (N_10484,N_10344,N_10315);
nand U10485 (N_10485,N_10346,N_10268);
xnor U10486 (N_10486,N_10246,N_10247);
xnor U10487 (N_10487,N_10336,N_10222);
and U10488 (N_10488,N_10285,N_10271);
or U10489 (N_10489,N_10303,N_10317);
nand U10490 (N_10490,N_10218,N_10282);
xnor U10491 (N_10491,N_10237,N_10211);
nor U10492 (N_10492,N_10227,N_10247);
nor U10493 (N_10493,N_10292,N_10274);
xor U10494 (N_10494,N_10252,N_10323);
xor U10495 (N_10495,N_10319,N_10324);
xor U10496 (N_10496,N_10336,N_10337);
nand U10497 (N_10497,N_10308,N_10276);
and U10498 (N_10498,N_10236,N_10319);
or U10499 (N_10499,N_10311,N_10303);
and U10500 (N_10500,N_10492,N_10432);
xor U10501 (N_10501,N_10479,N_10374);
or U10502 (N_10502,N_10389,N_10480);
xor U10503 (N_10503,N_10392,N_10360);
and U10504 (N_10504,N_10354,N_10399);
xor U10505 (N_10505,N_10458,N_10387);
nor U10506 (N_10506,N_10459,N_10496);
xor U10507 (N_10507,N_10351,N_10465);
nor U10508 (N_10508,N_10355,N_10420);
nand U10509 (N_10509,N_10365,N_10372);
or U10510 (N_10510,N_10486,N_10402);
nand U10511 (N_10511,N_10424,N_10472);
xnor U10512 (N_10512,N_10474,N_10401);
or U10513 (N_10513,N_10370,N_10356);
xnor U10514 (N_10514,N_10476,N_10388);
nand U10515 (N_10515,N_10437,N_10383);
or U10516 (N_10516,N_10469,N_10357);
nand U10517 (N_10517,N_10380,N_10483);
or U10518 (N_10518,N_10410,N_10470);
nand U10519 (N_10519,N_10413,N_10381);
nand U10520 (N_10520,N_10448,N_10439);
or U10521 (N_10521,N_10428,N_10426);
and U10522 (N_10522,N_10433,N_10361);
and U10523 (N_10523,N_10404,N_10441);
nand U10524 (N_10524,N_10373,N_10416);
nor U10525 (N_10525,N_10450,N_10452);
xor U10526 (N_10526,N_10394,N_10406);
and U10527 (N_10527,N_10430,N_10369);
nor U10528 (N_10528,N_10478,N_10386);
or U10529 (N_10529,N_10417,N_10379);
xnor U10530 (N_10530,N_10384,N_10421);
xor U10531 (N_10531,N_10471,N_10449);
xnor U10532 (N_10532,N_10414,N_10396);
xnor U10533 (N_10533,N_10422,N_10456);
xnor U10534 (N_10534,N_10425,N_10440);
or U10535 (N_10535,N_10451,N_10444);
nor U10536 (N_10536,N_10412,N_10475);
nor U10537 (N_10537,N_10467,N_10455);
or U10538 (N_10538,N_10435,N_10484);
nand U10539 (N_10539,N_10443,N_10353);
nand U10540 (N_10540,N_10385,N_10453);
and U10541 (N_10541,N_10495,N_10371);
and U10542 (N_10542,N_10442,N_10481);
nor U10543 (N_10543,N_10391,N_10382);
nor U10544 (N_10544,N_10364,N_10415);
and U10545 (N_10545,N_10407,N_10434);
nand U10546 (N_10546,N_10487,N_10362);
nand U10547 (N_10547,N_10462,N_10490);
xnor U10548 (N_10548,N_10411,N_10419);
or U10549 (N_10549,N_10427,N_10494);
nand U10550 (N_10550,N_10431,N_10423);
and U10551 (N_10551,N_10377,N_10446);
or U10552 (N_10552,N_10403,N_10499);
nand U10553 (N_10553,N_10390,N_10482);
nand U10554 (N_10554,N_10473,N_10352);
nor U10555 (N_10555,N_10429,N_10408);
and U10556 (N_10556,N_10477,N_10366);
xor U10557 (N_10557,N_10464,N_10497);
and U10558 (N_10558,N_10350,N_10375);
nand U10559 (N_10559,N_10498,N_10463);
nor U10560 (N_10560,N_10493,N_10418);
and U10561 (N_10561,N_10378,N_10398);
xnor U10562 (N_10562,N_10405,N_10368);
and U10563 (N_10563,N_10457,N_10436);
nor U10564 (N_10564,N_10489,N_10397);
nor U10565 (N_10565,N_10485,N_10367);
nor U10566 (N_10566,N_10438,N_10376);
nand U10567 (N_10567,N_10395,N_10358);
xor U10568 (N_10568,N_10363,N_10393);
xor U10569 (N_10569,N_10460,N_10409);
and U10570 (N_10570,N_10400,N_10488);
xor U10571 (N_10571,N_10468,N_10454);
nor U10572 (N_10572,N_10466,N_10445);
nor U10573 (N_10573,N_10447,N_10461);
nand U10574 (N_10574,N_10491,N_10359);
or U10575 (N_10575,N_10436,N_10414);
and U10576 (N_10576,N_10425,N_10454);
xor U10577 (N_10577,N_10396,N_10421);
or U10578 (N_10578,N_10384,N_10382);
nor U10579 (N_10579,N_10424,N_10461);
nand U10580 (N_10580,N_10497,N_10420);
or U10581 (N_10581,N_10485,N_10415);
or U10582 (N_10582,N_10472,N_10373);
or U10583 (N_10583,N_10499,N_10419);
or U10584 (N_10584,N_10402,N_10465);
nor U10585 (N_10585,N_10421,N_10481);
or U10586 (N_10586,N_10487,N_10484);
or U10587 (N_10587,N_10490,N_10441);
xnor U10588 (N_10588,N_10405,N_10430);
nor U10589 (N_10589,N_10398,N_10371);
nor U10590 (N_10590,N_10434,N_10466);
xnor U10591 (N_10591,N_10414,N_10358);
xor U10592 (N_10592,N_10457,N_10444);
nand U10593 (N_10593,N_10405,N_10434);
nand U10594 (N_10594,N_10486,N_10487);
and U10595 (N_10595,N_10466,N_10400);
nor U10596 (N_10596,N_10379,N_10434);
nor U10597 (N_10597,N_10400,N_10496);
nor U10598 (N_10598,N_10429,N_10372);
nand U10599 (N_10599,N_10374,N_10481);
and U10600 (N_10600,N_10423,N_10415);
nand U10601 (N_10601,N_10362,N_10490);
nand U10602 (N_10602,N_10458,N_10356);
nor U10603 (N_10603,N_10407,N_10480);
or U10604 (N_10604,N_10362,N_10410);
or U10605 (N_10605,N_10410,N_10479);
and U10606 (N_10606,N_10496,N_10482);
xor U10607 (N_10607,N_10420,N_10421);
and U10608 (N_10608,N_10415,N_10368);
nand U10609 (N_10609,N_10449,N_10443);
or U10610 (N_10610,N_10364,N_10454);
nand U10611 (N_10611,N_10453,N_10496);
nor U10612 (N_10612,N_10387,N_10421);
nor U10613 (N_10613,N_10395,N_10492);
and U10614 (N_10614,N_10377,N_10410);
xor U10615 (N_10615,N_10373,N_10359);
and U10616 (N_10616,N_10441,N_10395);
or U10617 (N_10617,N_10411,N_10444);
and U10618 (N_10618,N_10464,N_10358);
or U10619 (N_10619,N_10354,N_10475);
nand U10620 (N_10620,N_10490,N_10407);
nor U10621 (N_10621,N_10467,N_10408);
xnor U10622 (N_10622,N_10360,N_10394);
or U10623 (N_10623,N_10499,N_10495);
nor U10624 (N_10624,N_10396,N_10386);
and U10625 (N_10625,N_10370,N_10410);
nor U10626 (N_10626,N_10367,N_10457);
and U10627 (N_10627,N_10401,N_10495);
xnor U10628 (N_10628,N_10420,N_10370);
nand U10629 (N_10629,N_10435,N_10402);
nand U10630 (N_10630,N_10429,N_10406);
nand U10631 (N_10631,N_10456,N_10477);
and U10632 (N_10632,N_10396,N_10457);
nand U10633 (N_10633,N_10367,N_10427);
or U10634 (N_10634,N_10469,N_10432);
nand U10635 (N_10635,N_10393,N_10355);
xnor U10636 (N_10636,N_10360,N_10448);
nor U10637 (N_10637,N_10498,N_10483);
and U10638 (N_10638,N_10418,N_10491);
nor U10639 (N_10639,N_10464,N_10450);
nand U10640 (N_10640,N_10445,N_10382);
and U10641 (N_10641,N_10478,N_10496);
and U10642 (N_10642,N_10423,N_10381);
xnor U10643 (N_10643,N_10439,N_10470);
or U10644 (N_10644,N_10368,N_10438);
nor U10645 (N_10645,N_10486,N_10365);
or U10646 (N_10646,N_10396,N_10425);
xor U10647 (N_10647,N_10414,N_10408);
and U10648 (N_10648,N_10443,N_10427);
or U10649 (N_10649,N_10436,N_10440);
or U10650 (N_10650,N_10647,N_10576);
nor U10651 (N_10651,N_10502,N_10579);
nor U10652 (N_10652,N_10611,N_10519);
xnor U10653 (N_10653,N_10541,N_10500);
xor U10654 (N_10654,N_10572,N_10625);
nor U10655 (N_10655,N_10559,N_10548);
xor U10656 (N_10656,N_10609,N_10531);
nand U10657 (N_10657,N_10526,N_10538);
or U10658 (N_10658,N_10584,N_10577);
xor U10659 (N_10659,N_10567,N_10648);
nor U10660 (N_10660,N_10558,N_10529);
xnor U10661 (N_10661,N_10503,N_10602);
xor U10662 (N_10662,N_10616,N_10540);
xnor U10663 (N_10663,N_10597,N_10610);
or U10664 (N_10664,N_10588,N_10598);
and U10665 (N_10665,N_10596,N_10628);
xor U10666 (N_10666,N_10574,N_10507);
or U10667 (N_10667,N_10600,N_10593);
and U10668 (N_10668,N_10537,N_10509);
nor U10669 (N_10669,N_10641,N_10520);
nand U10670 (N_10670,N_10517,N_10514);
nand U10671 (N_10671,N_10606,N_10586);
and U10672 (N_10672,N_10630,N_10644);
or U10673 (N_10673,N_10512,N_10624);
xor U10674 (N_10674,N_10605,N_10532);
xor U10675 (N_10675,N_10561,N_10632);
xor U10676 (N_10676,N_10542,N_10578);
and U10677 (N_10677,N_10642,N_10634);
nand U10678 (N_10678,N_10560,N_10621);
xor U10679 (N_10679,N_10543,N_10562);
and U10680 (N_10680,N_10518,N_10568);
nor U10681 (N_10681,N_10516,N_10508);
and U10682 (N_10682,N_10501,N_10554);
xnor U10683 (N_10683,N_10613,N_10637);
xor U10684 (N_10684,N_10585,N_10645);
xor U10685 (N_10685,N_10544,N_10612);
nor U10686 (N_10686,N_10591,N_10510);
nand U10687 (N_10687,N_10513,N_10607);
nor U10688 (N_10688,N_10608,N_10525);
or U10689 (N_10689,N_10618,N_10549);
xor U10690 (N_10690,N_10617,N_10601);
nor U10691 (N_10691,N_10627,N_10569);
or U10692 (N_10692,N_10629,N_10594);
nor U10693 (N_10693,N_10563,N_10527);
xnor U10694 (N_10694,N_10557,N_10649);
nand U10695 (N_10695,N_10515,N_10590);
xor U10696 (N_10696,N_10603,N_10631);
or U10697 (N_10697,N_10522,N_10580);
nand U10698 (N_10698,N_10546,N_10564);
and U10699 (N_10699,N_10511,N_10599);
and U10700 (N_10700,N_10622,N_10555);
xnor U10701 (N_10701,N_10619,N_10589);
nand U10702 (N_10702,N_10573,N_10553);
or U10703 (N_10703,N_10550,N_10533);
xnor U10704 (N_10704,N_10626,N_10639);
nand U10705 (N_10705,N_10504,N_10552);
xor U10706 (N_10706,N_10582,N_10638);
or U10707 (N_10707,N_10566,N_10534);
and U10708 (N_10708,N_10521,N_10530);
xnor U10709 (N_10709,N_10636,N_10640);
or U10710 (N_10710,N_10536,N_10581);
nor U10711 (N_10711,N_10623,N_10583);
or U10712 (N_10712,N_10523,N_10575);
or U10713 (N_10713,N_10505,N_10595);
and U10714 (N_10714,N_10551,N_10633);
xnor U10715 (N_10715,N_10646,N_10570);
xor U10716 (N_10716,N_10535,N_10614);
or U10717 (N_10717,N_10556,N_10545);
or U10718 (N_10718,N_10565,N_10615);
and U10719 (N_10719,N_10643,N_10547);
or U10720 (N_10720,N_10571,N_10528);
or U10721 (N_10721,N_10604,N_10592);
nor U10722 (N_10722,N_10506,N_10635);
nand U10723 (N_10723,N_10620,N_10524);
nand U10724 (N_10724,N_10539,N_10587);
nand U10725 (N_10725,N_10546,N_10513);
xor U10726 (N_10726,N_10621,N_10528);
xor U10727 (N_10727,N_10531,N_10631);
xnor U10728 (N_10728,N_10540,N_10517);
and U10729 (N_10729,N_10584,N_10563);
nand U10730 (N_10730,N_10640,N_10547);
xor U10731 (N_10731,N_10630,N_10605);
xor U10732 (N_10732,N_10623,N_10555);
or U10733 (N_10733,N_10589,N_10572);
or U10734 (N_10734,N_10506,N_10510);
nor U10735 (N_10735,N_10525,N_10523);
xor U10736 (N_10736,N_10605,N_10646);
and U10737 (N_10737,N_10612,N_10525);
or U10738 (N_10738,N_10510,N_10631);
nor U10739 (N_10739,N_10607,N_10527);
xnor U10740 (N_10740,N_10604,N_10589);
xor U10741 (N_10741,N_10631,N_10574);
nand U10742 (N_10742,N_10617,N_10635);
nand U10743 (N_10743,N_10562,N_10555);
nand U10744 (N_10744,N_10552,N_10635);
xor U10745 (N_10745,N_10630,N_10538);
nand U10746 (N_10746,N_10508,N_10555);
or U10747 (N_10747,N_10536,N_10579);
and U10748 (N_10748,N_10512,N_10565);
or U10749 (N_10749,N_10567,N_10592);
nor U10750 (N_10750,N_10512,N_10540);
and U10751 (N_10751,N_10564,N_10601);
or U10752 (N_10752,N_10641,N_10589);
or U10753 (N_10753,N_10563,N_10578);
nor U10754 (N_10754,N_10556,N_10503);
and U10755 (N_10755,N_10553,N_10546);
xor U10756 (N_10756,N_10589,N_10585);
nor U10757 (N_10757,N_10584,N_10554);
or U10758 (N_10758,N_10578,N_10604);
nor U10759 (N_10759,N_10612,N_10629);
xor U10760 (N_10760,N_10531,N_10638);
and U10761 (N_10761,N_10538,N_10540);
and U10762 (N_10762,N_10568,N_10649);
or U10763 (N_10763,N_10588,N_10534);
and U10764 (N_10764,N_10617,N_10609);
or U10765 (N_10765,N_10574,N_10560);
nand U10766 (N_10766,N_10542,N_10599);
nor U10767 (N_10767,N_10527,N_10552);
nand U10768 (N_10768,N_10548,N_10606);
xor U10769 (N_10769,N_10613,N_10550);
or U10770 (N_10770,N_10580,N_10581);
or U10771 (N_10771,N_10647,N_10555);
and U10772 (N_10772,N_10608,N_10603);
nand U10773 (N_10773,N_10535,N_10522);
xor U10774 (N_10774,N_10588,N_10634);
or U10775 (N_10775,N_10593,N_10624);
and U10776 (N_10776,N_10581,N_10589);
nand U10777 (N_10777,N_10635,N_10536);
or U10778 (N_10778,N_10584,N_10566);
xor U10779 (N_10779,N_10511,N_10594);
nor U10780 (N_10780,N_10542,N_10552);
nand U10781 (N_10781,N_10586,N_10545);
and U10782 (N_10782,N_10552,N_10513);
and U10783 (N_10783,N_10606,N_10519);
and U10784 (N_10784,N_10594,N_10592);
and U10785 (N_10785,N_10620,N_10639);
nand U10786 (N_10786,N_10626,N_10614);
nor U10787 (N_10787,N_10627,N_10635);
and U10788 (N_10788,N_10505,N_10602);
or U10789 (N_10789,N_10547,N_10512);
xor U10790 (N_10790,N_10580,N_10551);
or U10791 (N_10791,N_10589,N_10536);
or U10792 (N_10792,N_10630,N_10571);
xnor U10793 (N_10793,N_10604,N_10631);
nand U10794 (N_10794,N_10565,N_10632);
xnor U10795 (N_10795,N_10558,N_10540);
or U10796 (N_10796,N_10577,N_10606);
or U10797 (N_10797,N_10503,N_10521);
xor U10798 (N_10798,N_10509,N_10535);
xor U10799 (N_10799,N_10542,N_10568);
or U10800 (N_10800,N_10786,N_10669);
and U10801 (N_10801,N_10701,N_10672);
nor U10802 (N_10802,N_10761,N_10658);
or U10803 (N_10803,N_10792,N_10706);
nor U10804 (N_10804,N_10754,N_10710);
and U10805 (N_10805,N_10678,N_10712);
or U10806 (N_10806,N_10675,N_10770);
nor U10807 (N_10807,N_10795,N_10724);
nand U10808 (N_10808,N_10788,N_10680);
or U10809 (N_10809,N_10749,N_10682);
nand U10810 (N_10810,N_10773,N_10717);
or U10811 (N_10811,N_10711,N_10751);
nor U10812 (N_10812,N_10699,N_10777);
xnor U10813 (N_10813,N_10767,N_10796);
nand U10814 (N_10814,N_10787,N_10685);
nor U10815 (N_10815,N_10654,N_10657);
nor U10816 (N_10816,N_10698,N_10764);
xor U10817 (N_10817,N_10737,N_10691);
nand U10818 (N_10818,N_10772,N_10771);
nand U10819 (N_10819,N_10695,N_10671);
xnor U10820 (N_10820,N_10728,N_10719);
nor U10821 (N_10821,N_10731,N_10718);
and U10822 (N_10822,N_10650,N_10756);
nand U10823 (N_10823,N_10727,N_10743);
xor U10824 (N_10824,N_10709,N_10708);
nor U10825 (N_10825,N_10759,N_10704);
and U10826 (N_10826,N_10655,N_10730);
and U10827 (N_10827,N_10668,N_10740);
and U10828 (N_10828,N_10747,N_10664);
and U10829 (N_10829,N_10652,N_10790);
nand U10830 (N_10830,N_10694,N_10666);
or U10831 (N_10831,N_10752,N_10679);
nand U10832 (N_10832,N_10779,N_10793);
nor U10833 (N_10833,N_10681,N_10662);
nand U10834 (N_10834,N_10721,N_10738);
xor U10835 (N_10835,N_10765,N_10775);
xnor U10836 (N_10836,N_10656,N_10739);
or U10837 (N_10837,N_10726,N_10748);
and U10838 (N_10838,N_10746,N_10791);
nor U10839 (N_10839,N_10692,N_10688);
nor U10840 (N_10840,N_10735,N_10663);
or U10841 (N_10841,N_10673,N_10689);
nand U10842 (N_10842,N_10741,N_10729);
nand U10843 (N_10843,N_10677,N_10774);
nor U10844 (N_10844,N_10716,N_10742);
nand U10845 (N_10845,N_10794,N_10697);
or U10846 (N_10846,N_10782,N_10784);
xnor U10847 (N_10847,N_10653,N_10705);
xnor U10848 (N_10848,N_10769,N_10723);
nand U10849 (N_10849,N_10744,N_10783);
nor U10850 (N_10850,N_10667,N_10660);
xnor U10851 (N_10851,N_10725,N_10722);
nor U10852 (N_10852,N_10713,N_10651);
or U10853 (N_10853,N_10693,N_10707);
or U10854 (N_10854,N_10674,N_10676);
nor U10855 (N_10855,N_10715,N_10750);
or U10856 (N_10856,N_10781,N_10763);
xor U10857 (N_10857,N_10687,N_10714);
nor U10858 (N_10858,N_10799,N_10661);
xnor U10859 (N_10859,N_10659,N_10798);
and U10860 (N_10860,N_10757,N_10736);
nor U10861 (N_10861,N_10745,N_10797);
nand U10862 (N_10862,N_10734,N_10785);
or U10863 (N_10863,N_10702,N_10778);
or U10864 (N_10864,N_10684,N_10683);
and U10865 (N_10865,N_10762,N_10733);
xnor U10866 (N_10866,N_10700,N_10758);
xnor U10867 (N_10867,N_10690,N_10665);
and U10868 (N_10868,N_10755,N_10789);
nor U10869 (N_10869,N_10732,N_10768);
or U10870 (N_10870,N_10720,N_10780);
or U10871 (N_10871,N_10753,N_10686);
nor U10872 (N_10872,N_10760,N_10766);
nand U10873 (N_10873,N_10776,N_10703);
and U10874 (N_10874,N_10670,N_10696);
and U10875 (N_10875,N_10706,N_10795);
nor U10876 (N_10876,N_10749,N_10712);
and U10877 (N_10877,N_10717,N_10725);
xnor U10878 (N_10878,N_10738,N_10720);
xnor U10879 (N_10879,N_10688,N_10650);
nand U10880 (N_10880,N_10694,N_10769);
or U10881 (N_10881,N_10678,N_10654);
nor U10882 (N_10882,N_10782,N_10726);
nand U10883 (N_10883,N_10723,N_10721);
nand U10884 (N_10884,N_10777,N_10729);
and U10885 (N_10885,N_10786,N_10737);
and U10886 (N_10886,N_10685,N_10794);
or U10887 (N_10887,N_10756,N_10799);
and U10888 (N_10888,N_10777,N_10687);
nand U10889 (N_10889,N_10777,N_10745);
and U10890 (N_10890,N_10694,N_10681);
nor U10891 (N_10891,N_10683,N_10661);
nor U10892 (N_10892,N_10748,N_10686);
nand U10893 (N_10893,N_10652,N_10783);
xnor U10894 (N_10894,N_10671,N_10745);
nor U10895 (N_10895,N_10711,N_10681);
or U10896 (N_10896,N_10740,N_10714);
or U10897 (N_10897,N_10770,N_10702);
nor U10898 (N_10898,N_10661,N_10672);
and U10899 (N_10899,N_10773,N_10690);
nand U10900 (N_10900,N_10794,N_10775);
xor U10901 (N_10901,N_10793,N_10788);
or U10902 (N_10902,N_10774,N_10721);
xnor U10903 (N_10903,N_10758,N_10756);
nor U10904 (N_10904,N_10745,N_10664);
nor U10905 (N_10905,N_10703,N_10706);
xor U10906 (N_10906,N_10787,N_10761);
or U10907 (N_10907,N_10768,N_10679);
xnor U10908 (N_10908,N_10676,N_10671);
and U10909 (N_10909,N_10675,N_10781);
or U10910 (N_10910,N_10732,N_10713);
or U10911 (N_10911,N_10769,N_10733);
and U10912 (N_10912,N_10797,N_10701);
nand U10913 (N_10913,N_10731,N_10764);
nor U10914 (N_10914,N_10777,N_10796);
or U10915 (N_10915,N_10689,N_10701);
xnor U10916 (N_10916,N_10766,N_10745);
or U10917 (N_10917,N_10707,N_10740);
or U10918 (N_10918,N_10711,N_10652);
nand U10919 (N_10919,N_10716,N_10709);
nand U10920 (N_10920,N_10753,N_10731);
nor U10921 (N_10921,N_10782,N_10796);
nor U10922 (N_10922,N_10676,N_10723);
nor U10923 (N_10923,N_10657,N_10696);
and U10924 (N_10924,N_10792,N_10688);
xnor U10925 (N_10925,N_10718,N_10661);
or U10926 (N_10926,N_10666,N_10674);
nand U10927 (N_10927,N_10705,N_10652);
or U10928 (N_10928,N_10768,N_10718);
nand U10929 (N_10929,N_10667,N_10717);
nand U10930 (N_10930,N_10714,N_10726);
nand U10931 (N_10931,N_10662,N_10795);
nor U10932 (N_10932,N_10728,N_10681);
xnor U10933 (N_10933,N_10693,N_10789);
nand U10934 (N_10934,N_10723,N_10737);
nand U10935 (N_10935,N_10696,N_10764);
nand U10936 (N_10936,N_10679,N_10694);
nand U10937 (N_10937,N_10743,N_10748);
and U10938 (N_10938,N_10765,N_10770);
or U10939 (N_10939,N_10688,N_10694);
or U10940 (N_10940,N_10745,N_10792);
xnor U10941 (N_10941,N_10674,N_10702);
xnor U10942 (N_10942,N_10699,N_10664);
nand U10943 (N_10943,N_10778,N_10714);
xnor U10944 (N_10944,N_10785,N_10791);
xor U10945 (N_10945,N_10788,N_10672);
or U10946 (N_10946,N_10653,N_10760);
nor U10947 (N_10947,N_10715,N_10794);
nand U10948 (N_10948,N_10744,N_10756);
or U10949 (N_10949,N_10654,N_10673);
or U10950 (N_10950,N_10846,N_10809);
nor U10951 (N_10951,N_10817,N_10899);
or U10952 (N_10952,N_10833,N_10849);
and U10953 (N_10953,N_10828,N_10907);
and U10954 (N_10954,N_10879,N_10826);
nor U10955 (N_10955,N_10818,N_10893);
nor U10956 (N_10956,N_10883,N_10896);
xor U10957 (N_10957,N_10909,N_10916);
xor U10958 (N_10958,N_10811,N_10800);
or U10959 (N_10959,N_10816,N_10812);
nand U10960 (N_10960,N_10930,N_10802);
xnor U10961 (N_10961,N_10865,N_10923);
nor U10962 (N_10962,N_10924,N_10917);
and U10963 (N_10963,N_10884,N_10860);
or U10964 (N_10964,N_10840,N_10868);
and U10965 (N_10965,N_10844,N_10837);
xor U10966 (N_10966,N_10827,N_10903);
xor U10967 (N_10967,N_10820,N_10841);
xnor U10968 (N_10968,N_10932,N_10901);
and U10969 (N_10969,N_10929,N_10919);
or U10970 (N_10970,N_10880,N_10904);
or U10971 (N_10971,N_10898,N_10823);
nand U10972 (N_10972,N_10870,N_10854);
or U10973 (N_10973,N_10829,N_10825);
nand U10974 (N_10974,N_10861,N_10848);
xnor U10975 (N_10975,N_10830,N_10937);
xnor U10976 (N_10976,N_10871,N_10892);
and U10977 (N_10977,N_10872,N_10857);
or U10978 (N_10978,N_10882,N_10863);
and U10979 (N_10979,N_10845,N_10851);
nor U10980 (N_10980,N_10824,N_10918);
or U10981 (N_10981,N_10887,N_10834);
and U10982 (N_10982,N_10921,N_10821);
nor U10983 (N_10983,N_10835,N_10910);
or U10984 (N_10984,N_10843,N_10886);
nor U10985 (N_10985,N_10933,N_10922);
nor U10986 (N_10986,N_10869,N_10867);
and U10987 (N_10987,N_10913,N_10808);
nand U10988 (N_10988,N_10873,N_10934);
or U10989 (N_10989,N_10912,N_10850);
or U10990 (N_10990,N_10945,N_10928);
and U10991 (N_10991,N_10925,N_10931);
and U10992 (N_10992,N_10856,N_10819);
nor U10993 (N_10993,N_10832,N_10949);
and U10994 (N_10994,N_10822,N_10814);
nand U10995 (N_10995,N_10878,N_10842);
and U10996 (N_10996,N_10946,N_10885);
nor U10997 (N_10997,N_10935,N_10938);
xnor U10998 (N_10998,N_10915,N_10889);
xnor U10999 (N_10999,N_10847,N_10894);
or U11000 (N_11000,N_10911,N_10864);
nand U11001 (N_11001,N_10862,N_10900);
nand U11002 (N_11002,N_10941,N_10853);
nor U11003 (N_11003,N_10891,N_10948);
and U11004 (N_11004,N_10888,N_10804);
xor U11005 (N_11005,N_10803,N_10908);
and U11006 (N_11006,N_10914,N_10943);
nand U11007 (N_11007,N_10813,N_10942);
nor U11008 (N_11008,N_10902,N_10936);
nand U11009 (N_11009,N_10805,N_10897);
and U11010 (N_11010,N_10895,N_10855);
xor U11011 (N_11011,N_10944,N_10874);
xor U11012 (N_11012,N_10939,N_10876);
nor U11013 (N_11013,N_10836,N_10839);
xor U11014 (N_11014,N_10858,N_10926);
and U11015 (N_11015,N_10810,N_10838);
nor U11016 (N_11016,N_10927,N_10920);
or U11017 (N_11017,N_10852,N_10881);
or U11018 (N_11018,N_10906,N_10890);
and U11019 (N_11019,N_10947,N_10807);
and U11020 (N_11020,N_10905,N_10806);
or U11021 (N_11021,N_10815,N_10875);
xor U11022 (N_11022,N_10877,N_10940);
nor U11023 (N_11023,N_10866,N_10859);
nor U11024 (N_11024,N_10831,N_10801);
or U11025 (N_11025,N_10833,N_10924);
xor U11026 (N_11026,N_10909,N_10922);
nor U11027 (N_11027,N_10926,N_10865);
nand U11028 (N_11028,N_10888,N_10930);
nor U11029 (N_11029,N_10824,N_10935);
and U11030 (N_11030,N_10886,N_10807);
nand U11031 (N_11031,N_10931,N_10835);
and U11032 (N_11032,N_10875,N_10854);
nor U11033 (N_11033,N_10808,N_10934);
xor U11034 (N_11034,N_10934,N_10898);
and U11035 (N_11035,N_10916,N_10895);
or U11036 (N_11036,N_10832,N_10881);
nor U11037 (N_11037,N_10917,N_10811);
and U11038 (N_11038,N_10831,N_10855);
nand U11039 (N_11039,N_10808,N_10837);
or U11040 (N_11040,N_10820,N_10853);
nor U11041 (N_11041,N_10926,N_10842);
and U11042 (N_11042,N_10873,N_10846);
xnor U11043 (N_11043,N_10824,N_10862);
and U11044 (N_11044,N_10803,N_10858);
and U11045 (N_11045,N_10905,N_10827);
nor U11046 (N_11046,N_10880,N_10890);
or U11047 (N_11047,N_10841,N_10801);
nand U11048 (N_11048,N_10842,N_10833);
and U11049 (N_11049,N_10815,N_10837);
xnor U11050 (N_11050,N_10926,N_10903);
nand U11051 (N_11051,N_10871,N_10878);
nand U11052 (N_11052,N_10868,N_10831);
nor U11053 (N_11053,N_10823,N_10831);
nor U11054 (N_11054,N_10859,N_10823);
or U11055 (N_11055,N_10827,N_10900);
and U11056 (N_11056,N_10897,N_10823);
xor U11057 (N_11057,N_10892,N_10908);
or U11058 (N_11058,N_10878,N_10933);
or U11059 (N_11059,N_10870,N_10851);
nor U11060 (N_11060,N_10862,N_10921);
nand U11061 (N_11061,N_10899,N_10873);
or U11062 (N_11062,N_10922,N_10928);
nor U11063 (N_11063,N_10944,N_10806);
and U11064 (N_11064,N_10911,N_10808);
xnor U11065 (N_11065,N_10935,N_10811);
xor U11066 (N_11066,N_10942,N_10823);
xor U11067 (N_11067,N_10883,N_10803);
or U11068 (N_11068,N_10868,N_10833);
nand U11069 (N_11069,N_10894,N_10927);
nand U11070 (N_11070,N_10853,N_10936);
or U11071 (N_11071,N_10921,N_10891);
and U11072 (N_11072,N_10824,N_10819);
and U11073 (N_11073,N_10852,N_10925);
nand U11074 (N_11074,N_10867,N_10948);
and U11075 (N_11075,N_10854,N_10805);
and U11076 (N_11076,N_10877,N_10810);
nand U11077 (N_11077,N_10849,N_10855);
and U11078 (N_11078,N_10808,N_10945);
and U11079 (N_11079,N_10873,N_10800);
xor U11080 (N_11080,N_10902,N_10819);
nand U11081 (N_11081,N_10938,N_10829);
or U11082 (N_11082,N_10846,N_10906);
and U11083 (N_11083,N_10913,N_10838);
or U11084 (N_11084,N_10896,N_10892);
and U11085 (N_11085,N_10835,N_10823);
xnor U11086 (N_11086,N_10909,N_10925);
nor U11087 (N_11087,N_10836,N_10881);
and U11088 (N_11088,N_10846,N_10890);
nor U11089 (N_11089,N_10930,N_10918);
nor U11090 (N_11090,N_10868,N_10879);
or U11091 (N_11091,N_10908,N_10828);
or U11092 (N_11092,N_10914,N_10916);
xor U11093 (N_11093,N_10902,N_10814);
nor U11094 (N_11094,N_10803,N_10831);
nor U11095 (N_11095,N_10918,N_10833);
xnor U11096 (N_11096,N_10912,N_10914);
nand U11097 (N_11097,N_10863,N_10874);
nand U11098 (N_11098,N_10908,N_10830);
nor U11099 (N_11099,N_10870,N_10934);
nor U11100 (N_11100,N_11056,N_10979);
or U11101 (N_11101,N_11054,N_11097);
or U11102 (N_11102,N_11057,N_11073);
nand U11103 (N_11103,N_10984,N_11087);
nand U11104 (N_11104,N_11096,N_11027);
nand U11105 (N_11105,N_11006,N_11005);
xnor U11106 (N_11106,N_11064,N_11048);
or U11107 (N_11107,N_11044,N_10983);
nor U11108 (N_11108,N_10950,N_10953);
or U11109 (N_11109,N_11013,N_11059);
xnor U11110 (N_11110,N_11039,N_11034);
or U11111 (N_11111,N_10977,N_11038);
xnor U11112 (N_11112,N_11007,N_10981);
or U11113 (N_11113,N_11015,N_11098);
nand U11114 (N_11114,N_10956,N_11080);
nor U11115 (N_11115,N_11071,N_10985);
xnor U11116 (N_11116,N_10975,N_11042);
nor U11117 (N_11117,N_11070,N_11051);
xor U11118 (N_11118,N_11084,N_11011);
nor U11119 (N_11119,N_11018,N_11076);
xor U11120 (N_11120,N_11092,N_10995);
nand U11121 (N_11121,N_11090,N_11031);
or U11122 (N_11122,N_10962,N_11021);
and U11123 (N_11123,N_11058,N_11060);
and U11124 (N_11124,N_10992,N_10997);
and U11125 (N_11125,N_11086,N_11037);
nor U11126 (N_11126,N_10993,N_10967);
or U11127 (N_11127,N_11068,N_11000);
and U11128 (N_11128,N_11049,N_10959);
nor U11129 (N_11129,N_11026,N_11043);
nor U11130 (N_11130,N_11099,N_10980);
nor U11131 (N_11131,N_10961,N_10982);
or U11132 (N_11132,N_10973,N_11033);
or U11133 (N_11133,N_11062,N_11074);
or U11134 (N_11134,N_10969,N_11032);
and U11135 (N_11135,N_11065,N_10954);
xnor U11136 (N_11136,N_11095,N_10987);
and U11137 (N_11137,N_11017,N_11066);
nor U11138 (N_11138,N_11078,N_11008);
and U11139 (N_11139,N_11036,N_10990);
and U11140 (N_11140,N_11081,N_10968);
xnor U11141 (N_11141,N_11061,N_11055);
nand U11142 (N_11142,N_10974,N_11041);
nor U11143 (N_11143,N_10991,N_11077);
nand U11144 (N_11144,N_11046,N_11019);
and U11145 (N_11145,N_11075,N_11085);
or U11146 (N_11146,N_10960,N_10952);
and U11147 (N_11147,N_11091,N_11022);
nor U11148 (N_11148,N_11050,N_11072);
or U11149 (N_11149,N_11004,N_11030);
xnor U11150 (N_11150,N_11012,N_11014);
nor U11151 (N_11151,N_10951,N_11063);
nand U11152 (N_11152,N_11003,N_11020);
nand U11153 (N_11153,N_11009,N_10971);
nand U11154 (N_11154,N_11052,N_11024);
nand U11155 (N_11155,N_11082,N_11069);
and U11156 (N_11156,N_11001,N_11088);
nor U11157 (N_11157,N_10955,N_10958);
nand U11158 (N_11158,N_11016,N_11029);
nor U11159 (N_11159,N_11053,N_10957);
or U11160 (N_11160,N_10965,N_10986);
nand U11161 (N_11161,N_10998,N_10966);
or U11162 (N_11162,N_11025,N_11079);
and U11163 (N_11163,N_11083,N_11010);
nand U11164 (N_11164,N_10994,N_11067);
nor U11165 (N_11165,N_10989,N_10963);
nand U11166 (N_11166,N_11094,N_11093);
nand U11167 (N_11167,N_10999,N_11035);
or U11168 (N_11168,N_11089,N_10988);
xor U11169 (N_11169,N_10972,N_10978);
nor U11170 (N_11170,N_10976,N_11028);
and U11171 (N_11171,N_11040,N_11002);
and U11172 (N_11172,N_10996,N_10964);
and U11173 (N_11173,N_11047,N_10970);
nor U11174 (N_11174,N_11023,N_11045);
and U11175 (N_11175,N_10973,N_10983);
nand U11176 (N_11176,N_11067,N_11074);
nor U11177 (N_11177,N_11092,N_11035);
and U11178 (N_11178,N_10975,N_10992);
nand U11179 (N_11179,N_11091,N_11003);
nand U11180 (N_11180,N_11008,N_10962);
nor U11181 (N_11181,N_11008,N_11053);
and U11182 (N_11182,N_11028,N_10956);
nand U11183 (N_11183,N_11051,N_11083);
nor U11184 (N_11184,N_11073,N_10960);
or U11185 (N_11185,N_11095,N_11073);
nor U11186 (N_11186,N_11067,N_10959);
xnor U11187 (N_11187,N_11035,N_10989);
xnor U11188 (N_11188,N_11063,N_11050);
and U11189 (N_11189,N_11034,N_11078);
nor U11190 (N_11190,N_11083,N_11012);
nand U11191 (N_11191,N_10968,N_10969);
xnor U11192 (N_11192,N_10994,N_11071);
nand U11193 (N_11193,N_10980,N_11062);
nand U11194 (N_11194,N_11074,N_10965);
or U11195 (N_11195,N_11039,N_10981);
xor U11196 (N_11196,N_11028,N_11059);
and U11197 (N_11197,N_11001,N_11020);
and U11198 (N_11198,N_11061,N_10964);
nand U11199 (N_11199,N_11083,N_11020);
nand U11200 (N_11200,N_10958,N_11083);
or U11201 (N_11201,N_11024,N_11044);
and U11202 (N_11202,N_10951,N_11016);
nand U11203 (N_11203,N_11067,N_11033);
or U11204 (N_11204,N_10957,N_11021);
nor U11205 (N_11205,N_11020,N_11012);
nor U11206 (N_11206,N_11059,N_11084);
nand U11207 (N_11207,N_10990,N_11082);
or U11208 (N_11208,N_10960,N_10981);
xnor U11209 (N_11209,N_10953,N_10995);
xor U11210 (N_11210,N_11063,N_11044);
or U11211 (N_11211,N_11085,N_11005);
or U11212 (N_11212,N_11099,N_10954);
or U11213 (N_11213,N_11088,N_11012);
nand U11214 (N_11214,N_11088,N_11034);
or U11215 (N_11215,N_11073,N_11034);
xor U11216 (N_11216,N_11049,N_11025);
or U11217 (N_11217,N_10974,N_11081);
or U11218 (N_11218,N_11088,N_11018);
xor U11219 (N_11219,N_11078,N_10972);
or U11220 (N_11220,N_11020,N_11027);
nand U11221 (N_11221,N_10954,N_10969);
or U11222 (N_11222,N_10990,N_10996);
nor U11223 (N_11223,N_11007,N_10979);
and U11224 (N_11224,N_11019,N_10966);
xnor U11225 (N_11225,N_11037,N_11015);
and U11226 (N_11226,N_10988,N_10970);
and U11227 (N_11227,N_11004,N_10982);
nand U11228 (N_11228,N_11035,N_11027);
nand U11229 (N_11229,N_10987,N_10979);
xnor U11230 (N_11230,N_11003,N_10972);
or U11231 (N_11231,N_11036,N_11044);
nand U11232 (N_11232,N_11010,N_11061);
nand U11233 (N_11233,N_10965,N_10998);
nand U11234 (N_11234,N_10972,N_11070);
or U11235 (N_11235,N_11009,N_10972);
xor U11236 (N_11236,N_11028,N_11043);
nand U11237 (N_11237,N_11083,N_11047);
and U11238 (N_11238,N_10991,N_10982);
xnor U11239 (N_11239,N_10999,N_10984);
or U11240 (N_11240,N_11066,N_11081);
nor U11241 (N_11241,N_11073,N_11068);
xor U11242 (N_11242,N_11089,N_11092);
nand U11243 (N_11243,N_11027,N_11014);
xnor U11244 (N_11244,N_10993,N_11043);
and U11245 (N_11245,N_11031,N_11063);
or U11246 (N_11246,N_10989,N_10977);
or U11247 (N_11247,N_11070,N_11092);
and U11248 (N_11248,N_11012,N_11017);
nor U11249 (N_11249,N_10976,N_10978);
and U11250 (N_11250,N_11110,N_11100);
and U11251 (N_11251,N_11236,N_11202);
or U11252 (N_11252,N_11221,N_11126);
xor U11253 (N_11253,N_11164,N_11226);
nor U11254 (N_11254,N_11129,N_11181);
and U11255 (N_11255,N_11134,N_11186);
or U11256 (N_11256,N_11238,N_11157);
or U11257 (N_11257,N_11116,N_11227);
nor U11258 (N_11258,N_11172,N_11224);
and U11259 (N_11259,N_11203,N_11122);
and U11260 (N_11260,N_11111,N_11103);
and U11261 (N_11261,N_11117,N_11171);
xnor U11262 (N_11262,N_11218,N_11245);
and U11263 (N_11263,N_11200,N_11127);
and U11264 (N_11264,N_11213,N_11178);
nor U11265 (N_11265,N_11188,N_11152);
or U11266 (N_11266,N_11174,N_11248);
xor U11267 (N_11267,N_11151,N_11191);
nor U11268 (N_11268,N_11131,N_11140);
nor U11269 (N_11269,N_11101,N_11220);
nor U11270 (N_11270,N_11231,N_11139);
nor U11271 (N_11271,N_11225,N_11158);
xor U11272 (N_11272,N_11168,N_11179);
or U11273 (N_11273,N_11135,N_11201);
xor U11274 (N_11274,N_11229,N_11118);
or U11275 (N_11275,N_11176,N_11109);
nand U11276 (N_11276,N_11119,N_11165);
nor U11277 (N_11277,N_11185,N_11183);
xor U11278 (N_11278,N_11195,N_11177);
or U11279 (N_11279,N_11156,N_11246);
and U11280 (N_11280,N_11237,N_11233);
nand U11281 (N_11281,N_11192,N_11137);
or U11282 (N_11282,N_11204,N_11147);
xnor U11283 (N_11283,N_11159,N_11124);
xor U11284 (N_11284,N_11113,N_11193);
xnor U11285 (N_11285,N_11241,N_11211);
xor U11286 (N_11286,N_11121,N_11136);
nand U11287 (N_11287,N_11115,N_11104);
or U11288 (N_11288,N_11112,N_11198);
nand U11289 (N_11289,N_11130,N_11120);
xnor U11290 (N_11290,N_11142,N_11215);
nor U11291 (N_11291,N_11228,N_11210);
and U11292 (N_11292,N_11209,N_11230);
xnor U11293 (N_11293,N_11128,N_11180);
and U11294 (N_11294,N_11235,N_11163);
and U11295 (N_11295,N_11167,N_11216);
nor U11296 (N_11296,N_11107,N_11239);
xnor U11297 (N_11297,N_11240,N_11123);
or U11298 (N_11298,N_11175,N_11214);
nor U11299 (N_11299,N_11196,N_11194);
nand U11300 (N_11300,N_11184,N_11125);
or U11301 (N_11301,N_11169,N_11199);
and U11302 (N_11302,N_11144,N_11219);
nand U11303 (N_11303,N_11173,N_11161);
xor U11304 (N_11304,N_11170,N_11222);
or U11305 (N_11305,N_11132,N_11190);
nand U11306 (N_11306,N_11145,N_11133);
nor U11307 (N_11307,N_11189,N_11149);
nand U11308 (N_11308,N_11102,N_11197);
or U11309 (N_11309,N_11143,N_11108);
nor U11310 (N_11310,N_11232,N_11155);
nor U11311 (N_11311,N_11162,N_11243);
and U11312 (N_11312,N_11223,N_11153);
nand U11313 (N_11313,N_11217,N_11205);
nand U11314 (N_11314,N_11106,N_11249);
xnor U11315 (N_11315,N_11212,N_11105);
nor U11316 (N_11316,N_11187,N_11160);
or U11317 (N_11317,N_11247,N_11206);
xor U11318 (N_11318,N_11166,N_11182);
or U11319 (N_11319,N_11114,N_11146);
nor U11320 (N_11320,N_11207,N_11234);
nand U11321 (N_11321,N_11150,N_11244);
xor U11322 (N_11322,N_11138,N_11141);
and U11323 (N_11323,N_11148,N_11208);
xnor U11324 (N_11324,N_11154,N_11242);
nand U11325 (N_11325,N_11198,N_11223);
or U11326 (N_11326,N_11156,N_11181);
and U11327 (N_11327,N_11212,N_11237);
and U11328 (N_11328,N_11102,N_11149);
or U11329 (N_11329,N_11173,N_11239);
nor U11330 (N_11330,N_11167,N_11243);
xnor U11331 (N_11331,N_11151,N_11199);
and U11332 (N_11332,N_11212,N_11215);
xnor U11333 (N_11333,N_11200,N_11112);
nor U11334 (N_11334,N_11101,N_11118);
nand U11335 (N_11335,N_11189,N_11225);
nor U11336 (N_11336,N_11191,N_11241);
xnor U11337 (N_11337,N_11139,N_11134);
or U11338 (N_11338,N_11187,N_11222);
nand U11339 (N_11339,N_11175,N_11136);
xnor U11340 (N_11340,N_11153,N_11230);
nor U11341 (N_11341,N_11220,N_11110);
nor U11342 (N_11342,N_11143,N_11211);
nand U11343 (N_11343,N_11195,N_11242);
nand U11344 (N_11344,N_11212,N_11203);
nand U11345 (N_11345,N_11134,N_11104);
or U11346 (N_11346,N_11213,N_11160);
nor U11347 (N_11347,N_11124,N_11156);
xor U11348 (N_11348,N_11230,N_11156);
xnor U11349 (N_11349,N_11118,N_11123);
nor U11350 (N_11350,N_11109,N_11181);
or U11351 (N_11351,N_11146,N_11154);
or U11352 (N_11352,N_11185,N_11235);
or U11353 (N_11353,N_11131,N_11210);
and U11354 (N_11354,N_11106,N_11201);
nand U11355 (N_11355,N_11118,N_11144);
and U11356 (N_11356,N_11132,N_11177);
nand U11357 (N_11357,N_11205,N_11168);
nor U11358 (N_11358,N_11109,N_11133);
xor U11359 (N_11359,N_11191,N_11116);
xnor U11360 (N_11360,N_11121,N_11175);
xnor U11361 (N_11361,N_11240,N_11192);
nor U11362 (N_11362,N_11195,N_11249);
xnor U11363 (N_11363,N_11184,N_11143);
and U11364 (N_11364,N_11175,N_11153);
nor U11365 (N_11365,N_11173,N_11123);
xnor U11366 (N_11366,N_11161,N_11162);
xnor U11367 (N_11367,N_11200,N_11237);
nand U11368 (N_11368,N_11243,N_11125);
and U11369 (N_11369,N_11107,N_11236);
nor U11370 (N_11370,N_11224,N_11137);
xnor U11371 (N_11371,N_11213,N_11228);
and U11372 (N_11372,N_11240,N_11229);
nor U11373 (N_11373,N_11230,N_11215);
and U11374 (N_11374,N_11233,N_11153);
xnor U11375 (N_11375,N_11220,N_11128);
xor U11376 (N_11376,N_11155,N_11108);
or U11377 (N_11377,N_11135,N_11160);
and U11378 (N_11378,N_11175,N_11201);
and U11379 (N_11379,N_11214,N_11100);
and U11380 (N_11380,N_11125,N_11235);
nand U11381 (N_11381,N_11154,N_11150);
nand U11382 (N_11382,N_11130,N_11221);
and U11383 (N_11383,N_11122,N_11179);
nor U11384 (N_11384,N_11192,N_11246);
and U11385 (N_11385,N_11187,N_11132);
and U11386 (N_11386,N_11145,N_11103);
and U11387 (N_11387,N_11212,N_11214);
xor U11388 (N_11388,N_11176,N_11105);
nor U11389 (N_11389,N_11182,N_11194);
or U11390 (N_11390,N_11100,N_11104);
nor U11391 (N_11391,N_11238,N_11146);
and U11392 (N_11392,N_11145,N_11172);
and U11393 (N_11393,N_11168,N_11125);
and U11394 (N_11394,N_11191,N_11164);
or U11395 (N_11395,N_11146,N_11161);
or U11396 (N_11396,N_11102,N_11249);
nor U11397 (N_11397,N_11216,N_11209);
and U11398 (N_11398,N_11115,N_11132);
nand U11399 (N_11399,N_11185,N_11207);
or U11400 (N_11400,N_11279,N_11292);
xnor U11401 (N_11401,N_11280,N_11300);
or U11402 (N_11402,N_11352,N_11291);
or U11403 (N_11403,N_11255,N_11378);
nor U11404 (N_11404,N_11281,N_11328);
xor U11405 (N_11405,N_11339,N_11285);
or U11406 (N_11406,N_11346,N_11350);
or U11407 (N_11407,N_11394,N_11298);
or U11408 (N_11408,N_11264,N_11327);
or U11409 (N_11409,N_11348,N_11276);
and U11410 (N_11410,N_11267,N_11286);
nor U11411 (N_11411,N_11322,N_11257);
nand U11412 (N_11412,N_11289,N_11368);
nand U11413 (N_11413,N_11284,N_11295);
xor U11414 (N_11414,N_11338,N_11376);
and U11415 (N_11415,N_11260,N_11333);
and U11416 (N_11416,N_11393,N_11335);
nor U11417 (N_11417,N_11358,N_11347);
nor U11418 (N_11418,N_11382,N_11366);
or U11419 (N_11419,N_11329,N_11282);
and U11420 (N_11420,N_11362,N_11306);
and U11421 (N_11421,N_11301,N_11251);
xnor U11422 (N_11422,N_11297,N_11356);
nor U11423 (N_11423,N_11321,N_11370);
nand U11424 (N_11424,N_11315,N_11367);
nand U11425 (N_11425,N_11363,N_11399);
and U11426 (N_11426,N_11360,N_11271);
or U11427 (N_11427,N_11256,N_11349);
nor U11428 (N_11428,N_11299,N_11277);
nand U11429 (N_11429,N_11354,N_11263);
or U11430 (N_11430,N_11381,N_11384);
or U11431 (N_11431,N_11269,N_11371);
or U11432 (N_11432,N_11364,N_11383);
and U11433 (N_11433,N_11325,N_11392);
xnor U11434 (N_11434,N_11397,N_11375);
and U11435 (N_11435,N_11357,N_11340);
xnor U11436 (N_11436,N_11307,N_11293);
or U11437 (N_11437,N_11254,N_11262);
nor U11438 (N_11438,N_11261,N_11305);
or U11439 (N_11439,N_11334,N_11396);
or U11440 (N_11440,N_11345,N_11250);
and U11441 (N_11441,N_11351,N_11309);
nor U11442 (N_11442,N_11341,N_11388);
and U11443 (N_11443,N_11353,N_11294);
xor U11444 (N_11444,N_11390,N_11374);
nand U11445 (N_11445,N_11296,N_11302);
and U11446 (N_11446,N_11389,N_11324);
nand U11447 (N_11447,N_11336,N_11318);
nor U11448 (N_11448,N_11359,N_11319);
nand U11449 (N_11449,N_11278,N_11310);
or U11450 (N_11450,N_11303,N_11268);
nand U11451 (N_11451,N_11273,N_11323);
and U11452 (N_11452,N_11283,N_11258);
or U11453 (N_11453,N_11337,N_11386);
and U11454 (N_11454,N_11343,N_11395);
nor U11455 (N_11455,N_11288,N_11365);
xnor U11456 (N_11456,N_11259,N_11377);
nor U11457 (N_11457,N_11253,N_11272);
or U11458 (N_11458,N_11373,N_11266);
nor U11459 (N_11459,N_11385,N_11311);
nor U11460 (N_11460,N_11331,N_11330);
nand U11461 (N_11461,N_11344,N_11379);
xnor U11462 (N_11462,N_11313,N_11265);
nor U11463 (N_11463,N_11275,N_11369);
xnor U11464 (N_11464,N_11372,N_11380);
nand U11465 (N_11465,N_11361,N_11398);
nand U11466 (N_11466,N_11320,N_11308);
and U11467 (N_11467,N_11314,N_11326);
and U11468 (N_11468,N_11342,N_11304);
and U11469 (N_11469,N_11391,N_11274);
nor U11470 (N_11470,N_11290,N_11355);
nor U11471 (N_11471,N_11387,N_11317);
or U11472 (N_11472,N_11270,N_11287);
xnor U11473 (N_11473,N_11316,N_11252);
or U11474 (N_11474,N_11332,N_11312);
and U11475 (N_11475,N_11319,N_11288);
and U11476 (N_11476,N_11268,N_11384);
xnor U11477 (N_11477,N_11329,N_11288);
nor U11478 (N_11478,N_11373,N_11338);
or U11479 (N_11479,N_11304,N_11394);
nand U11480 (N_11480,N_11294,N_11355);
or U11481 (N_11481,N_11398,N_11263);
nor U11482 (N_11482,N_11390,N_11395);
nand U11483 (N_11483,N_11287,N_11294);
or U11484 (N_11484,N_11353,N_11365);
nand U11485 (N_11485,N_11324,N_11332);
or U11486 (N_11486,N_11323,N_11284);
and U11487 (N_11487,N_11340,N_11303);
nand U11488 (N_11488,N_11395,N_11350);
nand U11489 (N_11489,N_11370,N_11263);
and U11490 (N_11490,N_11386,N_11297);
nand U11491 (N_11491,N_11368,N_11277);
nor U11492 (N_11492,N_11349,N_11281);
and U11493 (N_11493,N_11373,N_11366);
nand U11494 (N_11494,N_11285,N_11362);
and U11495 (N_11495,N_11263,N_11333);
nor U11496 (N_11496,N_11281,N_11278);
nor U11497 (N_11497,N_11350,N_11376);
and U11498 (N_11498,N_11356,N_11337);
and U11499 (N_11499,N_11339,N_11363);
or U11500 (N_11500,N_11300,N_11367);
and U11501 (N_11501,N_11373,N_11276);
xnor U11502 (N_11502,N_11394,N_11272);
nand U11503 (N_11503,N_11385,N_11299);
nand U11504 (N_11504,N_11354,N_11265);
and U11505 (N_11505,N_11310,N_11382);
or U11506 (N_11506,N_11294,N_11346);
and U11507 (N_11507,N_11261,N_11384);
or U11508 (N_11508,N_11344,N_11318);
and U11509 (N_11509,N_11269,N_11385);
or U11510 (N_11510,N_11348,N_11277);
or U11511 (N_11511,N_11279,N_11297);
nor U11512 (N_11512,N_11282,N_11298);
nor U11513 (N_11513,N_11284,N_11305);
or U11514 (N_11514,N_11258,N_11392);
nor U11515 (N_11515,N_11297,N_11288);
nor U11516 (N_11516,N_11290,N_11294);
xnor U11517 (N_11517,N_11292,N_11318);
nand U11518 (N_11518,N_11330,N_11256);
nor U11519 (N_11519,N_11335,N_11273);
nor U11520 (N_11520,N_11371,N_11299);
or U11521 (N_11521,N_11311,N_11277);
nand U11522 (N_11522,N_11325,N_11256);
xor U11523 (N_11523,N_11266,N_11342);
xnor U11524 (N_11524,N_11303,N_11293);
or U11525 (N_11525,N_11257,N_11253);
xnor U11526 (N_11526,N_11288,N_11306);
nand U11527 (N_11527,N_11298,N_11356);
xor U11528 (N_11528,N_11289,N_11257);
and U11529 (N_11529,N_11313,N_11364);
nor U11530 (N_11530,N_11352,N_11309);
nand U11531 (N_11531,N_11366,N_11290);
and U11532 (N_11532,N_11364,N_11332);
xnor U11533 (N_11533,N_11366,N_11272);
nor U11534 (N_11534,N_11302,N_11359);
and U11535 (N_11535,N_11370,N_11342);
xnor U11536 (N_11536,N_11290,N_11303);
xnor U11537 (N_11537,N_11261,N_11284);
nand U11538 (N_11538,N_11301,N_11297);
and U11539 (N_11539,N_11289,N_11323);
nor U11540 (N_11540,N_11298,N_11269);
and U11541 (N_11541,N_11331,N_11353);
nor U11542 (N_11542,N_11262,N_11263);
xnor U11543 (N_11543,N_11311,N_11319);
and U11544 (N_11544,N_11332,N_11276);
xnor U11545 (N_11545,N_11255,N_11263);
and U11546 (N_11546,N_11303,N_11253);
or U11547 (N_11547,N_11271,N_11371);
and U11548 (N_11548,N_11367,N_11349);
nor U11549 (N_11549,N_11361,N_11344);
nand U11550 (N_11550,N_11545,N_11433);
nor U11551 (N_11551,N_11504,N_11499);
or U11552 (N_11552,N_11420,N_11447);
nor U11553 (N_11553,N_11404,N_11413);
nand U11554 (N_11554,N_11489,N_11517);
nor U11555 (N_11555,N_11491,N_11459);
and U11556 (N_11556,N_11479,N_11511);
xor U11557 (N_11557,N_11414,N_11466);
or U11558 (N_11558,N_11529,N_11518);
and U11559 (N_11559,N_11541,N_11512);
or U11560 (N_11560,N_11448,N_11467);
nor U11561 (N_11561,N_11457,N_11549);
or U11562 (N_11562,N_11439,N_11493);
nor U11563 (N_11563,N_11417,N_11535);
nand U11564 (N_11564,N_11408,N_11488);
nand U11565 (N_11565,N_11484,N_11468);
or U11566 (N_11566,N_11492,N_11476);
and U11567 (N_11567,N_11515,N_11526);
and U11568 (N_11568,N_11410,N_11427);
xnor U11569 (N_11569,N_11415,N_11431);
xnor U11570 (N_11570,N_11537,N_11421);
or U11571 (N_11571,N_11501,N_11463);
or U11572 (N_11572,N_11542,N_11486);
nand U11573 (N_11573,N_11442,N_11543);
xor U11574 (N_11574,N_11498,N_11490);
nor U11575 (N_11575,N_11483,N_11422);
and U11576 (N_11576,N_11412,N_11524);
nand U11577 (N_11577,N_11530,N_11536);
nand U11578 (N_11578,N_11425,N_11438);
or U11579 (N_11579,N_11485,N_11465);
or U11580 (N_11580,N_11450,N_11528);
xor U11581 (N_11581,N_11435,N_11436);
xor U11582 (N_11582,N_11540,N_11520);
or U11583 (N_11583,N_11474,N_11470);
xnor U11584 (N_11584,N_11456,N_11445);
or U11585 (N_11585,N_11516,N_11471);
or U11586 (N_11586,N_11527,N_11453);
xor U11587 (N_11587,N_11482,N_11481);
and U11588 (N_11588,N_11429,N_11407);
or U11589 (N_11589,N_11444,N_11531);
nor U11590 (N_11590,N_11503,N_11454);
nand U11591 (N_11591,N_11525,N_11544);
or U11592 (N_11592,N_11405,N_11437);
or U11593 (N_11593,N_11514,N_11546);
nor U11594 (N_11594,N_11446,N_11478);
nand U11595 (N_11595,N_11547,N_11473);
nor U11596 (N_11596,N_11455,N_11495);
and U11597 (N_11597,N_11423,N_11521);
nor U11598 (N_11598,N_11548,N_11523);
and U11599 (N_11599,N_11502,N_11510);
and U11600 (N_11600,N_11452,N_11522);
and U11601 (N_11601,N_11507,N_11449);
and U11602 (N_11602,N_11508,N_11538);
xnor U11603 (N_11603,N_11406,N_11428);
and U11604 (N_11604,N_11461,N_11460);
nor U11605 (N_11605,N_11519,N_11539);
or U11606 (N_11606,N_11472,N_11430);
xnor U11607 (N_11607,N_11496,N_11400);
nor U11608 (N_11608,N_11440,N_11434);
and U11609 (N_11609,N_11416,N_11469);
xor U11610 (N_11610,N_11462,N_11506);
nor U11611 (N_11611,N_11419,N_11411);
xor U11612 (N_11612,N_11513,N_11487);
and U11613 (N_11613,N_11424,N_11480);
or U11614 (N_11614,N_11401,N_11509);
or U11615 (N_11615,N_11494,N_11477);
or U11616 (N_11616,N_11402,N_11426);
and U11617 (N_11617,N_11532,N_11451);
nor U11618 (N_11618,N_11500,N_11497);
nand U11619 (N_11619,N_11418,N_11409);
nand U11620 (N_11620,N_11505,N_11441);
or U11621 (N_11621,N_11443,N_11464);
and U11622 (N_11622,N_11432,N_11458);
and U11623 (N_11623,N_11403,N_11534);
and U11624 (N_11624,N_11475,N_11533);
xor U11625 (N_11625,N_11493,N_11490);
or U11626 (N_11626,N_11507,N_11444);
nor U11627 (N_11627,N_11477,N_11493);
and U11628 (N_11628,N_11531,N_11447);
xnor U11629 (N_11629,N_11525,N_11546);
nor U11630 (N_11630,N_11502,N_11471);
and U11631 (N_11631,N_11439,N_11540);
nor U11632 (N_11632,N_11425,N_11511);
nand U11633 (N_11633,N_11510,N_11454);
xnor U11634 (N_11634,N_11400,N_11429);
or U11635 (N_11635,N_11405,N_11445);
or U11636 (N_11636,N_11459,N_11546);
nor U11637 (N_11637,N_11410,N_11400);
or U11638 (N_11638,N_11504,N_11502);
nor U11639 (N_11639,N_11444,N_11469);
nor U11640 (N_11640,N_11410,N_11537);
nand U11641 (N_11641,N_11417,N_11434);
nand U11642 (N_11642,N_11407,N_11511);
xnor U11643 (N_11643,N_11513,N_11496);
nor U11644 (N_11644,N_11504,N_11473);
nor U11645 (N_11645,N_11400,N_11428);
or U11646 (N_11646,N_11533,N_11456);
nor U11647 (N_11647,N_11459,N_11446);
nand U11648 (N_11648,N_11545,N_11526);
nor U11649 (N_11649,N_11431,N_11500);
xnor U11650 (N_11650,N_11534,N_11532);
and U11651 (N_11651,N_11420,N_11410);
nand U11652 (N_11652,N_11498,N_11424);
nor U11653 (N_11653,N_11518,N_11544);
or U11654 (N_11654,N_11479,N_11454);
and U11655 (N_11655,N_11474,N_11489);
nor U11656 (N_11656,N_11432,N_11460);
and U11657 (N_11657,N_11521,N_11438);
nor U11658 (N_11658,N_11538,N_11442);
xor U11659 (N_11659,N_11537,N_11525);
and U11660 (N_11660,N_11491,N_11519);
xor U11661 (N_11661,N_11448,N_11483);
nor U11662 (N_11662,N_11518,N_11505);
xnor U11663 (N_11663,N_11482,N_11463);
and U11664 (N_11664,N_11455,N_11449);
nand U11665 (N_11665,N_11425,N_11539);
and U11666 (N_11666,N_11405,N_11491);
xnor U11667 (N_11667,N_11487,N_11542);
or U11668 (N_11668,N_11465,N_11410);
xnor U11669 (N_11669,N_11539,N_11474);
nor U11670 (N_11670,N_11544,N_11507);
xnor U11671 (N_11671,N_11475,N_11473);
nor U11672 (N_11672,N_11504,N_11538);
or U11673 (N_11673,N_11515,N_11546);
or U11674 (N_11674,N_11511,N_11540);
or U11675 (N_11675,N_11548,N_11455);
or U11676 (N_11676,N_11444,N_11450);
and U11677 (N_11677,N_11504,N_11440);
xnor U11678 (N_11678,N_11519,N_11508);
nor U11679 (N_11679,N_11419,N_11494);
nand U11680 (N_11680,N_11416,N_11535);
xnor U11681 (N_11681,N_11424,N_11503);
nor U11682 (N_11682,N_11438,N_11443);
xnor U11683 (N_11683,N_11470,N_11490);
nand U11684 (N_11684,N_11506,N_11500);
and U11685 (N_11685,N_11435,N_11424);
and U11686 (N_11686,N_11538,N_11529);
xor U11687 (N_11687,N_11456,N_11434);
or U11688 (N_11688,N_11458,N_11469);
and U11689 (N_11689,N_11542,N_11435);
xnor U11690 (N_11690,N_11407,N_11491);
nand U11691 (N_11691,N_11431,N_11438);
or U11692 (N_11692,N_11548,N_11415);
xnor U11693 (N_11693,N_11532,N_11433);
and U11694 (N_11694,N_11487,N_11449);
and U11695 (N_11695,N_11454,N_11481);
nor U11696 (N_11696,N_11460,N_11532);
nor U11697 (N_11697,N_11453,N_11450);
xnor U11698 (N_11698,N_11438,N_11444);
or U11699 (N_11699,N_11481,N_11450);
and U11700 (N_11700,N_11686,N_11669);
nor U11701 (N_11701,N_11668,N_11553);
xnor U11702 (N_11702,N_11578,N_11619);
nand U11703 (N_11703,N_11635,N_11621);
and U11704 (N_11704,N_11685,N_11646);
nand U11705 (N_11705,N_11630,N_11628);
xor U11706 (N_11706,N_11693,N_11594);
nand U11707 (N_11707,N_11580,N_11556);
nor U11708 (N_11708,N_11682,N_11656);
or U11709 (N_11709,N_11555,N_11609);
xnor U11710 (N_11710,N_11651,N_11625);
and U11711 (N_11711,N_11613,N_11590);
and U11712 (N_11712,N_11640,N_11652);
nor U11713 (N_11713,N_11627,N_11602);
xnor U11714 (N_11714,N_11551,N_11579);
xor U11715 (N_11715,N_11636,N_11573);
or U11716 (N_11716,N_11644,N_11643);
and U11717 (N_11717,N_11557,N_11661);
xnor U11718 (N_11718,N_11637,N_11663);
or U11719 (N_11719,N_11692,N_11695);
nor U11720 (N_11720,N_11599,N_11697);
and U11721 (N_11721,N_11698,N_11615);
xnor U11722 (N_11722,N_11670,N_11575);
and U11723 (N_11723,N_11563,N_11588);
nand U11724 (N_11724,N_11587,N_11649);
xor U11725 (N_11725,N_11560,N_11593);
or U11726 (N_11726,N_11632,N_11645);
or U11727 (N_11727,N_11567,N_11675);
nand U11728 (N_11728,N_11604,N_11659);
nor U11729 (N_11729,N_11654,N_11681);
nor U11730 (N_11730,N_11584,N_11606);
or U11731 (N_11731,N_11565,N_11629);
or U11732 (N_11732,N_11616,N_11673);
nand U11733 (N_11733,N_11631,N_11550);
and U11734 (N_11734,N_11634,N_11559);
nand U11735 (N_11735,N_11664,N_11660);
xnor U11736 (N_11736,N_11623,N_11591);
nand U11737 (N_11737,N_11603,N_11592);
or U11738 (N_11738,N_11564,N_11576);
xor U11739 (N_11739,N_11699,N_11566);
and U11740 (N_11740,N_11583,N_11679);
nor U11741 (N_11741,N_11595,N_11585);
nor U11742 (N_11742,N_11586,N_11624);
nor U11743 (N_11743,N_11689,N_11666);
nand U11744 (N_11744,N_11642,N_11650);
and U11745 (N_11745,N_11696,N_11600);
nand U11746 (N_11746,N_11648,N_11552);
or U11747 (N_11747,N_11598,N_11554);
and U11748 (N_11748,N_11607,N_11620);
or U11749 (N_11749,N_11687,N_11577);
or U11750 (N_11750,N_11562,N_11561);
nand U11751 (N_11751,N_11667,N_11655);
nor U11752 (N_11752,N_11572,N_11694);
and U11753 (N_11753,N_11683,N_11684);
or U11754 (N_11754,N_11653,N_11581);
nand U11755 (N_11755,N_11601,N_11690);
nor U11756 (N_11756,N_11626,N_11672);
or U11757 (N_11757,N_11612,N_11688);
nor U11758 (N_11758,N_11622,N_11676);
nand U11759 (N_11759,N_11597,N_11691);
nor U11760 (N_11760,N_11589,N_11558);
nor U11761 (N_11761,N_11618,N_11678);
xor U11762 (N_11762,N_11569,N_11570);
and U11763 (N_11763,N_11617,N_11639);
nor U11764 (N_11764,N_11568,N_11671);
nor U11765 (N_11765,N_11680,N_11574);
nor U11766 (N_11766,N_11665,N_11674);
nand U11767 (N_11767,N_11657,N_11610);
xnor U11768 (N_11768,N_11633,N_11571);
nand U11769 (N_11769,N_11582,N_11611);
or U11770 (N_11770,N_11605,N_11638);
xor U11771 (N_11771,N_11677,N_11608);
nand U11772 (N_11772,N_11662,N_11658);
or U11773 (N_11773,N_11641,N_11596);
or U11774 (N_11774,N_11614,N_11647);
xnor U11775 (N_11775,N_11652,N_11649);
or U11776 (N_11776,N_11582,N_11696);
nor U11777 (N_11777,N_11632,N_11677);
xor U11778 (N_11778,N_11578,N_11583);
nor U11779 (N_11779,N_11568,N_11577);
nor U11780 (N_11780,N_11610,N_11623);
or U11781 (N_11781,N_11633,N_11562);
and U11782 (N_11782,N_11566,N_11582);
and U11783 (N_11783,N_11552,N_11668);
nand U11784 (N_11784,N_11674,N_11598);
or U11785 (N_11785,N_11613,N_11621);
or U11786 (N_11786,N_11594,N_11677);
or U11787 (N_11787,N_11596,N_11680);
or U11788 (N_11788,N_11600,N_11639);
nand U11789 (N_11789,N_11664,N_11676);
or U11790 (N_11790,N_11661,N_11690);
and U11791 (N_11791,N_11692,N_11641);
or U11792 (N_11792,N_11645,N_11656);
nand U11793 (N_11793,N_11663,N_11595);
or U11794 (N_11794,N_11672,N_11610);
and U11795 (N_11795,N_11659,N_11657);
or U11796 (N_11796,N_11632,N_11691);
nor U11797 (N_11797,N_11668,N_11694);
and U11798 (N_11798,N_11582,N_11589);
and U11799 (N_11799,N_11665,N_11580);
nor U11800 (N_11800,N_11666,N_11589);
nor U11801 (N_11801,N_11574,N_11592);
nand U11802 (N_11802,N_11694,N_11675);
or U11803 (N_11803,N_11575,N_11657);
nand U11804 (N_11804,N_11604,N_11617);
xor U11805 (N_11805,N_11678,N_11622);
nand U11806 (N_11806,N_11601,N_11598);
and U11807 (N_11807,N_11606,N_11677);
nor U11808 (N_11808,N_11625,N_11668);
nand U11809 (N_11809,N_11630,N_11624);
nor U11810 (N_11810,N_11636,N_11569);
nand U11811 (N_11811,N_11635,N_11586);
nor U11812 (N_11812,N_11636,N_11633);
nand U11813 (N_11813,N_11605,N_11590);
or U11814 (N_11814,N_11561,N_11620);
nor U11815 (N_11815,N_11640,N_11635);
xor U11816 (N_11816,N_11614,N_11580);
and U11817 (N_11817,N_11554,N_11680);
nand U11818 (N_11818,N_11651,N_11552);
or U11819 (N_11819,N_11574,N_11663);
nand U11820 (N_11820,N_11625,N_11678);
nand U11821 (N_11821,N_11598,N_11614);
and U11822 (N_11822,N_11600,N_11622);
and U11823 (N_11823,N_11684,N_11580);
and U11824 (N_11824,N_11674,N_11595);
nor U11825 (N_11825,N_11689,N_11564);
xor U11826 (N_11826,N_11594,N_11685);
nor U11827 (N_11827,N_11570,N_11644);
or U11828 (N_11828,N_11564,N_11659);
and U11829 (N_11829,N_11609,N_11688);
or U11830 (N_11830,N_11556,N_11594);
nor U11831 (N_11831,N_11627,N_11673);
xnor U11832 (N_11832,N_11630,N_11572);
and U11833 (N_11833,N_11627,N_11639);
nor U11834 (N_11834,N_11610,N_11686);
nor U11835 (N_11835,N_11557,N_11554);
nor U11836 (N_11836,N_11567,N_11563);
nand U11837 (N_11837,N_11692,N_11682);
nand U11838 (N_11838,N_11575,N_11570);
nand U11839 (N_11839,N_11576,N_11587);
nor U11840 (N_11840,N_11679,N_11650);
and U11841 (N_11841,N_11666,N_11587);
or U11842 (N_11842,N_11683,N_11628);
nor U11843 (N_11843,N_11610,N_11693);
xnor U11844 (N_11844,N_11664,N_11585);
nor U11845 (N_11845,N_11637,N_11598);
or U11846 (N_11846,N_11609,N_11624);
or U11847 (N_11847,N_11666,N_11694);
nand U11848 (N_11848,N_11608,N_11620);
and U11849 (N_11849,N_11644,N_11684);
nand U11850 (N_11850,N_11838,N_11800);
nor U11851 (N_11851,N_11818,N_11725);
nand U11852 (N_11852,N_11828,N_11735);
or U11853 (N_11853,N_11746,N_11714);
and U11854 (N_11854,N_11719,N_11762);
or U11855 (N_11855,N_11738,N_11755);
xor U11856 (N_11856,N_11842,N_11841);
nand U11857 (N_11857,N_11777,N_11802);
or U11858 (N_11858,N_11748,N_11705);
or U11859 (N_11859,N_11816,N_11731);
xor U11860 (N_11860,N_11791,N_11712);
xnor U11861 (N_11861,N_11744,N_11811);
nand U11862 (N_11862,N_11826,N_11785);
and U11863 (N_11863,N_11837,N_11814);
xnor U11864 (N_11864,N_11703,N_11830);
nor U11865 (N_11865,N_11804,N_11779);
xor U11866 (N_11866,N_11722,N_11724);
nand U11867 (N_11867,N_11708,N_11789);
nor U11868 (N_11868,N_11780,N_11761);
nor U11869 (N_11869,N_11775,N_11817);
and U11870 (N_11870,N_11812,N_11803);
nand U11871 (N_11871,N_11786,N_11793);
nand U11872 (N_11872,N_11784,N_11776);
or U11873 (N_11873,N_11796,N_11706);
or U11874 (N_11874,N_11717,N_11824);
xor U11875 (N_11875,N_11726,N_11749);
and U11876 (N_11876,N_11745,N_11750);
xor U11877 (N_11877,N_11768,N_11741);
nor U11878 (N_11878,N_11711,N_11778);
or U11879 (N_11879,N_11718,N_11707);
or U11880 (N_11880,N_11773,N_11760);
nor U11881 (N_11881,N_11813,N_11821);
and U11882 (N_11882,N_11742,N_11835);
and U11883 (N_11883,N_11801,N_11831);
or U11884 (N_11884,N_11747,N_11700);
nor U11885 (N_11885,N_11765,N_11774);
nor U11886 (N_11886,N_11790,N_11763);
and U11887 (N_11887,N_11805,N_11819);
xnor U11888 (N_11888,N_11728,N_11729);
nand U11889 (N_11889,N_11716,N_11721);
nand U11890 (N_11890,N_11820,N_11736);
xnor U11891 (N_11891,N_11807,N_11815);
or U11892 (N_11892,N_11730,N_11848);
nand U11893 (N_11893,N_11734,N_11798);
nand U11894 (N_11894,N_11737,N_11701);
or U11895 (N_11895,N_11769,N_11733);
and U11896 (N_11896,N_11723,N_11727);
nor U11897 (N_11897,N_11836,N_11709);
and U11898 (N_11898,N_11756,N_11792);
nand U11899 (N_11899,N_11752,N_11839);
nand U11900 (N_11900,N_11758,N_11739);
or U11901 (N_11901,N_11787,N_11844);
xnor U11902 (N_11902,N_11766,N_11806);
nand U11903 (N_11903,N_11827,N_11770);
or U11904 (N_11904,N_11822,N_11751);
nor U11905 (N_11905,N_11767,N_11753);
or U11906 (N_11906,N_11832,N_11833);
and U11907 (N_11907,N_11715,N_11713);
nor U11908 (N_11908,N_11840,N_11757);
and U11909 (N_11909,N_11704,N_11710);
nand U11910 (N_11910,N_11771,N_11847);
nand U11911 (N_11911,N_11732,N_11834);
or U11912 (N_11912,N_11782,N_11794);
and U11913 (N_11913,N_11702,N_11799);
xnor U11914 (N_11914,N_11846,N_11788);
or U11915 (N_11915,N_11781,N_11849);
and U11916 (N_11916,N_11823,N_11795);
nand U11917 (N_11917,N_11797,N_11809);
or U11918 (N_11918,N_11829,N_11759);
or U11919 (N_11919,N_11740,N_11772);
and U11920 (N_11920,N_11845,N_11808);
xnor U11921 (N_11921,N_11764,N_11843);
xor U11922 (N_11922,N_11720,N_11754);
and U11923 (N_11923,N_11783,N_11743);
and U11924 (N_11924,N_11825,N_11810);
nand U11925 (N_11925,N_11818,N_11804);
nand U11926 (N_11926,N_11763,N_11720);
nor U11927 (N_11927,N_11831,N_11809);
or U11928 (N_11928,N_11703,N_11821);
nand U11929 (N_11929,N_11739,N_11837);
nand U11930 (N_11930,N_11790,N_11739);
and U11931 (N_11931,N_11758,N_11777);
nand U11932 (N_11932,N_11820,N_11785);
or U11933 (N_11933,N_11810,N_11813);
nor U11934 (N_11934,N_11813,N_11717);
or U11935 (N_11935,N_11812,N_11764);
and U11936 (N_11936,N_11719,N_11808);
nand U11937 (N_11937,N_11807,N_11738);
xnor U11938 (N_11938,N_11740,N_11825);
or U11939 (N_11939,N_11788,N_11789);
or U11940 (N_11940,N_11703,N_11705);
nand U11941 (N_11941,N_11815,N_11762);
nor U11942 (N_11942,N_11759,N_11827);
and U11943 (N_11943,N_11826,N_11782);
or U11944 (N_11944,N_11834,N_11703);
nor U11945 (N_11945,N_11761,N_11773);
or U11946 (N_11946,N_11706,N_11715);
xnor U11947 (N_11947,N_11820,N_11844);
xor U11948 (N_11948,N_11761,N_11803);
nand U11949 (N_11949,N_11800,N_11725);
xnor U11950 (N_11950,N_11718,N_11772);
or U11951 (N_11951,N_11759,N_11812);
or U11952 (N_11952,N_11730,N_11754);
xor U11953 (N_11953,N_11748,N_11713);
nand U11954 (N_11954,N_11780,N_11730);
xnor U11955 (N_11955,N_11802,N_11844);
and U11956 (N_11956,N_11817,N_11836);
or U11957 (N_11957,N_11738,N_11794);
nor U11958 (N_11958,N_11714,N_11767);
nand U11959 (N_11959,N_11743,N_11754);
and U11960 (N_11960,N_11836,N_11728);
xor U11961 (N_11961,N_11771,N_11785);
nand U11962 (N_11962,N_11756,N_11771);
or U11963 (N_11963,N_11794,N_11773);
nand U11964 (N_11964,N_11839,N_11800);
and U11965 (N_11965,N_11710,N_11846);
xnor U11966 (N_11966,N_11705,N_11808);
or U11967 (N_11967,N_11818,N_11755);
and U11968 (N_11968,N_11752,N_11815);
xor U11969 (N_11969,N_11766,N_11701);
nor U11970 (N_11970,N_11746,N_11720);
nor U11971 (N_11971,N_11839,N_11846);
and U11972 (N_11972,N_11747,N_11780);
and U11973 (N_11973,N_11826,N_11801);
nand U11974 (N_11974,N_11735,N_11821);
and U11975 (N_11975,N_11835,N_11707);
nor U11976 (N_11976,N_11748,N_11776);
xor U11977 (N_11977,N_11791,N_11754);
nand U11978 (N_11978,N_11785,N_11794);
and U11979 (N_11979,N_11702,N_11845);
nand U11980 (N_11980,N_11803,N_11747);
and U11981 (N_11981,N_11761,N_11718);
nand U11982 (N_11982,N_11786,N_11723);
xor U11983 (N_11983,N_11763,N_11819);
or U11984 (N_11984,N_11762,N_11807);
or U11985 (N_11985,N_11767,N_11821);
and U11986 (N_11986,N_11836,N_11751);
xnor U11987 (N_11987,N_11799,N_11792);
nand U11988 (N_11988,N_11738,N_11707);
xor U11989 (N_11989,N_11701,N_11731);
and U11990 (N_11990,N_11765,N_11798);
and U11991 (N_11991,N_11715,N_11801);
nand U11992 (N_11992,N_11736,N_11839);
or U11993 (N_11993,N_11771,N_11721);
or U11994 (N_11994,N_11837,N_11777);
xor U11995 (N_11995,N_11840,N_11790);
and U11996 (N_11996,N_11810,N_11712);
and U11997 (N_11997,N_11705,N_11732);
nand U11998 (N_11998,N_11780,N_11754);
xnor U11999 (N_11999,N_11759,N_11728);
nand U12000 (N_12000,N_11855,N_11921);
nand U12001 (N_12001,N_11945,N_11896);
nand U12002 (N_12002,N_11881,N_11906);
xnor U12003 (N_12003,N_11891,N_11926);
nand U12004 (N_12004,N_11866,N_11859);
nor U12005 (N_12005,N_11902,N_11877);
or U12006 (N_12006,N_11925,N_11898);
xnor U12007 (N_12007,N_11939,N_11951);
nand U12008 (N_12008,N_11999,N_11982);
and U12009 (N_12009,N_11934,N_11966);
nand U12010 (N_12010,N_11911,N_11989);
nand U12011 (N_12011,N_11930,N_11972);
nand U12012 (N_12012,N_11886,N_11947);
or U12013 (N_12013,N_11884,N_11998);
nor U12014 (N_12014,N_11956,N_11981);
nand U12015 (N_12015,N_11949,N_11927);
and U12016 (N_12016,N_11900,N_11991);
nor U12017 (N_12017,N_11931,N_11903);
nand U12018 (N_12018,N_11853,N_11978);
xor U12019 (N_12019,N_11996,N_11909);
nor U12020 (N_12020,N_11988,N_11916);
and U12021 (N_12021,N_11882,N_11852);
or U12022 (N_12022,N_11851,N_11917);
and U12023 (N_12023,N_11899,N_11987);
xnor U12024 (N_12024,N_11858,N_11980);
xnor U12025 (N_12025,N_11863,N_11983);
nand U12026 (N_12026,N_11936,N_11923);
nor U12027 (N_12027,N_11912,N_11963);
or U12028 (N_12028,N_11942,N_11967);
nor U12029 (N_12029,N_11965,N_11935);
nand U12030 (N_12030,N_11890,N_11862);
nor U12031 (N_12031,N_11889,N_11955);
nand U12032 (N_12032,N_11910,N_11893);
nand U12033 (N_12033,N_11958,N_11959);
nor U12034 (N_12034,N_11856,N_11997);
and U12035 (N_12035,N_11973,N_11854);
nor U12036 (N_12036,N_11888,N_11979);
and U12037 (N_12037,N_11977,N_11860);
nor U12038 (N_12038,N_11994,N_11929);
and U12039 (N_12039,N_11985,N_11897);
xnor U12040 (N_12040,N_11960,N_11915);
or U12041 (N_12041,N_11880,N_11894);
xor U12042 (N_12042,N_11957,N_11895);
and U12043 (N_12043,N_11976,N_11948);
nand U12044 (N_12044,N_11924,N_11943);
or U12045 (N_12045,N_11887,N_11940);
xnor U12046 (N_12046,N_11986,N_11938);
and U12047 (N_12047,N_11876,N_11969);
nand U12048 (N_12048,N_11964,N_11870);
xnor U12049 (N_12049,N_11954,N_11933);
xor U12050 (N_12050,N_11953,N_11868);
nor U12051 (N_12051,N_11920,N_11984);
nor U12052 (N_12052,N_11904,N_11992);
or U12053 (N_12053,N_11919,N_11908);
or U12054 (N_12054,N_11993,N_11914);
nand U12055 (N_12055,N_11922,N_11901);
or U12056 (N_12056,N_11869,N_11928);
nand U12057 (N_12057,N_11913,N_11875);
xor U12058 (N_12058,N_11865,N_11995);
nor U12059 (N_12059,N_11879,N_11905);
nand U12060 (N_12060,N_11990,N_11944);
nor U12061 (N_12061,N_11962,N_11970);
and U12062 (N_12062,N_11861,N_11892);
or U12063 (N_12063,N_11918,N_11975);
and U12064 (N_12064,N_11950,N_11850);
or U12065 (N_12065,N_11872,N_11946);
or U12066 (N_12066,N_11907,N_11867);
nand U12067 (N_12067,N_11873,N_11968);
nand U12068 (N_12068,N_11974,N_11878);
nor U12069 (N_12069,N_11857,N_11864);
and U12070 (N_12070,N_11937,N_11971);
nand U12071 (N_12071,N_11871,N_11885);
nand U12072 (N_12072,N_11961,N_11952);
xnor U12073 (N_12073,N_11941,N_11932);
and U12074 (N_12074,N_11874,N_11883);
nor U12075 (N_12075,N_11939,N_11921);
or U12076 (N_12076,N_11883,N_11972);
xnor U12077 (N_12077,N_11970,N_11885);
nand U12078 (N_12078,N_11907,N_11884);
xor U12079 (N_12079,N_11999,N_11918);
nand U12080 (N_12080,N_11963,N_11890);
and U12081 (N_12081,N_11997,N_11889);
and U12082 (N_12082,N_11923,N_11951);
and U12083 (N_12083,N_11943,N_11866);
and U12084 (N_12084,N_11925,N_11924);
nand U12085 (N_12085,N_11967,N_11885);
xnor U12086 (N_12086,N_11935,N_11980);
or U12087 (N_12087,N_11863,N_11909);
and U12088 (N_12088,N_11959,N_11892);
xor U12089 (N_12089,N_11924,N_11984);
nand U12090 (N_12090,N_11958,N_11851);
xnor U12091 (N_12091,N_11981,N_11966);
nor U12092 (N_12092,N_11975,N_11954);
and U12093 (N_12093,N_11967,N_11890);
or U12094 (N_12094,N_11935,N_11969);
and U12095 (N_12095,N_11860,N_11886);
and U12096 (N_12096,N_11958,N_11996);
xor U12097 (N_12097,N_11896,N_11871);
nand U12098 (N_12098,N_11936,N_11860);
xor U12099 (N_12099,N_11985,N_11931);
and U12100 (N_12100,N_11914,N_11922);
or U12101 (N_12101,N_11999,N_11969);
and U12102 (N_12102,N_11931,N_11892);
and U12103 (N_12103,N_11955,N_11871);
xor U12104 (N_12104,N_11862,N_11872);
nor U12105 (N_12105,N_11877,N_11966);
or U12106 (N_12106,N_11865,N_11936);
xor U12107 (N_12107,N_11881,N_11852);
and U12108 (N_12108,N_11851,N_11884);
xnor U12109 (N_12109,N_11943,N_11948);
or U12110 (N_12110,N_11946,N_11922);
nor U12111 (N_12111,N_11934,N_11868);
nor U12112 (N_12112,N_11876,N_11930);
nor U12113 (N_12113,N_11993,N_11866);
nand U12114 (N_12114,N_11963,N_11989);
and U12115 (N_12115,N_11852,N_11971);
and U12116 (N_12116,N_11865,N_11926);
nand U12117 (N_12117,N_11922,N_11962);
nor U12118 (N_12118,N_11863,N_11958);
xnor U12119 (N_12119,N_11992,N_11967);
nand U12120 (N_12120,N_11974,N_11958);
and U12121 (N_12121,N_11967,N_11857);
nand U12122 (N_12122,N_11976,N_11985);
or U12123 (N_12123,N_11936,N_11932);
xnor U12124 (N_12124,N_11956,N_11959);
or U12125 (N_12125,N_11936,N_11900);
xor U12126 (N_12126,N_11974,N_11990);
nand U12127 (N_12127,N_11912,N_11997);
and U12128 (N_12128,N_11883,N_11985);
xor U12129 (N_12129,N_11871,N_11898);
and U12130 (N_12130,N_11941,N_11897);
nand U12131 (N_12131,N_11966,N_11967);
nor U12132 (N_12132,N_11998,N_11893);
nor U12133 (N_12133,N_11888,N_11908);
and U12134 (N_12134,N_11936,N_11853);
xor U12135 (N_12135,N_11907,N_11962);
or U12136 (N_12136,N_11993,N_11979);
or U12137 (N_12137,N_11920,N_11864);
or U12138 (N_12138,N_11988,N_11922);
nor U12139 (N_12139,N_11858,N_11983);
or U12140 (N_12140,N_11913,N_11984);
xor U12141 (N_12141,N_11926,N_11987);
xnor U12142 (N_12142,N_11953,N_11857);
or U12143 (N_12143,N_11943,N_11908);
nor U12144 (N_12144,N_11918,N_11878);
xor U12145 (N_12145,N_11876,N_11970);
or U12146 (N_12146,N_11947,N_11885);
or U12147 (N_12147,N_11912,N_11928);
nor U12148 (N_12148,N_11892,N_11858);
and U12149 (N_12149,N_11941,N_11987);
and U12150 (N_12150,N_12113,N_12079);
and U12151 (N_12151,N_12008,N_12017);
xor U12152 (N_12152,N_12144,N_12028);
xor U12153 (N_12153,N_12085,N_12145);
nand U12154 (N_12154,N_12125,N_12015);
nand U12155 (N_12155,N_12050,N_12071);
xor U12156 (N_12156,N_12116,N_12078);
and U12157 (N_12157,N_12140,N_12060);
nor U12158 (N_12158,N_12056,N_12018);
nand U12159 (N_12159,N_12039,N_12112);
xnor U12160 (N_12160,N_12029,N_12124);
or U12161 (N_12161,N_12062,N_12073);
nand U12162 (N_12162,N_12033,N_12141);
xor U12163 (N_12163,N_12143,N_12107);
and U12164 (N_12164,N_12146,N_12005);
nand U12165 (N_12165,N_12032,N_12048);
and U12166 (N_12166,N_12076,N_12031);
nand U12167 (N_12167,N_12099,N_12069);
nand U12168 (N_12168,N_12109,N_12100);
and U12169 (N_12169,N_12058,N_12007);
and U12170 (N_12170,N_12128,N_12034);
xnor U12171 (N_12171,N_12023,N_12129);
or U12172 (N_12172,N_12096,N_12054);
nand U12173 (N_12173,N_12045,N_12091);
nor U12174 (N_12174,N_12021,N_12013);
xnor U12175 (N_12175,N_12094,N_12043);
or U12176 (N_12176,N_12011,N_12010);
or U12177 (N_12177,N_12119,N_12092);
nor U12178 (N_12178,N_12006,N_12088);
and U12179 (N_12179,N_12000,N_12135);
and U12180 (N_12180,N_12089,N_12072);
nor U12181 (N_12181,N_12123,N_12081);
nand U12182 (N_12182,N_12103,N_12070);
and U12183 (N_12183,N_12022,N_12003);
and U12184 (N_12184,N_12147,N_12019);
nand U12185 (N_12185,N_12049,N_12040);
nor U12186 (N_12186,N_12038,N_12042);
and U12187 (N_12187,N_12114,N_12097);
nand U12188 (N_12188,N_12142,N_12084);
xor U12189 (N_12189,N_12130,N_12064);
nand U12190 (N_12190,N_12044,N_12047);
nand U12191 (N_12191,N_12108,N_12137);
xnor U12192 (N_12192,N_12051,N_12012);
nand U12193 (N_12193,N_12035,N_12121);
xor U12194 (N_12194,N_12118,N_12061);
nand U12195 (N_12195,N_12009,N_12087);
nand U12196 (N_12196,N_12052,N_12041);
nor U12197 (N_12197,N_12075,N_12063);
nor U12198 (N_12198,N_12134,N_12046);
and U12199 (N_12199,N_12104,N_12068);
nand U12200 (N_12200,N_12066,N_12057);
nor U12201 (N_12201,N_12132,N_12106);
nand U12202 (N_12202,N_12037,N_12055);
or U12203 (N_12203,N_12082,N_12110);
nor U12204 (N_12204,N_12139,N_12020);
or U12205 (N_12205,N_12101,N_12086);
or U12206 (N_12206,N_12077,N_12053);
or U12207 (N_12207,N_12102,N_12080);
and U12208 (N_12208,N_12117,N_12027);
nor U12209 (N_12209,N_12093,N_12126);
and U12210 (N_12210,N_12122,N_12036);
nand U12211 (N_12211,N_12115,N_12065);
and U12212 (N_12212,N_12030,N_12059);
xor U12213 (N_12213,N_12025,N_12024);
xor U12214 (N_12214,N_12083,N_12149);
xnor U12215 (N_12215,N_12004,N_12026);
nor U12216 (N_12216,N_12014,N_12016);
nor U12217 (N_12217,N_12067,N_12098);
nand U12218 (N_12218,N_12111,N_12127);
nand U12219 (N_12219,N_12105,N_12133);
xor U12220 (N_12220,N_12120,N_12138);
nor U12221 (N_12221,N_12002,N_12001);
or U12222 (N_12222,N_12148,N_12074);
xor U12223 (N_12223,N_12131,N_12136);
nor U12224 (N_12224,N_12090,N_12095);
xnor U12225 (N_12225,N_12026,N_12103);
and U12226 (N_12226,N_12080,N_12118);
and U12227 (N_12227,N_12033,N_12051);
nand U12228 (N_12228,N_12119,N_12088);
and U12229 (N_12229,N_12023,N_12094);
nor U12230 (N_12230,N_12117,N_12024);
nand U12231 (N_12231,N_12027,N_12108);
and U12232 (N_12232,N_12109,N_12072);
xor U12233 (N_12233,N_12122,N_12144);
or U12234 (N_12234,N_12008,N_12033);
xnor U12235 (N_12235,N_12100,N_12043);
nand U12236 (N_12236,N_12119,N_12057);
nand U12237 (N_12237,N_12046,N_12075);
nand U12238 (N_12238,N_12117,N_12088);
or U12239 (N_12239,N_12080,N_12067);
nor U12240 (N_12240,N_12029,N_12059);
xor U12241 (N_12241,N_12029,N_12140);
and U12242 (N_12242,N_12054,N_12109);
nor U12243 (N_12243,N_12072,N_12086);
and U12244 (N_12244,N_12024,N_12129);
nand U12245 (N_12245,N_12104,N_12008);
nor U12246 (N_12246,N_12107,N_12101);
or U12247 (N_12247,N_12024,N_12074);
nand U12248 (N_12248,N_12066,N_12021);
and U12249 (N_12249,N_12091,N_12001);
or U12250 (N_12250,N_12065,N_12137);
or U12251 (N_12251,N_12112,N_12015);
xor U12252 (N_12252,N_12010,N_12138);
xnor U12253 (N_12253,N_12024,N_12128);
nand U12254 (N_12254,N_12005,N_12096);
nor U12255 (N_12255,N_12001,N_12010);
or U12256 (N_12256,N_12011,N_12089);
or U12257 (N_12257,N_12127,N_12041);
nand U12258 (N_12258,N_12131,N_12043);
nor U12259 (N_12259,N_12006,N_12130);
and U12260 (N_12260,N_12064,N_12093);
and U12261 (N_12261,N_12046,N_12042);
nand U12262 (N_12262,N_12139,N_12103);
and U12263 (N_12263,N_12116,N_12033);
nand U12264 (N_12264,N_12020,N_12119);
and U12265 (N_12265,N_12100,N_12005);
or U12266 (N_12266,N_12135,N_12125);
nor U12267 (N_12267,N_12059,N_12049);
and U12268 (N_12268,N_12029,N_12000);
or U12269 (N_12269,N_12089,N_12023);
nand U12270 (N_12270,N_12140,N_12051);
and U12271 (N_12271,N_12055,N_12124);
and U12272 (N_12272,N_12032,N_12025);
or U12273 (N_12273,N_12115,N_12079);
nor U12274 (N_12274,N_12054,N_12000);
or U12275 (N_12275,N_12120,N_12136);
nor U12276 (N_12276,N_12082,N_12044);
xnor U12277 (N_12277,N_12045,N_12141);
and U12278 (N_12278,N_12094,N_12120);
nand U12279 (N_12279,N_12096,N_12149);
or U12280 (N_12280,N_12053,N_12001);
nor U12281 (N_12281,N_12073,N_12145);
and U12282 (N_12282,N_12025,N_12100);
or U12283 (N_12283,N_12125,N_12045);
nand U12284 (N_12284,N_12041,N_12147);
nor U12285 (N_12285,N_12080,N_12041);
and U12286 (N_12286,N_12008,N_12060);
or U12287 (N_12287,N_12070,N_12040);
xnor U12288 (N_12288,N_12020,N_12064);
or U12289 (N_12289,N_12096,N_12114);
or U12290 (N_12290,N_12138,N_12093);
and U12291 (N_12291,N_12098,N_12108);
nand U12292 (N_12292,N_12082,N_12008);
xor U12293 (N_12293,N_12076,N_12138);
xnor U12294 (N_12294,N_12000,N_12067);
nor U12295 (N_12295,N_12125,N_12035);
and U12296 (N_12296,N_12143,N_12062);
xnor U12297 (N_12297,N_12126,N_12031);
or U12298 (N_12298,N_12076,N_12018);
or U12299 (N_12299,N_12109,N_12081);
nor U12300 (N_12300,N_12200,N_12258);
and U12301 (N_12301,N_12234,N_12191);
xor U12302 (N_12302,N_12266,N_12195);
nand U12303 (N_12303,N_12248,N_12214);
nand U12304 (N_12304,N_12196,N_12286);
or U12305 (N_12305,N_12172,N_12165);
nor U12306 (N_12306,N_12187,N_12203);
or U12307 (N_12307,N_12219,N_12282);
or U12308 (N_12308,N_12238,N_12185);
nand U12309 (N_12309,N_12295,N_12288);
and U12310 (N_12310,N_12184,N_12163);
and U12311 (N_12311,N_12161,N_12181);
nor U12312 (N_12312,N_12298,N_12299);
and U12313 (N_12313,N_12227,N_12255);
nand U12314 (N_12314,N_12267,N_12242);
nand U12315 (N_12315,N_12249,N_12275);
nor U12316 (N_12316,N_12157,N_12152);
or U12317 (N_12317,N_12269,N_12209);
nor U12318 (N_12318,N_12228,N_12220);
nand U12319 (N_12319,N_12287,N_12291);
nand U12320 (N_12320,N_12233,N_12174);
xnor U12321 (N_12321,N_12192,N_12237);
or U12322 (N_12322,N_12198,N_12271);
nor U12323 (N_12323,N_12178,N_12188);
or U12324 (N_12324,N_12221,N_12225);
nand U12325 (N_12325,N_12285,N_12229);
nor U12326 (N_12326,N_12205,N_12206);
nand U12327 (N_12327,N_12284,N_12189);
xor U12328 (N_12328,N_12171,N_12289);
and U12329 (N_12329,N_12263,N_12254);
nor U12330 (N_12330,N_12268,N_12247);
xnor U12331 (N_12331,N_12179,N_12273);
or U12332 (N_12332,N_12150,N_12186);
nand U12333 (N_12333,N_12283,N_12296);
nand U12334 (N_12334,N_12177,N_12158);
nand U12335 (N_12335,N_12217,N_12162);
nor U12336 (N_12336,N_12215,N_12155);
nor U12337 (N_12337,N_12256,N_12223);
and U12338 (N_12338,N_12252,N_12166);
or U12339 (N_12339,N_12243,N_12201);
nor U12340 (N_12340,N_12160,N_12204);
or U12341 (N_12341,N_12183,N_12167);
nor U12342 (N_12342,N_12182,N_12281);
nor U12343 (N_12343,N_12226,N_12224);
xnor U12344 (N_12344,N_12169,N_12239);
or U12345 (N_12345,N_12159,N_12262);
or U12346 (N_12346,N_12251,N_12272);
xnor U12347 (N_12347,N_12213,N_12168);
or U12348 (N_12348,N_12170,N_12290);
xor U12349 (N_12349,N_12277,N_12208);
xnor U12350 (N_12350,N_12297,N_12202);
nand U12351 (N_12351,N_12175,N_12207);
or U12352 (N_12352,N_12250,N_12278);
or U12353 (N_12353,N_12173,N_12199);
nand U12354 (N_12354,N_12294,N_12230);
xor U12355 (N_12355,N_12246,N_12218);
or U12356 (N_12356,N_12274,N_12292);
or U12357 (N_12357,N_12151,N_12253);
xor U12358 (N_12358,N_12279,N_12265);
or U12359 (N_12359,N_12211,N_12261);
xor U12360 (N_12360,N_12293,N_12241);
nand U12361 (N_12361,N_12232,N_12276);
xor U12362 (N_12362,N_12270,N_12280);
and U12363 (N_12363,N_12180,N_12231);
nand U12364 (N_12364,N_12240,N_12193);
nor U12365 (N_12365,N_12259,N_12222);
nand U12366 (N_12366,N_12244,N_12164);
nor U12367 (N_12367,N_12156,N_12245);
nand U12368 (N_12368,N_12236,N_12257);
nor U12369 (N_12369,N_12190,N_12235);
xnor U12370 (N_12370,N_12194,N_12197);
xor U12371 (N_12371,N_12176,N_12210);
and U12372 (N_12372,N_12154,N_12264);
xnor U12373 (N_12373,N_12216,N_12260);
nor U12374 (N_12374,N_12153,N_12212);
nor U12375 (N_12375,N_12189,N_12258);
nor U12376 (N_12376,N_12235,N_12284);
or U12377 (N_12377,N_12293,N_12195);
nor U12378 (N_12378,N_12170,N_12183);
xnor U12379 (N_12379,N_12155,N_12214);
nand U12380 (N_12380,N_12278,N_12225);
nand U12381 (N_12381,N_12152,N_12257);
and U12382 (N_12382,N_12229,N_12209);
or U12383 (N_12383,N_12184,N_12218);
xnor U12384 (N_12384,N_12218,N_12201);
xnor U12385 (N_12385,N_12297,N_12157);
or U12386 (N_12386,N_12286,N_12264);
xor U12387 (N_12387,N_12275,N_12176);
nand U12388 (N_12388,N_12263,N_12241);
or U12389 (N_12389,N_12213,N_12192);
nor U12390 (N_12390,N_12154,N_12220);
and U12391 (N_12391,N_12189,N_12201);
xor U12392 (N_12392,N_12265,N_12261);
or U12393 (N_12393,N_12176,N_12280);
xor U12394 (N_12394,N_12187,N_12201);
xor U12395 (N_12395,N_12206,N_12254);
nand U12396 (N_12396,N_12284,N_12224);
nor U12397 (N_12397,N_12214,N_12165);
and U12398 (N_12398,N_12220,N_12192);
nor U12399 (N_12399,N_12199,N_12152);
xnor U12400 (N_12400,N_12270,N_12168);
nor U12401 (N_12401,N_12285,N_12169);
or U12402 (N_12402,N_12238,N_12280);
or U12403 (N_12403,N_12193,N_12280);
or U12404 (N_12404,N_12185,N_12265);
xnor U12405 (N_12405,N_12178,N_12162);
xnor U12406 (N_12406,N_12236,N_12192);
or U12407 (N_12407,N_12167,N_12289);
or U12408 (N_12408,N_12157,N_12196);
nand U12409 (N_12409,N_12270,N_12264);
nor U12410 (N_12410,N_12279,N_12203);
and U12411 (N_12411,N_12214,N_12291);
or U12412 (N_12412,N_12278,N_12258);
xnor U12413 (N_12413,N_12174,N_12216);
nor U12414 (N_12414,N_12229,N_12240);
nor U12415 (N_12415,N_12178,N_12176);
and U12416 (N_12416,N_12182,N_12285);
or U12417 (N_12417,N_12235,N_12282);
or U12418 (N_12418,N_12158,N_12247);
xnor U12419 (N_12419,N_12237,N_12232);
xnor U12420 (N_12420,N_12293,N_12152);
and U12421 (N_12421,N_12194,N_12228);
xnor U12422 (N_12422,N_12254,N_12270);
or U12423 (N_12423,N_12278,N_12227);
nand U12424 (N_12424,N_12200,N_12256);
nor U12425 (N_12425,N_12258,N_12276);
nor U12426 (N_12426,N_12275,N_12278);
nand U12427 (N_12427,N_12256,N_12237);
or U12428 (N_12428,N_12185,N_12216);
and U12429 (N_12429,N_12226,N_12266);
xnor U12430 (N_12430,N_12180,N_12265);
or U12431 (N_12431,N_12265,N_12167);
nor U12432 (N_12432,N_12167,N_12290);
xnor U12433 (N_12433,N_12215,N_12202);
and U12434 (N_12434,N_12224,N_12252);
and U12435 (N_12435,N_12287,N_12215);
nor U12436 (N_12436,N_12283,N_12279);
or U12437 (N_12437,N_12294,N_12176);
or U12438 (N_12438,N_12236,N_12227);
or U12439 (N_12439,N_12202,N_12250);
xor U12440 (N_12440,N_12207,N_12256);
nor U12441 (N_12441,N_12184,N_12270);
or U12442 (N_12442,N_12237,N_12204);
and U12443 (N_12443,N_12182,N_12276);
or U12444 (N_12444,N_12285,N_12266);
nand U12445 (N_12445,N_12257,N_12286);
and U12446 (N_12446,N_12170,N_12271);
or U12447 (N_12447,N_12161,N_12274);
xnor U12448 (N_12448,N_12166,N_12233);
xnor U12449 (N_12449,N_12200,N_12271);
xor U12450 (N_12450,N_12398,N_12378);
xor U12451 (N_12451,N_12355,N_12405);
xor U12452 (N_12452,N_12396,N_12410);
xnor U12453 (N_12453,N_12430,N_12408);
nor U12454 (N_12454,N_12349,N_12389);
and U12455 (N_12455,N_12361,N_12354);
and U12456 (N_12456,N_12432,N_12309);
nand U12457 (N_12457,N_12395,N_12330);
or U12458 (N_12458,N_12304,N_12314);
or U12459 (N_12459,N_12318,N_12424);
nand U12460 (N_12460,N_12417,N_12436);
nand U12461 (N_12461,N_12365,N_12353);
or U12462 (N_12462,N_12350,N_12357);
or U12463 (N_12463,N_12306,N_12431);
nand U12464 (N_12464,N_12401,N_12352);
or U12465 (N_12465,N_12390,N_12356);
xnor U12466 (N_12466,N_12391,N_12428);
xor U12467 (N_12467,N_12383,N_12439);
nor U12468 (N_12468,N_12360,N_12308);
nand U12469 (N_12469,N_12399,N_12443);
xnor U12470 (N_12470,N_12363,N_12386);
nand U12471 (N_12471,N_12348,N_12415);
nor U12472 (N_12472,N_12420,N_12394);
and U12473 (N_12473,N_12406,N_12377);
or U12474 (N_12474,N_12444,N_12440);
nand U12475 (N_12475,N_12328,N_12336);
nand U12476 (N_12476,N_12324,N_12400);
nand U12477 (N_12477,N_12332,N_12435);
nor U12478 (N_12478,N_12445,N_12372);
nand U12479 (N_12479,N_12307,N_12313);
and U12480 (N_12480,N_12425,N_12423);
nor U12481 (N_12481,N_12376,N_12337);
and U12482 (N_12482,N_12421,N_12319);
nand U12483 (N_12483,N_12320,N_12333);
and U12484 (N_12484,N_12447,N_12413);
nor U12485 (N_12485,N_12414,N_12342);
or U12486 (N_12486,N_12416,N_12388);
nand U12487 (N_12487,N_12335,N_12317);
and U12488 (N_12488,N_12305,N_12323);
nor U12489 (N_12489,N_12334,N_12418);
and U12490 (N_12490,N_12446,N_12341);
and U12491 (N_12491,N_12409,N_12429);
xor U12492 (N_12492,N_12449,N_12382);
and U12493 (N_12493,N_12433,N_12301);
nor U12494 (N_12494,N_12427,N_12300);
and U12495 (N_12495,N_12325,N_12371);
nor U12496 (N_12496,N_12397,N_12404);
and U12497 (N_12497,N_12339,N_12366);
nand U12498 (N_12498,N_12434,N_12411);
xor U12499 (N_12499,N_12387,N_12422);
xnor U12500 (N_12500,N_12437,N_12385);
and U12501 (N_12501,N_12322,N_12327);
nor U12502 (N_12502,N_12346,N_12407);
nor U12503 (N_12503,N_12344,N_12331);
or U12504 (N_12504,N_12302,N_12329);
xor U12505 (N_12505,N_12379,N_12374);
nand U12506 (N_12506,N_12359,N_12438);
xnor U12507 (N_12507,N_12310,N_12362);
xor U12508 (N_12508,N_12351,N_12380);
and U12509 (N_12509,N_12381,N_12426);
or U12510 (N_12510,N_12311,N_12347);
nor U12511 (N_12511,N_12367,N_12338);
xnor U12512 (N_12512,N_12316,N_12448);
nor U12513 (N_12513,N_12315,N_12368);
nand U12514 (N_12514,N_12321,N_12392);
nand U12515 (N_12515,N_12303,N_12358);
and U12516 (N_12516,N_12345,N_12393);
or U12517 (N_12517,N_12419,N_12312);
and U12518 (N_12518,N_12442,N_12373);
and U12519 (N_12519,N_12340,N_12384);
or U12520 (N_12520,N_12369,N_12370);
or U12521 (N_12521,N_12402,N_12403);
or U12522 (N_12522,N_12364,N_12375);
xor U12523 (N_12523,N_12343,N_12412);
or U12524 (N_12524,N_12326,N_12441);
nor U12525 (N_12525,N_12336,N_12419);
and U12526 (N_12526,N_12319,N_12375);
and U12527 (N_12527,N_12356,N_12363);
xnor U12528 (N_12528,N_12340,N_12412);
nand U12529 (N_12529,N_12303,N_12377);
and U12530 (N_12530,N_12443,N_12428);
or U12531 (N_12531,N_12447,N_12346);
xnor U12532 (N_12532,N_12433,N_12425);
and U12533 (N_12533,N_12405,N_12447);
nand U12534 (N_12534,N_12409,N_12309);
xnor U12535 (N_12535,N_12334,N_12437);
xor U12536 (N_12536,N_12337,N_12404);
and U12537 (N_12537,N_12313,N_12417);
xnor U12538 (N_12538,N_12371,N_12443);
nor U12539 (N_12539,N_12428,N_12449);
nor U12540 (N_12540,N_12375,N_12449);
xor U12541 (N_12541,N_12352,N_12377);
nor U12542 (N_12542,N_12355,N_12371);
or U12543 (N_12543,N_12304,N_12306);
nor U12544 (N_12544,N_12423,N_12334);
nand U12545 (N_12545,N_12309,N_12408);
nor U12546 (N_12546,N_12379,N_12304);
nor U12547 (N_12547,N_12401,N_12380);
and U12548 (N_12548,N_12398,N_12304);
or U12549 (N_12549,N_12417,N_12364);
or U12550 (N_12550,N_12396,N_12431);
or U12551 (N_12551,N_12334,N_12395);
or U12552 (N_12552,N_12320,N_12434);
xor U12553 (N_12553,N_12449,N_12319);
xor U12554 (N_12554,N_12341,N_12376);
or U12555 (N_12555,N_12416,N_12350);
or U12556 (N_12556,N_12354,N_12444);
and U12557 (N_12557,N_12369,N_12314);
xor U12558 (N_12558,N_12340,N_12337);
xnor U12559 (N_12559,N_12355,N_12435);
xnor U12560 (N_12560,N_12418,N_12318);
nand U12561 (N_12561,N_12365,N_12370);
xor U12562 (N_12562,N_12418,N_12346);
and U12563 (N_12563,N_12361,N_12318);
and U12564 (N_12564,N_12376,N_12356);
nand U12565 (N_12565,N_12431,N_12301);
and U12566 (N_12566,N_12310,N_12316);
or U12567 (N_12567,N_12340,N_12372);
nand U12568 (N_12568,N_12365,N_12357);
nand U12569 (N_12569,N_12350,N_12445);
and U12570 (N_12570,N_12433,N_12375);
or U12571 (N_12571,N_12318,N_12415);
or U12572 (N_12572,N_12373,N_12302);
xor U12573 (N_12573,N_12342,N_12382);
and U12574 (N_12574,N_12371,N_12423);
nand U12575 (N_12575,N_12377,N_12329);
xnor U12576 (N_12576,N_12344,N_12391);
nor U12577 (N_12577,N_12438,N_12301);
nor U12578 (N_12578,N_12399,N_12307);
nor U12579 (N_12579,N_12308,N_12396);
xnor U12580 (N_12580,N_12383,N_12376);
nor U12581 (N_12581,N_12438,N_12335);
nand U12582 (N_12582,N_12417,N_12440);
nand U12583 (N_12583,N_12316,N_12377);
nor U12584 (N_12584,N_12319,N_12324);
nor U12585 (N_12585,N_12431,N_12318);
or U12586 (N_12586,N_12375,N_12437);
and U12587 (N_12587,N_12428,N_12366);
nand U12588 (N_12588,N_12322,N_12396);
or U12589 (N_12589,N_12329,N_12321);
nand U12590 (N_12590,N_12366,N_12418);
xor U12591 (N_12591,N_12349,N_12328);
xnor U12592 (N_12592,N_12325,N_12326);
xor U12593 (N_12593,N_12328,N_12350);
nand U12594 (N_12594,N_12434,N_12385);
or U12595 (N_12595,N_12423,N_12352);
xnor U12596 (N_12596,N_12437,N_12412);
xor U12597 (N_12597,N_12435,N_12344);
nand U12598 (N_12598,N_12366,N_12393);
or U12599 (N_12599,N_12306,N_12342);
nor U12600 (N_12600,N_12458,N_12578);
nor U12601 (N_12601,N_12525,N_12540);
and U12602 (N_12602,N_12488,N_12482);
nor U12603 (N_12603,N_12499,N_12541);
nand U12604 (N_12604,N_12536,N_12455);
xnor U12605 (N_12605,N_12465,N_12580);
and U12606 (N_12606,N_12514,N_12564);
or U12607 (N_12607,N_12461,N_12583);
xor U12608 (N_12608,N_12577,N_12464);
or U12609 (N_12609,N_12467,N_12593);
and U12610 (N_12610,N_12599,N_12506);
nand U12611 (N_12611,N_12556,N_12576);
nand U12612 (N_12612,N_12598,N_12551);
nand U12613 (N_12613,N_12498,N_12463);
nand U12614 (N_12614,N_12567,N_12517);
nor U12615 (N_12615,N_12454,N_12470);
nand U12616 (N_12616,N_12516,N_12574);
nor U12617 (N_12617,N_12459,N_12476);
nand U12618 (N_12618,N_12469,N_12535);
xnor U12619 (N_12619,N_12584,N_12460);
xnor U12620 (N_12620,N_12529,N_12594);
nor U12621 (N_12621,N_12552,N_12518);
nor U12622 (N_12622,N_12592,N_12542);
or U12623 (N_12623,N_12565,N_12489);
or U12624 (N_12624,N_12575,N_12477);
xnor U12625 (N_12625,N_12495,N_12504);
nor U12626 (N_12626,N_12558,N_12543);
and U12627 (N_12627,N_12490,N_12555);
xnor U12628 (N_12628,N_12595,N_12480);
nand U12629 (N_12629,N_12501,N_12472);
or U12630 (N_12630,N_12452,N_12523);
nand U12631 (N_12631,N_12557,N_12471);
nand U12632 (N_12632,N_12513,N_12561);
and U12633 (N_12633,N_12515,N_12596);
nor U12634 (N_12634,N_12533,N_12487);
or U12635 (N_12635,N_12481,N_12534);
nor U12636 (N_12636,N_12597,N_12586);
and U12637 (N_12637,N_12451,N_12473);
nand U12638 (N_12638,N_12522,N_12579);
and U12639 (N_12639,N_12563,N_12548);
nand U12640 (N_12640,N_12491,N_12478);
nor U12641 (N_12641,N_12483,N_12573);
nand U12642 (N_12642,N_12507,N_12520);
nand U12643 (N_12643,N_12512,N_12474);
xor U12644 (N_12644,N_12475,N_12545);
or U12645 (N_12645,N_12547,N_12485);
nand U12646 (N_12646,N_12570,N_12505);
nor U12647 (N_12647,N_12509,N_12496);
or U12648 (N_12648,N_12546,N_12486);
xor U12649 (N_12649,N_12553,N_12511);
or U12650 (N_12650,N_12560,N_12569);
and U12651 (N_12651,N_12559,N_12589);
nand U12652 (N_12652,N_12585,N_12493);
and U12653 (N_12653,N_12500,N_12554);
nor U12654 (N_12654,N_12562,N_12503);
and U12655 (N_12655,N_12591,N_12549);
or U12656 (N_12656,N_12571,N_12538);
nand U12657 (N_12657,N_12531,N_12590);
and U12658 (N_12658,N_12527,N_12468);
and U12659 (N_12659,N_12588,N_12537);
and U12660 (N_12660,N_12497,N_12526);
xor U12661 (N_12661,N_12456,N_12521);
xnor U12662 (N_12662,N_12453,N_12582);
or U12663 (N_12663,N_12568,N_12550);
and U12664 (N_12664,N_12530,N_12587);
nand U12665 (N_12665,N_12581,N_12466);
or U12666 (N_12666,N_12524,N_12519);
nand U12667 (N_12667,N_12508,N_12450);
or U12668 (N_12668,N_12484,N_12544);
and U12669 (N_12669,N_12572,N_12539);
or U12670 (N_12670,N_12510,N_12457);
or U12671 (N_12671,N_12502,N_12492);
nand U12672 (N_12672,N_12528,N_12494);
xor U12673 (N_12673,N_12532,N_12566);
or U12674 (N_12674,N_12462,N_12479);
nor U12675 (N_12675,N_12566,N_12455);
xor U12676 (N_12676,N_12494,N_12455);
nor U12677 (N_12677,N_12551,N_12532);
and U12678 (N_12678,N_12547,N_12524);
or U12679 (N_12679,N_12468,N_12530);
nand U12680 (N_12680,N_12539,N_12573);
nand U12681 (N_12681,N_12468,N_12561);
xor U12682 (N_12682,N_12499,N_12513);
xnor U12683 (N_12683,N_12581,N_12594);
nor U12684 (N_12684,N_12521,N_12583);
xor U12685 (N_12685,N_12573,N_12595);
or U12686 (N_12686,N_12565,N_12495);
nor U12687 (N_12687,N_12519,N_12571);
nand U12688 (N_12688,N_12531,N_12543);
xnor U12689 (N_12689,N_12589,N_12595);
nand U12690 (N_12690,N_12534,N_12460);
or U12691 (N_12691,N_12526,N_12560);
nand U12692 (N_12692,N_12578,N_12489);
nor U12693 (N_12693,N_12488,N_12490);
nand U12694 (N_12694,N_12565,N_12594);
nand U12695 (N_12695,N_12583,N_12573);
xnor U12696 (N_12696,N_12542,N_12467);
or U12697 (N_12697,N_12584,N_12513);
nand U12698 (N_12698,N_12492,N_12458);
nor U12699 (N_12699,N_12541,N_12562);
nand U12700 (N_12700,N_12544,N_12476);
and U12701 (N_12701,N_12580,N_12516);
nand U12702 (N_12702,N_12577,N_12481);
nor U12703 (N_12703,N_12477,N_12517);
nor U12704 (N_12704,N_12466,N_12451);
xor U12705 (N_12705,N_12465,N_12543);
nor U12706 (N_12706,N_12569,N_12487);
nand U12707 (N_12707,N_12468,N_12493);
nand U12708 (N_12708,N_12569,N_12464);
and U12709 (N_12709,N_12499,N_12528);
nand U12710 (N_12710,N_12454,N_12545);
and U12711 (N_12711,N_12484,N_12496);
nand U12712 (N_12712,N_12585,N_12581);
xor U12713 (N_12713,N_12517,N_12458);
and U12714 (N_12714,N_12498,N_12593);
nor U12715 (N_12715,N_12521,N_12518);
nor U12716 (N_12716,N_12564,N_12505);
and U12717 (N_12717,N_12544,N_12473);
nand U12718 (N_12718,N_12486,N_12489);
nand U12719 (N_12719,N_12596,N_12589);
and U12720 (N_12720,N_12509,N_12561);
nand U12721 (N_12721,N_12534,N_12496);
and U12722 (N_12722,N_12546,N_12466);
and U12723 (N_12723,N_12502,N_12491);
xnor U12724 (N_12724,N_12553,N_12480);
xor U12725 (N_12725,N_12558,N_12488);
nand U12726 (N_12726,N_12503,N_12517);
nor U12727 (N_12727,N_12467,N_12512);
xor U12728 (N_12728,N_12465,N_12574);
and U12729 (N_12729,N_12574,N_12594);
and U12730 (N_12730,N_12483,N_12526);
nand U12731 (N_12731,N_12523,N_12465);
nor U12732 (N_12732,N_12536,N_12469);
and U12733 (N_12733,N_12557,N_12453);
or U12734 (N_12734,N_12476,N_12484);
nor U12735 (N_12735,N_12469,N_12482);
nand U12736 (N_12736,N_12495,N_12515);
or U12737 (N_12737,N_12452,N_12546);
or U12738 (N_12738,N_12470,N_12542);
or U12739 (N_12739,N_12519,N_12539);
or U12740 (N_12740,N_12498,N_12499);
or U12741 (N_12741,N_12505,N_12511);
xnor U12742 (N_12742,N_12527,N_12510);
xnor U12743 (N_12743,N_12483,N_12477);
or U12744 (N_12744,N_12578,N_12523);
xnor U12745 (N_12745,N_12505,N_12552);
or U12746 (N_12746,N_12508,N_12574);
xnor U12747 (N_12747,N_12459,N_12569);
or U12748 (N_12748,N_12578,N_12536);
xnor U12749 (N_12749,N_12525,N_12465);
nand U12750 (N_12750,N_12749,N_12627);
and U12751 (N_12751,N_12636,N_12602);
nor U12752 (N_12752,N_12679,N_12666);
or U12753 (N_12753,N_12635,N_12641);
and U12754 (N_12754,N_12722,N_12659);
and U12755 (N_12755,N_12710,N_12611);
nor U12756 (N_12756,N_12681,N_12614);
and U12757 (N_12757,N_12733,N_12704);
xnor U12758 (N_12758,N_12654,N_12663);
and U12759 (N_12759,N_12615,N_12625);
nand U12760 (N_12760,N_12617,N_12739);
nor U12761 (N_12761,N_12737,N_12688);
nand U12762 (N_12762,N_12667,N_12683);
nor U12763 (N_12763,N_12656,N_12677);
nor U12764 (N_12764,N_12632,N_12622);
nand U12765 (N_12765,N_12670,N_12680);
xor U12766 (N_12766,N_12669,N_12660);
and U12767 (N_12767,N_12628,N_12673);
and U12768 (N_12768,N_12735,N_12716);
xnor U12769 (N_12769,N_12682,N_12706);
xor U12770 (N_12770,N_12631,N_12742);
nor U12771 (N_12771,N_12694,N_12606);
or U12772 (N_12772,N_12601,N_12637);
nand U12773 (N_12773,N_12623,N_12701);
nand U12774 (N_12774,N_12639,N_12674);
or U12775 (N_12775,N_12745,N_12638);
nand U12776 (N_12776,N_12652,N_12678);
or U12777 (N_12777,N_12715,N_12608);
nor U12778 (N_12778,N_12610,N_12721);
xnor U12779 (N_12779,N_12621,N_12668);
xnor U12780 (N_12780,N_12696,N_12643);
nand U12781 (N_12781,N_12714,N_12723);
and U12782 (N_12782,N_12671,N_12734);
nand U12783 (N_12783,N_12736,N_12703);
xnor U12784 (N_12784,N_12647,N_12743);
xnor U12785 (N_12785,N_12709,N_12740);
or U12786 (N_12786,N_12653,N_12729);
xnor U12787 (N_12787,N_12612,N_12690);
or U12788 (N_12788,N_12613,N_12619);
xor U12789 (N_12789,N_12665,N_12676);
and U12790 (N_12790,N_12747,N_12725);
nand U12791 (N_12791,N_12689,N_12720);
or U12792 (N_12792,N_12648,N_12616);
nor U12793 (N_12793,N_12717,N_12713);
xor U12794 (N_12794,N_12603,N_12630);
or U12795 (N_12795,N_12728,N_12726);
nor U12796 (N_12796,N_12711,N_12744);
nor U12797 (N_12797,N_12691,N_12732);
xor U12798 (N_12798,N_12708,N_12604);
or U12799 (N_12799,N_12664,N_12675);
and U12800 (N_12800,N_12730,N_12651);
and U12801 (N_12801,N_12657,N_12684);
and U12802 (N_12802,N_12646,N_12634);
nor U12803 (N_12803,N_12658,N_12697);
nor U12804 (N_12804,N_12633,N_12693);
nor U12805 (N_12805,N_12655,N_12609);
xor U12806 (N_12806,N_12738,N_12692);
or U12807 (N_12807,N_12605,N_12644);
nor U12808 (N_12808,N_12649,N_12662);
or U12809 (N_12809,N_12702,N_12642);
xor U12810 (N_12810,N_12724,N_12707);
xnor U12811 (N_12811,N_12727,N_12624);
and U12812 (N_12812,N_12607,N_12748);
nand U12813 (N_12813,N_12618,N_12705);
xnor U12814 (N_12814,N_12686,N_12687);
or U12815 (N_12815,N_12626,N_12718);
or U12816 (N_12816,N_12746,N_12712);
nor U12817 (N_12817,N_12640,N_12741);
nand U12818 (N_12818,N_12650,N_12672);
and U12819 (N_12819,N_12685,N_12731);
and U12820 (N_12820,N_12699,N_12661);
or U12821 (N_12821,N_12700,N_12719);
nand U12822 (N_12822,N_12629,N_12698);
xor U12823 (N_12823,N_12645,N_12695);
and U12824 (N_12824,N_12620,N_12600);
or U12825 (N_12825,N_12637,N_12728);
xnor U12826 (N_12826,N_12652,N_12613);
nor U12827 (N_12827,N_12614,N_12714);
or U12828 (N_12828,N_12749,N_12714);
and U12829 (N_12829,N_12707,N_12686);
xor U12830 (N_12830,N_12739,N_12665);
xor U12831 (N_12831,N_12678,N_12729);
or U12832 (N_12832,N_12614,N_12660);
nand U12833 (N_12833,N_12690,N_12699);
nand U12834 (N_12834,N_12697,N_12723);
xnor U12835 (N_12835,N_12650,N_12734);
nand U12836 (N_12836,N_12618,N_12697);
xor U12837 (N_12837,N_12674,N_12602);
or U12838 (N_12838,N_12692,N_12655);
nand U12839 (N_12839,N_12630,N_12606);
xor U12840 (N_12840,N_12742,N_12724);
xor U12841 (N_12841,N_12715,N_12697);
xor U12842 (N_12842,N_12615,N_12676);
xnor U12843 (N_12843,N_12675,N_12659);
and U12844 (N_12844,N_12730,N_12664);
xnor U12845 (N_12845,N_12747,N_12716);
or U12846 (N_12846,N_12640,N_12642);
nor U12847 (N_12847,N_12730,N_12706);
nand U12848 (N_12848,N_12718,N_12602);
nand U12849 (N_12849,N_12660,N_12687);
nor U12850 (N_12850,N_12719,N_12603);
nand U12851 (N_12851,N_12638,N_12604);
and U12852 (N_12852,N_12662,N_12745);
nand U12853 (N_12853,N_12628,N_12611);
and U12854 (N_12854,N_12692,N_12700);
and U12855 (N_12855,N_12711,N_12634);
nand U12856 (N_12856,N_12614,N_12662);
and U12857 (N_12857,N_12657,N_12676);
nor U12858 (N_12858,N_12675,N_12701);
or U12859 (N_12859,N_12635,N_12693);
or U12860 (N_12860,N_12665,N_12603);
and U12861 (N_12861,N_12706,N_12658);
nor U12862 (N_12862,N_12726,N_12659);
and U12863 (N_12863,N_12649,N_12722);
xnor U12864 (N_12864,N_12740,N_12747);
and U12865 (N_12865,N_12618,N_12698);
nand U12866 (N_12866,N_12727,N_12678);
or U12867 (N_12867,N_12700,N_12639);
nor U12868 (N_12868,N_12640,N_12643);
nand U12869 (N_12869,N_12709,N_12631);
or U12870 (N_12870,N_12635,N_12723);
nor U12871 (N_12871,N_12612,N_12675);
xnor U12872 (N_12872,N_12670,N_12745);
nand U12873 (N_12873,N_12711,N_12679);
nand U12874 (N_12874,N_12658,N_12714);
nor U12875 (N_12875,N_12600,N_12714);
and U12876 (N_12876,N_12734,N_12600);
nor U12877 (N_12877,N_12615,N_12645);
xnor U12878 (N_12878,N_12637,N_12685);
and U12879 (N_12879,N_12657,N_12733);
nand U12880 (N_12880,N_12724,N_12614);
nand U12881 (N_12881,N_12713,N_12745);
xnor U12882 (N_12882,N_12659,N_12740);
nor U12883 (N_12883,N_12672,N_12691);
nor U12884 (N_12884,N_12707,N_12671);
or U12885 (N_12885,N_12691,N_12685);
nor U12886 (N_12886,N_12604,N_12678);
nor U12887 (N_12887,N_12710,N_12730);
or U12888 (N_12888,N_12693,N_12617);
nor U12889 (N_12889,N_12735,N_12646);
or U12890 (N_12890,N_12657,N_12736);
or U12891 (N_12891,N_12659,N_12703);
and U12892 (N_12892,N_12638,N_12681);
xor U12893 (N_12893,N_12645,N_12613);
or U12894 (N_12894,N_12649,N_12602);
or U12895 (N_12895,N_12619,N_12728);
or U12896 (N_12896,N_12725,N_12661);
nand U12897 (N_12897,N_12703,N_12699);
and U12898 (N_12898,N_12656,N_12626);
or U12899 (N_12899,N_12718,N_12652);
nand U12900 (N_12900,N_12885,N_12798);
nand U12901 (N_12901,N_12837,N_12768);
nand U12902 (N_12902,N_12751,N_12802);
or U12903 (N_12903,N_12832,N_12822);
nand U12904 (N_12904,N_12894,N_12772);
xnor U12905 (N_12905,N_12897,N_12783);
nand U12906 (N_12906,N_12807,N_12784);
nor U12907 (N_12907,N_12826,N_12834);
or U12908 (N_12908,N_12895,N_12818);
or U12909 (N_12909,N_12876,N_12759);
and U12910 (N_12910,N_12854,N_12849);
nor U12911 (N_12911,N_12753,N_12887);
xnor U12912 (N_12912,N_12874,N_12760);
nor U12913 (N_12913,N_12840,N_12812);
nand U12914 (N_12914,N_12757,N_12843);
xor U12915 (N_12915,N_12884,N_12820);
xnor U12916 (N_12916,N_12765,N_12755);
xor U12917 (N_12917,N_12841,N_12786);
and U12918 (N_12918,N_12814,N_12882);
or U12919 (N_12919,N_12782,N_12819);
nand U12920 (N_12920,N_12808,N_12867);
and U12921 (N_12921,N_12830,N_12764);
xor U12922 (N_12922,N_12756,N_12868);
nand U12923 (N_12923,N_12898,N_12796);
and U12924 (N_12924,N_12869,N_12865);
nor U12925 (N_12925,N_12870,N_12770);
nand U12926 (N_12926,N_12766,N_12758);
xnor U12927 (N_12927,N_12763,N_12853);
nor U12928 (N_12928,N_12776,N_12813);
nand U12929 (N_12929,N_12785,N_12821);
nand U12930 (N_12930,N_12892,N_12899);
or U12931 (N_12931,N_12888,N_12815);
xnor U12932 (N_12932,N_12788,N_12787);
nand U12933 (N_12933,N_12825,N_12848);
xnor U12934 (N_12934,N_12752,N_12875);
xor U12935 (N_12935,N_12890,N_12835);
xnor U12936 (N_12936,N_12789,N_12817);
or U12937 (N_12937,N_12833,N_12851);
nand U12938 (N_12938,N_12855,N_12880);
nand U12939 (N_12939,N_12852,N_12891);
nand U12940 (N_12940,N_12750,N_12779);
xnor U12941 (N_12941,N_12836,N_12803);
and U12942 (N_12942,N_12767,N_12778);
or U12943 (N_12943,N_12777,N_12842);
nor U12944 (N_12944,N_12774,N_12864);
nand U12945 (N_12945,N_12847,N_12797);
and U12946 (N_12946,N_12791,N_12861);
nor U12947 (N_12947,N_12754,N_12863);
or U12948 (N_12948,N_12889,N_12775);
and U12949 (N_12949,N_12856,N_12883);
or U12950 (N_12950,N_12800,N_12877);
and U12951 (N_12951,N_12804,N_12860);
nor U12952 (N_12952,N_12773,N_12858);
xnor U12953 (N_12953,N_12793,N_12806);
nand U12954 (N_12954,N_12871,N_12771);
or U12955 (N_12955,N_12801,N_12886);
nor U12956 (N_12956,N_12829,N_12823);
or U12957 (N_12957,N_12790,N_12792);
xor U12958 (N_12958,N_12873,N_12831);
and U12959 (N_12959,N_12799,N_12810);
or U12960 (N_12960,N_12846,N_12795);
xnor U12961 (N_12961,N_12809,N_12794);
or U12962 (N_12962,N_12762,N_12828);
and U12963 (N_12963,N_12845,N_12872);
xnor U12964 (N_12964,N_12881,N_12780);
or U12965 (N_12965,N_12824,N_12805);
nand U12966 (N_12966,N_12850,N_12816);
xnor U12967 (N_12967,N_12761,N_12839);
nand U12968 (N_12968,N_12827,N_12878);
or U12969 (N_12969,N_12879,N_12859);
xnor U12970 (N_12970,N_12838,N_12811);
xnor U12971 (N_12971,N_12862,N_12893);
xnor U12972 (N_12972,N_12896,N_12781);
xor U12973 (N_12973,N_12769,N_12857);
nand U12974 (N_12974,N_12866,N_12844);
xor U12975 (N_12975,N_12825,N_12766);
nand U12976 (N_12976,N_12772,N_12797);
nand U12977 (N_12977,N_12765,N_12752);
nor U12978 (N_12978,N_12858,N_12783);
and U12979 (N_12979,N_12772,N_12861);
nor U12980 (N_12980,N_12896,N_12838);
and U12981 (N_12981,N_12770,N_12856);
or U12982 (N_12982,N_12882,N_12768);
nor U12983 (N_12983,N_12878,N_12765);
and U12984 (N_12984,N_12751,N_12836);
nand U12985 (N_12985,N_12754,N_12843);
and U12986 (N_12986,N_12871,N_12870);
xor U12987 (N_12987,N_12763,N_12795);
xnor U12988 (N_12988,N_12855,N_12845);
and U12989 (N_12989,N_12756,N_12768);
or U12990 (N_12990,N_12876,N_12881);
or U12991 (N_12991,N_12811,N_12752);
or U12992 (N_12992,N_12869,N_12755);
nor U12993 (N_12993,N_12776,N_12807);
or U12994 (N_12994,N_12830,N_12825);
nand U12995 (N_12995,N_12780,N_12751);
xnor U12996 (N_12996,N_12874,N_12859);
or U12997 (N_12997,N_12750,N_12892);
and U12998 (N_12998,N_12798,N_12823);
nand U12999 (N_12999,N_12800,N_12801);
xnor U13000 (N_13000,N_12750,N_12855);
xnor U13001 (N_13001,N_12890,N_12866);
or U13002 (N_13002,N_12862,N_12871);
nor U13003 (N_13003,N_12790,N_12767);
nand U13004 (N_13004,N_12825,N_12792);
xnor U13005 (N_13005,N_12874,N_12818);
xnor U13006 (N_13006,N_12868,N_12825);
xnor U13007 (N_13007,N_12839,N_12774);
nand U13008 (N_13008,N_12882,N_12848);
nand U13009 (N_13009,N_12809,N_12795);
or U13010 (N_13010,N_12836,N_12816);
xor U13011 (N_13011,N_12796,N_12811);
nor U13012 (N_13012,N_12836,N_12848);
and U13013 (N_13013,N_12755,N_12867);
or U13014 (N_13014,N_12837,N_12895);
nor U13015 (N_13015,N_12818,N_12821);
nor U13016 (N_13016,N_12780,N_12771);
xor U13017 (N_13017,N_12777,N_12873);
xor U13018 (N_13018,N_12834,N_12882);
nor U13019 (N_13019,N_12869,N_12886);
nand U13020 (N_13020,N_12786,N_12819);
nand U13021 (N_13021,N_12827,N_12887);
nor U13022 (N_13022,N_12874,N_12789);
or U13023 (N_13023,N_12768,N_12857);
nand U13024 (N_13024,N_12880,N_12877);
or U13025 (N_13025,N_12799,N_12874);
nor U13026 (N_13026,N_12864,N_12802);
or U13027 (N_13027,N_12809,N_12880);
nand U13028 (N_13028,N_12819,N_12894);
nand U13029 (N_13029,N_12895,N_12822);
or U13030 (N_13030,N_12803,N_12847);
and U13031 (N_13031,N_12760,N_12755);
xnor U13032 (N_13032,N_12851,N_12814);
nand U13033 (N_13033,N_12889,N_12811);
nor U13034 (N_13034,N_12840,N_12804);
nor U13035 (N_13035,N_12752,N_12881);
xnor U13036 (N_13036,N_12862,N_12784);
nor U13037 (N_13037,N_12815,N_12772);
nor U13038 (N_13038,N_12789,N_12773);
nor U13039 (N_13039,N_12898,N_12773);
nor U13040 (N_13040,N_12753,N_12824);
and U13041 (N_13041,N_12795,N_12899);
nor U13042 (N_13042,N_12754,N_12787);
xnor U13043 (N_13043,N_12869,N_12752);
xnor U13044 (N_13044,N_12805,N_12840);
nand U13045 (N_13045,N_12899,N_12779);
xnor U13046 (N_13046,N_12858,N_12849);
nand U13047 (N_13047,N_12846,N_12784);
or U13048 (N_13048,N_12782,N_12854);
xor U13049 (N_13049,N_12885,N_12838);
xnor U13050 (N_13050,N_12949,N_12959);
and U13051 (N_13051,N_12948,N_12932);
and U13052 (N_13052,N_13012,N_12905);
or U13053 (N_13053,N_12940,N_12922);
nand U13054 (N_13054,N_12986,N_12909);
or U13055 (N_13055,N_12925,N_13048);
xnor U13056 (N_13056,N_12979,N_13038);
nor U13057 (N_13057,N_13034,N_13020);
xnor U13058 (N_13058,N_13007,N_13037);
nor U13059 (N_13059,N_13035,N_12964);
and U13060 (N_13060,N_13049,N_12966);
xnor U13061 (N_13061,N_13029,N_12911);
or U13062 (N_13062,N_12950,N_13045);
nand U13063 (N_13063,N_12912,N_13043);
nand U13064 (N_13064,N_12938,N_13027);
and U13065 (N_13065,N_13018,N_12963);
nand U13066 (N_13066,N_12985,N_12976);
and U13067 (N_13067,N_13015,N_12998);
or U13068 (N_13068,N_12980,N_12951);
nand U13069 (N_13069,N_13016,N_12996);
nand U13070 (N_13070,N_12920,N_12945);
nor U13071 (N_13071,N_12946,N_12943);
xnor U13072 (N_13072,N_13047,N_12958);
or U13073 (N_13073,N_12960,N_12982);
xnor U13074 (N_13074,N_12901,N_13000);
and U13075 (N_13075,N_12962,N_12990);
nand U13076 (N_13076,N_13031,N_12965);
nand U13077 (N_13077,N_13028,N_13041);
nand U13078 (N_13078,N_13005,N_12937);
and U13079 (N_13079,N_13022,N_13023);
or U13080 (N_13080,N_12910,N_13004);
and U13081 (N_13081,N_12917,N_12955);
and U13082 (N_13082,N_13001,N_13039);
xor U13083 (N_13083,N_13026,N_12921);
nand U13084 (N_13084,N_12995,N_12947);
or U13085 (N_13085,N_13002,N_12939);
nand U13086 (N_13086,N_13040,N_12993);
xor U13087 (N_13087,N_12942,N_12929);
nand U13088 (N_13088,N_13032,N_12944);
nand U13089 (N_13089,N_12935,N_12904);
xnor U13090 (N_13090,N_12928,N_12997);
or U13091 (N_13091,N_12975,N_12903);
and U13092 (N_13092,N_12908,N_13003);
xor U13093 (N_13093,N_12907,N_12914);
or U13094 (N_13094,N_12926,N_12900);
and U13095 (N_13095,N_13036,N_12973);
nor U13096 (N_13096,N_12931,N_12927);
xnor U13097 (N_13097,N_12930,N_13046);
nor U13098 (N_13098,N_12934,N_12924);
nor U13099 (N_13099,N_12992,N_12936);
and U13100 (N_13100,N_13009,N_12915);
and U13101 (N_13101,N_12978,N_12918);
or U13102 (N_13102,N_12961,N_13021);
nand U13103 (N_13103,N_12954,N_13025);
nor U13104 (N_13104,N_13006,N_12977);
and U13105 (N_13105,N_13019,N_12981);
nand U13106 (N_13106,N_12972,N_12969);
nor U13107 (N_13107,N_12906,N_13033);
xnor U13108 (N_13108,N_12974,N_12967);
xor U13109 (N_13109,N_13014,N_13017);
nor U13110 (N_13110,N_12956,N_12983);
nand U13111 (N_13111,N_13011,N_12902);
and U13112 (N_13112,N_12988,N_12984);
nor U13113 (N_13113,N_12994,N_12987);
or U13114 (N_13114,N_12919,N_12989);
and U13115 (N_13115,N_12991,N_12913);
xor U13116 (N_13116,N_13013,N_12952);
nand U13117 (N_13117,N_12971,N_13024);
nand U13118 (N_13118,N_13042,N_12933);
nor U13119 (N_13119,N_12970,N_12916);
nand U13120 (N_13120,N_12953,N_13008);
nand U13121 (N_13121,N_12999,N_13030);
or U13122 (N_13122,N_12957,N_13010);
xnor U13123 (N_13123,N_12968,N_13044);
or U13124 (N_13124,N_12941,N_12923);
and U13125 (N_13125,N_13021,N_12914);
nor U13126 (N_13126,N_12914,N_12993);
nand U13127 (N_13127,N_12932,N_12994);
or U13128 (N_13128,N_12918,N_12981);
or U13129 (N_13129,N_13018,N_12966);
and U13130 (N_13130,N_12977,N_12953);
or U13131 (N_13131,N_12931,N_12995);
nor U13132 (N_13132,N_12948,N_12955);
nor U13133 (N_13133,N_12993,N_12959);
and U13134 (N_13134,N_12961,N_12992);
nand U13135 (N_13135,N_12926,N_12948);
xnor U13136 (N_13136,N_12999,N_12912);
and U13137 (N_13137,N_12960,N_12980);
xnor U13138 (N_13138,N_12959,N_12902);
and U13139 (N_13139,N_12975,N_13040);
xor U13140 (N_13140,N_12966,N_13029);
xor U13141 (N_13141,N_13001,N_12995);
nor U13142 (N_13142,N_13008,N_12958);
nor U13143 (N_13143,N_12976,N_13032);
or U13144 (N_13144,N_13035,N_12966);
nand U13145 (N_13145,N_12979,N_13043);
and U13146 (N_13146,N_13037,N_12974);
and U13147 (N_13147,N_12965,N_12904);
xnor U13148 (N_13148,N_13031,N_12905);
and U13149 (N_13149,N_13044,N_12970);
nand U13150 (N_13150,N_13047,N_13023);
nor U13151 (N_13151,N_12940,N_13036);
nand U13152 (N_13152,N_12943,N_12967);
nor U13153 (N_13153,N_13028,N_13043);
and U13154 (N_13154,N_12904,N_12931);
nor U13155 (N_13155,N_12932,N_12936);
or U13156 (N_13156,N_12968,N_13001);
nand U13157 (N_13157,N_12901,N_12903);
xnor U13158 (N_13158,N_12979,N_13031);
or U13159 (N_13159,N_12908,N_12977);
or U13160 (N_13160,N_12926,N_12951);
nand U13161 (N_13161,N_13012,N_12998);
xnor U13162 (N_13162,N_13035,N_12943);
xor U13163 (N_13163,N_12909,N_12956);
nand U13164 (N_13164,N_13025,N_13001);
nand U13165 (N_13165,N_13044,N_13003);
and U13166 (N_13166,N_13015,N_12987);
or U13167 (N_13167,N_12930,N_12952);
xnor U13168 (N_13168,N_12904,N_13014);
nor U13169 (N_13169,N_12975,N_13027);
nor U13170 (N_13170,N_12960,N_12969);
nand U13171 (N_13171,N_13048,N_12931);
nand U13172 (N_13172,N_12938,N_13011);
or U13173 (N_13173,N_13002,N_12955);
and U13174 (N_13174,N_12959,N_12974);
xor U13175 (N_13175,N_13048,N_13030);
or U13176 (N_13176,N_12910,N_12953);
or U13177 (N_13177,N_12912,N_13029);
and U13178 (N_13178,N_12921,N_12906);
or U13179 (N_13179,N_13002,N_13020);
nor U13180 (N_13180,N_13035,N_12921);
nand U13181 (N_13181,N_13032,N_12950);
nor U13182 (N_13182,N_12905,N_12973);
or U13183 (N_13183,N_12983,N_12982);
xnor U13184 (N_13184,N_13008,N_12905);
or U13185 (N_13185,N_13044,N_13030);
xor U13186 (N_13186,N_13014,N_12994);
nor U13187 (N_13187,N_12909,N_13026);
xor U13188 (N_13188,N_13025,N_13000);
nor U13189 (N_13189,N_12904,N_12959);
nor U13190 (N_13190,N_13036,N_12991);
nor U13191 (N_13191,N_13000,N_12934);
nand U13192 (N_13192,N_13035,N_12933);
xnor U13193 (N_13193,N_12963,N_12973);
xnor U13194 (N_13194,N_12954,N_12985);
nor U13195 (N_13195,N_12922,N_12928);
or U13196 (N_13196,N_12980,N_13029);
or U13197 (N_13197,N_13018,N_13011);
nor U13198 (N_13198,N_13031,N_12935);
nand U13199 (N_13199,N_12981,N_13044);
xnor U13200 (N_13200,N_13127,N_13161);
or U13201 (N_13201,N_13108,N_13198);
or U13202 (N_13202,N_13163,N_13117);
or U13203 (N_13203,N_13164,N_13134);
and U13204 (N_13204,N_13133,N_13146);
or U13205 (N_13205,N_13082,N_13067);
and U13206 (N_13206,N_13130,N_13055);
nand U13207 (N_13207,N_13183,N_13083);
nand U13208 (N_13208,N_13195,N_13053);
or U13209 (N_13209,N_13096,N_13184);
xor U13210 (N_13210,N_13078,N_13116);
nand U13211 (N_13211,N_13187,N_13099);
xnor U13212 (N_13212,N_13160,N_13132);
xnor U13213 (N_13213,N_13137,N_13106);
nor U13214 (N_13214,N_13169,N_13176);
and U13215 (N_13215,N_13181,N_13077);
xor U13216 (N_13216,N_13170,N_13168);
or U13217 (N_13217,N_13052,N_13136);
nor U13218 (N_13218,N_13050,N_13126);
or U13219 (N_13219,N_13144,N_13063);
nor U13220 (N_13220,N_13121,N_13084);
nand U13221 (N_13221,N_13149,N_13167);
nor U13222 (N_13222,N_13115,N_13141);
or U13223 (N_13223,N_13089,N_13192);
and U13224 (N_13224,N_13186,N_13062);
xnor U13225 (N_13225,N_13085,N_13147);
nand U13226 (N_13226,N_13102,N_13175);
or U13227 (N_13227,N_13190,N_13113);
nand U13228 (N_13228,N_13171,N_13079);
or U13229 (N_13229,N_13092,N_13066);
xor U13230 (N_13230,N_13093,N_13140);
nor U13231 (N_13231,N_13185,N_13142);
xnor U13232 (N_13232,N_13135,N_13087);
nor U13233 (N_13233,N_13097,N_13120);
nor U13234 (N_13234,N_13151,N_13157);
xor U13235 (N_13235,N_13155,N_13060);
nand U13236 (N_13236,N_13124,N_13178);
xnor U13237 (N_13237,N_13061,N_13103);
or U13238 (N_13238,N_13174,N_13112);
or U13239 (N_13239,N_13158,N_13098);
nor U13240 (N_13240,N_13086,N_13191);
nor U13241 (N_13241,N_13177,N_13091);
and U13242 (N_13242,N_13156,N_13165);
nand U13243 (N_13243,N_13145,N_13166);
nand U13244 (N_13244,N_13114,N_13090);
nor U13245 (N_13245,N_13069,N_13095);
and U13246 (N_13246,N_13122,N_13076);
and U13247 (N_13247,N_13159,N_13162);
nor U13248 (N_13248,N_13125,N_13197);
nand U13249 (N_13249,N_13110,N_13104);
nor U13250 (N_13250,N_13080,N_13094);
and U13251 (N_13251,N_13109,N_13129);
nor U13252 (N_13252,N_13070,N_13199);
and U13253 (N_13253,N_13107,N_13073);
and U13254 (N_13254,N_13100,N_13064);
nand U13255 (N_13255,N_13189,N_13138);
and U13256 (N_13256,N_13059,N_13057);
or U13257 (N_13257,N_13182,N_13071);
xnor U13258 (N_13258,N_13154,N_13196);
nor U13259 (N_13259,N_13118,N_13051);
nor U13260 (N_13260,N_13180,N_13131);
and U13261 (N_13261,N_13074,N_13143);
xnor U13262 (N_13262,N_13072,N_13188);
nand U13263 (N_13263,N_13065,N_13123);
xnor U13264 (N_13264,N_13088,N_13101);
and U13265 (N_13265,N_13173,N_13148);
and U13266 (N_13266,N_13111,N_13081);
nor U13267 (N_13267,N_13075,N_13193);
nand U13268 (N_13268,N_13054,N_13150);
and U13269 (N_13269,N_13068,N_13105);
or U13270 (N_13270,N_13194,N_13139);
or U13271 (N_13271,N_13179,N_13153);
and U13272 (N_13272,N_13152,N_13172);
nor U13273 (N_13273,N_13056,N_13128);
or U13274 (N_13274,N_13058,N_13119);
nand U13275 (N_13275,N_13121,N_13051);
nor U13276 (N_13276,N_13173,N_13127);
or U13277 (N_13277,N_13134,N_13075);
nor U13278 (N_13278,N_13086,N_13161);
nor U13279 (N_13279,N_13091,N_13149);
nand U13280 (N_13280,N_13196,N_13060);
and U13281 (N_13281,N_13135,N_13156);
nor U13282 (N_13282,N_13165,N_13180);
xnor U13283 (N_13283,N_13166,N_13194);
and U13284 (N_13284,N_13090,N_13104);
and U13285 (N_13285,N_13096,N_13094);
nor U13286 (N_13286,N_13198,N_13144);
nand U13287 (N_13287,N_13082,N_13083);
nor U13288 (N_13288,N_13168,N_13084);
nor U13289 (N_13289,N_13096,N_13100);
nand U13290 (N_13290,N_13184,N_13139);
xnor U13291 (N_13291,N_13050,N_13096);
nand U13292 (N_13292,N_13104,N_13116);
nand U13293 (N_13293,N_13155,N_13183);
nand U13294 (N_13294,N_13052,N_13189);
nor U13295 (N_13295,N_13176,N_13134);
and U13296 (N_13296,N_13078,N_13178);
nor U13297 (N_13297,N_13093,N_13183);
nand U13298 (N_13298,N_13065,N_13163);
xor U13299 (N_13299,N_13150,N_13050);
xnor U13300 (N_13300,N_13052,N_13181);
nand U13301 (N_13301,N_13154,N_13147);
and U13302 (N_13302,N_13102,N_13070);
or U13303 (N_13303,N_13180,N_13168);
nor U13304 (N_13304,N_13162,N_13061);
nor U13305 (N_13305,N_13174,N_13156);
nand U13306 (N_13306,N_13099,N_13053);
and U13307 (N_13307,N_13153,N_13050);
nand U13308 (N_13308,N_13095,N_13177);
nor U13309 (N_13309,N_13100,N_13147);
nand U13310 (N_13310,N_13050,N_13102);
or U13311 (N_13311,N_13065,N_13088);
or U13312 (N_13312,N_13079,N_13167);
and U13313 (N_13313,N_13133,N_13140);
or U13314 (N_13314,N_13109,N_13062);
or U13315 (N_13315,N_13118,N_13194);
xnor U13316 (N_13316,N_13138,N_13157);
nor U13317 (N_13317,N_13126,N_13081);
nand U13318 (N_13318,N_13155,N_13107);
or U13319 (N_13319,N_13126,N_13171);
and U13320 (N_13320,N_13085,N_13198);
xor U13321 (N_13321,N_13165,N_13050);
nor U13322 (N_13322,N_13157,N_13086);
and U13323 (N_13323,N_13133,N_13120);
nand U13324 (N_13324,N_13164,N_13104);
xnor U13325 (N_13325,N_13072,N_13092);
and U13326 (N_13326,N_13149,N_13081);
xnor U13327 (N_13327,N_13084,N_13055);
nand U13328 (N_13328,N_13059,N_13165);
nor U13329 (N_13329,N_13076,N_13126);
nor U13330 (N_13330,N_13131,N_13063);
and U13331 (N_13331,N_13194,N_13107);
and U13332 (N_13332,N_13080,N_13076);
and U13333 (N_13333,N_13142,N_13137);
xor U13334 (N_13334,N_13157,N_13097);
xnor U13335 (N_13335,N_13157,N_13127);
nand U13336 (N_13336,N_13168,N_13183);
xnor U13337 (N_13337,N_13168,N_13179);
or U13338 (N_13338,N_13072,N_13152);
and U13339 (N_13339,N_13136,N_13114);
xor U13340 (N_13340,N_13101,N_13160);
or U13341 (N_13341,N_13161,N_13124);
nand U13342 (N_13342,N_13079,N_13132);
nor U13343 (N_13343,N_13068,N_13079);
nor U13344 (N_13344,N_13182,N_13192);
and U13345 (N_13345,N_13162,N_13168);
nor U13346 (N_13346,N_13181,N_13129);
xnor U13347 (N_13347,N_13188,N_13191);
nor U13348 (N_13348,N_13089,N_13170);
and U13349 (N_13349,N_13175,N_13079);
nor U13350 (N_13350,N_13318,N_13277);
xnor U13351 (N_13351,N_13317,N_13319);
and U13352 (N_13352,N_13262,N_13344);
or U13353 (N_13353,N_13330,N_13289);
nor U13354 (N_13354,N_13327,N_13297);
or U13355 (N_13355,N_13258,N_13234);
and U13356 (N_13356,N_13214,N_13211);
or U13357 (N_13357,N_13250,N_13310);
nor U13358 (N_13358,N_13298,N_13336);
nand U13359 (N_13359,N_13240,N_13229);
or U13360 (N_13360,N_13343,N_13328);
xor U13361 (N_13361,N_13293,N_13307);
or U13362 (N_13362,N_13206,N_13255);
nor U13363 (N_13363,N_13228,N_13221);
nand U13364 (N_13364,N_13236,N_13210);
or U13365 (N_13365,N_13216,N_13225);
nor U13366 (N_13366,N_13347,N_13275);
xnor U13367 (N_13367,N_13242,N_13268);
nor U13368 (N_13368,N_13282,N_13299);
nand U13369 (N_13369,N_13323,N_13270);
xnor U13370 (N_13370,N_13278,N_13271);
xnor U13371 (N_13371,N_13230,N_13348);
and U13372 (N_13372,N_13224,N_13254);
or U13373 (N_13373,N_13219,N_13266);
xor U13374 (N_13374,N_13204,N_13263);
and U13375 (N_13375,N_13265,N_13260);
nor U13376 (N_13376,N_13329,N_13200);
or U13377 (N_13377,N_13202,N_13283);
and U13378 (N_13378,N_13291,N_13207);
or U13379 (N_13379,N_13295,N_13340);
and U13380 (N_13380,N_13239,N_13303);
and U13381 (N_13381,N_13209,N_13290);
xnor U13382 (N_13382,N_13201,N_13222);
or U13383 (N_13383,N_13237,N_13212);
and U13384 (N_13384,N_13247,N_13244);
or U13385 (N_13385,N_13304,N_13346);
and U13386 (N_13386,N_13243,N_13312);
xor U13387 (N_13387,N_13321,N_13253);
and U13388 (N_13388,N_13223,N_13241);
nand U13389 (N_13389,N_13300,N_13339);
xnor U13390 (N_13390,N_13285,N_13203);
nand U13391 (N_13391,N_13337,N_13231);
xor U13392 (N_13392,N_13256,N_13316);
xnor U13393 (N_13393,N_13334,N_13233);
or U13394 (N_13394,N_13306,N_13284);
nand U13395 (N_13395,N_13309,N_13322);
xnor U13396 (N_13396,N_13311,N_13314);
and U13397 (N_13397,N_13287,N_13248);
nand U13398 (N_13398,N_13269,N_13217);
nand U13399 (N_13399,N_13215,N_13259);
and U13400 (N_13400,N_13338,N_13341);
or U13401 (N_13401,N_13325,N_13245);
nand U13402 (N_13402,N_13274,N_13235);
nand U13403 (N_13403,N_13281,N_13331);
nand U13404 (N_13404,N_13301,N_13315);
nand U13405 (N_13405,N_13320,N_13273);
nand U13406 (N_13406,N_13246,N_13335);
nor U13407 (N_13407,N_13249,N_13261);
or U13408 (N_13408,N_13342,N_13349);
xnor U13409 (N_13409,N_13332,N_13305);
nand U13410 (N_13410,N_13302,N_13308);
nor U13411 (N_13411,N_13296,N_13294);
or U13412 (N_13412,N_13208,N_13252);
and U13413 (N_13413,N_13326,N_13313);
or U13414 (N_13414,N_13205,N_13324);
or U13415 (N_13415,N_13218,N_13232);
and U13416 (N_13416,N_13257,N_13292);
nor U13417 (N_13417,N_13280,N_13227);
nand U13418 (N_13418,N_13286,N_13333);
and U13419 (N_13419,N_13226,N_13238);
nor U13420 (N_13420,N_13276,N_13220);
or U13421 (N_13421,N_13288,N_13267);
xor U13422 (N_13422,N_13272,N_13345);
nor U13423 (N_13423,N_13264,N_13213);
nand U13424 (N_13424,N_13251,N_13279);
nand U13425 (N_13425,N_13319,N_13219);
nand U13426 (N_13426,N_13271,N_13226);
or U13427 (N_13427,N_13261,N_13327);
and U13428 (N_13428,N_13319,N_13208);
and U13429 (N_13429,N_13224,N_13243);
nand U13430 (N_13430,N_13290,N_13295);
xor U13431 (N_13431,N_13228,N_13303);
nand U13432 (N_13432,N_13256,N_13236);
or U13433 (N_13433,N_13334,N_13336);
nor U13434 (N_13434,N_13224,N_13225);
xnor U13435 (N_13435,N_13344,N_13283);
xnor U13436 (N_13436,N_13330,N_13309);
xnor U13437 (N_13437,N_13303,N_13261);
or U13438 (N_13438,N_13251,N_13249);
xor U13439 (N_13439,N_13224,N_13282);
or U13440 (N_13440,N_13264,N_13205);
nor U13441 (N_13441,N_13234,N_13319);
nor U13442 (N_13442,N_13255,N_13346);
and U13443 (N_13443,N_13346,N_13256);
xnor U13444 (N_13444,N_13300,N_13293);
xor U13445 (N_13445,N_13316,N_13289);
xnor U13446 (N_13446,N_13305,N_13238);
or U13447 (N_13447,N_13290,N_13289);
and U13448 (N_13448,N_13336,N_13348);
nand U13449 (N_13449,N_13212,N_13338);
xnor U13450 (N_13450,N_13282,N_13271);
nand U13451 (N_13451,N_13331,N_13210);
nand U13452 (N_13452,N_13280,N_13328);
xor U13453 (N_13453,N_13250,N_13206);
and U13454 (N_13454,N_13314,N_13263);
nand U13455 (N_13455,N_13273,N_13310);
nor U13456 (N_13456,N_13276,N_13248);
xnor U13457 (N_13457,N_13335,N_13205);
and U13458 (N_13458,N_13249,N_13305);
nor U13459 (N_13459,N_13284,N_13231);
nand U13460 (N_13460,N_13269,N_13310);
and U13461 (N_13461,N_13312,N_13237);
nor U13462 (N_13462,N_13204,N_13312);
or U13463 (N_13463,N_13202,N_13304);
nor U13464 (N_13464,N_13315,N_13269);
nor U13465 (N_13465,N_13294,N_13283);
nor U13466 (N_13466,N_13288,N_13225);
nand U13467 (N_13467,N_13312,N_13233);
nor U13468 (N_13468,N_13344,N_13290);
nor U13469 (N_13469,N_13203,N_13214);
or U13470 (N_13470,N_13284,N_13223);
nand U13471 (N_13471,N_13344,N_13336);
or U13472 (N_13472,N_13243,N_13261);
nor U13473 (N_13473,N_13232,N_13238);
or U13474 (N_13474,N_13314,N_13255);
nor U13475 (N_13475,N_13203,N_13297);
and U13476 (N_13476,N_13225,N_13274);
nand U13477 (N_13477,N_13249,N_13307);
nand U13478 (N_13478,N_13276,N_13262);
or U13479 (N_13479,N_13250,N_13323);
xnor U13480 (N_13480,N_13206,N_13201);
nor U13481 (N_13481,N_13262,N_13315);
xnor U13482 (N_13482,N_13255,N_13318);
and U13483 (N_13483,N_13342,N_13321);
nand U13484 (N_13484,N_13331,N_13301);
or U13485 (N_13485,N_13316,N_13315);
or U13486 (N_13486,N_13286,N_13290);
nand U13487 (N_13487,N_13346,N_13234);
and U13488 (N_13488,N_13323,N_13260);
or U13489 (N_13489,N_13278,N_13262);
nor U13490 (N_13490,N_13259,N_13289);
or U13491 (N_13491,N_13267,N_13296);
nor U13492 (N_13492,N_13202,N_13221);
and U13493 (N_13493,N_13202,N_13294);
nand U13494 (N_13494,N_13319,N_13258);
nand U13495 (N_13495,N_13287,N_13265);
nor U13496 (N_13496,N_13323,N_13246);
nor U13497 (N_13497,N_13273,N_13337);
nor U13498 (N_13498,N_13285,N_13230);
nor U13499 (N_13499,N_13262,N_13336);
and U13500 (N_13500,N_13393,N_13378);
xnor U13501 (N_13501,N_13400,N_13496);
and U13502 (N_13502,N_13491,N_13368);
xnor U13503 (N_13503,N_13359,N_13433);
nand U13504 (N_13504,N_13461,N_13424);
xor U13505 (N_13505,N_13481,N_13390);
nand U13506 (N_13506,N_13467,N_13463);
nand U13507 (N_13507,N_13401,N_13466);
xor U13508 (N_13508,N_13438,N_13361);
xnor U13509 (N_13509,N_13372,N_13404);
and U13510 (N_13510,N_13499,N_13374);
nor U13511 (N_13511,N_13470,N_13354);
nand U13512 (N_13512,N_13462,N_13385);
xnor U13513 (N_13513,N_13441,N_13488);
xor U13514 (N_13514,N_13376,N_13408);
or U13515 (N_13515,N_13432,N_13373);
or U13516 (N_13516,N_13449,N_13490);
and U13517 (N_13517,N_13483,N_13495);
xnor U13518 (N_13518,N_13356,N_13451);
nor U13519 (N_13519,N_13497,N_13492);
xnor U13520 (N_13520,N_13362,N_13429);
or U13521 (N_13521,N_13428,N_13389);
nor U13522 (N_13522,N_13425,N_13369);
or U13523 (N_13523,N_13448,N_13444);
nand U13524 (N_13524,N_13382,N_13353);
nor U13525 (N_13525,N_13399,N_13403);
and U13526 (N_13526,N_13405,N_13468);
xor U13527 (N_13527,N_13445,N_13427);
xnor U13528 (N_13528,N_13366,N_13419);
and U13529 (N_13529,N_13406,N_13358);
nor U13530 (N_13530,N_13457,N_13409);
nor U13531 (N_13531,N_13380,N_13471);
or U13532 (N_13532,N_13450,N_13446);
and U13533 (N_13533,N_13453,N_13398);
nand U13534 (N_13534,N_13485,N_13482);
nor U13535 (N_13535,N_13421,N_13402);
nor U13536 (N_13536,N_13469,N_13435);
nand U13537 (N_13537,N_13434,N_13377);
or U13538 (N_13538,N_13413,N_13464);
nand U13539 (N_13539,N_13375,N_13426);
nor U13540 (N_13540,N_13360,N_13414);
nor U13541 (N_13541,N_13364,N_13477);
or U13542 (N_13542,N_13420,N_13476);
nor U13543 (N_13543,N_13365,N_13447);
xnor U13544 (N_13544,N_13478,N_13473);
or U13545 (N_13545,N_13394,N_13392);
xor U13546 (N_13546,N_13396,N_13379);
and U13547 (N_13547,N_13363,N_13498);
xnor U13548 (N_13548,N_13381,N_13479);
or U13549 (N_13549,N_13371,N_13439);
xnor U13550 (N_13550,N_13475,N_13422);
and U13551 (N_13551,N_13487,N_13489);
xor U13552 (N_13552,N_13386,N_13350);
nor U13553 (N_13553,N_13387,N_13410);
xor U13554 (N_13554,N_13383,N_13388);
or U13555 (N_13555,N_13416,N_13458);
xor U13556 (N_13556,N_13493,N_13440);
xor U13557 (N_13557,N_13418,N_13411);
or U13558 (N_13558,N_13357,N_13412);
or U13559 (N_13559,N_13460,N_13456);
or U13560 (N_13560,N_13370,N_13395);
nor U13561 (N_13561,N_13352,N_13351);
or U13562 (N_13562,N_13423,N_13397);
xor U13563 (N_13563,N_13430,N_13455);
or U13564 (N_13564,N_13486,N_13431);
nand U13565 (N_13565,N_13474,N_13417);
xor U13566 (N_13566,N_13384,N_13459);
nor U13567 (N_13567,N_13443,N_13367);
nor U13568 (N_13568,N_13391,N_13415);
nand U13569 (N_13569,N_13436,N_13484);
nand U13570 (N_13570,N_13442,N_13437);
and U13571 (N_13571,N_13407,N_13472);
xnor U13572 (N_13572,N_13480,N_13465);
and U13573 (N_13573,N_13494,N_13355);
xnor U13574 (N_13574,N_13452,N_13454);
nor U13575 (N_13575,N_13429,N_13375);
and U13576 (N_13576,N_13471,N_13474);
or U13577 (N_13577,N_13457,N_13402);
xnor U13578 (N_13578,N_13371,N_13395);
nand U13579 (N_13579,N_13401,N_13375);
and U13580 (N_13580,N_13468,N_13417);
nand U13581 (N_13581,N_13381,N_13376);
or U13582 (N_13582,N_13382,N_13397);
nor U13583 (N_13583,N_13408,N_13427);
and U13584 (N_13584,N_13441,N_13374);
or U13585 (N_13585,N_13444,N_13479);
xor U13586 (N_13586,N_13368,N_13448);
nand U13587 (N_13587,N_13350,N_13353);
nand U13588 (N_13588,N_13369,N_13440);
and U13589 (N_13589,N_13387,N_13431);
xnor U13590 (N_13590,N_13452,N_13476);
nor U13591 (N_13591,N_13441,N_13402);
nor U13592 (N_13592,N_13351,N_13496);
nor U13593 (N_13593,N_13356,N_13366);
xor U13594 (N_13594,N_13416,N_13380);
or U13595 (N_13595,N_13392,N_13370);
nor U13596 (N_13596,N_13397,N_13400);
nand U13597 (N_13597,N_13384,N_13492);
xor U13598 (N_13598,N_13378,N_13363);
nand U13599 (N_13599,N_13384,N_13374);
and U13600 (N_13600,N_13360,N_13492);
nand U13601 (N_13601,N_13369,N_13399);
or U13602 (N_13602,N_13469,N_13426);
and U13603 (N_13603,N_13382,N_13461);
and U13604 (N_13604,N_13391,N_13375);
or U13605 (N_13605,N_13434,N_13362);
xor U13606 (N_13606,N_13481,N_13453);
xnor U13607 (N_13607,N_13458,N_13406);
or U13608 (N_13608,N_13399,N_13465);
xnor U13609 (N_13609,N_13445,N_13476);
or U13610 (N_13610,N_13481,N_13443);
nor U13611 (N_13611,N_13494,N_13373);
nor U13612 (N_13612,N_13461,N_13425);
and U13613 (N_13613,N_13432,N_13425);
nor U13614 (N_13614,N_13364,N_13468);
xnor U13615 (N_13615,N_13473,N_13368);
nor U13616 (N_13616,N_13478,N_13443);
or U13617 (N_13617,N_13419,N_13393);
or U13618 (N_13618,N_13442,N_13367);
xnor U13619 (N_13619,N_13444,N_13416);
xnor U13620 (N_13620,N_13367,N_13397);
nand U13621 (N_13621,N_13494,N_13352);
xor U13622 (N_13622,N_13395,N_13392);
nor U13623 (N_13623,N_13389,N_13382);
or U13624 (N_13624,N_13379,N_13404);
and U13625 (N_13625,N_13446,N_13497);
nand U13626 (N_13626,N_13459,N_13440);
nand U13627 (N_13627,N_13463,N_13495);
and U13628 (N_13628,N_13460,N_13432);
xnor U13629 (N_13629,N_13415,N_13466);
xor U13630 (N_13630,N_13354,N_13379);
or U13631 (N_13631,N_13423,N_13402);
nand U13632 (N_13632,N_13407,N_13427);
nor U13633 (N_13633,N_13479,N_13424);
nor U13634 (N_13634,N_13367,N_13473);
xnor U13635 (N_13635,N_13400,N_13403);
nor U13636 (N_13636,N_13483,N_13489);
nand U13637 (N_13637,N_13382,N_13381);
nor U13638 (N_13638,N_13376,N_13357);
or U13639 (N_13639,N_13396,N_13464);
and U13640 (N_13640,N_13422,N_13400);
xnor U13641 (N_13641,N_13403,N_13474);
and U13642 (N_13642,N_13473,N_13431);
nor U13643 (N_13643,N_13405,N_13360);
nand U13644 (N_13644,N_13401,N_13432);
and U13645 (N_13645,N_13439,N_13385);
nand U13646 (N_13646,N_13460,N_13449);
xor U13647 (N_13647,N_13485,N_13468);
xor U13648 (N_13648,N_13416,N_13490);
and U13649 (N_13649,N_13452,N_13451);
or U13650 (N_13650,N_13640,N_13536);
and U13651 (N_13651,N_13619,N_13508);
nor U13652 (N_13652,N_13579,N_13636);
and U13653 (N_13653,N_13639,N_13592);
and U13654 (N_13654,N_13598,N_13513);
xnor U13655 (N_13655,N_13567,N_13593);
xor U13656 (N_13656,N_13510,N_13591);
or U13657 (N_13657,N_13526,N_13525);
nand U13658 (N_13658,N_13546,N_13589);
or U13659 (N_13659,N_13607,N_13643);
nand U13660 (N_13660,N_13511,N_13558);
nor U13661 (N_13661,N_13524,N_13624);
xor U13662 (N_13662,N_13547,N_13646);
nand U13663 (N_13663,N_13527,N_13500);
nor U13664 (N_13664,N_13532,N_13577);
xnor U13665 (N_13665,N_13584,N_13630);
and U13666 (N_13666,N_13551,N_13585);
or U13667 (N_13667,N_13610,N_13556);
and U13668 (N_13668,N_13635,N_13520);
and U13669 (N_13669,N_13569,N_13620);
and U13670 (N_13670,N_13634,N_13538);
or U13671 (N_13671,N_13590,N_13506);
xor U13672 (N_13672,N_13563,N_13514);
and U13673 (N_13673,N_13565,N_13509);
nor U13674 (N_13674,N_13580,N_13537);
xnor U13675 (N_13675,N_13649,N_13517);
xor U13676 (N_13676,N_13564,N_13642);
nand U13677 (N_13677,N_13534,N_13632);
or U13678 (N_13678,N_13574,N_13605);
or U13679 (N_13679,N_13609,N_13600);
nand U13680 (N_13680,N_13612,N_13512);
nand U13681 (N_13681,N_13516,N_13638);
and U13682 (N_13682,N_13641,N_13622);
nor U13683 (N_13683,N_13608,N_13542);
or U13684 (N_13684,N_13614,N_13501);
and U13685 (N_13685,N_13587,N_13544);
or U13686 (N_13686,N_13596,N_13621);
nand U13687 (N_13687,N_13504,N_13644);
or U13688 (N_13688,N_13555,N_13616);
and U13689 (N_13689,N_13539,N_13535);
and U13690 (N_13690,N_13629,N_13515);
xnor U13691 (N_13691,N_13505,N_13571);
nand U13692 (N_13692,N_13531,N_13645);
and U13693 (N_13693,N_13543,N_13541);
and U13694 (N_13694,N_13548,N_13557);
xnor U13695 (N_13695,N_13560,N_13623);
nor U13696 (N_13696,N_13631,N_13637);
or U13697 (N_13697,N_13583,N_13528);
nor U13698 (N_13698,N_13562,N_13529);
xor U13699 (N_13699,N_13626,N_13599);
nand U13700 (N_13700,N_13595,N_13594);
nor U13701 (N_13701,N_13613,N_13572);
nor U13702 (N_13702,N_13597,N_13586);
or U13703 (N_13703,N_13518,N_13549);
xnor U13704 (N_13704,N_13573,N_13533);
nand U13705 (N_13705,N_13601,N_13627);
nand U13706 (N_13706,N_13617,N_13603);
and U13707 (N_13707,N_13602,N_13553);
xor U13708 (N_13708,N_13582,N_13575);
or U13709 (N_13709,N_13615,N_13604);
or U13710 (N_13710,N_13568,N_13522);
xor U13711 (N_13711,N_13559,N_13519);
or U13712 (N_13712,N_13570,N_13540);
nor U13713 (N_13713,N_13554,N_13550);
or U13714 (N_13714,N_13545,N_13588);
nand U13715 (N_13715,N_13507,N_13581);
nand U13716 (N_13716,N_13503,N_13523);
and U13717 (N_13717,N_13502,N_13633);
or U13718 (N_13718,N_13530,N_13566);
or U13719 (N_13719,N_13576,N_13618);
nand U13720 (N_13720,N_13625,N_13647);
nor U13721 (N_13721,N_13561,N_13611);
or U13722 (N_13722,N_13552,N_13521);
nand U13723 (N_13723,N_13606,N_13578);
nand U13724 (N_13724,N_13648,N_13628);
and U13725 (N_13725,N_13522,N_13544);
or U13726 (N_13726,N_13527,N_13637);
and U13727 (N_13727,N_13588,N_13532);
nor U13728 (N_13728,N_13501,N_13592);
nor U13729 (N_13729,N_13611,N_13536);
nor U13730 (N_13730,N_13542,N_13605);
nand U13731 (N_13731,N_13594,N_13635);
nand U13732 (N_13732,N_13571,N_13556);
nand U13733 (N_13733,N_13599,N_13598);
or U13734 (N_13734,N_13615,N_13585);
and U13735 (N_13735,N_13648,N_13603);
nand U13736 (N_13736,N_13530,N_13568);
xnor U13737 (N_13737,N_13548,N_13628);
xor U13738 (N_13738,N_13640,N_13546);
xnor U13739 (N_13739,N_13542,N_13576);
xor U13740 (N_13740,N_13570,N_13596);
xor U13741 (N_13741,N_13618,N_13635);
xor U13742 (N_13742,N_13563,N_13646);
nand U13743 (N_13743,N_13645,N_13633);
xor U13744 (N_13744,N_13609,N_13576);
and U13745 (N_13745,N_13594,N_13500);
nor U13746 (N_13746,N_13545,N_13504);
nor U13747 (N_13747,N_13628,N_13620);
nand U13748 (N_13748,N_13550,N_13634);
or U13749 (N_13749,N_13604,N_13570);
or U13750 (N_13750,N_13639,N_13595);
or U13751 (N_13751,N_13593,N_13548);
nor U13752 (N_13752,N_13544,N_13569);
nand U13753 (N_13753,N_13641,N_13596);
nor U13754 (N_13754,N_13520,N_13634);
xor U13755 (N_13755,N_13605,N_13636);
nand U13756 (N_13756,N_13647,N_13541);
nor U13757 (N_13757,N_13601,N_13596);
and U13758 (N_13758,N_13548,N_13649);
nor U13759 (N_13759,N_13516,N_13578);
xnor U13760 (N_13760,N_13548,N_13527);
nand U13761 (N_13761,N_13523,N_13551);
nand U13762 (N_13762,N_13583,N_13523);
xnor U13763 (N_13763,N_13575,N_13601);
nand U13764 (N_13764,N_13533,N_13537);
nand U13765 (N_13765,N_13517,N_13501);
nor U13766 (N_13766,N_13601,N_13604);
nor U13767 (N_13767,N_13507,N_13577);
or U13768 (N_13768,N_13537,N_13643);
and U13769 (N_13769,N_13597,N_13554);
nor U13770 (N_13770,N_13624,N_13584);
xnor U13771 (N_13771,N_13576,N_13616);
nor U13772 (N_13772,N_13531,N_13542);
and U13773 (N_13773,N_13517,N_13561);
nor U13774 (N_13774,N_13501,N_13506);
nor U13775 (N_13775,N_13597,N_13512);
or U13776 (N_13776,N_13566,N_13526);
nand U13777 (N_13777,N_13507,N_13596);
xor U13778 (N_13778,N_13611,N_13505);
nand U13779 (N_13779,N_13596,N_13512);
xor U13780 (N_13780,N_13549,N_13566);
and U13781 (N_13781,N_13560,N_13518);
or U13782 (N_13782,N_13544,N_13523);
or U13783 (N_13783,N_13506,N_13512);
and U13784 (N_13784,N_13504,N_13629);
xor U13785 (N_13785,N_13527,N_13516);
nand U13786 (N_13786,N_13551,N_13611);
and U13787 (N_13787,N_13571,N_13612);
and U13788 (N_13788,N_13601,N_13543);
and U13789 (N_13789,N_13534,N_13508);
nor U13790 (N_13790,N_13587,N_13567);
xnor U13791 (N_13791,N_13640,N_13517);
or U13792 (N_13792,N_13532,N_13614);
nand U13793 (N_13793,N_13581,N_13614);
nand U13794 (N_13794,N_13594,N_13618);
xor U13795 (N_13795,N_13534,N_13536);
nand U13796 (N_13796,N_13587,N_13525);
or U13797 (N_13797,N_13528,N_13546);
and U13798 (N_13798,N_13538,N_13589);
and U13799 (N_13799,N_13529,N_13592);
or U13800 (N_13800,N_13770,N_13698);
nand U13801 (N_13801,N_13797,N_13764);
xor U13802 (N_13802,N_13726,N_13684);
xor U13803 (N_13803,N_13717,N_13686);
nor U13804 (N_13804,N_13775,N_13734);
or U13805 (N_13805,N_13712,N_13679);
nand U13806 (N_13806,N_13733,N_13796);
and U13807 (N_13807,N_13784,N_13765);
or U13808 (N_13808,N_13740,N_13705);
nand U13809 (N_13809,N_13693,N_13776);
or U13810 (N_13810,N_13651,N_13745);
nor U13811 (N_13811,N_13773,N_13751);
and U13812 (N_13812,N_13655,N_13683);
and U13813 (N_13813,N_13700,N_13708);
nor U13814 (N_13814,N_13680,N_13779);
nand U13815 (N_13815,N_13676,N_13694);
nor U13816 (N_13816,N_13721,N_13695);
or U13817 (N_13817,N_13711,N_13743);
xnor U13818 (N_13818,N_13752,N_13750);
xor U13819 (N_13819,N_13774,N_13736);
xor U13820 (N_13820,N_13709,N_13656);
nand U13821 (N_13821,N_13672,N_13760);
nor U13822 (N_13822,N_13701,N_13744);
nor U13823 (N_13823,N_13718,N_13681);
xor U13824 (N_13824,N_13771,N_13790);
xnor U13825 (N_13825,N_13722,N_13691);
nand U13826 (N_13826,N_13769,N_13723);
xnor U13827 (N_13827,N_13737,N_13728);
xnor U13828 (N_13828,N_13696,N_13665);
nor U13829 (N_13829,N_13732,N_13714);
xor U13830 (N_13830,N_13677,N_13664);
xor U13831 (N_13831,N_13657,N_13731);
and U13832 (N_13832,N_13759,N_13725);
nand U13833 (N_13833,N_13652,N_13682);
and U13834 (N_13834,N_13762,N_13707);
and U13835 (N_13835,N_13670,N_13703);
xnor U13836 (N_13836,N_13787,N_13788);
nand U13837 (N_13837,N_13669,N_13650);
and U13838 (N_13838,N_13710,N_13793);
nand U13839 (N_13839,N_13742,N_13663);
nand U13840 (N_13840,N_13781,N_13795);
and U13841 (N_13841,N_13719,N_13791);
and U13842 (N_13842,N_13727,N_13706);
nand U13843 (N_13843,N_13689,N_13766);
nor U13844 (N_13844,N_13697,N_13778);
nand U13845 (N_13845,N_13756,N_13757);
or U13846 (N_13846,N_13768,N_13688);
xnor U13847 (N_13847,N_13799,N_13749);
xor U13848 (N_13848,N_13687,N_13747);
nor U13849 (N_13849,N_13748,N_13658);
xor U13850 (N_13850,N_13673,N_13685);
xnor U13851 (N_13851,N_13753,N_13716);
xnor U13852 (N_13852,N_13654,N_13661);
nand U13853 (N_13853,N_13675,N_13746);
or U13854 (N_13854,N_13720,N_13662);
nor U13855 (N_13855,N_13789,N_13729);
or U13856 (N_13856,N_13763,N_13735);
nand U13857 (N_13857,N_13702,N_13761);
and U13858 (N_13858,N_13782,N_13667);
and U13859 (N_13859,N_13767,N_13715);
xnor U13860 (N_13860,N_13792,N_13653);
xor U13861 (N_13861,N_13713,N_13666);
nor U13862 (N_13862,N_13739,N_13786);
or U13863 (N_13863,N_13772,N_13678);
xnor U13864 (N_13864,N_13692,N_13671);
and U13865 (N_13865,N_13755,N_13738);
and U13866 (N_13866,N_13785,N_13783);
and U13867 (N_13867,N_13668,N_13674);
and U13868 (N_13868,N_13730,N_13704);
and U13869 (N_13869,N_13798,N_13777);
nor U13870 (N_13870,N_13780,N_13660);
and U13871 (N_13871,N_13659,N_13741);
xnor U13872 (N_13872,N_13794,N_13699);
or U13873 (N_13873,N_13754,N_13724);
nor U13874 (N_13874,N_13690,N_13758);
xnor U13875 (N_13875,N_13732,N_13677);
or U13876 (N_13876,N_13796,N_13714);
xnor U13877 (N_13877,N_13697,N_13721);
or U13878 (N_13878,N_13758,N_13685);
nor U13879 (N_13879,N_13741,N_13777);
and U13880 (N_13880,N_13713,N_13753);
nor U13881 (N_13881,N_13725,N_13736);
or U13882 (N_13882,N_13788,N_13767);
and U13883 (N_13883,N_13797,N_13716);
nor U13884 (N_13884,N_13791,N_13713);
xor U13885 (N_13885,N_13712,N_13698);
nand U13886 (N_13886,N_13674,N_13725);
nor U13887 (N_13887,N_13763,N_13657);
nand U13888 (N_13888,N_13784,N_13697);
or U13889 (N_13889,N_13766,N_13781);
nand U13890 (N_13890,N_13752,N_13713);
or U13891 (N_13891,N_13767,N_13672);
nand U13892 (N_13892,N_13757,N_13768);
nor U13893 (N_13893,N_13684,N_13683);
nor U13894 (N_13894,N_13780,N_13682);
nor U13895 (N_13895,N_13702,N_13748);
nand U13896 (N_13896,N_13732,N_13776);
and U13897 (N_13897,N_13661,N_13727);
and U13898 (N_13898,N_13676,N_13675);
nor U13899 (N_13899,N_13795,N_13672);
or U13900 (N_13900,N_13729,N_13724);
nand U13901 (N_13901,N_13774,N_13761);
xnor U13902 (N_13902,N_13693,N_13775);
or U13903 (N_13903,N_13717,N_13769);
xnor U13904 (N_13904,N_13681,N_13710);
xnor U13905 (N_13905,N_13650,N_13742);
nor U13906 (N_13906,N_13744,N_13698);
xnor U13907 (N_13907,N_13665,N_13685);
and U13908 (N_13908,N_13660,N_13674);
and U13909 (N_13909,N_13780,N_13684);
or U13910 (N_13910,N_13659,N_13778);
xor U13911 (N_13911,N_13666,N_13787);
and U13912 (N_13912,N_13741,N_13698);
and U13913 (N_13913,N_13679,N_13696);
and U13914 (N_13914,N_13695,N_13671);
nand U13915 (N_13915,N_13661,N_13658);
xor U13916 (N_13916,N_13651,N_13787);
xor U13917 (N_13917,N_13727,N_13700);
nor U13918 (N_13918,N_13654,N_13741);
and U13919 (N_13919,N_13750,N_13702);
and U13920 (N_13920,N_13799,N_13697);
and U13921 (N_13921,N_13661,N_13663);
or U13922 (N_13922,N_13706,N_13736);
nor U13923 (N_13923,N_13722,N_13705);
xor U13924 (N_13924,N_13695,N_13747);
nand U13925 (N_13925,N_13677,N_13657);
or U13926 (N_13926,N_13767,N_13670);
xnor U13927 (N_13927,N_13760,N_13673);
and U13928 (N_13928,N_13661,N_13788);
nand U13929 (N_13929,N_13682,N_13705);
and U13930 (N_13930,N_13697,N_13764);
nand U13931 (N_13931,N_13795,N_13742);
xor U13932 (N_13932,N_13701,N_13780);
or U13933 (N_13933,N_13790,N_13692);
or U13934 (N_13934,N_13675,N_13747);
or U13935 (N_13935,N_13652,N_13727);
and U13936 (N_13936,N_13743,N_13740);
nand U13937 (N_13937,N_13657,N_13793);
or U13938 (N_13938,N_13780,N_13706);
nor U13939 (N_13939,N_13718,N_13677);
nand U13940 (N_13940,N_13728,N_13778);
and U13941 (N_13941,N_13710,N_13745);
and U13942 (N_13942,N_13694,N_13757);
nor U13943 (N_13943,N_13755,N_13677);
and U13944 (N_13944,N_13673,N_13790);
xnor U13945 (N_13945,N_13740,N_13677);
xor U13946 (N_13946,N_13666,N_13756);
xnor U13947 (N_13947,N_13789,N_13660);
nor U13948 (N_13948,N_13699,N_13750);
nand U13949 (N_13949,N_13682,N_13694);
nor U13950 (N_13950,N_13879,N_13908);
and U13951 (N_13951,N_13942,N_13903);
nand U13952 (N_13952,N_13815,N_13931);
nand U13953 (N_13953,N_13887,N_13829);
nor U13954 (N_13954,N_13926,N_13809);
and U13955 (N_13955,N_13873,N_13900);
nor U13956 (N_13956,N_13822,N_13823);
xor U13957 (N_13957,N_13919,N_13835);
nor U13958 (N_13958,N_13914,N_13867);
nand U13959 (N_13959,N_13834,N_13848);
or U13960 (N_13960,N_13875,N_13880);
nor U13961 (N_13961,N_13906,N_13806);
nand U13962 (N_13962,N_13925,N_13853);
nand U13963 (N_13963,N_13830,N_13858);
nand U13964 (N_13964,N_13932,N_13832);
nor U13965 (N_13965,N_13826,N_13939);
nand U13966 (N_13966,N_13840,N_13907);
nor U13967 (N_13967,N_13802,N_13947);
xor U13968 (N_13968,N_13821,N_13876);
or U13969 (N_13969,N_13898,N_13807);
and U13970 (N_13970,N_13850,N_13904);
and U13971 (N_13971,N_13837,N_13816);
nor U13972 (N_13972,N_13863,N_13843);
and U13973 (N_13973,N_13805,N_13937);
or U13974 (N_13974,N_13871,N_13888);
nand U13975 (N_13975,N_13921,N_13868);
xnor U13976 (N_13976,N_13943,N_13846);
xor U13977 (N_13977,N_13874,N_13804);
nand U13978 (N_13978,N_13899,N_13940);
nor U13979 (N_13979,N_13842,N_13841);
nand U13980 (N_13980,N_13866,N_13909);
or U13981 (N_13981,N_13844,N_13882);
and U13982 (N_13982,N_13810,N_13890);
xor U13983 (N_13983,N_13859,N_13820);
nor U13984 (N_13984,N_13905,N_13861);
and U13985 (N_13985,N_13941,N_13916);
or U13986 (N_13986,N_13845,N_13860);
or U13987 (N_13987,N_13948,N_13901);
or U13988 (N_13988,N_13895,N_13930);
or U13989 (N_13989,N_13819,N_13938);
nor U13990 (N_13990,N_13878,N_13949);
or U13991 (N_13991,N_13894,N_13920);
nor U13992 (N_13992,N_13865,N_13884);
xnor U13993 (N_13993,N_13902,N_13881);
or U13994 (N_13994,N_13801,N_13913);
and U13995 (N_13995,N_13849,N_13813);
or U13996 (N_13996,N_13944,N_13927);
nand U13997 (N_13997,N_13883,N_13855);
xor U13998 (N_13998,N_13862,N_13872);
nand U13999 (N_13999,N_13933,N_13818);
and U14000 (N_14000,N_13893,N_13812);
nor U14001 (N_14001,N_13817,N_13857);
and U14002 (N_14002,N_13897,N_13828);
or U14003 (N_14003,N_13833,N_13936);
xnor U14004 (N_14004,N_13869,N_13854);
or U14005 (N_14005,N_13827,N_13811);
nand U14006 (N_14006,N_13928,N_13839);
nor U14007 (N_14007,N_13847,N_13929);
xnor U14008 (N_14008,N_13838,N_13891);
and U14009 (N_14009,N_13924,N_13808);
and U14010 (N_14010,N_13852,N_13889);
or U14011 (N_14011,N_13912,N_13935);
nand U14012 (N_14012,N_13886,N_13923);
or U14013 (N_14013,N_13946,N_13831);
or U14014 (N_14014,N_13945,N_13803);
xnor U14015 (N_14015,N_13911,N_13851);
nor U14016 (N_14016,N_13824,N_13922);
nand U14017 (N_14017,N_13918,N_13800);
nor U14018 (N_14018,N_13885,N_13825);
nand U14019 (N_14019,N_13896,N_13856);
xnor U14020 (N_14020,N_13814,N_13877);
and U14021 (N_14021,N_13917,N_13915);
nand U14022 (N_14022,N_13870,N_13910);
nand U14023 (N_14023,N_13892,N_13864);
or U14024 (N_14024,N_13934,N_13836);
nand U14025 (N_14025,N_13841,N_13807);
nand U14026 (N_14026,N_13800,N_13910);
nor U14027 (N_14027,N_13876,N_13942);
nand U14028 (N_14028,N_13820,N_13915);
and U14029 (N_14029,N_13845,N_13883);
xor U14030 (N_14030,N_13856,N_13867);
and U14031 (N_14031,N_13903,N_13835);
xnor U14032 (N_14032,N_13841,N_13869);
nor U14033 (N_14033,N_13802,N_13837);
or U14034 (N_14034,N_13921,N_13880);
and U14035 (N_14035,N_13913,N_13946);
nor U14036 (N_14036,N_13864,N_13943);
or U14037 (N_14037,N_13817,N_13822);
nand U14038 (N_14038,N_13813,N_13840);
or U14039 (N_14039,N_13801,N_13823);
nor U14040 (N_14040,N_13927,N_13899);
and U14041 (N_14041,N_13852,N_13833);
and U14042 (N_14042,N_13900,N_13802);
and U14043 (N_14043,N_13853,N_13907);
and U14044 (N_14044,N_13806,N_13856);
and U14045 (N_14045,N_13898,N_13842);
nand U14046 (N_14046,N_13818,N_13805);
or U14047 (N_14047,N_13870,N_13847);
nor U14048 (N_14048,N_13840,N_13930);
nor U14049 (N_14049,N_13876,N_13949);
nor U14050 (N_14050,N_13848,N_13888);
xor U14051 (N_14051,N_13912,N_13886);
or U14052 (N_14052,N_13928,N_13872);
nor U14053 (N_14053,N_13937,N_13918);
nand U14054 (N_14054,N_13829,N_13881);
and U14055 (N_14055,N_13831,N_13815);
or U14056 (N_14056,N_13899,N_13882);
nor U14057 (N_14057,N_13897,N_13840);
xor U14058 (N_14058,N_13856,N_13801);
nor U14059 (N_14059,N_13911,N_13935);
or U14060 (N_14060,N_13879,N_13895);
or U14061 (N_14061,N_13853,N_13932);
nor U14062 (N_14062,N_13854,N_13946);
nand U14063 (N_14063,N_13815,N_13947);
or U14064 (N_14064,N_13821,N_13878);
nor U14065 (N_14065,N_13865,N_13888);
nor U14066 (N_14066,N_13815,N_13850);
xnor U14067 (N_14067,N_13874,N_13816);
or U14068 (N_14068,N_13939,N_13930);
nand U14069 (N_14069,N_13834,N_13915);
or U14070 (N_14070,N_13869,N_13914);
xor U14071 (N_14071,N_13936,N_13824);
nor U14072 (N_14072,N_13831,N_13923);
xor U14073 (N_14073,N_13930,N_13818);
and U14074 (N_14074,N_13879,N_13816);
nor U14075 (N_14075,N_13886,N_13887);
or U14076 (N_14076,N_13882,N_13800);
nor U14077 (N_14077,N_13851,N_13940);
and U14078 (N_14078,N_13895,N_13938);
or U14079 (N_14079,N_13914,N_13905);
xnor U14080 (N_14080,N_13841,N_13905);
nand U14081 (N_14081,N_13858,N_13942);
xor U14082 (N_14082,N_13837,N_13908);
nand U14083 (N_14083,N_13916,N_13866);
xnor U14084 (N_14084,N_13943,N_13858);
nand U14085 (N_14085,N_13855,N_13877);
and U14086 (N_14086,N_13941,N_13835);
nand U14087 (N_14087,N_13930,N_13948);
or U14088 (N_14088,N_13919,N_13839);
nand U14089 (N_14089,N_13867,N_13911);
and U14090 (N_14090,N_13908,N_13810);
and U14091 (N_14091,N_13949,N_13870);
xor U14092 (N_14092,N_13927,N_13808);
nand U14093 (N_14093,N_13873,N_13926);
nor U14094 (N_14094,N_13828,N_13946);
nand U14095 (N_14095,N_13832,N_13934);
and U14096 (N_14096,N_13828,N_13949);
and U14097 (N_14097,N_13820,N_13831);
or U14098 (N_14098,N_13822,N_13804);
and U14099 (N_14099,N_13886,N_13826);
and U14100 (N_14100,N_13958,N_13962);
nand U14101 (N_14101,N_14086,N_14073);
nand U14102 (N_14102,N_14035,N_14023);
or U14103 (N_14103,N_13986,N_14070);
or U14104 (N_14104,N_14002,N_14080);
nor U14105 (N_14105,N_13994,N_14043);
or U14106 (N_14106,N_13951,N_14007);
nand U14107 (N_14107,N_14029,N_14089);
or U14108 (N_14108,N_13999,N_14099);
nor U14109 (N_14109,N_14095,N_14049);
xor U14110 (N_14110,N_14090,N_13971);
or U14111 (N_14111,N_14097,N_14079);
nand U14112 (N_14112,N_13974,N_14085);
nor U14113 (N_14113,N_13970,N_13953);
nor U14114 (N_14114,N_14062,N_14059);
or U14115 (N_14115,N_14005,N_14056);
nor U14116 (N_14116,N_14014,N_14075);
nor U14117 (N_14117,N_14036,N_13976);
or U14118 (N_14118,N_14091,N_14016);
and U14119 (N_14119,N_14067,N_14017);
nor U14120 (N_14120,N_14001,N_13969);
xnor U14121 (N_14121,N_13961,N_14046);
or U14122 (N_14122,N_14011,N_14064);
nand U14123 (N_14123,N_14032,N_14088);
or U14124 (N_14124,N_14030,N_13979);
and U14125 (N_14125,N_13952,N_13988);
nor U14126 (N_14126,N_13960,N_14050);
nand U14127 (N_14127,N_14081,N_13998);
xor U14128 (N_14128,N_14092,N_14024);
or U14129 (N_14129,N_13984,N_14060);
nor U14130 (N_14130,N_13954,N_13997);
or U14131 (N_14131,N_14031,N_13967);
xor U14132 (N_14132,N_14010,N_14026);
and U14133 (N_14133,N_14068,N_13995);
xor U14134 (N_14134,N_14012,N_13992);
nor U14135 (N_14135,N_14055,N_14034);
nand U14136 (N_14136,N_14093,N_14074);
and U14137 (N_14137,N_14069,N_14000);
and U14138 (N_14138,N_14048,N_14072);
and U14139 (N_14139,N_13989,N_14096);
and U14140 (N_14140,N_13963,N_14071);
nand U14141 (N_14141,N_14018,N_14022);
nor U14142 (N_14142,N_14027,N_14057);
or U14143 (N_14143,N_14020,N_14051);
xnor U14144 (N_14144,N_13955,N_14041);
xnor U14145 (N_14145,N_14077,N_14052);
and U14146 (N_14146,N_14028,N_14042);
nand U14147 (N_14147,N_13987,N_13957);
nor U14148 (N_14148,N_14054,N_14076);
nand U14149 (N_14149,N_13981,N_13996);
nand U14150 (N_14150,N_14004,N_14094);
nor U14151 (N_14151,N_14058,N_14084);
nor U14152 (N_14152,N_14082,N_14040);
nor U14153 (N_14153,N_13977,N_14039);
and U14154 (N_14154,N_14008,N_14053);
nor U14155 (N_14155,N_14021,N_14087);
nor U14156 (N_14156,N_14098,N_13985);
nand U14157 (N_14157,N_13950,N_14066);
or U14158 (N_14158,N_14038,N_13959);
xnor U14159 (N_14159,N_13968,N_14037);
nor U14160 (N_14160,N_14047,N_13965);
nor U14161 (N_14161,N_13972,N_14045);
nand U14162 (N_14162,N_13991,N_13956);
xor U14163 (N_14163,N_14033,N_13980);
xnor U14164 (N_14164,N_14009,N_14015);
nor U14165 (N_14165,N_14078,N_13964);
nor U14166 (N_14166,N_13983,N_14065);
nor U14167 (N_14167,N_14063,N_13966);
nor U14168 (N_14168,N_13978,N_13982);
xor U14169 (N_14169,N_14006,N_13993);
xnor U14170 (N_14170,N_14025,N_13973);
or U14171 (N_14171,N_14083,N_14061);
xor U14172 (N_14172,N_13975,N_14019);
nand U14173 (N_14173,N_14003,N_14044);
or U14174 (N_14174,N_14013,N_13990);
and U14175 (N_14175,N_13966,N_14088);
or U14176 (N_14176,N_13981,N_13989);
nor U14177 (N_14177,N_14020,N_13972);
and U14178 (N_14178,N_14015,N_13980);
and U14179 (N_14179,N_13981,N_13976);
nand U14180 (N_14180,N_14058,N_14076);
and U14181 (N_14181,N_14030,N_14007);
nand U14182 (N_14182,N_13985,N_14030);
nor U14183 (N_14183,N_14014,N_13963);
nor U14184 (N_14184,N_14033,N_13962);
nand U14185 (N_14185,N_13985,N_14008);
xnor U14186 (N_14186,N_14027,N_14058);
nand U14187 (N_14187,N_14061,N_13981);
xor U14188 (N_14188,N_14031,N_13991);
xnor U14189 (N_14189,N_14015,N_14008);
and U14190 (N_14190,N_14022,N_13977);
or U14191 (N_14191,N_14034,N_13993);
nand U14192 (N_14192,N_14070,N_14021);
nor U14193 (N_14193,N_14090,N_13979);
nand U14194 (N_14194,N_14034,N_14064);
or U14195 (N_14195,N_14063,N_14015);
and U14196 (N_14196,N_13969,N_13962);
and U14197 (N_14197,N_13966,N_13996);
nand U14198 (N_14198,N_14069,N_14041);
or U14199 (N_14199,N_14014,N_14074);
xor U14200 (N_14200,N_14039,N_14099);
xnor U14201 (N_14201,N_14089,N_14087);
xnor U14202 (N_14202,N_14027,N_14084);
and U14203 (N_14203,N_14017,N_14057);
nand U14204 (N_14204,N_14033,N_13971);
and U14205 (N_14205,N_14080,N_13985);
xor U14206 (N_14206,N_13960,N_14090);
and U14207 (N_14207,N_13976,N_14096);
nand U14208 (N_14208,N_14022,N_14069);
and U14209 (N_14209,N_14066,N_14085);
or U14210 (N_14210,N_14063,N_14031);
or U14211 (N_14211,N_14091,N_13999);
xor U14212 (N_14212,N_14073,N_14000);
xnor U14213 (N_14213,N_13973,N_14036);
or U14214 (N_14214,N_14083,N_14034);
or U14215 (N_14215,N_13987,N_14083);
xnor U14216 (N_14216,N_14090,N_13959);
xnor U14217 (N_14217,N_14075,N_13988);
and U14218 (N_14218,N_13966,N_13962);
and U14219 (N_14219,N_14047,N_14059);
nand U14220 (N_14220,N_13962,N_14034);
or U14221 (N_14221,N_13978,N_14014);
or U14222 (N_14222,N_13973,N_13970);
nand U14223 (N_14223,N_14099,N_13977);
nand U14224 (N_14224,N_13997,N_14012);
or U14225 (N_14225,N_13964,N_14055);
or U14226 (N_14226,N_14050,N_13971);
nand U14227 (N_14227,N_14054,N_13961);
nor U14228 (N_14228,N_14004,N_14063);
xnor U14229 (N_14229,N_13984,N_13958);
nand U14230 (N_14230,N_14047,N_13999);
xor U14231 (N_14231,N_14070,N_14063);
xor U14232 (N_14232,N_14060,N_14089);
and U14233 (N_14233,N_14055,N_14024);
and U14234 (N_14234,N_13963,N_14064);
or U14235 (N_14235,N_14007,N_13972);
and U14236 (N_14236,N_14032,N_13996);
nor U14237 (N_14237,N_14064,N_14048);
or U14238 (N_14238,N_13954,N_13964);
and U14239 (N_14239,N_13989,N_14042);
nor U14240 (N_14240,N_14030,N_14014);
and U14241 (N_14241,N_13984,N_14058);
and U14242 (N_14242,N_14029,N_13959);
xor U14243 (N_14243,N_13984,N_14086);
and U14244 (N_14244,N_14049,N_14075);
xnor U14245 (N_14245,N_13988,N_14000);
xnor U14246 (N_14246,N_13958,N_14032);
or U14247 (N_14247,N_14086,N_14094);
xor U14248 (N_14248,N_13984,N_13968);
and U14249 (N_14249,N_13968,N_14065);
nor U14250 (N_14250,N_14104,N_14195);
nor U14251 (N_14251,N_14246,N_14191);
and U14252 (N_14252,N_14207,N_14154);
xnor U14253 (N_14253,N_14202,N_14166);
or U14254 (N_14254,N_14220,N_14144);
xor U14255 (N_14255,N_14152,N_14175);
xor U14256 (N_14256,N_14223,N_14233);
nand U14257 (N_14257,N_14117,N_14174);
nor U14258 (N_14258,N_14176,N_14214);
and U14259 (N_14259,N_14222,N_14188);
nand U14260 (N_14260,N_14146,N_14213);
xnor U14261 (N_14261,N_14189,N_14249);
nor U14262 (N_14262,N_14196,N_14122);
xnor U14263 (N_14263,N_14192,N_14147);
and U14264 (N_14264,N_14161,N_14136);
or U14265 (N_14265,N_14138,N_14100);
and U14266 (N_14266,N_14225,N_14140);
xor U14267 (N_14267,N_14108,N_14148);
nor U14268 (N_14268,N_14157,N_14141);
xor U14269 (N_14269,N_14105,N_14119);
nor U14270 (N_14270,N_14211,N_14245);
nand U14271 (N_14271,N_14242,N_14165);
and U14272 (N_14272,N_14215,N_14127);
nand U14273 (N_14273,N_14109,N_14184);
or U14274 (N_14274,N_14118,N_14145);
xnor U14275 (N_14275,N_14143,N_14179);
nor U14276 (N_14276,N_14111,N_14230);
or U14277 (N_14277,N_14212,N_14234);
xnor U14278 (N_14278,N_14209,N_14125);
and U14279 (N_14279,N_14149,N_14208);
or U14280 (N_14280,N_14228,N_14126);
or U14281 (N_14281,N_14158,N_14240);
nor U14282 (N_14282,N_14150,N_14218);
xnor U14283 (N_14283,N_14133,N_14204);
nand U14284 (N_14284,N_14178,N_14112);
or U14285 (N_14285,N_14194,N_14200);
nor U14286 (N_14286,N_14137,N_14110);
xor U14287 (N_14287,N_14185,N_14227);
or U14288 (N_14288,N_14201,N_14183);
xor U14289 (N_14289,N_14160,N_14239);
and U14290 (N_14290,N_14226,N_14229);
nand U14291 (N_14291,N_14151,N_14219);
and U14292 (N_14292,N_14248,N_14162);
xnor U14293 (N_14293,N_14156,N_14221);
or U14294 (N_14294,N_14129,N_14244);
or U14295 (N_14295,N_14216,N_14113);
and U14296 (N_14296,N_14164,N_14210);
nor U14297 (N_14297,N_14224,N_14114);
nor U14298 (N_14298,N_14172,N_14155);
nor U14299 (N_14299,N_14131,N_14198);
nand U14300 (N_14300,N_14167,N_14168);
nor U14301 (N_14301,N_14170,N_14187);
or U14302 (N_14302,N_14190,N_14203);
nor U14303 (N_14303,N_14102,N_14128);
nor U14304 (N_14304,N_14232,N_14199);
nand U14305 (N_14305,N_14124,N_14132);
nand U14306 (N_14306,N_14134,N_14103);
xnor U14307 (N_14307,N_14153,N_14139);
nand U14308 (N_14308,N_14159,N_14135);
or U14309 (N_14309,N_14238,N_14101);
and U14310 (N_14310,N_14177,N_14241);
nor U14311 (N_14311,N_14186,N_14235);
nand U14312 (N_14312,N_14193,N_14247);
or U14313 (N_14313,N_14115,N_14169);
xor U14314 (N_14314,N_14237,N_14206);
xor U14315 (N_14315,N_14120,N_14197);
nor U14316 (N_14316,N_14107,N_14123);
or U14317 (N_14317,N_14243,N_14171);
xnor U14318 (N_14318,N_14106,N_14163);
or U14319 (N_14319,N_14236,N_14217);
nand U14320 (N_14320,N_14173,N_14180);
or U14321 (N_14321,N_14142,N_14116);
xor U14322 (N_14322,N_14182,N_14130);
nor U14323 (N_14323,N_14231,N_14121);
and U14324 (N_14324,N_14205,N_14181);
nand U14325 (N_14325,N_14161,N_14143);
and U14326 (N_14326,N_14166,N_14163);
nor U14327 (N_14327,N_14179,N_14172);
and U14328 (N_14328,N_14104,N_14233);
nand U14329 (N_14329,N_14158,N_14161);
and U14330 (N_14330,N_14114,N_14132);
or U14331 (N_14331,N_14158,N_14230);
nor U14332 (N_14332,N_14188,N_14186);
nor U14333 (N_14333,N_14215,N_14177);
nand U14334 (N_14334,N_14152,N_14172);
nor U14335 (N_14335,N_14170,N_14137);
nand U14336 (N_14336,N_14154,N_14127);
nand U14337 (N_14337,N_14107,N_14147);
nor U14338 (N_14338,N_14134,N_14104);
and U14339 (N_14339,N_14227,N_14178);
nor U14340 (N_14340,N_14216,N_14140);
xor U14341 (N_14341,N_14193,N_14103);
nand U14342 (N_14342,N_14148,N_14165);
and U14343 (N_14343,N_14208,N_14145);
and U14344 (N_14344,N_14209,N_14212);
and U14345 (N_14345,N_14222,N_14231);
and U14346 (N_14346,N_14212,N_14239);
xor U14347 (N_14347,N_14133,N_14101);
and U14348 (N_14348,N_14184,N_14134);
nand U14349 (N_14349,N_14184,N_14228);
or U14350 (N_14350,N_14228,N_14181);
or U14351 (N_14351,N_14231,N_14232);
xor U14352 (N_14352,N_14173,N_14199);
xor U14353 (N_14353,N_14179,N_14116);
nand U14354 (N_14354,N_14143,N_14112);
xnor U14355 (N_14355,N_14196,N_14168);
or U14356 (N_14356,N_14118,N_14124);
xor U14357 (N_14357,N_14142,N_14138);
and U14358 (N_14358,N_14120,N_14224);
nor U14359 (N_14359,N_14194,N_14159);
xnor U14360 (N_14360,N_14202,N_14206);
nor U14361 (N_14361,N_14105,N_14187);
or U14362 (N_14362,N_14111,N_14160);
nor U14363 (N_14363,N_14118,N_14148);
nand U14364 (N_14364,N_14194,N_14186);
and U14365 (N_14365,N_14133,N_14165);
nand U14366 (N_14366,N_14113,N_14150);
xnor U14367 (N_14367,N_14112,N_14120);
or U14368 (N_14368,N_14165,N_14177);
or U14369 (N_14369,N_14185,N_14187);
and U14370 (N_14370,N_14233,N_14116);
nand U14371 (N_14371,N_14128,N_14191);
nand U14372 (N_14372,N_14245,N_14199);
and U14373 (N_14373,N_14111,N_14223);
xnor U14374 (N_14374,N_14203,N_14118);
xnor U14375 (N_14375,N_14160,N_14195);
nor U14376 (N_14376,N_14228,N_14127);
and U14377 (N_14377,N_14133,N_14156);
nand U14378 (N_14378,N_14196,N_14104);
xnor U14379 (N_14379,N_14177,N_14147);
nor U14380 (N_14380,N_14135,N_14148);
nand U14381 (N_14381,N_14230,N_14215);
nand U14382 (N_14382,N_14156,N_14106);
nand U14383 (N_14383,N_14107,N_14135);
nand U14384 (N_14384,N_14104,N_14146);
nor U14385 (N_14385,N_14177,N_14237);
or U14386 (N_14386,N_14122,N_14213);
or U14387 (N_14387,N_14159,N_14187);
nand U14388 (N_14388,N_14112,N_14124);
or U14389 (N_14389,N_14218,N_14204);
xor U14390 (N_14390,N_14232,N_14181);
or U14391 (N_14391,N_14186,N_14202);
and U14392 (N_14392,N_14104,N_14107);
or U14393 (N_14393,N_14223,N_14163);
nand U14394 (N_14394,N_14238,N_14221);
nand U14395 (N_14395,N_14169,N_14154);
xor U14396 (N_14396,N_14236,N_14133);
nor U14397 (N_14397,N_14245,N_14222);
and U14398 (N_14398,N_14233,N_14129);
or U14399 (N_14399,N_14134,N_14219);
nand U14400 (N_14400,N_14392,N_14316);
and U14401 (N_14401,N_14372,N_14260);
and U14402 (N_14402,N_14391,N_14349);
nand U14403 (N_14403,N_14329,N_14394);
nor U14404 (N_14404,N_14359,N_14283);
nand U14405 (N_14405,N_14333,N_14309);
nor U14406 (N_14406,N_14293,N_14371);
and U14407 (N_14407,N_14250,N_14263);
nor U14408 (N_14408,N_14279,N_14314);
and U14409 (N_14409,N_14258,N_14286);
or U14410 (N_14410,N_14395,N_14261);
nor U14411 (N_14411,N_14291,N_14327);
nor U14412 (N_14412,N_14312,N_14364);
or U14413 (N_14413,N_14362,N_14301);
or U14414 (N_14414,N_14389,N_14383);
and U14415 (N_14415,N_14397,N_14377);
nand U14416 (N_14416,N_14320,N_14318);
nor U14417 (N_14417,N_14340,N_14262);
or U14418 (N_14418,N_14330,N_14325);
nor U14419 (N_14419,N_14398,N_14310);
nand U14420 (N_14420,N_14302,N_14341);
or U14421 (N_14421,N_14277,N_14305);
xor U14422 (N_14422,N_14284,N_14274);
nor U14423 (N_14423,N_14254,N_14361);
xor U14424 (N_14424,N_14294,N_14350);
nor U14425 (N_14425,N_14342,N_14307);
and U14426 (N_14426,N_14355,N_14317);
nor U14427 (N_14427,N_14381,N_14255);
xor U14428 (N_14428,N_14267,N_14282);
nand U14429 (N_14429,N_14337,N_14370);
or U14430 (N_14430,N_14272,N_14299);
and U14431 (N_14431,N_14303,N_14360);
nand U14432 (N_14432,N_14311,N_14386);
xor U14433 (N_14433,N_14313,N_14288);
and U14434 (N_14434,N_14353,N_14266);
and U14435 (N_14435,N_14259,N_14376);
nor U14436 (N_14436,N_14382,N_14368);
or U14437 (N_14437,N_14369,N_14332);
nor U14438 (N_14438,N_14315,N_14363);
nand U14439 (N_14439,N_14326,N_14396);
xor U14440 (N_14440,N_14351,N_14345);
or U14441 (N_14441,N_14328,N_14253);
or U14442 (N_14442,N_14264,N_14304);
xor U14443 (N_14443,N_14390,N_14346);
nor U14444 (N_14444,N_14280,N_14335);
xnor U14445 (N_14445,N_14285,N_14297);
or U14446 (N_14446,N_14352,N_14344);
or U14447 (N_14447,N_14324,N_14268);
xnor U14448 (N_14448,N_14323,N_14354);
and U14449 (N_14449,N_14378,N_14269);
and U14450 (N_14450,N_14252,N_14347);
nor U14451 (N_14451,N_14365,N_14290);
nor U14452 (N_14452,N_14399,N_14373);
nor U14453 (N_14453,N_14338,N_14331);
or U14454 (N_14454,N_14256,N_14322);
or U14455 (N_14455,N_14308,N_14393);
xnor U14456 (N_14456,N_14388,N_14380);
and U14457 (N_14457,N_14296,N_14387);
nand U14458 (N_14458,N_14374,N_14357);
and U14459 (N_14459,N_14375,N_14281);
or U14460 (N_14460,N_14343,N_14321);
or U14461 (N_14461,N_14278,N_14379);
or U14462 (N_14462,N_14348,N_14251);
and U14463 (N_14463,N_14384,N_14339);
or U14464 (N_14464,N_14257,N_14273);
xor U14465 (N_14465,N_14271,N_14275);
and U14466 (N_14466,N_14367,N_14358);
or U14467 (N_14467,N_14287,N_14270);
or U14468 (N_14468,N_14265,N_14276);
nor U14469 (N_14469,N_14298,N_14300);
or U14470 (N_14470,N_14319,N_14292);
and U14471 (N_14471,N_14336,N_14295);
or U14472 (N_14472,N_14366,N_14289);
nand U14473 (N_14473,N_14385,N_14334);
and U14474 (N_14474,N_14306,N_14356);
nand U14475 (N_14475,N_14289,N_14365);
or U14476 (N_14476,N_14308,N_14387);
nand U14477 (N_14477,N_14290,N_14278);
nand U14478 (N_14478,N_14362,N_14377);
nand U14479 (N_14479,N_14352,N_14364);
and U14480 (N_14480,N_14266,N_14364);
nand U14481 (N_14481,N_14394,N_14368);
or U14482 (N_14482,N_14330,N_14348);
nand U14483 (N_14483,N_14272,N_14283);
or U14484 (N_14484,N_14356,N_14320);
and U14485 (N_14485,N_14396,N_14392);
nor U14486 (N_14486,N_14319,N_14277);
or U14487 (N_14487,N_14344,N_14295);
and U14488 (N_14488,N_14367,N_14257);
xnor U14489 (N_14489,N_14390,N_14325);
nand U14490 (N_14490,N_14252,N_14281);
xnor U14491 (N_14491,N_14341,N_14373);
nand U14492 (N_14492,N_14395,N_14324);
nand U14493 (N_14493,N_14313,N_14372);
and U14494 (N_14494,N_14399,N_14302);
nor U14495 (N_14495,N_14394,N_14305);
nand U14496 (N_14496,N_14252,N_14304);
and U14497 (N_14497,N_14298,N_14349);
nor U14498 (N_14498,N_14365,N_14338);
or U14499 (N_14499,N_14272,N_14298);
or U14500 (N_14500,N_14335,N_14327);
or U14501 (N_14501,N_14350,N_14348);
xor U14502 (N_14502,N_14295,N_14391);
nor U14503 (N_14503,N_14269,N_14270);
or U14504 (N_14504,N_14325,N_14297);
and U14505 (N_14505,N_14283,N_14260);
and U14506 (N_14506,N_14300,N_14330);
nand U14507 (N_14507,N_14391,N_14252);
nand U14508 (N_14508,N_14326,N_14392);
nand U14509 (N_14509,N_14317,N_14369);
nand U14510 (N_14510,N_14339,N_14281);
or U14511 (N_14511,N_14376,N_14306);
xnor U14512 (N_14512,N_14349,N_14263);
nand U14513 (N_14513,N_14382,N_14285);
and U14514 (N_14514,N_14310,N_14344);
nor U14515 (N_14515,N_14251,N_14325);
and U14516 (N_14516,N_14392,N_14397);
xor U14517 (N_14517,N_14250,N_14271);
nand U14518 (N_14518,N_14308,N_14352);
or U14519 (N_14519,N_14348,N_14311);
and U14520 (N_14520,N_14276,N_14293);
nand U14521 (N_14521,N_14373,N_14355);
xor U14522 (N_14522,N_14388,N_14282);
nand U14523 (N_14523,N_14250,N_14302);
nor U14524 (N_14524,N_14288,N_14300);
nor U14525 (N_14525,N_14302,N_14392);
and U14526 (N_14526,N_14393,N_14310);
or U14527 (N_14527,N_14283,N_14325);
xor U14528 (N_14528,N_14327,N_14348);
and U14529 (N_14529,N_14384,N_14358);
or U14530 (N_14530,N_14333,N_14335);
nand U14531 (N_14531,N_14293,N_14386);
xor U14532 (N_14532,N_14294,N_14290);
nor U14533 (N_14533,N_14386,N_14345);
or U14534 (N_14534,N_14309,N_14315);
nand U14535 (N_14535,N_14383,N_14322);
xnor U14536 (N_14536,N_14283,N_14270);
nor U14537 (N_14537,N_14331,N_14297);
nand U14538 (N_14538,N_14250,N_14379);
nor U14539 (N_14539,N_14266,N_14250);
and U14540 (N_14540,N_14254,N_14331);
nor U14541 (N_14541,N_14335,N_14385);
nor U14542 (N_14542,N_14284,N_14272);
xor U14543 (N_14543,N_14264,N_14259);
or U14544 (N_14544,N_14377,N_14331);
and U14545 (N_14545,N_14334,N_14257);
xnor U14546 (N_14546,N_14258,N_14349);
and U14547 (N_14547,N_14297,N_14373);
xor U14548 (N_14548,N_14367,N_14346);
xnor U14549 (N_14549,N_14391,N_14338);
or U14550 (N_14550,N_14492,N_14503);
nor U14551 (N_14551,N_14514,N_14445);
xor U14552 (N_14552,N_14466,N_14405);
or U14553 (N_14553,N_14528,N_14535);
xor U14554 (N_14554,N_14547,N_14404);
and U14555 (N_14555,N_14447,N_14462);
nand U14556 (N_14556,N_14494,N_14488);
or U14557 (N_14557,N_14434,N_14474);
xor U14558 (N_14558,N_14456,N_14433);
and U14559 (N_14559,N_14448,N_14517);
xnor U14560 (N_14560,N_14450,N_14424);
nor U14561 (N_14561,N_14439,N_14473);
nor U14562 (N_14562,N_14423,N_14435);
nor U14563 (N_14563,N_14507,N_14417);
xor U14564 (N_14564,N_14432,N_14459);
or U14565 (N_14565,N_14512,N_14463);
and U14566 (N_14566,N_14430,N_14486);
nor U14567 (N_14567,N_14478,N_14504);
nand U14568 (N_14568,N_14500,N_14541);
and U14569 (N_14569,N_14443,N_14421);
nor U14570 (N_14570,N_14455,N_14457);
nor U14571 (N_14571,N_14542,N_14436);
or U14572 (N_14572,N_14482,N_14539);
or U14573 (N_14573,N_14511,N_14544);
and U14574 (N_14574,N_14427,N_14526);
nor U14575 (N_14575,N_14529,N_14429);
nand U14576 (N_14576,N_14470,N_14520);
or U14577 (N_14577,N_14549,N_14483);
or U14578 (N_14578,N_14491,N_14468);
nor U14579 (N_14579,N_14460,N_14413);
or U14580 (N_14580,N_14442,N_14425);
nor U14581 (N_14581,N_14431,N_14505);
nor U14582 (N_14582,N_14506,N_14426);
xnor U14583 (N_14583,N_14400,N_14414);
and U14584 (N_14584,N_14411,N_14437);
or U14585 (N_14585,N_14537,N_14403);
and U14586 (N_14586,N_14522,N_14452);
nand U14587 (N_14587,N_14444,N_14484);
nor U14588 (N_14588,N_14408,N_14519);
nand U14589 (N_14589,N_14475,N_14489);
or U14590 (N_14590,N_14485,N_14471);
or U14591 (N_14591,N_14441,N_14438);
and U14592 (N_14592,N_14454,N_14536);
and U14593 (N_14593,N_14497,N_14451);
xor U14594 (N_14594,N_14458,N_14465);
nor U14595 (N_14595,N_14415,N_14487);
nor U14596 (N_14596,N_14513,N_14499);
xor U14597 (N_14597,N_14546,N_14518);
xnor U14598 (N_14598,N_14481,N_14498);
nand U14599 (N_14599,N_14496,N_14510);
nor U14600 (N_14600,N_14502,N_14446);
nand U14601 (N_14601,N_14516,N_14515);
and U14602 (N_14602,N_14472,N_14509);
and U14603 (N_14603,N_14490,N_14467);
nand U14604 (N_14604,N_14495,N_14407);
nor U14605 (N_14605,N_14412,N_14406);
xor U14606 (N_14606,N_14530,N_14538);
nand U14607 (N_14607,N_14480,N_14508);
and U14608 (N_14608,N_14410,N_14543);
xnor U14609 (N_14609,N_14409,N_14461);
nand U14610 (N_14610,N_14469,N_14416);
or U14611 (N_14611,N_14419,N_14476);
nand U14612 (N_14612,N_14453,N_14501);
xnor U14613 (N_14613,N_14428,N_14401);
nand U14614 (N_14614,N_14440,N_14493);
and U14615 (N_14615,N_14531,N_14548);
or U14616 (N_14616,N_14418,N_14479);
or U14617 (N_14617,N_14521,N_14545);
nand U14618 (N_14618,N_14402,N_14449);
nand U14619 (N_14619,N_14534,N_14523);
or U14620 (N_14620,N_14533,N_14525);
and U14621 (N_14621,N_14540,N_14477);
or U14622 (N_14622,N_14527,N_14422);
xnor U14623 (N_14623,N_14464,N_14532);
nor U14624 (N_14624,N_14524,N_14420);
or U14625 (N_14625,N_14488,N_14535);
or U14626 (N_14626,N_14485,N_14533);
nor U14627 (N_14627,N_14489,N_14431);
xnor U14628 (N_14628,N_14411,N_14496);
xor U14629 (N_14629,N_14501,N_14533);
and U14630 (N_14630,N_14491,N_14413);
and U14631 (N_14631,N_14547,N_14420);
and U14632 (N_14632,N_14462,N_14534);
and U14633 (N_14633,N_14521,N_14510);
and U14634 (N_14634,N_14518,N_14465);
nand U14635 (N_14635,N_14528,N_14452);
nor U14636 (N_14636,N_14525,N_14467);
xor U14637 (N_14637,N_14500,N_14548);
or U14638 (N_14638,N_14491,N_14428);
or U14639 (N_14639,N_14535,N_14426);
nor U14640 (N_14640,N_14537,N_14520);
and U14641 (N_14641,N_14466,N_14481);
nor U14642 (N_14642,N_14477,N_14486);
xnor U14643 (N_14643,N_14432,N_14497);
and U14644 (N_14644,N_14540,N_14451);
xnor U14645 (N_14645,N_14454,N_14418);
nand U14646 (N_14646,N_14428,N_14472);
nand U14647 (N_14647,N_14481,N_14530);
xnor U14648 (N_14648,N_14493,N_14535);
nor U14649 (N_14649,N_14412,N_14485);
nand U14650 (N_14650,N_14438,N_14541);
nor U14651 (N_14651,N_14528,N_14512);
or U14652 (N_14652,N_14544,N_14480);
nand U14653 (N_14653,N_14490,N_14481);
or U14654 (N_14654,N_14511,N_14512);
or U14655 (N_14655,N_14466,N_14424);
or U14656 (N_14656,N_14412,N_14454);
nand U14657 (N_14657,N_14528,N_14504);
nor U14658 (N_14658,N_14541,N_14489);
xor U14659 (N_14659,N_14423,N_14542);
xnor U14660 (N_14660,N_14454,N_14533);
and U14661 (N_14661,N_14402,N_14494);
nand U14662 (N_14662,N_14499,N_14474);
xnor U14663 (N_14663,N_14457,N_14438);
nand U14664 (N_14664,N_14528,N_14505);
or U14665 (N_14665,N_14404,N_14473);
or U14666 (N_14666,N_14425,N_14426);
or U14667 (N_14667,N_14450,N_14425);
nor U14668 (N_14668,N_14528,N_14405);
xor U14669 (N_14669,N_14541,N_14414);
nand U14670 (N_14670,N_14465,N_14489);
xor U14671 (N_14671,N_14446,N_14462);
xor U14672 (N_14672,N_14408,N_14452);
nor U14673 (N_14673,N_14487,N_14481);
xor U14674 (N_14674,N_14539,N_14461);
and U14675 (N_14675,N_14400,N_14517);
nand U14676 (N_14676,N_14463,N_14452);
xnor U14677 (N_14677,N_14435,N_14434);
or U14678 (N_14678,N_14474,N_14539);
nor U14679 (N_14679,N_14487,N_14515);
or U14680 (N_14680,N_14441,N_14546);
or U14681 (N_14681,N_14519,N_14545);
or U14682 (N_14682,N_14449,N_14521);
or U14683 (N_14683,N_14488,N_14418);
nand U14684 (N_14684,N_14451,N_14454);
or U14685 (N_14685,N_14410,N_14537);
or U14686 (N_14686,N_14519,N_14532);
nand U14687 (N_14687,N_14441,N_14425);
and U14688 (N_14688,N_14495,N_14489);
or U14689 (N_14689,N_14444,N_14538);
nor U14690 (N_14690,N_14530,N_14541);
xor U14691 (N_14691,N_14476,N_14543);
and U14692 (N_14692,N_14533,N_14497);
and U14693 (N_14693,N_14530,N_14413);
nor U14694 (N_14694,N_14403,N_14491);
and U14695 (N_14695,N_14459,N_14446);
nand U14696 (N_14696,N_14492,N_14531);
nor U14697 (N_14697,N_14527,N_14473);
xor U14698 (N_14698,N_14447,N_14533);
nor U14699 (N_14699,N_14452,N_14409);
or U14700 (N_14700,N_14662,N_14606);
xor U14701 (N_14701,N_14660,N_14692);
nand U14702 (N_14702,N_14690,N_14643);
xor U14703 (N_14703,N_14614,N_14580);
or U14704 (N_14704,N_14619,N_14584);
or U14705 (N_14705,N_14626,N_14563);
xnor U14706 (N_14706,N_14671,N_14616);
or U14707 (N_14707,N_14665,N_14551);
or U14708 (N_14708,N_14659,N_14674);
and U14709 (N_14709,N_14646,N_14586);
nor U14710 (N_14710,N_14581,N_14676);
or U14711 (N_14711,N_14603,N_14657);
nand U14712 (N_14712,N_14589,N_14558);
nand U14713 (N_14713,N_14684,N_14651);
nand U14714 (N_14714,N_14573,N_14639);
and U14715 (N_14715,N_14645,N_14661);
nor U14716 (N_14716,N_14695,N_14561);
nand U14717 (N_14717,N_14680,N_14585);
and U14718 (N_14718,N_14594,N_14569);
and U14719 (N_14719,N_14649,N_14673);
or U14720 (N_14720,N_14636,N_14620);
nand U14721 (N_14721,N_14608,N_14553);
xor U14722 (N_14722,N_14596,N_14679);
nor U14723 (N_14723,N_14567,N_14693);
and U14724 (N_14724,N_14562,N_14559);
and U14725 (N_14725,N_14611,N_14654);
nand U14726 (N_14726,N_14655,N_14642);
and U14727 (N_14727,N_14658,N_14622);
nand U14728 (N_14728,N_14572,N_14628);
nor U14729 (N_14729,N_14637,N_14688);
or U14730 (N_14730,N_14578,N_14554);
nand U14731 (N_14731,N_14579,N_14587);
or U14732 (N_14732,N_14564,N_14598);
or U14733 (N_14733,N_14550,N_14565);
xor U14734 (N_14734,N_14666,N_14650);
and U14735 (N_14735,N_14670,N_14597);
and U14736 (N_14736,N_14689,N_14566);
or U14737 (N_14737,N_14691,N_14610);
nor U14738 (N_14738,N_14568,N_14571);
nor U14739 (N_14739,N_14555,N_14678);
xnor U14740 (N_14740,N_14602,N_14683);
xnor U14741 (N_14741,N_14682,N_14618);
nor U14742 (N_14742,N_14648,N_14699);
nor U14743 (N_14743,N_14686,N_14574);
nor U14744 (N_14744,N_14604,N_14615);
nand U14745 (N_14745,N_14590,N_14640);
or U14746 (N_14746,N_14698,N_14656);
nand U14747 (N_14747,N_14599,N_14627);
and U14748 (N_14748,N_14576,N_14638);
and U14749 (N_14749,N_14623,N_14663);
xor U14750 (N_14750,N_14668,N_14644);
nor U14751 (N_14751,N_14633,N_14591);
nor U14752 (N_14752,N_14592,N_14617);
or U14753 (N_14753,N_14612,N_14630);
and U14754 (N_14754,N_14556,N_14647);
and U14755 (N_14755,N_14687,N_14607);
xor U14756 (N_14756,N_14557,N_14588);
or U14757 (N_14757,N_14624,N_14672);
nand U14758 (N_14758,N_14675,N_14583);
nand U14759 (N_14759,N_14696,N_14601);
or U14760 (N_14760,N_14664,N_14641);
xnor U14761 (N_14761,N_14582,N_14609);
xnor U14762 (N_14762,N_14575,N_14653);
and U14763 (N_14763,N_14694,N_14613);
and U14764 (N_14764,N_14667,N_14621);
nor U14765 (N_14765,N_14595,N_14570);
xor U14766 (N_14766,N_14697,N_14560);
xor U14767 (N_14767,N_14631,N_14634);
or U14768 (N_14768,N_14669,N_14593);
or U14769 (N_14769,N_14605,N_14552);
nor U14770 (N_14770,N_14685,N_14625);
nor U14771 (N_14771,N_14677,N_14652);
and U14772 (N_14772,N_14629,N_14600);
xor U14773 (N_14773,N_14577,N_14635);
nand U14774 (N_14774,N_14632,N_14681);
nor U14775 (N_14775,N_14612,N_14575);
nor U14776 (N_14776,N_14670,N_14666);
or U14777 (N_14777,N_14565,N_14606);
nor U14778 (N_14778,N_14583,N_14681);
nor U14779 (N_14779,N_14585,N_14554);
or U14780 (N_14780,N_14649,N_14590);
nand U14781 (N_14781,N_14688,N_14569);
nor U14782 (N_14782,N_14659,N_14633);
nor U14783 (N_14783,N_14658,N_14567);
xnor U14784 (N_14784,N_14686,N_14585);
nor U14785 (N_14785,N_14656,N_14663);
nor U14786 (N_14786,N_14659,N_14613);
nor U14787 (N_14787,N_14622,N_14580);
xnor U14788 (N_14788,N_14596,N_14604);
or U14789 (N_14789,N_14592,N_14650);
xor U14790 (N_14790,N_14632,N_14604);
xor U14791 (N_14791,N_14633,N_14558);
nor U14792 (N_14792,N_14603,N_14590);
nand U14793 (N_14793,N_14562,N_14659);
nor U14794 (N_14794,N_14608,N_14685);
xnor U14795 (N_14795,N_14667,N_14647);
nand U14796 (N_14796,N_14666,N_14602);
nor U14797 (N_14797,N_14630,N_14584);
and U14798 (N_14798,N_14564,N_14607);
nor U14799 (N_14799,N_14623,N_14560);
and U14800 (N_14800,N_14625,N_14658);
nand U14801 (N_14801,N_14676,N_14584);
and U14802 (N_14802,N_14574,N_14580);
nor U14803 (N_14803,N_14599,N_14682);
xnor U14804 (N_14804,N_14638,N_14697);
and U14805 (N_14805,N_14658,N_14615);
or U14806 (N_14806,N_14616,N_14591);
or U14807 (N_14807,N_14698,N_14610);
xor U14808 (N_14808,N_14690,N_14695);
nand U14809 (N_14809,N_14578,N_14584);
nor U14810 (N_14810,N_14625,N_14639);
or U14811 (N_14811,N_14565,N_14560);
xor U14812 (N_14812,N_14616,N_14643);
and U14813 (N_14813,N_14626,N_14650);
xor U14814 (N_14814,N_14663,N_14574);
or U14815 (N_14815,N_14601,N_14614);
xnor U14816 (N_14816,N_14632,N_14624);
xor U14817 (N_14817,N_14693,N_14564);
and U14818 (N_14818,N_14628,N_14588);
nor U14819 (N_14819,N_14675,N_14593);
nand U14820 (N_14820,N_14699,N_14665);
or U14821 (N_14821,N_14631,N_14598);
xnor U14822 (N_14822,N_14551,N_14614);
and U14823 (N_14823,N_14660,N_14583);
nor U14824 (N_14824,N_14616,N_14623);
xor U14825 (N_14825,N_14572,N_14583);
nand U14826 (N_14826,N_14664,N_14575);
and U14827 (N_14827,N_14576,N_14596);
nor U14828 (N_14828,N_14663,N_14622);
xnor U14829 (N_14829,N_14571,N_14666);
xor U14830 (N_14830,N_14568,N_14586);
or U14831 (N_14831,N_14616,N_14583);
xor U14832 (N_14832,N_14680,N_14608);
nand U14833 (N_14833,N_14573,N_14567);
or U14834 (N_14834,N_14656,N_14612);
xor U14835 (N_14835,N_14628,N_14664);
nor U14836 (N_14836,N_14552,N_14604);
or U14837 (N_14837,N_14603,N_14684);
nor U14838 (N_14838,N_14587,N_14588);
nand U14839 (N_14839,N_14628,N_14695);
nor U14840 (N_14840,N_14626,N_14555);
nor U14841 (N_14841,N_14691,N_14676);
nor U14842 (N_14842,N_14561,N_14577);
and U14843 (N_14843,N_14681,N_14697);
nor U14844 (N_14844,N_14640,N_14621);
nor U14845 (N_14845,N_14613,N_14550);
or U14846 (N_14846,N_14614,N_14637);
xor U14847 (N_14847,N_14659,N_14615);
and U14848 (N_14848,N_14567,N_14581);
nand U14849 (N_14849,N_14566,N_14635);
xnor U14850 (N_14850,N_14749,N_14755);
or U14851 (N_14851,N_14779,N_14747);
nor U14852 (N_14852,N_14744,N_14740);
and U14853 (N_14853,N_14772,N_14841);
nand U14854 (N_14854,N_14845,N_14806);
nor U14855 (N_14855,N_14801,N_14726);
and U14856 (N_14856,N_14708,N_14762);
and U14857 (N_14857,N_14736,N_14798);
and U14858 (N_14858,N_14847,N_14788);
or U14859 (N_14859,N_14713,N_14836);
and U14860 (N_14860,N_14700,N_14828);
and U14861 (N_14861,N_14840,N_14827);
nand U14862 (N_14862,N_14838,N_14730);
nand U14863 (N_14863,N_14725,N_14831);
and U14864 (N_14864,N_14712,N_14792);
and U14865 (N_14865,N_14705,N_14748);
nor U14866 (N_14866,N_14818,N_14820);
nor U14867 (N_14867,N_14751,N_14797);
nand U14868 (N_14868,N_14848,N_14727);
and U14869 (N_14869,N_14791,N_14701);
nor U14870 (N_14870,N_14724,N_14813);
nand U14871 (N_14871,N_14812,N_14821);
nand U14872 (N_14872,N_14750,N_14768);
and U14873 (N_14873,N_14711,N_14731);
and U14874 (N_14874,N_14834,N_14765);
nor U14875 (N_14875,N_14829,N_14769);
and U14876 (N_14876,N_14849,N_14719);
and U14877 (N_14877,N_14710,N_14810);
or U14878 (N_14878,N_14781,N_14787);
and U14879 (N_14879,N_14775,N_14824);
or U14880 (N_14880,N_14830,N_14763);
nor U14881 (N_14881,N_14739,N_14833);
xor U14882 (N_14882,N_14745,N_14837);
or U14883 (N_14883,N_14816,N_14702);
or U14884 (N_14884,N_14843,N_14716);
nor U14885 (N_14885,N_14799,N_14789);
or U14886 (N_14886,N_14814,N_14774);
nand U14887 (N_14887,N_14786,N_14709);
or U14888 (N_14888,N_14807,N_14790);
and U14889 (N_14889,N_14839,N_14728);
or U14890 (N_14890,N_14793,N_14796);
and U14891 (N_14891,N_14735,N_14817);
xnor U14892 (N_14892,N_14770,N_14720);
or U14893 (N_14893,N_14783,N_14771);
nor U14894 (N_14894,N_14723,N_14732);
or U14895 (N_14895,N_14803,N_14800);
nor U14896 (N_14896,N_14760,N_14844);
nand U14897 (N_14897,N_14707,N_14784);
nor U14898 (N_14898,N_14729,N_14823);
nor U14899 (N_14899,N_14756,N_14778);
xor U14900 (N_14900,N_14795,N_14822);
or U14901 (N_14901,N_14802,N_14846);
nor U14902 (N_14902,N_14804,N_14752);
and U14903 (N_14903,N_14805,N_14780);
or U14904 (N_14904,N_14815,N_14706);
nor U14905 (N_14905,N_14776,N_14741);
nand U14906 (N_14906,N_14826,N_14809);
xor U14907 (N_14907,N_14704,N_14754);
nor U14908 (N_14908,N_14773,N_14832);
nor U14909 (N_14909,N_14738,N_14718);
xor U14910 (N_14910,N_14764,N_14746);
and U14911 (N_14911,N_14766,N_14758);
xnor U14912 (N_14912,N_14722,N_14737);
or U14913 (N_14913,N_14703,N_14753);
nor U14914 (N_14914,N_14794,N_14825);
or U14915 (N_14915,N_14734,N_14742);
nand U14916 (N_14916,N_14819,N_14757);
xor U14917 (N_14917,N_14842,N_14759);
xor U14918 (N_14918,N_14714,N_14808);
nand U14919 (N_14919,N_14785,N_14767);
and U14920 (N_14920,N_14715,N_14733);
or U14921 (N_14921,N_14777,N_14761);
or U14922 (N_14922,N_14811,N_14721);
nor U14923 (N_14923,N_14743,N_14835);
and U14924 (N_14924,N_14717,N_14782);
and U14925 (N_14925,N_14706,N_14756);
nand U14926 (N_14926,N_14840,N_14708);
or U14927 (N_14927,N_14827,N_14730);
nand U14928 (N_14928,N_14797,N_14796);
nand U14929 (N_14929,N_14821,N_14700);
xor U14930 (N_14930,N_14716,N_14805);
nor U14931 (N_14931,N_14772,N_14760);
nor U14932 (N_14932,N_14781,N_14720);
or U14933 (N_14933,N_14831,N_14744);
and U14934 (N_14934,N_14830,N_14701);
nor U14935 (N_14935,N_14801,N_14838);
or U14936 (N_14936,N_14778,N_14847);
xor U14937 (N_14937,N_14742,N_14809);
or U14938 (N_14938,N_14805,N_14708);
xor U14939 (N_14939,N_14804,N_14763);
and U14940 (N_14940,N_14793,N_14783);
nand U14941 (N_14941,N_14792,N_14703);
nor U14942 (N_14942,N_14760,N_14804);
xor U14943 (N_14943,N_14788,N_14758);
or U14944 (N_14944,N_14741,N_14794);
or U14945 (N_14945,N_14824,N_14713);
or U14946 (N_14946,N_14807,N_14734);
or U14947 (N_14947,N_14776,N_14718);
xor U14948 (N_14948,N_14840,N_14742);
nand U14949 (N_14949,N_14766,N_14775);
xor U14950 (N_14950,N_14722,N_14787);
nor U14951 (N_14951,N_14715,N_14812);
or U14952 (N_14952,N_14829,N_14846);
nand U14953 (N_14953,N_14724,N_14799);
and U14954 (N_14954,N_14822,N_14826);
or U14955 (N_14955,N_14769,N_14726);
nand U14956 (N_14956,N_14825,N_14751);
or U14957 (N_14957,N_14822,N_14839);
or U14958 (N_14958,N_14776,N_14711);
or U14959 (N_14959,N_14757,N_14709);
nor U14960 (N_14960,N_14794,N_14728);
and U14961 (N_14961,N_14735,N_14700);
nor U14962 (N_14962,N_14716,N_14813);
nor U14963 (N_14963,N_14717,N_14768);
nor U14964 (N_14964,N_14718,N_14816);
or U14965 (N_14965,N_14825,N_14732);
xor U14966 (N_14966,N_14840,N_14716);
or U14967 (N_14967,N_14813,N_14814);
nor U14968 (N_14968,N_14749,N_14797);
nand U14969 (N_14969,N_14799,N_14759);
xor U14970 (N_14970,N_14839,N_14793);
nor U14971 (N_14971,N_14791,N_14798);
xnor U14972 (N_14972,N_14819,N_14738);
or U14973 (N_14973,N_14800,N_14830);
or U14974 (N_14974,N_14814,N_14810);
xnor U14975 (N_14975,N_14719,N_14724);
nand U14976 (N_14976,N_14807,N_14834);
or U14977 (N_14977,N_14811,N_14784);
xor U14978 (N_14978,N_14823,N_14812);
and U14979 (N_14979,N_14811,N_14749);
nand U14980 (N_14980,N_14735,N_14740);
nand U14981 (N_14981,N_14756,N_14745);
nand U14982 (N_14982,N_14759,N_14780);
nor U14983 (N_14983,N_14811,N_14782);
nor U14984 (N_14984,N_14778,N_14824);
xor U14985 (N_14985,N_14727,N_14833);
or U14986 (N_14986,N_14834,N_14791);
nor U14987 (N_14987,N_14784,N_14741);
xnor U14988 (N_14988,N_14754,N_14723);
or U14989 (N_14989,N_14710,N_14753);
xnor U14990 (N_14990,N_14736,N_14793);
or U14991 (N_14991,N_14727,N_14829);
or U14992 (N_14992,N_14759,N_14760);
nand U14993 (N_14993,N_14821,N_14785);
and U14994 (N_14994,N_14716,N_14812);
nand U14995 (N_14995,N_14711,N_14728);
and U14996 (N_14996,N_14714,N_14785);
nand U14997 (N_14997,N_14803,N_14819);
or U14998 (N_14998,N_14793,N_14823);
nor U14999 (N_14999,N_14751,N_14739);
xnor UO_0 (O_0,N_14917,N_14981);
nand UO_1 (O_1,N_14923,N_14915);
nor UO_2 (O_2,N_14999,N_14956);
nand UO_3 (O_3,N_14871,N_14980);
nor UO_4 (O_4,N_14870,N_14960);
nand UO_5 (O_5,N_14951,N_14899);
and UO_6 (O_6,N_14907,N_14931);
nand UO_7 (O_7,N_14942,N_14856);
and UO_8 (O_8,N_14912,N_14983);
and UO_9 (O_9,N_14932,N_14987);
and UO_10 (O_10,N_14922,N_14892);
nor UO_11 (O_11,N_14853,N_14862);
nand UO_12 (O_12,N_14945,N_14865);
or UO_13 (O_13,N_14860,N_14926);
or UO_14 (O_14,N_14969,N_14888);
nand UO_15 (O_15,N_14934,N_14995);
nand UO_16 (O_16,N_14974,N_14978);
nor UO_17 (O_17,N_14877,N_14894);
and UO_18 (O_18,N_14982,N_14873);
nor UO_19 (O_19,N_14906,N_14867);
nand UO_20 (O_20,N_14954,N_14971);
nor UO_21 (O_21,N_14891,N_14869);
or UO_22 (O_22,N_14903,N_14916);
and UO_23 (O_23,N_14927,N_14882);
nor UO_24 (O_24,N_14904,N_14879);
nor UO_25 (O_25,N_14959,N_14929);
and UO_26 (O_26,N_14878,N_14962);
xor UO_27 (O_27,N_14925,N_14943);
nand UO_28 (O_28,N_14985,N_14998);
and UO_29 (O_29,N_14898,N_14957);
nor UO_30 (O_30,N_14914,N_14857);
nor UO_31 (O_31,N_14941,N_14940);
or UO_32 (O_32,N_14970,N_14855);
nand UO_33 (O_33,N_14972,N_14893);
nor UO_34 (O_34,N_14852,N_14947);
nand UO_35 (O_35,N_14919,N_14868);
nand UO_36 (O_36,N_14949,N_14986);
or UO_37 (O_37,N_14886,N_14938);
xor UO_38 (O_38,N_14897,N_14890);
and UO_39 (O_39,N_14876,N_14953);
nor UO_40 (O_40,N_14885,N_14850);
or UO_41 (O_41,N_14968,N_14939);
and UO_42 (O_42,N_14920,N_14863);
nor UO_43 (O_43,N_14997,N_14921);
xor UO_44 (O_44,N_14875,N_14918);
nand UO_45 (O_45,N_14965,N_14859);
or UO_46 (O_46,N_14909,N_14900);
nand UO_47 (O_47,N_14889,N_14901);
nand UO_48 (O_48,N_14977,N_14988);
nor UO_49 (O_49,N_14861,N_14944);
or UO_50 (O_50,N_14880,N_14854);
and UO_51 (O_51,N_14866,N_14924);
or UO_52 (O_52,N_14884,N_14992);
nor UO_53 (O_53,N_14930,N_14973);
and UO_54 (O_54,N_14976,N_14896);
nor UO_55 (O_55,N_14955,N_14961);
nand UO_56 (O_56,N_14948,N_14887);
nand UO_57 (O_57,N_14958,N_14881);
xor UO_58 (O_58,N_14975,N_14883);
or UO_59 (O_59,N_14946,N_14990);
nor UO_60 (O_60,N_14911,N_14913);
nor UO_61 (O_61,N_14936,N_14935);
and UO_62 (O_62,N_14872,N_14864);
and UO_63 (O_63,N_14874,N_14908);
and UO_64 (O_64,N_14950,N_14905);
nor UO_65 (O_65,N_14964,N_14910);
nor UO_66 (O_66,N_14933,N_14996);
and UO_67 (O_67,N_14858,N_14994);
nor UO_68 (O_68,N_14902,N_14993);
nand UO_69 (O_69,N_14895,N_14991);
nor UO_70 (O_70,N_14851,N_14966);
and UO_71 (O_71,N_14967,N_14963);
or UO_72 (O_72,N_14984,N_14937);
xnor UO_73 (O_73,N_14928,N_14979);
nor UO_74 (O_74,N_14989,N_14952);
nor UO_75 (O_75,N_14853,N_14999);
and UO_76 (O_76,N_14887,N_14913);
and UO_77 (O_77,N_14970,N_14912);
or UO_78 (O_78,N_14888,N_14885);
or UO_79 (O_79,N_14931,N_14877);
xnor UO_80 (O_80,N_14892,N_14901);
xor UO_81 (O_81,N_14858,N_14936);
and UO_82 (O_82,N_14933,N_14926);
nand UO_83 (O_83,N_14953,N_14909);
nand UO_84 (O_84,N_14944,N_14924);
or UO_85 (O_85,N_14890,N_14886);
and UO_86 (O_86,N_14973,N_14881);
or UO_87 (O_87,N_14895,N_14933);
xnor UO_88 (O_88,N_14943,N_14890);
or UO_89 (O_89,N_14948,N_14860);
xnor UO_90 (O_90,N_14940,N_14926);
xor UO_91 (O_91,N_14966,N_14900);
nor UO_92 (O_92,N_14942,N_14935);
xnor UO_93 (O_93,N_14916,N_14973);
xnor UO_94 (O_94,N_14926,N_14886);
xnor UO_95 (O_95,N_14880,N_14970);
xor UO_96 (O_96,N_14877,N_14907);
nand UO_97 (O_97,N_14950,N_14855);
xor UO_98 (O_98,N_14872,N_14885);
or UO_99 (O_99,N_14914,N_14919);
and UO_100 (O_100,N_14897,N_14973);
nor UO_101 (O_101,N_14909,N_14884);
or UO_102 (O_102,N_14927,N_14938);
or UO_103 (O_103,N_14933,N_14976);
and UO_104 (O_104,N_14939,N_14938);
nand UO_105 (O_105,N_14946,N_14855);
nor UO_106 (O_106,N_14979,N_14927);
nand UO_107 (O_107,N_14868,N_14892);
or UO_108 (O_108,N_14896,N_14879);
xnor UO_109 (O_109,N_14997,N_14966);
and UO_110 (O_110,N_14919,N_14918);
or UO_111 (O_111,N_14998,N_14971);
nand UO_112 (O_112,N_14952,N_14945);
nand UO_113 (O_113,N_14890,N_14966);
xnor UO_114 (O_114,N_14967,N_14995);
xnor UO_115 (O_115,N_14881,N_14884);
nor UO_116 (O_116,N_14941,N_14993);
and UO_117 (O_117,N_14900,N_14919);
nor UO_118 (O_118,N_14915,N_14949);
xor UO_119 (O_119,N_14992,N_14909);
xnor UO_120 (O_120,N_14914,N_14931);
nand UO_121 (O_121,N_14985,N_14991);
nor UO_122 (O_122,N_14862,N_14978);
nor UO_123 (O_123,N_14947,N_14949);
and UO_124 (O_124,N_14897,N_14980);
nand UO_125 (O_125,N_14912,N_14879);
nand UO_126 (O_126,N_14916,N_14963);
and UO_127 (O_127,N_14893,N_14878);
xor UO_128 (O_128,N_14891,N_14996);
nor UO_129 (O_129,N_14924,N_14869);
or UO_130 (O_130,N_14951,N_14941);
or UO_131 (O_131,N_14875,N_14900);
or UO_132 (O_132,N_14881,N_14907);
nor UO_133 (O_133,N_14966,N_14930);
and UO_134 (O_134,N_14858,N_14953);
or UO_135 (O_135,N_14949,N_14858);
nor UO_136 (O_136,N_14989,N_14963);
or UO_137 (O_137,N_14879,N_14935);
xnor UO_138 (O_138,N_14909,N_14930);
or UO_139 (O_139,N_14928,N_14980);
or UO_140 (O_140,N_14990,N_14866);
and UO_141 (O_141,N_14897,N_14866);
xnor UO_142 (O_142,N_14880,N_14893);
or UO_143 (O_143,N_14881,N_14964);
and UO_144 (O_144,N_14985,N_14999);
xnor UO_145 (O_145,N_14976,N_14917);
xor UO_146 (O_146,N_14882,N_14946);
or UO_147 (O_147,N_14988,N_14950);
or UO_148 (O_148,N_14854,N_14863);
or UO_149 (O_149,N_14948,N_14933);
or UO_150 (O_150,N_14923,N_14940);
nand UO_151 (O_151,N_14956,N_14925);
nor UO_152 (O_152,N_14871,N_14885);
nor UO_153 (O_153,N_14989,N_14973);
xor UO_154 (O_154,N_14920,N_14861);
and UO_155 (O_155,N_14949,N_14860);
and UO_156 (O_156,N_14949,N_14981);
nand UO_157 (O_157,N_14994,N_14879);
nand UO_158 (O_158,N_14873,N_14891);
and UO_159 (O_159,N_14918,N_14923);
and UO_160 (O_160,N_14862,N_14901);
nand UO_161 (O_161,N_14991,N_14973);
xor UO_162 (O_162,N_14957,N_14964);
nor UO_163 (O_163,N_14870,N_14979);
or UO_164 (O_164,N_14935,N_14975);
or UO_165 (O_165,N_14995,N_14997);
xnor UO_166 (O_166,N_14890,N_14923);
nor UO_167 (O_167,N_14965,N_14870);
nand UO_168 (O_168,N_14861,N_14943);
nor UO_169 (O_169,N_14984,N_14919);
or UO_170 (O_170,N_14936,N_14954);
nand UO_171 (O_171,N_14899,N_14904);
and UO_172 (O_172,N_14879,N_14961);
and UO_173 (O_173,N_14891,N_14999);
nor UO_174 (O_174,N_14895,N_14988);
nor UO_175 (O_175,N_14974,N_14873);
xor UO_176 (O_176,N_14957,N_14877);
or UO_177 (O_177,N_14976,N_14975);
or UO_178 (O_178,N_14973,N_14867);
nor UO_179 (O_179,N_14896,N_14949);
and UO_180 (O_180,N_14936,N_14963);
xor UO_181 (O_181,N_14965,N_14856);
or UO_182 (O_182,N_14906,N_14925);
nand UO_183 (O_183,N_14906,N_14889);
or UO_184 (O_184,N_14919,N_14877);
or UO_185 (O_185,N_14853,N_14886);
xnor UO_186 (O_186,N_14986,N_14852);
nand UO_187 (O_187,N_14985,N_14883);
and UO_188 (O_188,N_14862,N_14924);
xor UO_189 (O_189,N_14992,N_14899);
nand UO_190 (O_190,N_14938,N_14903);
xnor UO_191 (O_191,N_14981,N_14979);
nand UO_192 (O_192,N_14896,N_14920);
xnor UO_193 (O_193,N_14932,N_14964);
nand UO_194 (O_194,N_14864,N_14970);
nand UO_195 (O_195,N_14914,N_14887);
nand UO_196 (O_196,N_14976,N_14993);
or UO_197 (O_197,N_14920,N_14901);
and UO_198 (O_198,N_14918,N_14880);
xnor UO_199 (O_199,N_14893,N_14886);
and UO_200 (O_200,N_14964,N_14959);
or UO_201 (O_201,N_14944,N_14936);
and UO_202 (O_202,N_14939,N_14995);
xor UO_203 (O_203,N_14872,N_14981);
nor UO_204 (O_204,N_14951,N_14908);
nand UO_205 (O_205,N_14934,N_14987);
and UO_206 (O_206,N_14892,N_14969);
xnor UO_207 (O_207,N_14889,N_14854);
or UO_208 (O_208,N_14978,N_14877);
nand UO_209 (O_209,N_14929,N_14967);
xor UO_210 (O_210,N_14966,N_14914);
or UO_211 (O_211,N_14939,N_14866);
and UO_212 (O_212,N_14981,N_14863);
xnor UO_213 (O_213,N_14963,N_14996);
and UO_214 (O_214,N_14939,N_14894);
xnor UO_215 (O_215,N_14861,N_14901);
xnor UO_216 (O_216,N_14860,N_14913);
xor UO_217 (O_217,N_14916,N_14930);
and UO_218 (O_218,N_14983,N_14953);
nor UO_219 (O_219,N_14861,N_14993);
and UO_220 (O_220,N_14930,N_14956);
nand UO_221 (O_221,N_14906,N_14880);
or UO_222 (O_222,N_14979,N_14942);
xnor UO_223 (O_223,N_14914,N_14869);
xnor UO_224 (O_224,N_14853,N_14952);
nor UO_225 (O_225,N_14911,N_14992);
and UO_226 (O_226,N_14942,N_14923);
nor UO_227 (O_227,N_14902,N_14956);
and UO_228 (O_228,N_14949,N_14926);
and UO_229 (O_229,N_14950,N_14963);
nand UO_230 (O_230,N_14949,N_14907);
or UO_231 (O_231,N_14905,N_14923);
nor UO_232 (O_232,N_14914,N_14970);
nor UO_233 (O_233,N_14926,N_14956);
nor UO_234 (O_234,N_14952,N_14997);
nand UO_235 (O_235,N_14900,N_14874);
xnor UO_236 (O_236,N_14865,N_14857);
and UO_237 (O_237,N_14953,N_14899);
nor UO_238 (O_238,N_14893,N_14990);
or UO_239 (O_239,N_14893,N_14966);
nand UO_240 (O_240,N_14866,N_14865);
nor UO_241 (O_241,N_14890,N_14972);
nor UO_242 (O_242,N_14995,N_14941);
nand UO_243 (O_243,N_14974,N_14979);
nand UO_244 (O_244,N_14905,N_14912);
nor UO_245 (O_245,N_14923,N_14999);
and UO_246 (O_246,N_14872,N_14994);
and UO_247 (O_247,N_14852,N_14856);
xor UO_248 (O_248,N_14984,N_14936);
nor UO_249 (O_249,N_14919,N_14983);
nand UO_250 (O_250,N_14850,N_14870);
nand UO_251 (O_251,N_14969,N_14883);
xor UO_252 (O_252,N_14870,N_14974);
or UO_253 (O_253,N_14909,N_14893);
nand UO_254 (O_254,N_14902,N_14863);
nand UO_255 (O_255,N_14898,N_14976);
xor UO_256 (O_256,N_14988,N_14931);
or UO_257 (O_257,N_14939,N_14914);
or UO_258 (O_258,N_14966,N_14905);
and UO_259 (O_259,N_14931,N_14985);
nor UO_260 (O_260,N_14851,N_14981);
and UO_261 (O_261,N_14928,N_14944);
or UO_262 (O_262,N_14984,N_14914);
and UO_263 (O_263,N_14925,N_14901);
nand UO_264 (O_264,N_14951,N_14853);
xor UO_265 (O_265,N_14994,N_14982);
and UO_266 (O_266,N_14911,N_14884);
and UO_267 (O_267,N_14987,N_14956);
xnor UO_268 (O_268,N_14987,N_14997);
and UO_269 (O_269,N_14859,N_14935);
xnor UO_270 (O_270,N_14891,N_14852);
nor UO_271 (O_271,N_14942,N_14851);
or UO_272 (O_272,N_14912,N_14951);
nand UO_273 (O_273,N_14868,N_14890);
nor UO_274 (O_274,N_14932,N_14851);
xor UO_275 (O_275,N_14884,N_14998);
xnor UO_276 (O_276,N_14997,N_14958);
nand UO_277 (O_277,N_14993,N_14874);
xor UO_278 (O_278,N_14969,N_14912);
and UO_279 (O_279,N_14860,N_14875);
nor UO_280 (O_280,N_14862,N_14982);
nand UO_281 (O_281,N_14877,N_14930);
and UO_282 (O_282,N_14911,N_14891);
and UO_283 (O_283,N_14890,N_14957);
nor UO_284 (O_284,N_14886,N_14900);
nand UO_285 (O_285,N_14998,N_14917);
xor UO_286 (O_286,N_14981,N_14980);
or UO_287 (O_287,N_14986,N_14895);
or UO_288 (O_288,N_14924,N_14945);
and UO_289 (O_289,N_14886,N_14915);
or UO_290 (O_290,N_14946,N_14889);
and UO_291 (O_291,N_14972,N_14958);
xor UO_292 (O_292,N_14962,N_14871);
nand UO_293 (O_293,N_14882,N_14856);
or UO_294 (O_294,N_14903,N_14904);
or UO_295 (O_295,N_14939,N_14870);
nor UO_296 (O_296,N_14908,N_14990);
nand UO_297 (O_297,N_14952,N_14983);
nor UO_298 (O_298,N_14991,N_14882);
nor UO_299 (O_299,N_14998,N_14898);
or UO_300 (O_300,N_14873,N_14958);
or UO_301 (O_301,N_14958,N_14940);
nor UO_302 (O_302,N_14852,N_14928);
xnor UO_303 (O_303,N_14850,N_14953);
nor UO_304 (O_304,N_14934,N_14938);
xor UO_305 (O_305,N_14900,N_14970);
nor UO_306 (O_306,N_14983,N_14972);
and UO_307 (O_307,N_14858,N_14950);
nand UO_308 (O_308,N_14961,N_14903);
or UO_309 (O_309,N_14975,N_14914);
and UO_310 (O_310,N_14893,N_14979);
and UO_311 (O_311,N_14885,N_14905);
nor UO_312 (O_312,N_14992,N_14960);
nand UO_313 (O_313,N_14951,N_14904);
or UO_314 (O_314,N_14920,N_14850);
or UO_315 (O_315,N_14982,N_14963);
nor UO_316 (O_316,N_14986,N_14870);
or UO_317 (O_317,N_14897,N_14921);
xnor UO_318 (O_318,N_14925,N_14870);
nor UO_319 (O_319,N_14998,N_14868);
nand UO_320 (O_320,N_14984,N_14888);
xor UO_321 (O_321,N_14918,N_14948);
or UO_322 (O_322,N_14862,N_14883);
or UO_323 (O_323,N_14854,N_14981);
xnor UO_324 (O_324,N_14930,N_14986);
xnor UO_325 (O_325,N_14969,N_14994);
or UO_326 (O_326,N_14925,N_14942);
xor UO_327 (O_327,N_14978,N_14963);
and UO_328 (O_328,N_14974,N_14852);
or UO_329 (O_329,N_14989,N_14868);
or UO_330 (O_330,N_14966,N_14860);
xnor UO_331 (O_331,N_14945,N_14936);
or UO_332 (O_332,N_14883,N_14909);
or UO_333 (O_333,N_14901,N_14979);
xor UO_334 (O_334,N_14976,N_14995);
nand UO_335 (O_335,N_14936,N_14871);
or UO_336 (O_336,N_14859,N_14867);
and UO_337 (O_337,N_14874,N_14865);
nor UO_338 (O_338,N_14898,N_14993);
nand UO_339 (O_339,N_14878,N_14879);
or UO_340 (O_340,N_14919,N_14902);
nor UO_341 (O_341,N_14905,N_14913);
or UO_342 (O_342,N_14902,N_14952);
nor UO_343 (O_343,N_14999,N_14992);
nor UO_344 (O_344,N_14913,N_14943);
nand UO_345 (O_345,N_14936,N_14970);
or UO_346 (O_346,N_14908,N_14897);
xnor UO_347 (O_347,N_14965,N_14894);
or UO_348 (O_348,N_14988,N_14941);
or UO_349 (O_349,N_14950,N_14977);
nand UO_350 (O_350,N_14902,N_14905);
nor UO_351 (O_351,N_14865,N_14980);
xor UO_352 (O_352,N_14877,N_14982);
or UO_353 (O_353,N_14971,N_14886);
nand UO_354 (O_354,N_14880,N_14926);
nand UO_355 (O_355,N_14932,N_14854);
or UO_356 (O_356,N_14859,N_14988);
and UO_357 (O_357,N_14948,N_14938);
and UO_358 (O_358,N_14976,N_14910);
nor UO_359 (O_359,N_14869,N_14993);
nand UO_360 (O_360,N_14859,N_14946);
xnor UO_361 (O_361,N_14903,N_14917);
or UO_362 (O_362,N_14867,N_14988);
or UO_363 (O_363,N_14852,N_14980);
xnor UO_364 (O_364,N_14859,N_14921);
nand UO_365 (O_365,N_14999,N_14880);
or UO_366 (O_366,N_14999,N_14944);
xnor UO_367 (O_367,N_14908,N_14943);
nor UO_368 (O_368,N_14900,N_14850);
xnor UO_369 (O_369,N_14948,N_14927);
or UO_370 (O_370,N_14870,N_14918);
nor UO_371 (O_371,N_14917,N_14983);
xor UO_372 (O_372,N_14944,N_14886);
or UO_373 (O_373,N_14863,N_14924);
or UO_374 (O_374,N_14929,N_14948);
and UO_375 (O_375,N_14919,N_14852);
or UO_376 (O_376,N_14883,N_14948);
and UO_377 (O_377,N_14929,N_14916);
nand UO_378 (O_378,N_14855,N_14910);
and UO_379 (O_379,N_14949,N_14877);
and UO_380 (O_380,N_14932,N_14945);
xnor UO_381 (O_381,N_14902,N_14851);
nor UO_382 (O_382,N_14981,N_14894);
xnor UO_383 (O_383,N_14874,N_14949);
nor UO_384 (O_384,N_14904,N_14870);
or UO_385 (O_385,N_14938,N_14987);
nand UO_386 (O_386,N_14913,N_14929);
nor UO_387 (O_387,N_14917,N_14972);
nor UO_388 (O_388,N_14980,N_14878);
nor UO_389 (O_389,N_14962,N_14943);
nor UO_390 (O_390,N_14968,N_14850);
or UO_391 (O_391,N_14890,N_14948);
and UO_392 (O_392,N_14862,N_14885);
xor UO_393 (O_393,N_14928,N_14853);
xnor UO_394 (O_394,N_14922,N_14961);
nor UO_395 (O_395,N_14859,N_14967);
nand UO_396 (O_396,N_14861,N_14937);
or UO_397 (O_397,N_14850,N_14950);
xor UO_398 (O_398,N_14880,N_14981);
and UO_399 (O_399,N_14979,N_14891);
nand UO_400 (O_400,N_14920,N_14893);
nor UO_401 (O_401,N_14965,N_14935);
nand UO_402 (O_402,N_14959,N_14882);
nand UO_403 (O_403,N_14983,N_14937);
or UO_404 (O_404,N_14870,N_14951);
nand UO_405 (O_405,N_14873,N_14852);
xor UO_406 (O_406,N_14855,N_14877);
xor UO_407 (O_407,N_14860,N_14929);
nor UO_408 (O_408,N_14959,N_14876);
nor UO_409 (O_409,N_14931,N_14998);
or UO_410 (O_410,N_14976,N_14897);
and UO_411 (O_411,N_14948,N_14971);
or UO_412 (O_412,N_14973,N_14882);
nand UO_413 (O_413,N_14963,N_14983);
or UO_414 (O_414,N_14901,N_14951);
nor UO_415 (O_415,N_14877,N_14853);
nand UO_416 (O_416,N_14896,N_14860);
or UO_417 (O_417,N_14855,N_14852);
or UO_418 (O_418,N_14946,N_14969);
nor UO_419 (O_419,N_14981,N_14972);
xor UO_420 (O_420,N_14940,N_14974);
xnor UO_421 (O_421,N_14892,N_14990);
or UO_422 (O_422,N_14894,N_14978);
nand UO_423 (O_423,N_14938,N_14936);
nor UO_424 (O_424,N_14861,N_14988);
or UO_425 (O_425,N_14883,N_14920);
or UO_426 (O_426,N_14877,N_14890);
and UO_427 (O_427,N_14861,N_14873);
nor UO_428 (O_428,N_14989,N_14969);
and UO_429 (O_429,N_14859,N_14891);
nand UO_430 (O_430,N_14990,N_14986);
or UO_431 (O_431,N_14898,N_14942);
nor UO_432 (O_432,N_14856,N_14905);
and UO_433 (O_433,N_14862,N_14887);
nor UO_434 (O_434,N_14927,N_14891);
nor UO_435 (O_435,N_14877,N_14927);
xor UO_436 (O_436,N_14937,N_14865);
and UO_437 (O_437,N_14998,N_14946);
and UO_438 (O_438,N_14928,N_14981);
or UO_439 (O_439,N_14993,N_14911);
nand UO_440 (O_440,N_14900,N_14995);
or UO_441 (O_441,N_14941,N_14969);
nand UO_442 (O_442,N_14881,N_14878);
and UO_443 (O_443,N_14913,N_14856);
xnor UO_444 (O_444,N_14853,N_14900);
nor UO_445 (O_445,N_14862,N_14983);
and UO_446 (O_446,N_14908,N_14939);
and UO_447 (O_447,N_14926,N_14894);
or UO_448 (O_448,N_14875,N_14851);
nor UO_449 (O_449,N_14863,N_14972);
nand UO_450 (O_450,N_14888,N_14905);
xnor UO_451 (O_451,N_14873,N_14858);
or UO_452 (O_452,N_14923,N_14977);
and UO_453 (O_453,N_14874,N_14902);
and UO_454 (O_454,N_14925,N_14963);
xor UO_455 (O_455,N_14916,N_14938);
nand UO_456 (O_456,N_14998,N_14922);
nand UO_457 (O_457,N_14856,N_14928);
xor UO_458 (O_458,N_14956,N_14916);
nor UO_459 (O_459,N_14891,N_14978);
and UO_460 (O_460,N_14852,N_14977);
xor UO_461 (O_461,N_14915,N_14974);
or UO_462 (O_462,N_14977,N_14924);
or UO_463 (O_463,N_14850,N_14863);
nor UO_464 (O_464,N_14988,N_14934);
nor UO_465 (O_465,N_14910,N_14873);
xor UO_466 (O_466,N_14876,N_14994);
or UO_467 (O_467,N_14922,N_14908);
nand UO_468 (O_468,N_14874,N_14850);
and UO_469 (O_469,N_14957,N_14989);
xor UO_470 (O_470,N_14858,N_14981);
xnor UO_471 (O_471,N_14868,N_14884);
and UO_472 (O_472,N_14876,N_14880);
or UO_473 (O_473,N_14991,N_14972);
xnor UO_474 (O_474,N_14923,N_14906);
or UO_475 (O_475,N_14891,N_14884);
xor UO_476 (O_476,N_14864,N_14888);
nand UO_477 (O_477,N_14893,N_14896);
xnor UO_478 (O_478,N_14879,N_14861);
or UO_479 (O_479,N_14888,N_14986);
or UO_480 (O_480,N_14872,N_14937);
nand UO_481 (O_481,N_14944,N_14913);
or UO_482 (O_482,N_14879,N_14868);
xnor UO_483 (O_483,N_14996,N_14982);
xor UO_484 (O_484,N_14902,N_14976);
and UO_485 (O_485,N_14965,N_14977);
or UO_486 (O_486,N_14877,N_14966);
xor UO_487 (O_487,N_14864,N_14907);
nand UO_488 (O_488,N_14939,N_14943);
xor UO_489 (O_489,N_14852,N_14982);
nand UO_490 (O_490,N_14993,N_14991);
nand UO_491 (O_491,N_14957,N_14970);
xor UO_492 (O_492,N_14890,N_14911);
xor UO_493 (O_493,N_14952,N_14893);
xnor UO_494 (O_494,N_14977,N_14969);
xnor UO_495 (O_495,N_14945,N_14851);
or UO_496 (O_496,N_14909,N_14889);
and UO_497 (O_497,N_14959,N_14923);
nor UO_498 (O_498,N_14945,N_14922);
nand UO_499 (O_499,N_14904,N_14920);
and UO_500 (O_500,N_14893,N_14945);
or UO_501 (O_501,N_14857,N_14995);
nand UO_502 (O_502,N_14946,N_14850);
and UO_503 (O_503,N_14947,N_14906);
and UO_504 (O_504,N_14945,N_14972);
xnor UO_505 (O_505,N_14906,N_14967);
or UO_506 (O_506,N_14894,N_14879);
nand UO_507 (O_507,N_14887,N_14856);
and UO_508 (O_508,N_14998,N_14916);
or UO_509 (O_509,N_14856,N_14922);
and UO_510 (O_510,N_14875,N_14869);
or UO_511 (O_511,N_14960,N_14955);
and UO_512 (O_512,N_14902,N_14894);
nand UO_513 (O_513,N_14987,N_14982);
xor UO_514 (O_514,N_14864,N_14877);
and UO_515 (O_515,N_14881,N_14927);
nor UO_516 (O_516,N_14866,N_14976);
xor UO_517 (O_517,N_14923,N_14980);
and UO_518 (O_518,N_14918,N_14852);
and UO_519 (O_519,N_14869,N_14989);
and UO_520 (O_520,N_14972,N_14925);
and UO_521 (O_521,N_14972,N_14913);
nor UO_522 (O_522,N_14865,N_14851);
or UO_523 (O_523,N_14948,N_14851);
nand UO_524 (O_524,N_14856,N_14921);
or UO_525 (O_525,N_14964,N_14927);
and UO_526 (O_526,N_14965,N_14956);
xnor UO_527 (O_527,N_14870,N_14877);
xnor UO_528 (O_528,N_14992,N_14949);
or UO_529 (O_529,N_14919,N_14879);
nor UO_530 (O_530,N_14886,N_14885);
and UO_531 (O_531,N_14916,N_14876);
xor UO_532 (O_532,N_14975,N_14981);
nor UO_533 (O_533,N_14931,N_14876);
or UO_534 (O_534,N_14890,N_14875);
nand UO_535 (O_535,N_14858,N_14865);
and UO_536 (O_536,N_14876,N_14862);
nor UO_537 (O_537,N_14925,N_14917);
or UO_538 (O_538,N_14988,N_14994);
nand UO_539 (O_539,N_14894,N_14969);
xor UO_540 (O_540,N_14991,N_14859);
nand UO_541 (O_541,N_14994,N_14943);
or UO_542 (O_542,N_14853,N_14901);
and UO_543 (O_543,N_14898,N_14938);
xor UO_544 (O_544,N_14934,N_14893);
and UO_545 (O_545,N_14927,N_14949);
nand UO_546 (O_546,N_14973,N_14959);
xor UO_547 (O_547,N_14938,N_14949);
xnor UO_548 (O_548,N_14908,N_14896);
nand UO_549 (O_549,N_14976,N_14972);
or UO_550 (O_550,N_14968,N_14945);
xnor UO_551 (O_551,N_14960,N_14908);
and UO_552 (O_552,N_14895,N_14946);
or UO_553 (O_553,N_14872,N_14883);
nand UO_554 (O_554,N_14894,N_14974);
nor UO_555 (O_555,N_14979,N_14940);
nor UO_556 (O_556,N_14862,N_14991);
or UO_557 (O_557,N_14858,N_14882);
and UO_558 (O_558,N_14862,N_14965);
or UO_559 (O_559,N_14947,N_14997);
or UO_560 (O_560,N_14950,N_14878);
nor UO_561 (O_561,N_14923,N_14869);
or UO_562 (O_562,N_14861,N_14987);
nor UO_563 (O_563,N_14870,N_14943);
and UO_564 (O_564,N_14957,N_14889);
or UO_565 (O_565,N_14921,N_14854);
nand UO_566 (O_566,N_14861,N_14996);
and UO_567 (O_567,N_14957,N_14897);
and UO_568 (O_568,N_14926,N_14936);
xor UO_569 (O_569,N_14871,N_14969);
or UO_570 (O_570,N_14920,N_14853);
and UO_571 (O_571,N_14865,N_14992);
xor UO_572 (O_572,N_14968,N_14924);
and UO_573 (O_573,N_14886,N_14984);
nand UO_574 (O_574,N_14879,N_14893);
or UO_575 (O_575,N_14871,N_14887);
nand UO_576 (O_576,N_14940,N_14956);
and UO_577 (O_577,N_14883,N_14954);
and UO_578 (O_578,N_14892,N_14895);
xnor UO_579 (O_579,N_14955,N_14973);
nor UO_580 (O_580,N_14856,N_14945);
nor UO_581 (O_581,N_14958,N_14882);
nand UO_582 (O_582,N_14982,N_14979);
xor UO_583 (O_583,N_14976,N_14929);
and UO_584 (O_584,N_14917,N_14882);
or UO_585 (O_585,N_14977,N_14963);
or UO_586 (O_586,N_14917,N_14916);
xnor UO_587 (O_587,N_14965,N_14853);
nor UO_588 (O_588,N_14985,N_14865);
nor UO_589 (O_589,N_14968,N_14928);
nor UO_590 (O_590,N_14967,N_14925);
nand UO_591 (O_591,N_14871,N_14925);
and UO_592 (O_592,N_14877,N_14941);
nor UO_593 (O_593,N_14850,N_14911);
nand UO_594 (O_594,N_14986,N_14924);
nand UO_595 (O_595,N_14885,N_14936);
or UO_596 (O_596,N_14964,N_14926);
xnor UO_597 (O_597,N_14998,N_14856);
xnor UO_598 (O_598,N_14912,N_14960);
xnor UO_599 (O_599,N_14967,N_14953);
nor UO_600 (O_600,N_14980,N_14964);
nor UO_601 (O_601,N_14878,N_14875);
nand UO_602 (O_602,N_14965,N_14950);
and UO_603 (O_603,N_14976,N_14885);
nor UO_604 (O_604,N_14984,N_14887);
or UO_605 (O_605,N_14986,N_14959);
or UO_606 (O_606,N_14981,N_14926);
and UO_607 (O_607,N_14943,N_14991);
nand UO_608 (O_608,N_14996,N_14859);
nand UO_609 (O_609,N_14905,N_14921);
and UO_610 (O_610,N_14880,N_14899);
nor UO_611 (O_611,N_14938,N_14913);
nor UO_612 (O_612,N_14877,N_14993);
or UO_613 (O_613,N_14978,N_14857);
and UO_614 (O_614,N_14992,N_14852);
nand UO_615 (O_615,N_14916,N_14883);
xor UO_616 (O_616,N_14939,N_14867);
and UO_617 (O_617,N_14862,N_14986);
xor UO_618 (O_618,N_14990,N_14913);
or UO_619 (O_619,N_14998,N_14907);
or UO_620 (O_620,N_14864,N_14869);
xor UO_621 (O_621,N_14983,N_14867);
and UO_622 (O_622,N_14879,N_14883);
nor UO_623 (O_623,N_14971,N_14873);
xor UO_624 (O_624,N_14860,N_14886);
xor UO_625 (O_625,N_14918,N_14873);
or UO_626 (O_626,N_14854,N_14850);
or UO_627 (O_627,N_14882,N_14984);
nand UO_628 (O_628,N_14877,N_14945);
nand UO_629 (O_629,N_14860,N_14942);
nand UO_630 (O_630,N_14917,N_14912);
and UO_631 (O_631,N_14956,N_14919);
and UO_632 (O_632,N_14919,N_14896);
nor UO_633 (O_633,N_14904,N_14882);
xnor UO_634 (O_634,N_14876,N_14913);
nor UO_635 (O_635,N_14901,N_14885);
and UO_636 (O_636,N_14876,N_14943);
nor UO_637 (O_637,N_14909,N_14967);
or UO_638 (O_638,N_14922,N_14866);
nor UO_639 (O_639,N_14980,N_14949);
nand UO_640 (O_640,N_14891,N_14904);
or UO_641 (O_641,N_14902,N_14940);
xnor UO_642 (O_642,N_14975,N_14924);
or UO_643 (O_643,N_14885,N_14968);
nand UO_644 (O_644,N_14953,N_14906);
xnor UO_645 (O_645,N_14986,N_14940);
nor UO_646 (O_646,N_14925,N_14872);
or UO_647 (O_647,N_14930,N_14977);
nand UO_648 (O_648,N_14959,N_14921);
nand UO_649 (O_649,N_14870,N_14944);
and UO_650 (O_650,N_14932,N_14925);
xnor UO_651 (O_651,N_14875,N_14963);
or UO_652 (O_652,N_14923,N_14867);
nand UO_653 (O_653,N_14884,N_14919);
nand UO_654 (O_654,N_14857,N_14904);
nand UO_655 (O_655,N_14994,N_14899);
nor UO_656 (O_656,N_14891,N_14909);
xnor UO_657 (O_657,N_14913,N_14893);
nand UO_658 (O_658,N_14928,N_14995);
and UO_659 (O_659,N_14972,N_14965);
nand UO_660 (O_660,N_14885,N_14913);
xor UO_661 (O_661,N_14990,N_14900);
and UO_662 (O_662,N_14870,N_14891);
nand UO_663 (O_663,N_14916,N_14954);
and UO_664 (O_664,N_14851,N_14926);
or UO_665 (O_665,N_14876,N_14924);
xnor UO_666 (O_666,N_14949,N_14942);
or UO_667 (O_667,N_14874,N_14995);
nand UO_668 (O_668,N_14907,N_14914);
xor UO_669 (O_669,N_14852,N_14949);
nor UO_670 (O_670,N_14940,N_14854);
or UO_671 (O_671,N_14892,N_14959);
and UO_672 (O_672,N_14854,N_14888);
xnor UO_673 (O_673,N_14944,N_14930);
nor UO_674 (O_674,N_14933,N_14990);
nand UO_675 (O_675,N_14865,N_14881);
xnor UO_676 (O_676,N_14916,N_14945);
and UO_677 (O_677,N_14933,N_14852);
nor UO_678 (O_678,N_14931,N_14990);
nor UO_679 (O_679,N_14851,N_14983);
nor UO_680 (O_680,N_14922,N_14884);
and UO_681 (O_681,N_14859,N_14931);
or UO_682 (O_682,N_14991,N_14890);
nand UO_683 (O_683,N_14951,N_14987);
and UO_684 (O_684,N_14915,N_14976);
or UO_685 (O_685,N_14917,N_14855);
and UO_686 (O_686,N_14893,N_14883);
and UO_687 (O_687,N_14917,N_14968);
and UO_688 (O_688,N_14974,N_14996);
xnor UO_689 (O_689,N_14937,N_14913);
nor UO_690 (O_690,N_14974,N_14890);
or UO_691 (O_691,N_14887,N_14925);
and UO_692 (O_692,N_14870,N_14855);
nand UO_693 (O_693,N_14907,N_14984);
xor UO_694 (O_694,N_14927,N_14913);
or UO_695 (O_695,N_14978,N_14912);
nand UO_696 (O_696,N_14986,N_14861);
nand UO_697 (O_697,N_14913,N_14908);
nor UO_698 (O_698,N_14866,N_14896);
or UO_699 (O_699,N_14912,N_14856);
or UO_700 (O_700,N_14894,N_14927);
nor UO_701 (O_701,N_14998,N_14979);
nor UO_702 (O_702,N_14935,N_14971);
nand UO_703 (O_703,N_14933,N_14868);
nand UO_704 (O_704,N_14964,N_14885);
and UO_705 (O_705,N_14932,N_14974);
and UO_706 (O_706,N_14971,N_14891);
and UO_707 (O_707,N_14988,N_14889);
xor UO_708 (O_708,N_14880,N_14979);
and UO_709 (O_709,N_14863,N_14919);
nand UO_710 (O_710,N_14927,N_14899);
and UO_711 (O_711,N_14974,N_14964);
nor UO_712 (O_712,N_14939,N_14912);
nor UO_713 (O_713,N_14860,N_14944);
or UO_714 (O_714,N_14962,N_14879);
nor UO_715 (O_715,N_14949,N_14996);
xor UO_716 (O_716,N_14887,N_14889);
or UO_717 (O_717,N_14857,N_14927);
or UO_718 (O_718,N_14994,N_14946);
nor UO_719 (O_719,N_14876,N_14935);
nand UO_720 (O_720,N_14910,N_14970);
or UO_721 (O_721,N_14966,N_14925);
nand UO_722 (O_722,N_14923,N_14963);
and UO_723 (O_723,N_14970,N_14872);
and UO_724 (O_724,N_14860,N_14979);
nor UO_725 (O_725,N_14962,N_14979);
or UO_726 (O_726,N_14988,N_14890);
and UO_727 (O_727,N_14857,N_14872);
nor UO_728 (O_728,N_14960,N_14957);
nand UO_729 (O_729,N_14943,N_14940);
nor UO_730 (O_730,N_14866,N_14964);
nor UO_731 (O_731,N_14954,N_14922);
nand UO_732 (O_732,N_14978,N_14927);
xor UO_733 (O_733,N_14957,N_14937);
nand UO_734 (O_734,N_14926,N_14861);
or UO_735 (O_735,N_14977,N_14902);
xnor UO_736 (O_736,N_14893,N_14877);
or UO_737 (O_737,N_14866,N_14917);
xor UO_738 (O_738,N_14877,N_14947);
nand UO_739 (O_739,N_14881,N_14891);
xor UO_740 (O_740,N_14859,N_14980);
nand UO_741 (O_741,N_14942,N_14867);
or UO_742 (O_742,N_14969,N_14897);
nand UO_743 (O_743,N_14881,N_14974);
xnor UO_744 (O_744,N_14970,N_14923);
nor UO_745 (O_745,N_14882,N_14878);
nand UO_746 (O_746,N_14974,N_14995);
nand UO_747 (O_747,N_14938,N_14888);
xor UO_748 (O_748,N_14939,N_14946);
nor UO_749 (O_749,N_14989,N_14931);
or UO_750 (O_750,N_14967,N_14924);
nand UO_751 (O_751,N_14876,N_14892);
nor UO_752 (O_752,N_14991,N_14997);
xor UO_753 (O_753,N_14956,N_14975);
xnor UO_754 (O_754,N_14980,N_14966);
or UO_755 (O_755,N_14918,N_14890);
xor UO_756 (O_756,N_14970,N_14898);
nor UO_757 (O_757,N_14895,N_14949);
nand UO_758 (O_758,N_14913,N_14872);
xnor UO_759 (O_759,N_14903,N_14870);
xnor UO_760 (O_760,N_14955,N_14944);
nor UO_761 (O_761,N_14980,N_14957);
nand UO_762 (O_762,N_14907,N_14905);
or UO_763 (O_763,N_14915,N_14932);
or UO_764 (O_764,N_14863,N_14940);
nand UO_765 (O_765,N_14963,N_14887);
and UO_766 (O_766,N_14900,N_14888);
nor UO_767 (O_767,N_14907,N_14923);
and UO_768 (O_768,N_14898,N_14929);
and UO_769 (O_769,N_14882,N_14851);
nor UO_770 (O_770,N_14992,N_14898);
or UO_771 (O_771,N_14917,N_14900);
and UO_772 (O_772,N_14868,N_14946);
xor UO_773 (O_773,N_14984,N_14941);
nor UO_774 (O_774,N_14936,N_14992);
nand UO_775 (O_775,N_14980,N_14967);
or UO_776 (O_776,N_14952,N_14926);
nand UO_777 (O_777,N_14915,N_14874);
or UO_778 (O_778,N_14865,N_14958);
or UO_779 (O_779,N_14915,N_14945);
or UO_780 (O_780,N_14891,N_14899);
and UO_781 (O_781,N_14901,N_14941);
nand UO_782 (O_782,N_14874,N_14873);
or UO_783 (O_783,N_14915,N_14972);
xnor UO_784 (O_784,N_14900,N_14931);
or UO_785 (O_785,N_14935,N_14926);
nand UO_786 (O_786,N_14867,N_14960);
xnor UO_787 (O_787,N_14940,N_14949);
or UO_788 (O_788,N_14930,N_14861);
and UO_789 (O_789,N_14880,N_14912);
nand UO_790 (O_790,N_14915,N_14927);
nand UO_791 (O_791,N_14932,N_14967);
nand UO_792 (O_792,N_14939,N_14910);
xor UO_793 (O_793,N_14934,N_14974);
nand UO_794 (O_794,N_14944,N_14967);
nor UO_795 (O_795,N_14940,N_14985);
nand UO_796 (O_796,N_14894,N_14914);
and UO_797 (O_797,N_14897,N_14900);
or UO_798 (O_798,N_14888,N_14855);
nor UO_799 (O_799,N_14972,N_14869);
xnor UO_800 (O_800,N_14984,N_14990);
nor UO_801 (O_801,N_14886,N_14999);
or UO_802 (O_802,N_14867,N_14951);
nor UO_803 (O_803,N_14972,N_14935);
and UO_804 (O_804,N_14913,N_14853);
and UO_805 (O_805,N_14965,N_14933);
xor UO_806 (O_806,N_14889,N_14867);
nand UO_807 (O_807,N_14866,N_14853);
xnor UO_808 (O_808,N_14879,N_14983);
xnor UO_809 (O_809,N_14925,N_14969);
or UO_810 (O_810,N_14974,N_14989);
nand UO_811 (O_811,N_14912,N_14946);
xnor UO_812 (O_812,N_14896,N_14875);
and UO_813 (O_813,N_14944,N_14977);
nor UO_814 (O_814,N_14985,N_14908);
and UO_815 (O_815,N_14883,N_14930);
and UO_816 (O_816,N_14967,N_14911);
nand UO_817 (O_817,N_14876,N_14982);
and UO_818 (O_818,N_14891,N_14882);
or UO_819 (O_819,N_14898,N_14999);
or UO_820 (O_820,N_14945,N_14933);
nand UO_821 (O_821,N_14913,N_14992);
or UO_822 (O_822,N_14850,N_14996);
or UO_823 (O_823,N_14891,N_14902);
xnor UO_824 (O_824,N_14903,N_14861);
or UO_825 (O_825,N_14879,N_14892);
nor UO_826 (O_826,N_14851,N_14925);
and UO_827 (O_827,N_14873,N_14947);
or UO_828 (O_828,N_14934,N_14979);
nor UO_829 (O_829,N_14926,N_14984);
nor UO_830 (O_830,N_14888,N_14939);
and UO_831 (O_831,N_14954,N_14862);
nor UO_832 (O_832,N_14887,N_14868);
nor UO_833 (O_833,N_14970,N_14984);
nor UO_834 (O_834,N_14929,N_14952);
or UO_835 (O_835,N_14918,N_14959);
or UO_836 (O_836,N_14962,N_14976);
nand UO_837 (O_837,N_14894,N_14916);
xnor UO_838 (O_838,N_14873,N_14977);
nand UO_839 (O_839,N_14966,N_14961);
xnor UO_840 (O_840,N_14910,N_14963);
and UO_841 (O_841,N_14948,N_14916);
nor UO_842 (O_842,N_14897,N_14860);
nor UO_843 (O_843,N_14948,N_14877);
nor UO_844 (O_844,N_14909,N_14959);
or UO_845 (O_845,N_14865,N_14951);
or UO_846 (O_846,N_14869,N_14893);
or UO_847 (O_847,N_14929,N_14994);
nand UO_848 (O_848,N_14957,N_14953);
nor UO_849 (O_849,N_14999,N_14984);
xor UO_850 (O_850,N_14924,N_14926);
and UO_851 (O_851,N_14881,N_14871);
or UO_852 (O_852,N_14868,N_14912);
nand UO_853 (O_853,N_14944,N_14880);
or UO_854 (O_854,N_14923,N_14948);
or UO_855 (O_855,N_14938,N_14893);
nand UO_856 (O_856,N_14960,N_14914);
or UO_857 (O_857,N_14970,N_14873);
nor UO_858 (O_858,N_14947,N_14981);
xor UO_859 (O_859,N_14895,N_14971);
and UO_860 (O_860,N_14881,N_14931);
nor UO_861 (O_861,N_14975,N_14884);
xnor UO_862 (O_862,N_14936,N_14862);
nand UO_863 (O_863,N_14968,N_14869);
xnor UO_864 (O_864,N_14989,N_14871);
nor UO_865 (O_865,N_14990,N_14867);
or UO_866 (O_866,N_14986,N_14864);
and UO_867 (O_867,N_14994,N_14875);
nor UO_868 (O_868,N_14895,N_14958);
nand UO_869 (O_869,N_14939,N_14982);
nor UO_870 (O_870,N_14855,N_14983);
xor UO_871 (O_871,N_14984,N_14910);
xnor UO_872 (O_872,N_14853,N_14991);
nor UO_873 (O_873,N_14860,N_14967);
or UO_874 (O_874,N_14893,N_14853);
nand UO_875 (O_875,N_14904,N_14912);
and UO_876 (O_876,N_14935,N_14869);
nor UO_877 (O_877,N_14938,N_14982);
xnor UO_878 (O_878,N_14991,N_14896);
nor UO_879 (O_879,N_14957,N_14985);
and UO_880 (O_880,N_14962,N_14892);
xnor UO_881 (O_881,N_14877,N_14954);
nor UO_882 (O_882,N_14905,N_14949);
nor UO_883 (O_883,N_14877,N_14943);
or UO_884 (O_884,N_14963,N_14942);
nor UO_885 (O_885,N_14927,N_14888);
xnor UO_886 (O_886,N_14853,N_14995);
and UO_887 (O_887,N_14871,N_14935);
nor UO_888 (O_888,N_14931,N_14895);
nor UO_889 (O_889,N_14858,N_14927);
and UO_890 (O_890,N_14885,N_14927);
nor UO_891 (O_891,N_14873,N_14909);
xor UO_892 (O_892,N_14858,N_14900);
and UO_893 (O_893,N_14904,N_14886);
and UO_894 (O_894,N_14911,N_14859);
nor UO_895 (O_895,N_14902,N_14990);
nand UO_896 (O_896,N_14874,N_14866);
nand UO_897 (O_897,N_14885,N_14895);
xnor UO_898 (O_898,N_14897,N_14924);
xor UO_899 (O_899,N_14927,N_14974);
and UO_900 (O_900,N_14912,N_14998);
nand UO_901 (O_901,N_14948,N_14885);
and UO_902 (O_902,N_14978,N_14976);
nor UO_903 (O_903,N_14880,N_14932);
or UO_904 (O_904,N_14879,N_14863);
nor UO_905 (O_905,N_14936,N_14933);
and UO_906 (O_906,N_14919,N_14992);
or UO_907 (O_907,N_14917,N_14994);
or UO_908 (O_908,N_14993,N_14944);
and UO_909 (O_909,N_14959,N_14874);
or UO_910 (O_910,N_14960,N_14926);
nand UO_911 (O_911,N_14989,N_14880);
xnor UO_912 (O_912,N_14851,N_14856);
nor UO_913 (O_913,N_14966,N_14992);
or UO_914 (O_914,N_14982,N_14978);
or UO_915 (O_915,N_14979,N_14920);
nor UO_916 (O_916,N_14860,N_14988);
or UO_917 (O_917,N_14993,N_14954);
or UO_918 (O_918,N_14866,N_14883);
nand UO_919 (O_919,N_14863,N_14973);
nand UO_920 (O_920,N_14943,N_14916);
nand UO_921 (O_921,N_14962,N_14950);
or UO_922 (O_922,N_14928,N_14999);
and UO_923 (O_923,N_14894,N_14857);
or UO_924 (O_924,N_14939,N_14992);
nand UO_925 (O_925,N_14980,N_14929);
and UO_926 (O_926,N_14911,N_14919);
and UO_927 (O_927,N_14880,N_14931);
xor UO_928 (O_928,N_14897,N_14889);
and UO_929 (O_929,N_14973,N_14856);
or UO_930 (O_930,N_14942,N_14877);
nor UO_931 (O_931,N_14873,N_14953);
xor UO_932 (O_932,N_14918,N_14958);
xor UO_933 (O_933,N_14871,N_14884);
xor UO_934 (O_934,N_14966,N_14864);
nand UO_935 (O_935,N_14877,N_14987);
nand UO_936 (O_936,N_14911,N_14917);
nor UO_937 (O_937,N_14945,N_14931);
and UO_938 (O_938,N_14948,N_14987);
and UO_939 (O_939,N_14958,N_14924);
and UO_940 (O_940,N_14922,N_14896);
xor UO_941 (O_941,N_14990,N_14856);
nand UO_942 (O_942,N_14882,N_14978);
or UO_943 (O_943,N_14979,N_14875);
and UO_944 (O_944,N_14934,N_14884);
xor UO_945 (O_945,N_14909,N_14907);
xnor UO_946 (O_946,N_14984,N_14899);
or UO_947 (O_947,N_14912,N_14891);
or UO_948 (O_948,N_14852,N_14969);
or UO_949 (O_949,N_14970,N_14884);
nand UO_950 (O_950,N_14975,N_14971);
xnor UO_951 (O_951,N_14939,N_14945);
or UO_952 (O_952,N_14878,N_14961);
and UO_953 (O_953,N_14984,N_14931);
nor UO_954 (O_954,N_14965,N_14860);
and UO_955 (O_955,N_14917,N_14884);
nor UO_956 (O_956,N_14998,N_14925);
or UO_957 (O_957,N_14880,N_14930);
nor UO_958 (O_958,N_14871,N_14877);
and UO_959 (O_959,N_14972,N_14992);
and UO_960 (O_960,N_14862,N_14851);
and UO_961 (O_961,N_14850,N_14867);
nand UO_962 (O_962,N_14901,N_14851);
nand UO_963 (O_963,N_14869,N_14936);
nor UO_964 (O_964,N_14854,N_14936);
nand UO_965 (O_965,N_14910,N_14864);
xnor UO_966 (O_966,N_14887,N_14991);
nand UO_967 (O_967,N_14987,N_14996);
nor UO_968 (O_968,N_14924,N_14997);
nand UO_969 (O_969,N_14993,N_14892);
or UO_970 (O_970,N_14924,N_14879);
xnor UO_971 (O_971,N_14997,N_14960);
nor UO_972 (O_972,N_14982,N_14961);
nor UO_973 (O_973,N_14936,N_14942);
nor UO_974 (O_974,N_14878,N_14931);
nand UO_975 (O_975,N_14939,N_14919);
or UO_976 (O_976,N_14874,N_14896);
nand UO_977 (O_977,N_14894,N_14977);
nor UO_978 (O_978,N_14912,N_14896);
or UO_979 (O_979,N_14920,N_14998);
nor UO_980 (O_980,N_14901,N_14978);
nand UO_981 (O_981,N_14963,N_14852);
nor UO_982 (O_982,N_14887,N_14867);
and UO_983 (O_983,N_14964,N_14861);
nor UO_984 (O_984,N_14931,N_14905);
xor UO_985 (O_985,N_14890,N_14987);
nor UO_986 (O_986,N_14943,N_14879);
xnor UO_987 (O_987,N_14868,N_14928);
and UO_988 (O_988,N_14931,N_14951);
nor UO_989 (O_989,N_14900,N_14955);
nand UO_990 (O_990,N_14956,N_14890);
nor UO_991 (O_991,N_14899,N_14869);
and UO_992 (O_992,N_14876,N_14927);
and UO_993 (O_993,N_14939,N_14973);
and UO_994 (O_994,N_14937,N_14870);
nand UO_995 (O_995,N_14886,N_14859);
nand UO_996 (O_996,N_14938,N_14937);
nor UO_997 (O_997,N_14991,N_14891);
or UO_998 (O_998,N_14977,N_14911);
nor UO_999 (O_999,N_14987,N_14855);
xnor UO_1000 (O_1000,N_14940,N_14862);
xor UO_1001 (O_1001,N_14998,N_14959);
nor UO_1002 (O_1002,N_14902,N_14870);
or UO_1003 (O_1003,N_14854,N_14875);
xnor UO_1004 (O_1004,N_14942,N_14983);
and UO_1005 (O_1005,N_14852,N_14871);
or UO_1006 (O_1006,N_14984,N_14876);
nor UO_1007 (O_1007,N_14973,N_14972);
and UO_1008 (O_1008,N_14952,N_14946);
nor UO_1009 (O_1009,N_14850,N_14954);
and UO_1010 (O_1010,N_14931,N_14983);
nor UO_1011 (O_1011,N_14915,N_14872);
nand UO_1012 (O_1012,N_14951,N_14972);
xnor UO_1013 (O_1013,N_14988,N_14917);
xnor UO_1014 (O_1014,N_14973,N_14888);
and UO_1015 (O_1015,N_14862,N_14879);
xor UO_1016 (O_1016,N_14887,N_14928);
and UO_1017 (O_1017,N_14905,N_14992);
or UO_1018 (O_1018,N_14899,N_14989);
and UO_1019 (O_1019,N_14902,N_14922);
nor UO_1020 (O_1020,N_14876,N_14934);
nor UO_1021 (O_1021,N_14920,N_14925);
and UO_1022 (O_1022,N_14913,N_14987);
xnor UO_1023 (O_1023,N_14850,N_14883);
nand UO_1024 (O_1024,N_14946,N_14922);
xor UO_1025 (O_1025,N_14865,N_14947);
and UO_1026 (O_1026,N_14955,N_14910);
and UO_1027 (O_1027,N_14943,N_14966);
and UO_1028 (O_1028,N_14883,N_14899);
nor UO_1029 (O_1029,N_14954,N_14892);
or UO_1030 (O_1030,N_14918,N_14944);
and UO_1031 (O_1031,N_14978,N_14884);
or UO_1032 (O_1032,N_14983,N_14986);
nand UO_1033 (O_1033,N_14888,N_14883);
nand UO_1034 (O_1034,N_14999,N_14991);
xnor UO_1035 (O_1035,N_14898,N_14904);
and UO_1036 (O_1036,N_14874,N_14857);
nor UO_1037 (O_1037,N_14914,N_14999);
or UO_1038 (O_1038,N_14872,N_14852);
nor UO_1039 (O_1039,N_14883,N_14877);
xor UO_1040 (O_1040,N_14866,N_14860);
nor UO_1041 (O_1041,N_14946,N_14999);
or UO_1042 (O_1042,N_14890,N_14869);
xnor UO_1043 (O_1043,N_14876,N_14978);
nor UO_1044 (O_1044,N_14938,N_14901);
xor UO_1045 (O_1045,N_14930,N_14981);
nor UO_1046 (O_1046,N_14908,N_14918);
xnor UO_1047 (O_1047,N_14954,N_14853);
or UO_1048 (O_1048,N_14852,N_14902);
nor UO_1049 (O_1049,N_14855,N_14994);
and UO_1050 (O_1050,N_14926,N_14944);
and UO_1051 (O_1051,N_14960,N_14900);
xor UO_1052 (O_1052,N_14998,N_14949);
nor UO_1053 (O_1053,N_14922,N_14951);
nand UO_1054 (O_1054,N_14852,N_14897);
xnor UO_1055 (O_1055,N_14874,N_14892);
and UO_1056 (O_1056,N_14932,N_14944);
and UO_1057 (O_1057,N_14986,N_14961);
xnor UO_1058 (O_1058,N_14928,N_14915);
xnor UO_1059 (O_1059,N_14946,N_14984);
and UO_1060 (O_1060,N_14884,N_14886);
xnor UO_1061 (O_1061,N_14952,N_14890);
nand UO_1062 (O_1062,N_14865,N_14915);
or UO_1063 (O_1063,N_14889,N_14959);
xnor UO_1064 (O_1064,N_14948,N_14910);
or UO_1065 (O_1065,N_14942,N_14953);
or UO_1066 (O_1066,N_14857,N_14966);
nor UO_1067 (O_1067,N_14976,N_14994);
nor UO_1068 (O_1068,N_14934,N_14930);
and UO_1069 (O_1069,N_14996,N_14990);
nand UO_1070 (O_1070,N_14909,N_14853);
or UO_1071 (O_1071,N_14947,N_14929);
or UO_1072 (O_1072,N_14952,N_14986);
or UO_1073 (O_1073,N_14925,N_14885);
nand UO_1074 (O_1074,N_14952,N_14988);
xor UO_1075 (O_1075,N_14980,N_14885);
nor UO_1076 (O_1076,N_14975,N_14943);
nand UO_1077 (O_1077,N_14893,N_14857);
xnor UO_1078 (O_1078,N_14930,N_14952);
nand UO_1079 (O_1079,N_14932,N_14963);
or UO_1080 (O_1080,N_14874,N_14955);
and UO_1081 (O_1081,N_14896,N_14990);
nor UO_1082 (O_1082,N_14898,N_14971);
nor UO_1083 (O_1083,N_14882,N_14875);
and UO_1084 (O_1084,N_14862,N_14996);
or UO_1085 (O_1085,N_14981,N_14866);
xor UO_1086 (O_1086,N_14975,N_14999);
nand UO_1087 (O_1087,N_14859,N_14870);
and UO_1088 (O_1088,N_14854,N_14982);
xnor UO_1089 (O_1089,N_14939,N_14978);
nor UO_1090 (O_1090,N_14938,N_14905);
nand UO_1091 (O_1091,N_14850,N_14969);
nand UO_1092 (O_1092,N_14983,N_14954);
and UO_1093 (O_1093,N_14903,N_14908);
nand UO_1094 (O_1094,N_14991,N_14986);
or UO_1095 (O_1095,N_14956,N_14988);
and UO_1096 (O_1096,N_14975,N_14996);
xnor UO_1097 (O_1097,N_14917,N_14919);
nand UO_1098 (O_1098,N_14956,N_14955);
or UO_1099 (O_1099,N_14887,N_14852);
xnor UO_1100 (O_1100,N_14970,N_14899);
nor UO_1101 (O_1101,N_14878,N_14949);
xnor UO_1102 (O_1102,N_14894,N_14962);
or UO_1103 (O_1103,N_14867,N_14977);
nand UO_1104 (O_1104,N_14916,N_14873);
nor UO_1105 (O_1105,N_14934,N_14926);
or UO_1106 (O_1106,N_14975,N_14968);
xor UO_1107 (O_1107,N_14860,N_14876);
nand UO_1108 (O_1108,N_14920,N_14940);
or UO_1109 (O_1109,N_14912,N_14945);
or UO_1110 (O_1110,N_14941,N_14943);
nor UO_1111 (O_1111,N_14924,N_14951);
xor UO_1112 (O_1112,N_14933,N_14960);
nor UO_1113 (O_1113,N_14856,N_14974);
nand UO_1114 (O_1114,N_14956,N_14891);
nor UO_1115 (O_1115,N_14931,N_14977);
and UO_1116 (O_1116,N_14853,N_14939);
and UO_1117 (O_1117,N_14942,N_14993);
xor UO_1118 (O_1118,N_14850,N_14864);
or UO_1119 (O_1119,N_14894,N_14970);
nor UO_1120 (O_1120,N_14870,N_14938);
nor UO_1121 (O_1121,N_14917,N_14987);
nor UO_1122 (O_1122,N_14958,N_14914);
nor UO_1123 (O_1123,N_14965,N_14916);
and UO_1124 (O_1124,N_14945,N_14885);
and UO_1125 (O_1125,N_14887,N_14886);
or UO_1126 (O_1126,N_14909,N_14854);
xnor UO_1127 (O_1127,N_14857,N_14990);
nor UO_1128 (O_1128,N_14961,N_14862);
xnor UO_1129 (O_1129,N_14899,N_14914);
nand UO_1130 (O_1130,N_14882,N_14989);
xor UO_1131 (O_1131,N_14926,N_14863);
nor UO_1132 (O_1132,N_14853,N_14937);
nand UO_1133 (O_1133,N_14951,N_14902);
nand UO_1134 (O_1134,N_14858,N_14972);
and UO_1135 (O_1135,N_14860,N_14936);
nor UO_1136 (O_1136,N_14882,N_14934);
or UO_1137 (O_1137,N_14854,N_14934);
nand UO_1138 (O_1138,N_14926,N_14975);
and UO_1139 (O_1139,N_14904,N_14965);
xnor UO_1140 (O_1140,N_14977,N_14957);
nand UO_1141 (O_1141,N_14993,N_14887);
and UO_1142 (O_1142,N_14971,N_14899);
xnor UO_1143 (O_1143,N_14953,N_14887);
and UO_1144 (O_1144,N_14945,N_14998);
or UO_1145 (O_1145,N_14909,N_14901);
nand UO_1146 (O_1146,N_14881,N_14982);
or UO_1147 (O_1147,N_14973,N_14866);
nor UO_1148 (O_1148,N_14999,N_14897);
xnor UO_1149 (O_1149,N_14887,N_14891);
xor UO_1150 (O_1150,N_14899,N_14876);
and UO_1151 (O_1151,N_14904,N_14856);
nor UO_1152 (O_1152,N_14936,N_14861);
nor UO_1153 (O_1153,N_14978,N_14897);
and UO_1154 (O_1154,N_14937,N_14945);
nand UO_1155 (O_1155,N_14977,N_14990);
nand UO_1156 (O_1156,N_14852,N_14940);
and UO_1157 (O_1157,N_14909,N_14990);
xor UO_1158 (O_1158,N_14864,N_14932);
xor UO_1159 (O_1159,N_14979,N_14924);
nor UO_1160 (O_1160,N_14898,N_14997);
nand UO_1161 (O_1161,N_14919,N_14862);
nor UO_1162 (O_1162,N_14902,N_14972);
or UO_1163 (O_1163,N_14965,N_14984);
nor UO_1164 (O_1164,N_14988,N_14999);
nor UO_1165 (O_1165,N_14882,N_14896);
nor UO_1166 (O_1166,N_14893,N_14860);
nor UO_1167 (O_1167,N_14937,N_14876);
nor UO_1168 (O_1168,N_14974,N_14859);
nor UO_1169 (O_1169,N_14939,N_14865);
nand UO_1170 (O_1170,N_14914,N_14920);
and UO_1171 (O_1171,N_14928,N_14860);
and UO_1172 (O_1172,N_14855,N_14963);
nand UO_1173 (O_1173,N_14884,N_14967);
nor UO_1174 (O_1174,N_14886,N_14939);
xor UO_1175 (O_1175,N_14921,N_14974);
nand UO_1176 (O_1176,N_14946,N_14919);
nor UO_1177 (O_1177,N_14875,N_14944);
and UO_1178 (O_1178,N_14955,N_14949);
or UO_1179 (O_1179,N_14992,N_14902);
xor UO_1180 (O_1180,N_14924,N_14933);
xor UO_1181 (O_1181,N_14936,N_14961);
and UO_1182 (O_1182,N_14916,N_14984);
nand UO_1183 (O_1183,N_14893,N_14866);
nor UO_1184 (O_1184,N_14921,N_14917);
and UO_1185 (O_1185,N_14917,N_14975);
xor UO_1186 (O_1186,N_14992,N_14892);
xnor UO_1187 (O_1187,N_14897,N_14944);
xnor UO_1188 (O_1188,N_14900,N_14943);
or UO_1189 (O_1189,N_14921,N_14939);
nor UO_1190 (O_1190,N_14876,N_14919);
nor UO_1191 (O_1191,N_14951,N_14862);
or UO_1192 (O_1192,N_14864,N_14897);
and UO_1193 (O_1193,N_14886,N_14928);
nor UO_1194 (O_1194,N_14895,N_14918);
xnor UO_1195 (O_1195,N_14998,N_14966);
nand UO_1196 (O_1196,N_14882,N_14964);
or UO_1197 (O_1197,N_14901,N_14879);
nor UO_1198 (O_1198,N_14936,N_14934);
or UO_1199 (O_1199,N_14907,N_14965);
and UO_1200 (O_1200,N_14870,N_14876);
or UO_1201 (O_1201,N_14859,N_14959);
and UO_1202 (O_1202,N_14944,N_14857);
nor UO_1203 (O_1203,N_14963,N_14975);
and UO_1204 (O_1204,N_14997,N_14990);
nor UO_1205 (O_1205,N_14969,N_14943);
xor UO_1206 (O_1206,N_14989,N_14903);
nand UO_1207 (O_1207,N_14983,N_14924);
and UO_1208 (O_1208,N_14987,N_14966);
xor UO_1209 (O_1209,N_14974,N_14953);
nand UO_1210 (O_1210,N_14909,N_14916);
and UO_1211 (O_1211,N_14894,N_14985);
or UO_1212 (O_1212,N_14885,N_14914);
nor UO_1213 (O_1213,N_14981,N_14870);
and UO_1214 (O_1214,N_14948,N_14991);
xor UO_1215 (O_1215,N_14882,N_14926);
nor UO_1216 (O_1216,N_14928,N_14989);
nand UO_1217 (O_1217,N_14897,N_14968);
nor UO_1218 (O_1218,N_14855,N_14933);
xnor UO_1219 (O_1219,N_14941,N_14918);
or UO_1220 (O_1220,N_14947,N_14879);
xnor UO_1221 (O_1221,N_14894,N_14854);
nand UO_1222 (O_1222,N_14902,N_14950);
or UO_1223 (O_1223,N_14911,N_14995);
nor UO_1224 (O_1224,N_14998,N_14951);
nor UO_1225 (O_1225,N_14929,N_14932);
xor UO_1226 (O_1226,N_14946,N_14900);
nand UO_1227 (O_1227,N_14975,N_14942);
nor UO_1228 (O_1228,N_14892,N_14863);
nand UO_1229 (O_1229,N_14949,N_14973);
xnor UO_1230 (O_1230,N_14971,N_14968);
or UO_1231 (O_1231,N_14850,N_14902);
and UO_1232 (O_1232,N_14923,N_14878);
xnor UO_1233 (O_1233,N_14935,N_14946);
or UO_1234 (O_1234,N_14938,N_14975);
and UO_1235 (O_1235,N_14858,N_14978);
or UO_1236 (O_1236,N_14998,N_14899);
or UO_1237 (O_1237,N_14925,N_14899);
and UO_1238 (O_1238,N_14972,N_14920);
nand UO_1239 (O_1239,N_14867,N_14949);
nand UO_1240 (O_1240,N_14914,N_14921);
nand UO_1241 (O_1241,N_14889,N_14990);
and UO_1242 (O_1242,N_14864,N_14871);
nand UO_1243 (O_1243,N_14920,N_14953);
nor UO_1244 (O_1244,N_14906,N_14970);
and UO_1245 (O_1245,N_14948,N_14957);
xor UO_1246 (O_1246,N_14900,N_14892);
and UO_1247 (O_1247,N_14934,N_14869);
and UO_1248 (O_1248,N_14932,N_14998);
nor UO_1249 (O_1249,N_14884,N_14953);
xnor UO_1250 (O_1250,N_14970,N_14981);
nor UO_1251 (O_1251,N_14945,N_14872);
nand UO_1252 (O_1252,N_14921,N_14964);
xor UO_1253 (O_1253,N_14906,N_14937);
or UO_1254 (O_1254,N_14947,N_14860);
nor UO_1255 (O_1255,N_14894,N_14941);
xor UO_1256 (O_1256,N_14918,N_14942);
or UO_1257 (O_1257,N_14950,N_14857);
xor UO_1258 (O_1258,N_14974,N_14948);
nor UO_1259 (O_1259,N_14929,N_14866);
xor UO_1260 (O_1260,N_14972,N_14851);
or UO_1261 (O_1261,N_14923,N_14950);
xnor UO_1262 (O_1262,N_14932,N_14930);
xor UO_1263 (O_1263,N_14953,N_14943);
or UO_1264 (O_1264,N_14954,N_14852);
or UO_1265 (O_1265,N_14929,N_14853);
and UO_1266 (O_1266,N_14899,N_14957);
nor UO_1267 (O_1267,N_14978,N_14896);
or UO_1268 (O_1268,N_14953,N_14903);
nand UO_1269 (O_1269,N_14902,N_14864);
or UO_1270 (O_1270,N_14942,N_14858);
nor UO_1271 (O_1271,N_14879,N_14914);
nand UO_1272 (O_1272,N_14878,N_14906);
or UO_1273 (O_1273,N_14961,N_14968);
or UO_1274 (O_1274,N_14998,N_14918);
or UO_1275 (O_1275,N_14852,N_14853);
and UO_1276 (O_1276,N_14905,N_14855);
and UO_1277 (O_1277,N_14938,N_14999);
and UO_1278 (O_1278,N_14923,N_14865);
or UO_1279 (O_1279,N_14868,N_14973);
and UO_1280 (O_1280,N_14992,N_14890);
nand UO_1281 (O_1281,N_14885,N_14918);
nand UO_1282 (O_1282,N_14966,N_14957);
and UO_1283 (O_1283,N_14891,N_14975);
nor UO_1284 (O_1284,N_14958,N_14855);
xor UO_1285 (O_1285,N_14957,N_14923);
and UO_1286 (O_1286,N_14889,N_14947);
and UO_1287 (O_1287,N_14986,N_14941);
or UO_1288 (O_1288,N_14956,N_14924);
xnor UO_1289 (O_1289,N_14969,N_14904);
and UO_1290 (O_1290,N_14983,N_14909);
nor UO_1291 (O_1291,N_14859,N_14885);
xnor UO_1292 (O_1292,N_14930,N_14898);
nor UO_1293 (O_1293,N_14990,N_14883);
nand UO_1294 (O_1294,N_14889,N_14864);
nor UO_1295 (O_1295,N_14851,N_14884);
nand UO_1296 (O_1296,N_14885,N_14981);
nor UO_1297 (O_1297,N_14865,N_14957);
and UO_1298 (O_1298,N_14997,N_14977);
xnor UO_1299 (O_1299,N_14968,N_14914);
and UO_1300 (O_1300,N_14872,N_14958);
and UO_1301 (O_1301,N_14940,N_14912);
nor UO_1302 (O_1302,N_14923,N_14927);
or UO_1303 (O_1303,N_14990,N_14884);
or UO_1304 (O_1304,N_14919,N_14882);
xnor UO_1305 (O_1305,N_14858,N_14878);
xnor UO_1306 (O_1306,N_14971,N_14970);
nand UO_1307 (O_1307,N_14852,N_14957);
nand UO_1308 (O_1308,N_14897,N_14861);
nor UO_1309 (O_1309,N_14989,N_14923);
xnor UO_1310 (O_1310,N_14917,N_14970);
nor UO_1311 (O_1311,N_14872,N_14999);
and UO_1312 (O_1312,N_14913,N_14955);
nand UO_1313 (O_1313,N_14877,N_14981);
or UO_1314 (O_1314,N_14954,N_14973);
nor UO_1315 (O_1315,N_14942,N_14991);
and UO_1316 (O_1316,N_14998,N_14957);
xor UO_1317 (O_1317,N_14942,N_14875);
xor UO_1318 (O_1318,N_14998,N_14972);
nor UO_1319 (O_1319,N_14990,N_14945);
or UO_1320 (O_1320,N_14943,N_14979);
and UO_1321 (O_1321,N_14850,N_14931);
or UO_1322 (O_1322,N_14906,N_14852);
xor UO_1323 (O_1323,N_14862,N_14974);
and UO_1324 (O_1324,N_14950,N_14932);
xor UO_1325 (O_1325,N_14979,N_14897);
nor UO_1326 (O_1326,N_14857,N_14938);
nor UO_1327 (O_1327,N_14976,N_14980);
nand UO_1328 (O_1328,N_14999,N_14963);
nor UO_1329 (O_1329,N_14925,N_14964);
nor UO_1330 (O_1330,N_14976,N_14884);
xnor UO_1331 (O_1331,N_14896,N_14915);
nand UO_1332 (O_1332,N_14917,N_14850);
nand UO_1333 (O_1333,N_14959,N_14947);
or UO_1334 (O_1334,N_14851,N_14914);
and UO_1335 (O_1335,N_14851,N_14946);
and UO_1336 (O_1336,N_14943,N_14921);
nand UO_1337 (O_1337,N_14874,N_14863);
nor UO_1338 (O_1338,N_14997,N_14975);
nand UO_1339 (O_1339,N_14994,N_14953);
or UO_1340 (O_1340,N_14852,N_14997);
and UO_1341 (O_1341,N_14990,N_14915);
nor UO_1342 (O_1342,N_14948,N_14996);
nand UO_1343 (O_1343,N_14853,N_14871);
xor UO_1344 (O_1344,N_14861,N_14927);
nand UO_1345 (O_1345,N_14969,N_14917);
or UO_1346 (O_1346,N_14997,N_14949);
nand UO_1347 (O_1347,N_14959,N_14955);
or UO_1348 (O_1348,N_14943,N_14896);
nand UO_1349 (O_1349,N_14941,N_14972);
nor UO_1350 (O_1350,N_14932,N_14901);
nand UO_1351 (O_1351,N_14977,N_14900);
or UO_1352 (O_1352,N_14907,N_14940);
or UO_1353 (O_1353,N_14895,N_14911);
nand UO_1354 (O_1354,N_14902,N_14862);
and UO_1355 (O_1355,N_14925,N_14910);
xnor UO_1356 (O_1356,N_14867,N_14893);
nor UO_1357 (O_1357,N_14999,N_14883);
nand UO_1358 (O_1358,N_14950,N_14854);
nor UO_1359 (O_1359,N_14962,N_14852);
and UO_1360 (O_1360,N_14990,N_14999);
or UO_1361 (O_1361,N_14956,N_14872);
nor UO_1362 (O_1362,N_14940,N_14873);
xnor UO_1363 (O_1363,N_14953,N_14910);
nor UO_1364 (O_1364,N_14907,N_14957);
nor UO_1365 (O_1365,N_14951,N_14965);
or UO_1366 (O_1366,N_14940,N_14915);
nand UO_1367 (O_1367,N_14871,N_14963);
nand UO_1368 (O_1368,N_14995,N_14937);
xor UO_1369 (O_1369,N_14993,N_14872);
or UO_1370 (O_1370,N_14918,N_14886);
nand UO_1371 (O_1371,N_14901,N_14940);
xor UO_1372 (O_1372,N_14976,N_14895);
or UO_1373 (O_1373,N_14906,N_14854);
and UO_1374 (O_1374,N_14892,N_14985);
and UO_1375 (O_1375,N_14887,N_14942);
and UO_1376 (O_1376,N_14922,N_14868);
and UO_1377 (O_1377,N_14883,N_14867);
nor UO_1378 (O_1378,N_14960,N_14938);
or UO_1379 (O_1379,N_14938,N_14859);
and UO_1380 (O_1380,N_14884,N_14944);
nor UO_1381 (O_1381,N_14863,N_14964);
nor UO_1382 (O_1382,N_14993,N_14970);
or UO_1383 (O_1383,N_14882,N_14852);
xor UO_1384 (O_1384,N_14965,N_14986);
and UO_1385 (O_1385,N_14879,N_14858);
nand UO_1386 (O_1386,N_14894,N_14958);
nor UO_1387 (O_1387,N_14914,N_14881);
nor UO_1388 (O_1388,N_14940,N_14925);
nor UO_1389 (O_1389,N_14936,N_14964);
nand UO_1390 (O_1390,N_14872,N_14928);
nor UO_1391 (O_1391,N_14869,N_14955);
nand UO_1392 (O_1392,N_14884,N_14954);
nand UO_1393 (O_1393,N_14908,N_14924);
or UO_1394 (O_1394,N_14975,N_14977);
and UO_1395 (O_1395,N_14906,N_14971);
nand UO_1396 (O_1396,N_14858,N_14977);
or UO_1397 (O_1397,N_14923,N_14960);
xnor UO_1398 (O_1398,N_14903,N_14996);
nand UO_1399 (O_1399,N_14971,N_14917);
and UO_1400 (O_1400,N_14995,N_14909);
xnor UO_1401 (O_1401,N_14865,N_14974);
xnor UO_1402 (O_1402,N_14921,N_14942);
nor UO_1403 (O_1403,N_14866,N_14890);
or UO_1404 (O_1404,N_14990,N_14991);
nor UO_1405 (O_1405,N_14912,N_14964);
xnor UO_1406 (O_1406,N_14864,N_14898);
nand UO_1407 (O_1407,N_14983,N_14899);
or UO_1408 (O_1408,N_14929,N_14851);
and UO_1409 (O_1409,N_14925,N_14949);
and UO_1410 (O_1410,N_14883,N_14874);
or UO_1411 (O_1411,N_14983,N_14872);
and UO_1412 (O_1412,N_14919,N_14858);
and UO_1413 (O_1413,N_14954,N_14975);
nand UO_1414 (O_1414,N_14969,N_14962);
nand UO_1415 (O_1415,N_14881,N_14967);
nor UO_1416 (O_1416,N_14951,N_14935);
nor UO_1417 (O_1417,N_14958,N_14995);
nor UO_1418 (O_1418,N_14963,N_14856);
or UO_1419 (O_1419,N_14991,N_14971);
nand UO_1420 (O_1420,N_14997,N_14961);
xnor UO_1421 (O_1421,N_14968,N_14907);
nor UO_1422 (O_1422,N_14979,N_14944);
xor UO_1423 (O_1423,N_14999,N_14881);
and UO_1424 (O_1424,N_14980,N_14936);
and UO_1425 (O_1425,N_14987,N_14874);
nand UO_1426 (O_1426,N_14987,N_14919);
and UO_1427 (O_1427,N_14954,N_14989);
and UO_1428 (O_1428,N_14948,N_14859);
nand UO_1429 (O_1429,N_14901,N_14860);
nor UO_1430 (O_1430,N_14971,N_14916);
and UO_1431 (O_1431,N_14909,N_14857);
nand UO_1432 (O_1432,N_14963,N_14903);
and UO_1433 (O_1433,N_14860,N_14878);
or UO_1434 (O_1434,N_14857,N_14986);
xnor UO_1435 (O_1435,N_14869,N_14970);
nand UO_1436 (O_1436,N_14961,N_14993);
xnor UO_1437 (O_1437,N_14879,N_14998);
or UO_1438 (O_1438,N_14952,N_14869);
and UO_1439 (O_1439,N_14995,N_14975);
or UO_1440 (O_1440,N_14975,N_14912);
or UO_1441 (O_1441,N_14862,N_14967);
and UO_1442 (O_1442,N_14885,N_14935);
nor UO_1443 (O_1443,N_14897,N_14884);
and UO_1444 (O_1444,N_14994,N_14863);
xor UO_1445 (O_1445,N_14988,N_14869);
nor UO_1446 (O_1446,N_14877,N_14990);
or UO_1447 (O_1447,N_14979,N_14912);
nand UO_1448 (O_1448,N_14921,N_14884);
xor UO_1449 (O_1449,N_14894,N_14915);
xnor UO_1450 (O_1450,N_14922,N_14882);
xnor UO_1451 (O_1451,N_14979,N_14907);
nand UO_1452 (O_1452,N_14880,N_14946);
xnor UO_1453 (O_1453,N_14957,N_14965);
or UO_1454 (O_1454,N_14978,N_14863);
and UO_1455 (O_1455,N_14931,N_14896);
and UO_1456 (O_1456,N_14872,N_14916);
xor UO_1457 (O_1457,N_14905,N_14875);
and UO_1458 (O_1458,N_14865,N_14948);
nand UO_1459 (O_1459,N_14954,N_14925);
and UO_1460 (O_1460,N_14856,N_14876);
or UO_1461 (O_1461,N_14905,N_14943);
nor UO_1462 (O_1462,N_14864,N_14955);
and UO_1463 (O_1463,N_14900,N_14934);
or UO_1464 (O_1464,N_14882,N_14994);
nor UO_1465 (O_1465,N_14889,N_14945);
xor UO_1466 (O_1466,N_14963,N_14919);
nor UO_1467 (O_1467,N_14955,N_14886);
nand UO_1468 (O_1468,N_14938,N_14947);
or UO_1469 (O_1469,N_14926,N_14858);
or UO_1470 (O_1470,N_14982,N_14967);
nor UO_1471 (O_1471,N_14969,N_14968);
xnor UO_1472 (O_1472,N_14889,N_14886);
nand UO_1473 (O_1473,N_14998,N_14965);
xnor UO_1474 (O_1474,N_14872,N_14858);
xor UO_1475 (O_1475,N_14855,N_14885);
and UO_1476 (O_1476,N_14935,N_14912);
xnor UO_1477 (O_1477,N_14884,N_14985);
and UO_1478 (O_1478,N_14994,N_14985);
nor UO_1479 (O_1479,N_14888,N_14974);
and UO_1480 (O_1480,N_14957,N_14994);
and UO_1481 (O_1481,N_14958,N_14884);
xor UO_1482 (O_1482,N_14899,N_14930);
or UO_1483 (O_1483,N_14921,N_14955);
nor UO_1484 (O_1484,N_14940,N_14950);
xor UO_1485 (O_1485,N_14957,N_14914);
nor UO_1486 (O_1486,N_14880,N_14961);
and UO_1487 (O_1487,N_14921,N_14919);
nand UO_1488 (O_1488,N_14893,N_14889);
nor UO_1489 (O_1489,N_14872,N_14953);
xor UO_1490 (O_1490,N_14992,N_14907);
xnor UO_1491 (O_1491,N_14889,N_14998);
nor UO_1492 (O_1492,N_14991,N_14880);
and UO_1493 (O_1493,N_14908,N_14917);
nor UO_1494 (O_1494,N_14880,N_14993);
and UO_1495 (O_1495,N_14893,N_14903);
xnor UO_1496 (O_1496,N_14916,N_14931);
or UO_1497 (O_1497,N_14867,N_14894);
or UO_1498 (O_1498,N_14892,N_14977);
nor UO_1499 (O_1499,N_14904,N_14877);
nand UO_1500 (O_1500,N_14894,N_14945);
xnor UO_1501 (O_1501,N_14944,N_14954);
and UO_1502 (O_1502,N_14892,N_14939);
nand UO_1503 (O_1503,N_14901,N_14965);
nand UO_1504 (O_1504,N_14903,N_14853);
and UO_1505 (O_1505,N_14866,N_14963);
nor UO_1506 (O_1506,N_14928,N_14927);
and UO_1507 (O_1507,N_14862,N_14968);
nor UO_1508 (O_1508,N_14955,N_14926);
or UO_1509 (O_1509,N_14888,N_14930);
nand UO_1510 (O_1510,N_14910,N_14954);
nand UO_1511 (O_1511,N_14896,N_14952);
nand UO_1512 (O_1512,N_14960,N_14980);
or UO_1513 (O_1513,N_14853,N_14896);
or UO_1514 (O_1514,N_14874,N_14858);
nand UO_1515 (O_1515,N_14950,N_14947);
nor UO_1516 (O_1516,N_14892,N_14940);
or UO_1517 (O_1517,N_14989,N_14914);
and UO_1518 (O_1518,N_14923,N_14902);
and UO_1519 (O_1519,N_14911,N_14956);
nor UO_1520 (O_1520,N_14861,N_14990);
nand UO_1521 (O_1521,N_14939,N_14997);
or UO_1522 (O_1522,N_14904,N_14917);
or UO_1523 (O_1523,N_14986,N_14899);
nand UO_1524 (O_1524,N_14930,N_14857);
or UO_1525 (O_1525,N_14933,N_14934);
and UO_1526 (O_1526,N_14881,N_14870);
nand UO_1527 (O_1527,N_14961,N_14992);
and UO_1528 (O_1528,N_14953,N_14969);
xnor UO_1529 (O_1529,N_14961,N_14981);
nand UO_1530 (O_1530,N_14992,N_14951);
or UO_1531 (O_1531,N_14994,N_14866);
nor UO_1532 (O_1532,N_14975,N_14967);
nor UO_1533 (O_1533,N_14883,N_14876);
nor UO_1534 (O_1534,N_14866,N_14926);
xor UO_1535 (O_1535,N_14905,N_14916);
xor UO_1536 (O_1536,N_14907,N_14974);
nor UO_1537 (O_1537,N_14908,N_14888);
nand UO_1538 (O_1538,N_14947,N_14940);
nor UO_1539 (O_1539,N_14929,N_14962);
nor UO_1540 (O_1540,N_14973,N_14957);
nand UO_1541 (O_1541,N_14970,N_14987);
nand UO_1542 (O_1542,N_14995,N_14969);
nand UO_1543 (O_1543,N_14935,N_14862);
nor UO_1544 (O_1544,N_14937,N_14991);
xor UO_1545 (O_1545,N_14873,N_14850);
nor UO_1546 (O_1546,N_14957,N_14858);
nor UO_1547 (O_1547,N_14977,N_14972);
nor UO_1548 (O_1548,N_14935,N_14908);
nor UO_1549 (O_1549,N_14921,N_14907);
xnor UO_1550 (O_1550,N_14871,N_14956);
or UO_1551 (O_1551,N_14961,N_14957);
nor UO_1552 (O_1552,N_14928,N_14877);
nand UO_1553 (O_1553,N_14924,N_14998);
nand UO_1554 (O_1554,N_14988,N_14974);
and UO_1555 (O_1555,N_14965,N_14884);
nand UO_1556 (O_1556,N_14937,N_14871);
or UO_1557 (O_1557,N_14867,N_14979);
and UO_1558 (O_1558,N_14989,N_14886);
or UO_1559 (O_1559,N_14944,N_14925);
and UO_1560 (O_1560,N_14905,N_14919);
xor UO_1561 (O_1561,N_14876,N_14991);
nor UO_1562 (O_1562,N_14991,N_14871);
xnor UO_1563 (O_1563,N_14911,N_14940);
nor UO_1564 (O_1564,N_14970,N_14874);
xnor UO_1565 (O_1565,N_14904,N_14895);
or UO_1566 (O_1566,N_14900,N_14936);
xnor UO_1567 (O_1567,N_14899,N_14973);
or UO_1568 (O_1568,N_14933,N_14889);
and UO_1569 (O_1569,N_14941,N_14921);
xor UO_1570 (O_1570,N_14934,N_14873);
nor UO_1571 (O_1571,N_14925,N_14912);
nor UO_1572 (O_1572,N_14937,N_14890);
xor UO_1573 (O_1573,N_14893,N_14894);
nor UO_1574 (O_1574,N_14903,N_14897);
xnor UO_1575 (O_1575,N_14894,N_14896);
or UO_1576 (O_1576,N_14982,N_14958);
xor UO_1577 (O_1577,N_14953,N_14949);
nor UO_1578 (O_1578,N_14867,N_14886);
xor UO_1579 (O_1579,N_14944,N_14901);
nor UO_1580 (O_1580,N_14940,N_14932);
nor UO_1581 (O_1581,N_14862,N_14938);
nand UO_1582 (O_1582,N_14977,N_14999);
and UO_1583 (O_1583,N_14930,N_14895);
nor UO_1584 (O_1584,N_14875,N_14980);
nor UO_1585 (O_1585,N_14926,N_14862);
nand UO_1586 (O_1586,N_14885,N_14917);
and UO_1587 (O_1587,N_14897,N_14997);
and UO_1588 (O_1588,N_14854,N_14979);
and UO_1589 (O_1589,N_14984,N_14854);
nor UO_1590 (O_1590,N_14935,N_14923);
nor UO_1591 (O_1591,N_14995,N_14914);
nand UO_1592 (O_1592,N_14964,N_14905);
nor UO_1593 (O_1593,N_14930,N_14951);
and UO_1594 (O_1594,N_14918,N_14898);
xor UO_1595 (O_1595,N_14917,N_14881);
nand UO_1596 (O_1596,N_14952,N_14972);
or UO_1597 (O_1597,N_14961,N_14921);
or UO_1598 (O_1598,N_14879,N_14882);
or UO_1599 (O_1599,N_14901,N_14964);
nor UO_1600 (O_1600,N_14940,N_14879);
nor UO_1601 (O_1601,N_14902,N_14892);
nand UO_1602 (O_1602,N_14979,N_14922);
nor UO_1603 (O_1603,N_14913,N_14984);
and UO_1604 (O_1604,N_14890,N_14910);
or UO_1605 (O_1605,N_14985,N_14853);
nand UO_1606 (O_1606,N_14925,N_14884);
nor UO_1607 (O_1607,N_14905,N_14887);
and UO_1608 (O_1608,N_14937,N_14859);
or UO_1609 (O_1609,N_14941,N_14992);
nand UO_1610 (O_1610,N_14860,N_14976);
or UO_1611 (O_1611,N_14875,N_14937);
nor UO_1612 (O_1612,N_14851,N_14994);
xnor UO_1613 (O_1613,N_14963,N_14930);
nand UO_1614 (O_1614,N_14864,N_14937);
nor UO_1615 (O_1615,N_14935,N_14875);
nor UO_1616 (O_1616,N_14887,N_14904);
and UO_1617 (O_1617,N_14963,N_14892);
and UO_1618 (O_1618,N_14854,N_14933);
nand UO_1619 (O_1619,N_14859,N_14944);
or UO_1620 (O_1620,N_14921,N_14935);
and UO_1621 (O_1621,N_14979,N_14968);
or UO_1622 (O_1622,N_14885,N_14867);
nor UO_1623 (O_1623,N_14897,N_14901);
and UO_1624 (O_1624,N_14855,N_14926);
and UO_1625 (O_1625,N_14994,N_14906);
or UO_1626 (O_1626,N_14951,N_14911);
and UO_1627 (O_1627,N_14850,N_14893);
nand UO_1628 (O_1628,N_14865,N_14906);
nor UO_1629 (O_1629,N_14886,N_14855);
nand UO_1630 (O_1630,N_14921,N_14909);
nand UO_1631 (O_1631,N_14959,N_14985);
xor UO_1632 (O_1632,N_14878,N_14960);
xor UO_1633 (O_1633,N_14921,N_14985);
nor UO_1634 (O_1634,N_14881,N_14970);
nand UO_1635 (O_1635,N_14984,N_14978);
nor UO_1636 (O_1636,N_14966,N_14981);
nand UO_1637 (O_1637,N_14955,N_14860);
nand UO_1638 (O_1638,N_14940,N_14900);
nor UO_1639 (O_1639,N_14927,N_14987);
and UO_1640 (O_1640,N_14988,N_14926);
xnor UO_1641 (O_1641,N_14883,N_14994);
and UO_1642 (O_1642,N_14877,N_14936);
and UO_1643 (O_1643,N_14938,N_14966);
or UO_1644 (O_1644,N_14889,N_14875);
or UO_1645 (O_1645,N_14931,N_14857);
or UO_1646 (O_1646,N_14919,N_14952);
nor UO_1647 (O_1647,N_14981,N_14971);
and UO_1648 (O_1648,N_14871,N_14950);
nand UO_1649 (O_1649,N_14990,N_14952);
nor UO_1650 (O_1650,N_14928,N_14914);
and UO_1651 (O_1651,N_14863,N_14941);
nor UO_1652 (O_1652,N_14930,N_14929);
nor UO_1653 (O_1653,N_14923,N_14971);
xnor UO_1654 (O_1654,N_14962,N_14872);
xor UO_1655 (O_1655,N_14873,N_14948);
or UO_1656 (O_1656,N_14968,N_14888);
xnor UO_1657 (O_1657,N_14935,N_14893);
xnor UO_1658 (O_1658,N_14910,N_14885);
nor UO_1659 (O_1659,N_14851,N_14920);
nor UO_1660 (O_1660,N_14988,N_14959);
or UO_1661 (O_1661,N_14850,N_14965);
and UO_1662 (O_1662,N_14918,N_14971);
and UO_1663 (O_1663,N_14987,N_14895);
and UO_1664 (O_1664,N_14931,N_14940);
or UO_1665 (O_1665,N_14976,N_14922);
xor UO_1666 (O_1666,N_14903,N_14902);
xor UO_1667 (O_1667,N_14867,N_14982);
nand UO_1668 (O_1668,N_14866,N_14856);
nor UO_1669 (O_1669,N_14954,N_14994);
nand UO_1670 (O_1670,N_14858,N_14997);
and UO_1671 (O_1671,N_14858,N_14895);
xor UO_1672 (O_1672,N_14856,N_14947);
xor UO_1673 (O_1673,N_14933,N_14857);
nand UO_1674 (O_1674,N_14964,N_14922);
or UO_1675 (O_1675,N_14948,N_14963);
or UO_1676 (O_1676,N_14977,N_14907);
or UO_1677 (O_1677,N_14995,N_14954);
nor UO_1678 (O_1678,N_14896,N_14929);
nor UO_1679 (O_1679,N_14994,N_14949);
xor UO_1680 (O_1680,N_14985,N_14863);
or UO_1681 (O_1681,N_14874,N_14884);
nand UO_1682 (O_1682,N_14995,N_14919);
and UO_1683 (O_1683,N_14878,N_14986);
xnor UO_1684 (O_1684,N_14984,N_14864);
nor UO_1685 (O_1685,N_14968,N_14896);
nor UO_1686 (O_1686,N_14998,N_14921);
nand UO_1687 (O_1687,N_14862,N_14892);
nor UO_1688 (O_1688,N_14937,N_14889);
nor UO_1689 (O_1689,N_14982,N_14962);
or UO_1690 (O_1690,N_14967,N_14890);
xnor UO_1691 (O_1691,N_14904,N_14851);
or UO_1692 (O_1692,N_14909,N_14934);
nand UO_1693 (O_1693,N_14852,N_14944);
nand UO_1694 (O_1694,N_14887,N_14983);
and UO_1695 (O_1695,N_14861,N_14971);
and UO_1696 (O_1696,N_14886,N_14854);
nand UO_1697 (O_1697,N_14933,N_14898);
or UO_1698 (O_1698,N_14890,N_14862);
nor UO_1699 (O_1699,N_14986,N_14931);
and UO_1700 (O_1700,N_14901,N_14937);
nand UO_1701 (O_1701,N_14851,N_14881);
or UO_1702 (O_1702,N_14981,N_14996);
and UO_1703 (O_1703,N_14855,N_14904);
nand UO_1704 (O_1704,N_14927,N_14950);
and UO_1705 (O_1705,N_14856,N_14962);
or UO_1706 (O_1706,N_14854,N_14939);
nor UO_1707 (O_1707,N_14927,N_14890);
or UO_1708 (O_1708,N_14854,N_14977);
or UO_1709 (O_1709,N_14989,N_14999);
xor UO_1710 (O_1710,N_14868,N_14927);
nand UO_1711 (O_1711,N_14872,N_14870);
or UO_1712 (O_1712,N_14887,N_14888);
xnor UO_1713 (O_1713,N_14970,N_14890);
or UO_1714 (O_1714,N_14940,N_14972);
nand UO_1715 (O_1715,N_14965,N_14867);
and UO_1716 (O_1716,N_14939,N_14971);
nor UO_1717 (O_1717,N_14895,N_14875);
and UO_1718 (O_1718,N_14939,N_14949);
xnor UO_1719 (O_1719,N_14863,N_14916);
nand UO_1720 (O_1720,N_14854,N_14964);
nand UO_1721 (O_1721,N_14930,N_14999);
and UO_1722 (O_1722,N_14944,N_14946);
nand UO_1723 (O_1723,N_14916,N_14992);
or UO_1724 (O_1724,N_14907,N_14898);
or UO_1725 (O_1725,N_14965,N_14873);
xnor UO_1726 (O_1726,N_14865,N_14876);
or UO_1727 (O_1727,N_14932,N_14979);
or UO_1728 (O_1728,N_14985,N_14919);
nand UO_1729 (O_1729,N_14858,N_14943);
and UO_1730 (O_1730,N_14869,N_14994);
xnor UO_1731 (O_1731,N_14902,N_14932);
xor UO_1732 (O_1732,N_14860,N_14870);
or UO_1733 (O_1733,N_14986,N_14962);
nor UO_1734 (O_1734,N_14885,N_14852);
nand UO_1735 (O_1735,N_14984,N_14952);
nand UO_1736 (O_1736,N_14946,N_14860);
nor UO_1737 (O_1737,N_14962,N_14884);
or UO_1738 (O_1738,N_14931,N_14888);
xnor UO_1739 (O_1739,N_14869,N_14888);
and UO_1740 (O_1740,N_14946,N_14878);
xor UO_1741 (O_1741,N_14944,N_14862);
nor UO_1742 (O_1742,N_14910,N_14998);
nor UO_1743 (O_1743,N_14985,N_14876);
nand UO_1744 (O_1744,N_14863,N_14925);
and UO_1745 (O_1745,N_14946,N_14865);
nand UO_1746 (O_1746,N_14979,N_14903);
xor UO_1747 (O_1747,N_14942,N_14913);
nor UO_1748 (O_1748,N_14958,N_14976);
and UO_1749 (O_1749,N_14863,N_14971);
xnor UO_1750 (O_1750,N_14904,N_14863);
and UO_1751 (O_1751,N_14886,N_14881);
nand UO_1752 (O_1752,N_14916,N_14924);
nor UO_1753 (O_1753,N_14882,N_14889);
or UO_1754 (O_1754,N_14915,N_14988);
xnor UO_1755 (O_1755,N_14902,N_14878);
and UO_1756 (O_1756,N_14982,N_14850);
nor UO_1757 (O_1757,N_14883,N_14992);
and UO_1758 (O_1758,N_14927,N_14908);
nor UO_1759 (O_1759,N_14995,N_14870);
and UO_1760 (O_1760,N_14993,N_14934);
and UO_1761 (O_1761,N_14968,N_14935);
nor UO_1762 (O_1762,N_14930,N_14996);
nor UO_1763 (O_1763,N_14931,N_14954);
nor UO_1764 (O_1764,N_14910,N_14926);
nand UO_1765 (O_1765,N_14930,N_14908);
or UO_1766 (O_1766,N_14936,N_14899);
nor UO_1767 (O_1767,N_14942,N_14999);
or UO_1768 (O_1768,N_14860,N_14917);
nor UO_1769 (O_1769,N_14867,N_14858);
nor UO_1770 (O_1770,N_14946,N_14958);
nand UO_1771 (O_1771,N_14900,N_14976);
and UO_1772 (O_1772,N_14899,N_14947);
or UO_1773 (O_1773,N_14937,N_14932);
nor UO_1774 (O_1774,N_14871,N_14899);
and UO_1775 (O_1775,N_14938,N_14863);
xor UO_1776 (O_1776,N_14857,N_14997);
xor UO_1777 (O_1777,N_14971,N_14961);
nor UO_1778 (O_1778,N_14940,N_14929);
nand UO_1779 (O_1779,N_14966,N_14923);
nor UO_1780 (O_1780,N_14870,N_14912);
and UO_1781 (O_1781,N_14919,N_14927);
nand UO_1782 (O_1782,N_14903,N_14922);
nand UO_1783 (O_1783,N_14870,N_14879);
xnor UO_1784 (O_1784,N_14945,N_14959);
nand UO_1785 (O_1785,N_14859,N_14940);
or UO_1786 (O_1786,N_14864,N_14967);
xor UO_1787 (O_1787,N_14926,N_14962);
xnor UO_1788 (O_1788,N_14946,N_14907);
nor UO_1789 (O_1789,N_14900,N_14912);
nand UO_1790 (O_1790,N_14932,N_14981);
and UO_1791 (O_1791,N_14853,N_14953);
or UO_1792 (O_1792,N_14989,N_14970);
xnor UO_1793 (O_1793,N_14858,N_14986);
nand UO_1794 (O_1794,N_14904,N_14873);
or UO_1795 (O_1795,N_14874,N_14860);
nor UO_1796 (O_1796,N_14886,N_14931);
or UO_1797 (O_1797,N_14981,N_14900);
nor UO_1798 (O_1798,N_14868,N_14920);
and UO_1799 (O_1799,N_14916,N_14927);
xnor UO_1800 (O_1800,N_14862,N_14864);
nand UO_1801 (O_1801,N_14977,N_14903);
nor UO_1802 (O_1802,N_14897,N_14963);
xnor UO_1803 (O_1803,N_14874,N_14942);
nor UO_1804 (O_1804,N_14910,N_14947);
nand UO_1805 (O_1805,N_14858,N_14889);
and UO_1806 (O_1806,N_14935,N_14976);
nor UO_1807 (O_1807,N_14998,N_14941);
nor UO_1808 (O_1808,N_14924,N_14855);
nor UO_1809 (O_1809,N_14912,N_14872);
nand UO_1810 (O_1810,N_14940,N_14906);
nor UO_1811 (O_1811,N_14933,N_14915);
nand UO_1812 (O_1812,N_14851,N_14922);
nor UO_1813 (O_1813,N_14944,N_14978);
nand UO_1814 (O_1814,N_14879,N_14925);
xor UO_1815 (O_1815,N_14981,N_14861);
nand UO_1816 (O_1816,N_14882,N_14871);
xor UO_1817 (O_1817,N_14851,N_14963);
nor UO_1818 (O_1818,N_14955,N_14946);
and UO_1819 (O_1819,N_14873,N_14878);
and UO_1820 (O_1820,N_14916,N_14870);
xor UO_1821 (O_1821,N_14889,N_14948);
nand UO_1822 (O_1822,N_14860,N_14890);
and UO_1823 (O_1823,N_14987,N_14981);
or UO_1824 (O_1824,N_14886,N_14861);
nor UO_1825 (O_1825,N_14970,N_14851);
and UO_1826 (O_1826,N_14885,N_14915);
nor UO_1827 (O_1827,N_14955,N_14980);
nor UO_1828 (O_1828,N_14950,N_14982);
xor UO_1829 (O_1829,N_14946,N_14947);
xor UO_1830 (O_1830,N_14986,N_14872);
and UO_1831 (O_1831,N_14987,N_14909);
xor UO_1832 (O_1832,N_14972,N_14852);
xnor UO_1833 (O_1833,N_14941,N_14991);
nand UO_1834 (O_1834,N_14935,N_14916);
xor UO_1835 (O_1835,N_14864,N_14854);
nand UO_1836 (O_1836,N_14915,N_14996);
nand UO_1837 (O_1837,N_14944,N_14887);
or UO_1838 (O_1838,N_14916,N_14901);
and UO_1839 (O_1839,N_14890,N_14872);
nand UO_1840 (O_1840,N_14957,N_14891);
nand UO_1841 (O_1841,N_14962,N_14941);
and UO_1842 (O_1842,N_14922,N_14854);
and UO_1843 (O_1843,N_14888,N_14972);
xnor UO_1844 (O_1844,N_14870,N_14867);
nand UO_1845 (O_1845,N_14961,N_14988);
xor UO_1846 (O_1846,N_14862,N_14912);
and UO_1847 (O_1847,N_14963,N_14940);
or UO_1848 (O_1848,N_14920,N_14941);
nand UO_1849 (O_1849,N_14939,N_14987);
nand UO_1850 (O_1850,N_14900,N_14972);
and UO_1851 (O_1851,N_14996,N_14934);
or UO_1852 (O_1852,N_14975,N_14879);
and UO_1853 (O_1853,N_14866,N_14968);
and UO_1854 (O_1854,N_14885,N_14874);
or UO_1855 (O_1855,N_14867,N_14980);
xor UO_1856 (O_1856,N_14856,N_14914);
and UO_1857 (O_1857,N_14904,N_14992);
or UO_1858 (O_1858,N_14956,N_14879);
xor UO_1859 (O_1859,N_14958,N_14915);
nand UO_1860 (O_1860,N_14940,N_14973);
xnor UO_1861 (O_1861,N_14881,N_14955);
nand UO_1862 (O_1862,N_14905,N_14952);
and UO_1863 (O_1863,N_14879,N_14905);
xor UO_1864 (O_1864,N_14862,N_14868);
nand UO_1865 (O_1865,N_14986,N_14939);
xnor UO_1866 (O_1866,N_14959,N_14867);
xnor UO_1867 (O_1867,N_14871,N_14954);
nor UO_1868 (O_1868,N_14952,N_14928);
or UO_1869 (O_1869,N_14981,N_14927);
xnor UO_1870 (O_1870,N_14855,N_14859);
or UO_1871 (O_1871,N_14990,N_14969);
and UO_1872 (O_1872,N_14959,N_14987);
or UO_1873 (O_1873,N_14936,N_14971);
nand UO_1874 (O_1874,N_14965,N_14896);
and UO_1875 (O_1875,N_14923,N_14988);
xnor UO_1876 (O_1876,N_14937,N_14921);
nor UO_1877 (O_1877,N_14971,N_14987);
and UO_1878 (O_1878,N_14998,N_14968);
nand UO_1879 (O_1879,N_14921,N_14949);
and UO_1880 (O_1880,N_14932,N_14995);
or UO_1881 (O_1881,N_14994,N_14932);
nor UO_1882 (O_1882,N_14872,N_14907);
nor UO_1883 (O_1883,N_14905,N_14963);
nand UO_1884 (O_1884,N_14984,N_14932);
and UO_1885 (O_1885,N_14860,N_14941);
and UO_1886 (O_1886,N_14865,N_14896);
and UO_1887 (O_1887,N_14868,N_14969);
and UO_1888 (O_1888,N_14960,N_14979);
nor UO_1889 (O_1889,N_14996,N_14871);
xnor UO_1890 (O_1890,N_14953,N_14958);
xor UO_1891 (O_1891,N_14919,N_14893);
and UO_1892 (O_1892,N_14871,N_14895);
xor UO_1893 (O_1893,N_14980,N_14939);
xnor UO_1894 (O_1894,N_14879,N_14890);
nand UO_1895 (O_1895,N_14856,N_14992);
nor UO_1896 (O_1896,N_14902,N_14928);
nand UO_1897 (O_1897,N_14911,N_14885);
nor UO_1898 (O_1898,N_14883,N_14980);
or UO_1899 (O_1899,N_14884,N_14966);
nand UO_1900 (O_1900,N_14855,N_14875);
nor UO_1901 (O_1901,N_14947,N_14986);
nor UO_1902 (O_1902,N_14987,N_14872);
nand UO_1903 (O_1903,N_14927,N_14870);
xnor UO_1904 (O_1904,N_14874,N_14972);
and UO_1905 (O_1905,N_14859,N_14973);
or UO_1906 (O_1906,N_14904,N_14864);
and UO_1907 (O_1907,N_14890,N_14905);
or UO_1908 (O_1908,N_14942,N_14992);
xnor UO_1909 (O_1909,N_14933,N_14866);
xnor UO_1910 (O_1910,N_14948,N_14902);
nor UO_1911 (O_1911,N_14948,N_14995);
nor UO_1912 (O_1912,N_14993,N_14923);
or UO_1913 (O_1913,N_14915,N_14953);
nor UO_1914 (O_1914,N_14922,N_14944);
or UO_1915 (O_1915,N_14998,N_14937);
or UO_1916 (O_1916,N_14964,N_14924);
nand UO_1917 (O_1917,N_14956,N_14895);
xnor UO_1918 (O_1918,N_14996,N_14969);
and UO_1919 (O_1919,N_14947,N_14900);
xor UO_1920 (O_1920,N_14999,N_14943);
nand UO_1921 (O_1921,N_14950,N_14890);
and UO_1922 (O_1922,N_14996,N_14916);
and UO_1923 (O_1923,N_14953,N_14947);
xnor UO_1924 (O_1924,N_14997,N_14978);
nor UO_1925 (O_1925,N_14900,N_14908);
and UO_1926 (O_1926,N_14920,N_14999);
nand UO_1927 (O_1927,N_14969,N_14987);
and UO_1928 (O_1928,N_14933,N_14911);
nand UO_1929 (O_1929,N_14963,N_14858);
and UO_1930 (O_1930,N_14989,N_14909);
or UO_1931 (O_1931,N_14959,N_14977);
or UO_1932 (O_1932,N_14862,N_14920);
or UO_1933 (O_1933,N_14963,N_14883);
or UO_1934 (O_1934,N_14988,N_14951);
or UO_1935 (O_1935,N_14863,N_14858);
or UO_1936 (O_1936,N_14866,N_14947);
or UO_1937 (O_1937,N_14943,N_14973);
xnor UO_1938 (O_1938,N_14988,N_14940);
and UO_1939 (O_1939,N_14970,N_14955);
nor UO_1940 (O_1940,N_14915,N_14889);
or UO_1941 (O_1941,N_14882,N_14948);
nand UO_1942 (O_1942,N_14897,N_14913);
and UO_1943 (O_1943,N_14917,N_14902);
nor UO_1944 (O_1944,N_14929,N_14942);
nor UO_1945 (O_1945,N_14949,N_14974);
nand UO_1946 (O_1946,N_14993,N_14988);
and UO_1947 (O_1947,N_14876,N_14942);
nor UO_1948 (O_1948,N_14909,N_14982);
nor UO_1949 (O_1949,N_14877,N_14996);
nor UO_1950 (O_1950,N_14988,N_14963);
and UO_1951 (O_1951,N_14995,N_14883);
or UO_1952 (O_1952,N_14860,N_14914);
nand UO_1953 (O_1953,N_14997,N_14896);
and UO_1954 (O_1954,N_14891,N_14867);
and UO_1955 (O_1955,N_14991,N_14979);
and UO_1956 (O_1956,N_14898,N_14850);
or UO_1957 (O_1957,N_14879,N_14875);
nor UO_1958 (O_1958,N_14916,N_14928);
or UO_1959 (O_1959,N_14999,N_14993);
nor UO_1960 (O_1960,N_14930,N_14925);
nand UO_1961 (O_1961,N_14882,N_14988);
and UO_1962 (O_1962,N_14867,N_14964);
and UO_1963 (O_1963,N_14994,N_14964);
and UO_1964 (O_1964,N_14906,N_14850);
nor UO_1965 (O_1965,N_14991,N_14872);
nor UO_1966 (O_1966,N_14935,N_14973);
xnor UO_1967 (O_1967,N_14947,N_14930);
or UO_1968 (O_1968,N_14969,N_14982);
or UO_1969 (O_1969,N_14994,N_14877);
xnor UO_1970 (O_1970,N_14990,N_14918);
xor UO_1971 (O_1971,N_14871,N_14916);
nand UO_1972 (O_1972,N_14948,N_14985);
and UO_1973 (O_1973,N_14884,N_14971);
nor UO_1974 (O_1974,N_14908,N_14968);
nor UO_1975 (O_1975,N_14855,N_14892);
or UO_1976 (O_1976,N_14959,N_14881);
or UO_1977 (O_1977,N_14953,N_14976);
xnor UO_1978 (O_1978,N_14913,N_14877);
nor UO_1979 (O_1979,N_14984,N_14917);
or UO_1980 (O_1980,N_14871,N_14960);
nand UO_1981 (O_1981,N_14965,N_14958);
and UO_1982 (O_1982,N_14980,N_14992);
nand UO_1983 (O_1983,N_14945,N_14942);
nor UO_1984 (O_1984,N_14919,N_14989);
nand UO_1985 (O_1985,N_14854,N_14976);
and UO_1986 (O_1986,N_14973,N_14942);
xor UO_1987 (O_1987,N_14876,N_14983);
nand UO_1988 (O_1988,N_14910,N_14893);
and UO_1989 (O_1989,N_14992,N_14965);
xnor UO_1990 (O_1990,N_14859,N_14875);
nor UO_1991 (O_1991,N_14969,N_14974);
and UO_1992 (O_1992,N_14874,N_14967);
nand UO_1993 (O_1993,N_14955,N_14915);
xnor UO_1994 (O_1994,N_14857,N_14915);
and UO_1995 (O_1995,N_14913,N_14952);
nand UO_1996 (O_1996,N_14951,N_14850);
or UO_1997 (O_1997,N_14905,N_14930);
and UO_1998 (O_1998,N_14863,N_14890);
xnor UO_1999 (O_1999,N_14943,N_14944);
endmodule