module basic_500_3000_500_60_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_67,In_273);
nor U1 (N_1,In_487,In_448);
nor U2 (N_2,In_355,In_155);
nand U3 (N_3,In_357,In_30);
xor U4 (N_4,In_331,In_211);
nand U5 (N_5,In_437,In_449);
or U6 (N_6,In_152,In_108);
or U7 (N_7,In_317,In_271);
nand U8 (N_8,In_176,In_324);
nand U9 (N_9,In_354,In_256);
xor U10 (N_10,In_353,In_378);
or U11 (N_11,In_148,In_164);
and U12 (N_12,In_304,In_62);
and U13 (N_13,In_165,In_139);
nand U14 (N_14,In_429,In_124);
nand U15 (N_15,In_370,In_20);
nand U16 (N_16,In_54,In_91);
or U17 (N_17,In_470,In_296);
and U18 (N_18,In_8,In_446);
nor U19 (N_19,In_434,In_102);
or U20 (N_20,In_258,In_371);
nor U21 (N_21,In_295,In_206);
nor U22 (N_22,In_74,In_68);
or U23 (N_23,In_178,In_478);
and U24 (N_24,In_460,In_229);
nor U25 (N_25,In_484,In_366);
nand U26 (N_26,In_40,In_336);
nand U27 (N_27,In_230,In_294);
and U28 (N_28,In_315,In_187);
nor U29 (N_29,In_472,In_406);
or U30 (N_30,In_392,In_220);
nand U31 (N_31,In_49,In_22);
nand U32 (N_32,In_466,In_32);
nand U33 (N_33,In_272,In_432);
nand U34 (N_34,In_401,In_403);
and U35 (N_35,In_42,In_408);
nand U36 (N_36,In_66,In_467);
nand U37 (N_37,In_239,In_480);
xor U38 (N_38,In_126,In_443);
xor U39 (N_39,In_6,In_377);
or U40 (N_40,In_435,In_422);
xor U41 (N_41,In_34,In_363);
nor U42 (N_42,In_56,In_426);
nand U43 (N_43,In_360,In_409);
or U44 (N_44,In_439,In_16);
nor U45 (N_45,In_402,In_495);
and U46 (N_46,In_85,In_87);
or U47 (N_47,In_29,In_395);
nor U48 (N_48,In_23,In_288);
nor U49 (N_49,In_468,In_337);
nand U50 (N_50,In_129,In_442);
and U51 (N_51,In_162,In_43);
nor U52 (N_52,In_151,In_398);
nand U53 (N_53,In_51,In_420);
or U54 (N_54,In_463,In_69);
and U55 (N_55,In_269,N_40);
and U56 (N_56,In_223,In_326);
or U57 (N_57,In_216,N_9);
and U58 (N_58,In_3,In_339);
nor U59 (N_59,In_209,In_356);
nor U60 (N_60,In_298,In_341);
nor U61 (N_61,In_416,In_334);
nand U62 (N_62,In_419,In_367);
nor U63 (N_63,In_455,In_184);
nor U64 (N_64,In_332,In_35);
nor U65 (N_65,In_219,N_34);
and U66 (N_66,In_33,In_14);
nand U67 (N_67,In_10,In_57);
or U68 (N_68,In_247,In_462);
nand U69 (N_69,In_405,In_465);
and U70 (N_70,In_103,In_143);
nor U71 (N_71,In_488,In_347);
nor U72 (N_72,In_414,In_375);
xor U73 (N_73,In_7,In_399);
nand U74 (N_74,In_425,In_179);
or U75 (N_75,In_44,In_485);
nand U76 (N_76,In_145,In_84);
and U77 (N_77,In_191,In_352);
nand U78 (N_78,In_415,In_246);
or U79 (N_79,In_170,In_167);
and U80 (N_80,In_474,In_438);
nand U81 (N_81,In_496,In_78);
and U82 (N_82,In_286,In_476);
nand U83 (N_83,In_88,In_413);
or U84 (N_84,N_1,In_127);
nor U85 (N_85,In_86,In_45);
nor U86 (N_86,In_380,In_492);
nor U87 (N_87,In_193,In_199);
and U88 (N_88,In_201,In_259);
nand U89 (N_89,In_106,In_115);
nand U90 (N_90,In_477,In_311);
xor U91 (N_91,In_77,In_257);
or U92 (N_92,In_335,In_323);
or U93 (N_93,In_329,In_25);
or U94 (N_94,In_140,In_365);
and U95 (N_95,In_109,N_25);
and U96 (N_96,In_96,In_190);
or U97 (N_97,In_278,In_58);
xor U98 (N_98,In_15,In_142);
or U99 (N_99,In_252,In_338);
nor U100 (N_100,In_130,In_79);
and U101 (N_101,In_359,In_279);
or U102 (N_102,In_100,N_83);
nand U103 (N_103,In_232,In_447);
or U104 (N_104,In_38,In_391);
or U105 (N_105,In_307,In_90);
nor U106 (N_106,In_224,N_70);
and U107 (N_107,N_49,In_228);
nand U108 (N_108,In_445,In_452);
nor U109 (N_109,In_430,In_168);
and U110 (N_110,In_404,In_469);
xnor U111 (N_111,In_372,In_111);
and U112 (N_112,In_348,In_458);
xor U113 (N_113,N_10,N_35);
nor U114 (N_114,In_301,In_237);
or U115 (N_115,In_154,In_158);
nor U116 (N_116,In_222,In_72);
and U117 (N_117,In_235,In_19);
and U118 (N_118,In_384,In_198);
or U119 (N_119,In_362,In_342);
or U120 (N_120,In_400,N_5);
and U121 (N_121,In_456,In_379);
nor U122 (N_122,N_54,N_47);
nor U123 (N_123,In_5,In_451);
or U124 (N_124,In_289,N_32);
nand U125 (N_125,In_11,In_489);
and U126 (N_126,In_9,In_61);
or U127 (N_127,In_188,In_159);
nor U128 (N_128,In_174,In_101);
nand U129 (N_129,In_350,In_284);
or U130 (N_130,In_241,In_1);
nand U131 (N_131,N_95,In_183);
and U132 (N_132,In_381,N_98);
nand U133 (N_133,In_459,N_57);
nor U134 (N_134,In_94,In_48);
nor U135 (N_135,In_128,In_24);
and U136 (N_136,In_196,In_475);
nor U137 (N_137,N_94,In_95);
and U138 (N_138,N_77,In_358);
nand U139 (N_139,In_441,N_7);
nor U140 (N_140,In_299,In_76);
or U141 (N_141,In_156,In_104);
nand U142 (N_142,In_177,In_316);
nand U143 (N_143,In_283,In_471);
nor U144 (N_144,In_412,N_62);
nor U145 (N_145,N_74,In_464);
and U146 (N_146,In_312,In_123);
nand U147 (N_147,In_134,In_208);
and U148 (N_148,In_75,In_138);
xnor U149 (N_149,In_189,In_262);
xnor U150 (N_150,N_0,N_36);
nor U151 (N_151,In_233,In_493);
nand U152 (N_152,N_79,N_96);
xor U153 (N_153,In_81,In_263);
nand U154 (N_154,In_248,In_93);
or U155 (N_155,In_393,In_265);
nand U156 (N_156,In_397,In_213);
nor U157 (N_157,N_91,In_36);
nand U158 (N_158,N_51,N_55);
nand U159 (N_159,In_110,In_97);
or U160 (N_160,N_100,In_65);
nand U161 (N_161,N_131,N_43);
nand U162 (N_162,N_128,N_133);
xor U163 (N_163,N_97,In_321);
xnor U164 (N_164,N_3,In_287);
nor U165 (N_165,In_306,N_132);
nand U166 (N_166,In_82,In_389);
or U167 (N_167,In_133,In_141);
and U168 (N_168,In_157,In_276);
and U169 (N_169,N_11,In_346);
nand U170 (N_170,N_56,In_116);
nand U171 (N_171,In_107,N_80);
or U172 (N_172,In_499,In_227);
or U173 (N_173,In_411,In_112);
and U174 (N_174,In_436,In_270);
or U175 (N_175,N_142,In_238);
or U176 (N_176,N_147,N_104);
or U177 (N_177,N_67,In_70);
or U178 (N_178,In_431,In_394);
nor U179 (N_179,In_345,In_310);
nor U180 (N_180,In_374,In_4);
nand U181 (N_181,In_264,In_105);
and U182 (N_182,N_24,N_105);
nor U183 (N_183,N_89,N_39);
nor U184 (N_184,In_234,In_386);
or U185 (N_185,In_266,In_173);
nor U186 (N_186,In_147,In_387);
nand U187 (N_187,N_134,In_433);
nor U188 (N_188,In_320,N_103);
or U189 (N_189,In_308,In_121);
or U190 (N_190,In_98,In_225);
or U191 (N_191,N_52,In_254);
nand U192 (N_192,In_285,In_59);
nor U193 (N_193,In_214,In_163);
nor U194 (N_194,In_71,N_26);
and U195 (N_195,N_108,In_39);
xor U196 (N_196,In_250,N_87);
nand U197 (N_197,In_125,In_309);
or U198 (N_198,In_146,N_85);
nor U199 (N_199,In_344,N_21);
or U200 (N_200,In_17,In_364);
xnor U201 (N_201,N_28,In_497);
or U202 (N_202,In_63,In_251);
nand U203 (N_203,In_131,In_55);
nor U204 (N_204,N_193,N_154);
or U205 (N_205,N_58,N_61);
or U206 (N_206,In_268,N_181);
nor U207 (N_207,In_203,N_149);
nor U208 (N_208,N_136,In_13);
nor U209 (N_209,In_114,In_473);
and U210 (N_210,In_382,N_164);
nor U211 (N_211,In_12,N_76);
nand U212 (N_212,In_150,N_41);
and U213 (N_213,N_153,In_275);
nor U214 (N_214,In_351,In_293);
and U215 (N_215,In_161,In_319);
nand U216 (N_216,In_169,N_152);
and U217 (N_217,N_110,N_185);
nor U218 (N_218,In_53,In_195);
and U219 (N_219,N_157,In_491);
and U220 (N_220,N_199,In_290);
and U221 (N_221,In_383,In_483);
and U222 (N_222,N_46,N_22);
or U223 (N_223,In_349,In_282);
and U224 (N_224,N_44,N_184);
and U225 (N_225,N_68,In_322);
xnor U226 (N_226,N_141,N_116);
or U227 (N_227,In_277,N_163);
or U228 (N_228,N_64,In_160);
nand U229 (N_229,N_50,N_107);
and U230 (N_230,In_424,In_255);
xnor U231 (N_231,N_135,In_80);
or U232 (N_232,N_146,In_457);
nor U233 (N_233,In_454,In_200);
and U234 (N_234,N_78,In_181);
nor U235 (N_235,N_59,In_2);
xor U236 (N_236,N_82,N_92);
and U237 (N_237,In_92,In_26);
and U238 (N_238,In_482,In_297);
nand U239 (N_239,In_204,In_328);
xor U240 (N_240,In_410,N_101);
and U241 (N_241,N_86,N_81);
and U242 (N_242,N_129,In_302);
and U243 (N_243,In_444,In_260);
or U244 (N_244,In_120,N_171);
and U245 (N_245,In_314,In_243);
nor U246 (N_246,N_45,In_253);
or U247 (N_247,In_361,N_126);
and U248 (N_248,In_99,N_48);
nor U249 (N_249,N_138,N_102);
xor U250 (N_250,In_421,N_20);
or U251 (N_251,In_194,In_292);
nand U252 (N_252,N_139,N_228);
nand U253 (N_253,N_167,N_183);
or U254 (N_254,N_188,In_135);
nand U255 (N_255,N_207,N_118);
nand U256 (N_256,In_407,N_214);
nor U257 (N_257,N_173,N_38);
nor U258 (N_258,N_195,N_209);
or U259 (N_259,N_14,N_166);
nor U260 (N_260,N_65,N_180);
nand U261 (N_261,N_224,In_368);
and U262 (N_262,N_120,N_53);
nand U263 (N_263,N_234,N_182);
or U264 (N_264,N_192,N_161);
or U265 (N_265,N_223,N_127);
nand U266 (N_266,In_83,In_153);
and U267 (N_267,N_75,N_169);
nand U268 (N_268,N_227,In_215);
and U269 (N_269,In_440,In_144);
nand U270 (N_270,N_114,In_31);
and U271 (N_271,N_29,N_66);
nor U272 (N_272,N_4,In_137);
nand U273 (N_273,In_305,N_143);
and U274 (N_274,N_230,In_333);
and U275 (N_275,N_179,N_244);
or U276 (N_276,N_148,In_369);
and U277 (N_277,N_201,In_50);
nor U278 (N_278,In_245,N_151);
nand U279 (N_279,In_267,In_180);
nor U280 (N_280,N_73,In_89);
and U281 (N_281,N_162,N_90);
or U282 (N_282,In_212,In_494);
and U283 (N_283,In_202,N_219);
nor U284 (N_284,In_481,In_52);
or U285 (N_285,In_291,N_93);
or U286 (N_286,In_244,N_177);
xnor U287 (N_287,N_248,In_175);
or U288 (N_288,In_390,In_166);
xnor U289 (N_289,In_325,N_145);
nand U290 (N_290,In_205,N_247);
nand U291 (N_291,In_236,In_318);
and U292 (N_292,N_150,N_235);
and U293 (N_293,In_281,In_327);
or U294 (N_294,N_196,N_190);
nor U295 (N_295,In_428,N_13);
and U296 (N_296,In_28,N_208);
and U297 (N_297,N_63,In_217);
nor U298 (N_298,In_18,In_274);
nand U299 (N_299,N_170,In_186);
or U300 (N_300,In_197,N_200);
nor U301 (N_301,In_60,N_88);
and U302 (N_302,N_299,N_243);
or U303 (N_303,In_122,N_175);
and U304 (N_304,In_185,N_187);
and U305 (N_305,In_218,N_19);
nand U306 (N_306,N_294,N_264);
nor U307 (N_307,In_343,N_254);
and U308 (N_308,N_123,N_269);
nor U309 (N_309,N_109,In_427);
nand U310 (N_310,N_226,In_73);
and U311 (N_311,N_160,In_41);
and U312 (N_312,N_267,N_191);
xnor U313 (N_313,N_111,N_178);
or U314 (N_314,N_241,N_15);
and U315 (N_315,In_226,In_132);
xnor U316 (N_316,In_396,In_261);
and U317 (N_317,N_237,N_176);
or U318 (N_318,N_198,In_453);
or U319 (N_319,N_194,In_388);
nor U320 (N_320,N_211,In_385);
nand U321 (N_321,In_486,N_202);
xor U322 (N_322,N_258,In_64);
xnor U323 (N_323,In_207,N_225);
or U324 (N_324,N_255,In_490);
nor U325 (N_325,In_313,In_21);
nand U326 (N_326,In_450,N_246);
nand U327 (N_327,N_159,N_220);
nor U328 (N_328,N_130,In_46);
nand U329 (N_329,In_242,N_156);
nand U330 (N_330,In_231,N_286);
nand U331 (N_331,N_245,N_275);
nand U332 (N_332,In_172,In_418);
and U333 (N_333,N_16,N_271);
nor U334 (N_334,N_229,N_213);
or U335 (N_335,N_298,N_204);
nand U336 (N_336,N_115,In_300);
or U337 (N_337,N_119,N_297);
xnor U338 (N_338,N_273,N_296);
and U339 (N_339,In_118,N_289);
or U340 (N_340,N_221,N_251);
or U341 (N_341,N_232,N_84);
nor U342 (N_342,N_242,N_33);
and U343 (N_343,N_282,N_290);
nand U344 (N_344,N_263,In_340);
nor U345 (N_345,N_288,N_293);
nand U346 (N_346,N_144,In_149);
xnor U347 (N_347,N_17,N_253);
nor U348 (N_348,N_295,N_233);
nor U349 (N_349,N_215,In_479);
nand U350 (N_350,N_340,N_283);
xor U351 (N_351,N_60,N_238);
xnor U352 (N_352,N_323,N_312);
or U353 (N_353,N_42,N_330);
or U354 (N_354,N_268,N_2);
nand U355 (N_355,N_31,N_333);
or U356 (N_356,N_222,In_210);
nor U357 (N_357,N_125,N_23);
or U358 (N_358,N_117,N_318);
nand U359 (N_359,In_376,In_192);
or U360 (N_360,In_280,In_47);
nand U361 (N_361,N_336,N_306);
nand U362 (N_362,N_328,N_218);
nand U363 (N_363,N_210,N_155);
nand U364 (N_364,In_27,N_343);
nand U365 (N_365,N_285,N_265);
or U366 (N_366,N_341,N_197);
xor U367 (N_367,N_276,N_310);
nor U368 (N_368,N_106,N_274);
nor U369 (N_369,N_345,N_280);
nor U370 (N_370,N_18,N_261);
and U371 (N_371,N_279,N_27);
or U372 (N_372,N_72,N_320);
nor U373 (N_373,N_257,N_347);
nand U374 (N_374,N_321,N_71);
nor U375 (N_375,N_205,N_329);
nor U376 (N_376,In_113,N_292);
nand U377 (N_377,N_332,N_314);
nor U378 (N_378,N_112,N_231);
or U379 (N_379,N_12,N_319);
nor U380 (N_380,N_313,N_311);
nand U381 (N_381,In_240,N_324);
nand U382 (N_382,N_337,N_301);
nand U383 (N_383,N_278,N_236);
nor U384 (N_384,N_316,In_136);
or U385 (N_385,N_334,N_277);
nor U386 (N_386,In_330,N_6);
nor U387 (N_387,In_171,N_259);
xor U388 (N_388,N_272,N_338);
nor U389 (N_389,N_342,N_326);
nand U390 (N_390,N_249,N_303);
and U391 (N_391,N_99,N_69);
nand U392 (N_392,In_221,N_291);
nand U393 (N_393,N_158,N_308);
nand U394 (N_394,N_317,N_203);
or U395 (N_395,N_335,N_140);
and U396 (N_396,N_284,N_37);
and U397 (N_397,N_124,N_239);
and U398 (N_398,N_260,N_300);
or U399 (N_399,N_287,N_348);
xor U400 (N_400,N_387,N_360);
or U401 (N_401,N_380,N_381);
and U402 (N_402,In_119,N_399);
nand U403 (N_403,N_206,N_376);
nand U404 (N_404,In_373,N_386);
nand U405 (N_405,N_217,N_256);
or U406 (N_406,N_396,N_240);
nor U407 (N_407,N_391,N_368);
nor U408 (N_408,N_358,N_379);
nand U409 (N_409,N_373,N_393);
nor U410 (N_410,N_383,N_388);
and U411 (N_411,In_37,N_370);
xor U412 (N_412,N_270,N_351);
xor U413 (N_413,N_137,N_395);
or U414 (N_414,N_216,In_461);
nor U415 (N_415,N_165,N_307);
nand U416 (N_416,In_182,N_354);
and U417 (N_417,N_353,N_168);
or U418 (N_418,N_315,N_378);
and U419 (N_419,N_377,N_355);
nor U420 (N_420,N_374,N_322);
and U421 (N_421,N_398,In_249);
nor U422 (N_422,N_362,N_352);
nand U423 (N_423,N_250,N_349);
or U424 (N_424,In_417,N_397);
or U425 (N_425,N_384,N_344);
and U426 (N_426,N_364,In_498);
and U427 (N_427,N_331,N_365);
xor U428 (N_428,N_325,N_382);
and U429 (N_429,N_212,In_303);
nor U430 (N_430,N_363,In_0);
nand U431 (N_431,N_366,N_359);
or U432 (N_432,N_189,N_186);
and U433 (N_433,In_117,N_356);
nor U434 (N_434,In_423,N_346);
and U435 (N_435,N_172,N_372);
nand U436 (N_436,N_339,N_305);
and U437 (N_437,N_367,N_369);
and U438 (N_438,N_262,N_304);
or U439 (N_439,N_309,N_357);
xor U440 (N_440,N_113,N_375);
nand U441 (N_441,N_174,N_385);
nand U442 (N_442,N_266,N_327);
and U443 (N_443,N_8,N_302);
and U444 (N_444,N_390,N_392);
nor U445 (N_445,N_389,N_30);
nand U446 (N_446,N_252,N_121);
or U447 (N_447,N_371,N_394);
or U448 (N_448,N_122,N_350);
nand U449 (N_449,N_361,N_281);
and U450 (N_450,N_421,N_423);
nor U451 (N_451,N_409,N_418);
nand U452 (N_452,N_447,N_442);
nand U453 (N_453,N_416,N_417);
nor U454 (N_454,N_410,N_431);
nand U455 (N_455,N_428,N_430);
nor U456 (N_456,N_405,N_422);
or U457 (N_457,N_426,N_407);
or U458 (N_458,N_425,N_411);
nand U459 (N_459,N_429,N_448);
and U460 (N_460,N_433,N_427);
nor U461 (N_461,N_436,N_400);
xor U462 (N_462,N_414,N_412);
and U463 (N_463,N_434,N_413);
and U464 (N_464,N_435,N_408);
or U465 (N_465,N_419,N_438);
and U466 (N_466,N_439,N_424);
or U467 (N_467,N_432,N_420);
or U468 (N_468,N_446,N_445);
nor U469 (N_469,N_401,N_415);
nand U470 (N_470,N_404,N_443);
nand U471 (N_471,N_406,N_441);
and U472 (N_472,N_437,N_402);
nor U473 (N_473,N_449,N_403);
and U474 (N_474,N_440,N_444);
or U475 (N_475,N_400,N_403);
xnor U476 (N_476,N_406,N_429);
nand U477 (N_477,N_420,N_426);
xor U478 (N_478,N_417,N_430);
and U479 (N_479,N_432,N_425);
nor U480 (N_480,N_414,N_403);
nor U481 (N_481,N_417,N_448);
and U482 (N_482,N_408,N_449);
nor U483 (N_483,N_446,N_449);
and U484 (N_484,N_417,N_435);
nand U485 (N_485,N_421,N_416);
nor U486 (N_486,N_436,N_406);
or U487 (N_487,N_423,N_407);
and U488 (N_488,N_404,N_418);
nor U489 (N_489,N_416,N_437);
or U490 (N_490,N_446,N_413);
nand U491 (N_491,N_441,N_435);
or U492 (N_492,N_423,N_419);
nor U493 (N_493,N_427,N_418);
nor U494 (N_494,N_428,N_425);
and U495 (N_495,N_440,N_435);
and U496 (N_496,N_432,N_409);
nand U497 (N_497,N_416,N_433);
and U498 (N_498,N_403,N_431);
nor U499 (N_499,N_408,N_432);
nand U500 (N_500,N_477,N_479);
nand U501 (N_501,N_474,N_457);
nand U502 (N_502,N_464,N_489);
and U503 (N_503,N_460,N_491);
nor U504 (N_504,N_485,N_492);
nand U505 (N_505,N_450,N_454);
nand U506 (N_506,N_470,N_467);
xor U507 (N_507,N_478,N_497);
or U508 (N_508,N_486,N_496);
nor U509 (N_509,N_475,N_461);
xor U510 (N_510,N_452,N_480);
and U511 (N_511,N_487,N_456);
nand U512 (N_512,N_459,N_488);
and U513 (N_513,N_494,N_472);
xor U514 (N_514,N_455,N_484);
xnor U515 (N_515,N_471,N_476);
or U516 (N_516,N_495,N_481);
or U517 (N_517,N_466,N_499);
nand U518 (N_518,N_453,N_482);
nand U519 (N_519,N_451,N_465);
or U520 (N_520,N_463,N_468);
nand U521 (N_521,N_462,N_469);
nand U522 (N_522,N_483,N_458);
nand U523 (N_523,N_473,N_493);
or U524 (N_524,N_498,N_490);
nand U525 (N_525,N_464,N_470);
nor U526 (N_526,N_485,N_461);
nand U527 (N_527,N_492,N_481);
nor U528 (N_528,N_478,N_466);
and U529 (N_529,N_495,N_467);
xor U530 (N_530,N_477,N_468);
or U531 (N_531,N_466,N_476);
nand U532 (N_532,N_451,N_487);
and U533 (N_533,N_497,N_477);
xnor U534 (N_534,N_478,N_461);
or U535 (N_535,N_493,N_458);
and U536 (N_536,N_465,N_485);
and U537 (N_537,N_459,N_495);
nand U538 (N_538,N_493,N_479);
nand U539 (N_539,N_474,N_486);
nand U540 (N_540,N_480,N_478);
or U541 (N_541,N_457,N_478);
nand U542 (N_542,N_499,N_464);
or U543 (N_543,N_479,N_460);
nand U544 (N_544,N_494,N_454);
or U545 (N_545,N_454,N_493);
and U546 (N_546,N_483,N_487);
nand U547 (N_547,N_467,N_491);
nor U548 (N_548,N_490,N_454);
or U549 (N_549,N_456,N_497);
xor U550 (N_550,N_516,N_538);
and U551 (N_551,N_505,N_523);
xnor U552 (N_552,N_527,N_515);
nor U553 (N_553,N_525,N_506);
nor U554 (N_554,N_536,N_510);
nand U555 (N_555,N_521,N_535);
and U556 (N_556,N_501,N_504);
or U557 (N_557,N_503,N_511);
and U558 (N_558,N_537,N_541);
or U559 (N_559,N_509,N_528);
nor U560 (N_560,N_540,N_546);
nor U561 (N_561,N_500,N_531);
or U562 (N_562,N_539,N_534);
or U563 (N_563,N_533,N_507);
nor U564 (N_564,N_513,N_514);
nor U565 (N_565,N_502,N_547);
or U566 (N_566,N_532,N_549);
nor U567 (N_567,N_530,N_543);
and U568 (N_568,N_512,N_520);
xnor U569 (N_569,N_548,N_522);
nand U570 (N_570,N_524,N_545);
and U571 (N_571,N_518,N_529);
nand U572 (N_572,N_519,N_517);
or U573 (N_573,N_544,N_542);
xor U574 (N_574,N_526,N_508);
and U575 (N_575,N_505,N_542);
and U576 (N_576,N_542,N_548);
nor U577 (N_577,N_530,N_503);
nand U578 (N_578,N_544,N_516);
or U579 (N_579,N_520,N_534);
nand U580 (N_580,N_525,N_507);
nand U581 (N_581,N_535,N_513);
nand U582 (N_582,N_522,N_536);
nor U583 (N_583,N_514,N_509);
or U584 (N_584,N_535,N_540);
nand U585 (N_585,N_519,N_520);
and U586 (N_586,N_529,N_520);
nand U587 (N_587,N_536,N_516);
or U588 (N_588,N_525,N_520);
and U589 (N_589,N_515,N_541);
nor U590 (N_590,N_536,N_540);
nor U591 (N_591,N_519,N_536);
or U592 (N_592,N_513,N_504);
nand U593 (N_593,N_533,N_535);
nand U594 (N_594,N_549,N_526);
and U595 (N_595,N_514,N_549);
and U596 (N_596,N_511,N_505);
or U597 (N_597,N_522,N_533);
and U598 (N_598,N_515,N_526);
xor U599 (N_599,N_519,N_510);
and U600 (N_600,N_553,N_560);
and U601 (N_601,N_552,N_584);
nand U602 (N_602,N_573,N_555);
and U603 (N_603,N_585,N_579);
or U604 (N_604,N_589,N_568);
nand U605 (N_605,N_598,N_566);
and U606 (N_606,N_551,N_561);
and U607 (N_607,N_580,N_587);
nand U608 (N_608,N_586,N_558);
or U609 (N_609,N_570,N_583);
nand U610 (N_610,N_588,N_571);
or U611 (N_611,N_593,N_563);
nand U612 (N_612,N_595,N_564);
nor U613 (N_613,N_574,N_576);
or U614 (N_614,N_594,N_550);
or U615 (N_615,N_569,N_578);
nand U616 (N_616,N_591,N_554);
or U617 (N_617,N_581,N_575);
or U618 (N_618,N_556,N_597);
and U619 (N_619,N_567,N_577);
nor U620 (N_620,N_557,N_582);
xor U621 (N_621,N_559,N_596);
and U622 (N_622,N_599,N_590);
or U623 (N_623,N_592,N_562);
nand U624 (N_624,N_565,N_572);
nand U625 (N_625,N_554,N_557);
nor U626 (N_626,N_567,N_584);
and U627 (N_627,N_560,N_585);
nand U628 (N_628,N_591,N_596);
nor U629 (N_629,N_571,N_564);
or U630 (N_630,N_584,N_568);
or U631 (N_631,N_555,N_598);
and U632 (N_632,N_550,N_591);
or U633 (N_633,N_585,N_557);
nand U634 (N_634,N_579,N_599);
nor U635 (N_635,N_560,N_561);
or U636 (N_636,N_557,N_574);
and U637 (N_637,N_572,N_585);
nand U638 (N_638,N_575,N_558);
and U639 (N_639,N_596,N_553);
nor U640 (N_640,N_589,N_587);
nand U641 (N_641,N_590,N_580);
nand U642 (N_642,N_569,N_562);
and U643 (N_643,N_591,N_557);
and U644 (N_644,N_563,N_570);
and U645 (N_645,N_593,N_598);
nor U646 (N_646,N_590,N_579);
or U647 (N_647,N_552,N_564);
nand U648 (N_648,N_583,N_574);
nor U649 (N_649,N_580,N_567);
nor U650 (N_650,N_637,N_619);
xor U651 (N_651,N_645,N_638);
nor U652 (N_652,N_620,N_602);
or U653 (N_653,N_610,N_631);
or U654 (N_654,N_604,N_624);
or U655 (N_655,N_630,N_625);
xor U656 (N_656,N_641,N_613);
and U657 (N_657,N_614,N_635);
or U658 (N_658,N_615,N_603);
or U659 (N_659,N_642,N_647);
and U660 (N_660,N_616,N_646);
or U661 (N_661,N_639,N_628);
nand U662 (N_662,N_626,N_612);
or U663 (N_663,N_621,N_618);
nand U664 (N_664,N_640,N_648);
nor U665 (N_665,N_636,N_622);
or U666 (N_666,N_623,N_644);
nand U667 (N_667,N_643,N_605);
nand U668 (N_668,N_632,N_629);
nand U669 (N_669,N_608,N_600);
nor U670 (N_670,N_627,N_607);
or U671 (N_671,N_649,N_634);
nand U672 (N_672,N_633,N_617);
or U673 (N_673,N_601,N_611);
nor U674 (N_674,N_606,N_609);
nor U675 (N_675,N_614,N_608);
nor U676 (N_676,N_645,N_620);
nor U677 (N_677,N_606,N_617);
nor U678 (N_678,N_609,N_601);
nand U679 (N_679,N_649,N_612);
xnor U680 (N_680,N_610,N_604);
nand U681 (N_681,N_624,N_647);
nor U682 (N_682,N_647,N_601);
nor U683 (N_683,N_624,N_600);
or U684 (N_684,N_608,N_623);
and U685 (N_685,N_606,N_614);
or U686 (N_686,N_626,N_606);
and U687 (N_687,N_615,N_613);
or U688 (N_688,N_646,N_628);
or U689 (N_689,N_614,N_602);
nor U690 (N_690,N_603,N_610);
nand U691 (N_691,N_616,N_621);
and U692 (N_692,N_621,N_625);
and U693 (N_693,N_634,N_608);
or U694 (N_694,N_622,N_630);
nor U695 (N_695,N_605,N_612);
nand U696 (N_696,N_644,N_632);
and U697 (N_697,N_610,N_614);
and U698 (N_698,N_620,N_638);
nand U699 (N_699,N_618,N_633);
and U700 (N_700,N_662,N_664);
nor U701 (N_701,N_691,N_696);
or U702 (N_702,N_698,N_659);
or U703 (N_703,N_681,N_655);
xnor U704 (N_704,N_690,N_692);
and U705 (N_705,N_667,N_653);
nor U706 (N_706,N_685,N_678);
nand U707 (N_707,N_680,N_657);
nand U708 (N_708,N_666,N_693);
nor U709 (N_709,N_670,N_668);
nand U710 (N_710,N_674,N_697);
and U711 (N_711,N_689,N_695);
nand U712 (N_712,N_658,N_660);
or U713 (N_713,N_677,N_651);
or U714 (N_714,N_652,N_672);
nor U715 (N_715,N_679,N_686);
nor U716 (N_716,N_665,N_663);
or U717 (N_717,N_675,N_656);
and U718 (N_718,N_661,N_682);
nor U719 (N_719,N_673,N_654);
and U720 (N_720,N_687,N_669);
or U721 (N_721,N_671,N_688);
nor U722 (N_722,N_694,N_650);
nor U723 (N_723,N_683,N_676);
or U724 (N_724,N_684,N_699);
or U725 (N_725,N_677,N_662);
and U726 (N_726,N_657,N_671);
nand U727 (N_727,N_677,N_663);
and U728 (N_728,N_661,N_656);
nor U729 (N_729,N_664,N_695);
nand U730 (N_730,N_657,N_686);
and U731 (N_731,N_664,N_678);
nor U732 (N_732,N_681,N_667);
xnor U733 (N_733,N_691,N_662);
nor U734 (N_734,N_660,N_657);
and U735 (N_735,N_688,N_678);
and U736 (N_736,N_668,N_654);
nand U737 (N_737,N_655,N_691);
and U738 (N_738,N_680,N_686);
or U739 (N_739,N_669,N_665);
nand U740 (N_740,N_653,N_665);
and U741 (N_741,N_674,N_673);
and U742 (N_742,N_683,N_668);
nor U743 (N_743,N_675,N_679);
nand U744 (N_744,N_686,N_685);
nor U745 (N_745,N_674,N_693);
nand U746 (N_746,N_684,N_667);
or U747 (N_747,N_654,N_663);
and U748 (N_748,N_663,N_683);
nor U749 (N_749,N_681,N_672);
xnor U750 (N_750,N_734,N_728);
and U751 (N_751,N_736,N_725);
nor U752 (N_752,N_703,N_700);
nand U753 (N_753,N_748,N_733);
nand U754 (N_754,N_701,N_735);
xnor U755 (N_755,N_715,N_737);
nor U756 (N_756,N_711,N_708);
nand U757 (N_757,N_732,N_706);
xnor U758 (N_758,N_740,N_718);
or U759 (N_759,N_719,N_720);
nor U760 (N_760,N_709,N_713);
or U761 (N_761,N_705,N_746);
and U762 (N_762,N_726,N_710);
or U763 (N_763,N_747,N_738);
nor U764 (N_764,N_739,N_742);
xor U765 (N_765,N_743,N_727);
xnor U766 (N_766,N_744,N_712);
nor U767 (N_767,N_722,N_730);
nand U768 (N_768,N_716,N_731);
or U769 (N_769,N_745,N_741);
and U770 (N_770,N_702,N_704);
nor U771 (N_771,N_721,N_707);
or U772 (N_772,N_749,N_717);
and U773 (N_773,N_723,N_724);
and U774 (N_774,N_714,N_729);
nor U775 (N_775,N_717,N_733);
nor U776 (N_776,N_705,N_736);
nor U777 (N_777,N_713,N_708);
nand U778 (N_778,N_704,N_742);
and U779 (N_779,N_708,N_740);
and U780 (N_780,N_732,N_714);
nor U781 (N_781,N_732,N_715);
nand U782 (N_782,N_700,N_736);
nand U783 (N_783,N_709,N_727);
or U784 (N_784,N_718,N_741);
nand U785 (N_785,N_730,N_744);
nor U786 (N_786,N_734,N_727);
nand U787 (N_787,N_714,N_712);
and U788 (N_788,N_742,N_724);
and U789 (N_789,N_723,N_746);
nor U790 (N_790,N_716,N_718);
nand U791 (N_791,N_731,N_704);
or U792 (N_792,N_728,N_730);
xnor U793 (N_793,N_719,N_730);
and U794 (N_794,N_736,N_714);
or U795 (N_795,N_723,N_704);
nand U796 (N_796,N_743,N_709);
and U797 (N_797,N_731,N_746);
or U798 (N_798,N_706,N_700);
or U799 (N_799,N_730,N_716);
or U800 (N_800,N_762,N_753);
xor U801 (N_801,N_752,N_760);
and U802 (N_802,N_792,N_790);
or U803 (N_803,N_769,N_776);
and U804 (N_804,N_751,N_756);
or U805 (N_805,N_785,N_770);
nor U806 (N_806,N_767,N_777);
nor U807 (N_807,N_755,N_791);
nand U808 (N_808,N_759,N_750);
and U809 (N_809,N_781,N_789);
and U810 (N_810,N_793,N_764);
and U811 (N_811,N_754,N_780);
and U812 (N_812,N_787,N_779);
nand U813 (N_813,N_772,N_797);
or U814 (N_814,N_788,N_796);
nor U815 (N_815,N_778,N_765);
nand U816 (N_816,N_795,N_766);
nand U817 (N_817,N_798,N_774);
nor U818 (N_818,N_782,N_763);
and U819 (N_819,N_773,N_786);
nand U820 (N_820,N_758,N_768);
nor U821 (N_821,N_794,N_761);
and U822 (N_822,N_799,N_783);
and U823 (N_823,N_775,N_771);
nand U824 (N_824,N_784,N_757);
nor U825 (N_825,N_792,N_779);
xor U826 (N_826,N_777,N_781);
nor U827 (N_827,N_776,N_761);
nor U828 (N_828,N_796,N_768);
nor U829 (N_829,N_788,N_784);
or U830 (N_830,N_759,N_778);
and U831 (N_831,N_792,N_793);
or U832 (N_832,N_766,N_788);
or U833 (N_833,N_784,N_762);
nand U834 (N_834,N_781,N_784);
nor U835 (N_835,N_784,N_756);
and U836 (N_836,N_757,N_771);
xor U837 (N_837,N_751,N_754);
nor U838 (N_838,N_793,N_761);
and U839 (N_839,N_780,N_785);
or U840 (N_840,N_760,N_773);
nor U841 (N_841,N_763,N_751);
and U842 (N_842,N_795,N_764);
nand U843 (N_843,N_750,N_774);
and U844 (N_844,N_774,N_785);
nand U845 (N_845,N_775,N_787);
nand U846 (N_846,N_779,N_782);
or U847 (N_847,N_750,N_754);
nor U848 (N_848,N_793,N_769);
xnor U849 (N_849,N_789,N_768);
nor U850 (N_850,N_812,N_815);
or U851 (N_851,N_804,N_811);
nor U852 (N_852,N_813,N_820);
nand U853 (N_853,N_840,N_816);
or U854 (N_854,N_848,N_833);
or U855 (N_855,N_822,N_827);
nand U856 (N_856,N_818,N_817);
nor U857 (N_857,N_837,N_802);
nand U858 (N_858,N_823,N_801);
xnor U859 (N_859,N_825,N_829);
or U860 (N_860,N_835,N_842);
nor U861 (N_861,N_843,N_805);
xnor U862 (N_862,N_824,N_830);
xor U863 (N_863,N_806,N_826);
xor U864 (N_864,N_845,N_807);
nor U865 (N_865,N_832,N_838);
nor U866 (N_866,N_814,N_836);
or U867 (N_867,N_844,N_819);
or U868 (N_868,N_841,N_839);
nor U869 (N_869,N_803,N_821);
nand U870 (N_870,N_800,N_831);
and U871 (N_871,N_847,N_849);
nor U872 (N_872,N_846,N_808);
and U873 (N_873,N_809,N_828);
or U874 (N_874,N_810,N_834);
nand U875 (N_875,N_812,N_825);
or U876 (N_876,N_833,N_814);
or U877 (N_877,N_849,N_806);
nor U878 (N_878,N_838,N_828);
xnor U879 (N_879,N_849,N_835);
nor U880 (N_880,N_830,N_811);
and U881 (N_881,N_825,N_802);
nand U882 (N_882,N_829,N_846);
and U883 (N_883,N_844,N_833);
nor U884 (N_884,N_821,N_841);
and U885 (N_885,N_815,N_825);
xnor U886 (N_886,N_824,N_801);
or U887 (N_887,N_838,N_845);
or U888 (N_888,N_805,N_808);
nand U889 (N_889,N_839,N_815);
or U890 (N_890,N_814,N_838);
nand U891 (N_891,N_849,N_813);
nor U892 (N_892,N_813,N_830);
nand U893 (N_893,N_840,N_803);
and U894 (N_894,N_816,N_807);
nor U895 (N_895,N_832,N_822);
nand U896 (N_896,N_837,N_801);
and U897 (N_897,N_820,N_804);
xor U898 (N_898,N_812,N_818);
and U899 (N_899,N_816,N_822);
or U900 (N_900,N_875,N_893);
or U901 (N_901,N_894,N_862);
or U902 (N_902,N_876,N_858);
nor U903 (N_903,N_860,N_867);
nor U904 (N_904,N_872,N_854);
nand U905 (N_905,N_882,N_852);
and U906 (N_906,N_889,N_866);
nand U907 (N_907,N_863,N_856);
nor U908 (N_908,N_884,N_892);
nor U909 (N_909,N_871,N_898);
xnor U910 (N_910,N_899,N_879);
and U911 (N_911,N_896,N_873);
and U912 (N_912,N_853,N_865);
nand U913 (N_913,N_861,N_891);
xor U914 (N_914,N_859,N_888);
nor U915 (N_915,N_890,N_878);
or U916 (N_916,N_886,N_877);
and U917 (N_917,N_851,N_880);
and U918 (N_918,N_864,N_869);
nand U919 (N_919,N_887,N_870);
nor U920 (N_920,N_874,N_855);
and U921 (N_921,N_857,N_881);
or U922 (N_922,N_897,N_895);
nor U923 (N_923,N_850,N_868);
nor U924 (N_924,N_885,N_883);
nand U925 (N_925,N_890,N_881);
or U926 (N_926,N_894,N_876);
or U927 (N_927,N_879,N_880);
or U928 (N_928,N_867,N_850);
nand U929 (N_929,N_875,N_876);
nand U930 (N_930,N_898,N_882);
or U931 (N_931,N_899,N_896);
nor U932 (N_932,N_891,N_872);
or U933 (N_933,N_871,N_884);
or U934 (N_934,N_854,N_856);
nand U935 (N_935,N_859,N_865);
nor U936 (N_936,N_861,N_872);
xnor U937 (N_937,N_878,N_881);
and U938 (N_938,N_864,N_873);
nand U939 (N_939,N_895,N_867);
xor U940 (N_940,N_871,N_851);
or U941 (N_941,N_877,N_880);
and U942 (N_942,N_890,N_887);
nand U943 (N_943,N_852,N_875);
nor U944 (N_944,N_859,N_868);
nand U945 (N_945,N_853,N_864);
nor U946 (N_946,N_894,N_857);
or U947 (N_947,N_872,N_874);
or U948 (N_948,N_853,N_880);
xor U949 (N_949,N_890,N_882);
or U950 (N_950,N_942,N_931);
nand U951 (N_951,N_948,N_927);
and U952 (N_952,N_923,N_947);
nand U953 (N_953,N_929,N_903);
or U954 (N_954,N_907,N_904);
or U955 (N_955,N_944,N_928);
nor U956 (N_956,N_938,N_943);
nor U957 (N_957,N_941,N_925);
or U958 (N_958,N_946,N_913);
nor U959 (N_959,N_912,N_930);
and U960 (N_960,N_902,N_924);
or U961 (N_961,N_920,N_926);
and U962 (N_962,N_901,N_940);
nand U963 (N_963,N_934,N_905);
nor U964 (N_964,N_922,N_911);
nor U965 (N_965,N_932,N_921);
nor U966 (N_966,N_945,N_939);
nand U967 (N_967,N_919,N_935);
nand U968 (N_968,N_936,N_915);
and U969 (N_969,N_917,N_914);
nor U970 (N_970,N_908,N_906);
nand U971 (N_971,N_916,N_949);
and U972 (N_972,N_909,N_918);
nand U973 (N_973,N_910,N_900);
and U974 (N_974,N_933,N_937);
nand U975 (N_975,N_938,N_924);
or U976 (N_976,N_948,N_946);
or U977 (N_977,N_907,N_926);
or U978 (N_978,N_939,N_900);
nor U979 (N_979,N_923,N_915);
or U980 (N_980,N_923,N_906);
nor U981 (N_981,N_937,N_906);
nand U982 (N_982,N_940,N_904);
or U983 (N_983,N_925,N_928);
nor U984 (N_984,N_948,N_914);
and U985 (N_985,N_915,N_944);
or U986 (N_986,N_931,N_909);
xnor U987 (N_987,N_917,N_934);
or U988 (N_988,N_906,N_901);
or U989 (N_989,N_910,N_938);
nor U990 (N_990,N_917,N_933);
nor U991 (N_991,N_906,N_925);
nand U992 (N_992,N_939,N_912);
nor U993 (N_993,N_922,N_901);
or U994 (N_994,N_933,N_945);
nand U995 (N_995,N_943,N_902);
and U996 (N_996,N_905,N_900);
nor U997 (N_997,N_942,N_915);
and U998 (N_998,N_909,N_942);
or U999 (N_999,N_917,N_949);
nand U1000 (N_1000,N_989,N_974);
nand U1001 (N_1001,N_982,N_970);
and U1002 (N_1002,N_986,N_973);
and U1003 (N_1003,N_964,N_976);
and U1004 (N_1004,N_953,N_967);
nand U1005 (N_1005,N_968,N_971);
nand U1006 (N_1006,N_951,N_979);
or U1007 (N_1007,N_981,N_999);
nand U1008 (N_1008,N_980,N_983);
or U1009 (N_1009,N_992,N_963);
nor U1010 (N_1010,N_965,N_952);
or U1011 (N_1011,N_997,N_960);
and U1012 (N_1012,N_985,N_996);
and U1013 (N_1013,N_984,N_969);
nand U1014 (N_1014,N_962,N_957);
nor U1015 (N_1015,N_958,N_995);
nand U1016 (N_1016,N_950,N_987);
and U1017 (N_1017,N_998,N_975);
nand U1018 (N_1018,N_977,N_994);
xor U1019 (N_1019,N_955,N_993);
and U1020 (N_1020,N_959,N_978);
nor U1021 (N_1021,N_956,N_961);
xor U1022 (N_1022,N_954,N_988);
nor U1023 (N_1023,N_990,N_966);
nor U1024 (N_1024,N_991,N_972);
nor U1025 (N_1025,N_990,N_991);
xnor U1026 (N_1026,N_959,N_972);
nand U1027 (N_1027,N_954,N_976);
xor U1028 (N_1028,N_952,N_975);
nand U1029 (N_1029,N_968,N_953);
xor U1030 (N_1030,N_982,N_992);
nor U1031 (N_1031,N_984,N_981);
and U1032 (N_1032,N_978,N_990);
or U1033 (N_1033,N_991,N_957);
and U1034 (N_1034,N_981,N_954);
nor U1035 (N_1035,N_965,N_998);
xor U1036 (N_1036,N_964,N_970);
nor U1037 (N_1037,N_992,N_995);
nand U1038 (N_1038,N_973,N_972);
nor U1039 (N_1039,N_993,N_976);
and U1040 (N_1040,N_951,N_997);
nor U1041 (N_1041,N_958,N_989);
and U1042 (N_1042,N_997,N_986);
or U1043 (N_1043,N_985,N_965);
nand U1044 (N_1044,N_956,N_996);
or U1045 (N_1045,N_992,N_985);
or U1046 (N_1046,N_962,N_976);
and U1047 (N_1047,N_951,N_999);
nand U1048 (N_1048,N_964,N_983);
xor U1049 (N_1049,N_967,N_969);
and U1050 (N_1050,N_1047,N_1019);
or U1051 (N_1051,N_1042,N_1005);
nand U1052 (N_1052,N_1046,N_1022);
or U1053 (N_1053,N_1012,N_1027);
and U1054 (N_1054,N_1006,N_1034);
nor U1055 (N_1055,N_1020,N_1040);
nor U1056 (N_1056,N_1045,N_1037);
nor U1057 (N_1057,N_1018,N_1010);
or U1058 (N_1058,N_1031,N_1025);
and U1059 (N_1059,N_1032,N_1028);
nor U1060 (N_1060,N_1039,N_1013);
or U1061 (N_1061,N_1035,N_1002);
or U1062 (N_1062,N_1041,N_1003);
nor U1063 (N_1063,N_1004,N_1008);
nor U1064 (N_1064,N_1043,N_1009);
nor U1065 (N_1065,N_1023,N_1007);
nor U1066 (N_1066,N_1036,N_1029);
or U1067 (N_1067,N_1021,N_1001);
nor U1068 (N_1068,N_1015,N_1049);
nor U1069 (N_1069,N_1024,N_1014);
and U1070 (N_1070,N_1016,N_1038);
or U1071 (N_1071,N_1033,N_1011);
and U1072 (N_1072,N_1030,N_1017);
nand U1073 (N_1073,N_1044,N_1026);
and U1074 (N_1074,N_1000,N_1048);
nor U1075 (N_1075,N_1021,N_1013);
and U1076 (N_1076,N_1035,N_1001);
nand U1077 (N_1077,N_1039,N_1016);
nand U1078 (N_1078,N_1035,N_1047);
nand U1079 (N_1079,N_1048,N_1037);
nor U1080 (N_1080,N_1042,N_1024);
and U1081 (N_1081,N_1010,N_1023);
or U1082 (N_1082,N_1040,N_1031);
xor U1083 (N_1083,N_1021,N_1009);
or U1084 (N_1084,N_1036,N_1005);
or U1085 (N_1085,N_1043,N_1024);
or U1086 (N_1086,N_1040,N_1003);
and U1087 (N_1087,N_1006,N_1017);
nand U1088 (N_1088,N_1012,N_1007);
nand U1089 (N_1089,N_1013,N_1049);
nor U1090 (N_1090,N_1014,N_1020);
nor U1091 (N_1091,N_1007,N_1044);
and U1092 (N_1092,N_1002,N_1014);
nor U1093 (N_1093,N_1003,N_1034);
nand U1094 (N_1094,N_1032,N_1009);
nand U1095 (N_1095,N_1020,N_1043);
nand U1096 (N_1096,N_1049,N_1035);
nor U1097 (N_1097,N_1045,N_1012);
nand U1098 (N_1098,N_1048,N_1031);
or U1099 (N_1099,N_1019,N_1045);
or U1100 (N_1100,N_1056,N_1070);
nor U1101 (N_1101,N_1059,N_1073);
xor U1102 (N_1102,N_1060,N_1051);
nand U1103 (N_1103,N_1058,N_1063);
nor U1104 (N_1104,N_1072,N_1062);
and U1105 (N_1105,N_1087,N_1089);
and U1106 (N_1106,N_1068,N_1077);
nor U1107 (N_1107,N_1071,N_1094);
and U1108 (N_1108,N_1092,N_1095);
and U1109 (N_1109,N_1076,N_1078);
nand U1110 (N_1110,N_1088,N_1064);
nor U1111 (N_1111,N_1090,N_1052);
or U1112 (N_1112,N_1054,N_1086);
and U1113 (N_1113,N_1075,N_1053);
nor U1114 (N_1114,N_1067,N_1066);
or U1115 (N_1115,N_1057,N_1050);
and U1116 (N_1116,N_1085,N_1074);
or U1117 (N_1117,N_1097,N_1081);
or U1118 (N_1118,N_1069,N_1093);
xor U1119 (N_1119,N_1061,N_1096);
nand U1120 (N_1120,N_1079,N_1080);
and U1121 (N_1121,N_1065,N_1083);
nand U1122 (N_1122,N_1084,N_1055);
and U1123 (N_1123,N_1091,N_1099);
or U1124 (N_1124,N_1098,N_1082);
nor U1125 (N_1125,N_1052,N_1063);
and U1126 (N_1126,N_1078,N_1074);
and U1127 (N_1127,N_1056,N_1087);
nand U1128 (N_1128,N_1068,N_1081);
nor U1129 (N_1129,N_1089,N_1096);
or U1130 (N_1130,N_1065,N_1051);
and U1131 (N_1131,N_1087,N_1098);
and U1132 (N_1132,N_1058,N_1096);
nor U1133 (N_1133,N_1062,N_1052);
or U1134 (N_1134,N_1093,N_1094);
nor U1135 (N_1135,N_1085,N_1083);
nand U1136 (N_1136,N_1055,N_1054);
or U1137 (N_1137,N_1096,N_1084);
nor U1138 (N_1138,N_1098,N_1065);
and U1139 (N_1139,N_1082,N_1066);
or U1140 (N_1140,N_1060,N_1078);
or U1141 (N_1141,N_1091,N_1084);
nor U1142 (N_1142,N_1077,N_1098);
xor U1143 (N_1143,N_1084,N_1089);
or U1144 (N_1144,N_1057,N_1093);
or U1145 (N_1145,N_1071,N_1078);
or U1146 (N_1146,N_1053,N_1098);
nand U1147 (N_1147,N_1070,N_1058);
nand U1148 (N_1148,N_1080,N_1075);
and U1149 (N_1149,N_1094,N_1063);
and U1150 (N_1150,N_1117,N_1149);
and U1151 (N_1151,N_1140,N_1111);
nor U1152 (N_1152,N_1120,N_1105);
and U1153 (N_1153,N_1138,N_1100);
nor U1154 (N_1154,N_1146,N_1125);
or U1155 (N_1155,N_1119,N_1127);
nor U1156 (N_1156,N_1137,N_1110);
xor U1157 (N_1157,N_1133,N_1107);
nand U1158 (N_1158,N_1102,N_1113);
or U1159 (N_1159,N_1101,N_1128);
nor U1160 (N_1160,N_1136,N_1148);
nor U1161 (N_1161,N_1106,N_1122);
and U1162 (N_1162,N_1124,N_1114);
nand U1163 (N_1163,N_1143,N_1131);
xnor U1164 (N_1164,N_1129,N_1121);
or U1165 (N_1165,N_1141,N_1130);
and U1166 (N_1166,N_1103,N_1135);
and U1167 (N_1167,N_1145,N_1144);
nand U1168 (N_1168,N_1126,N_1109);
or U1169 (N_1169,N_1118,N_1132);
nor U1170 (N_1170,N_1112,N_1123);
nor U1171 (N_1171,N_1108,N_1142);
nand U1172 (N_1172,N_1139,N_1116);
or U1173 (N_1173,N_1115,N_1104);
and U1174 (N_1174,N_1147,N_1134);
nand U1175 (N_1175,N_1141,N_1143);
xnor U1176 (N_1176,N_1108,N_1141);
and U1177 (N_1177,N_1110,N_1109);
or U1178 (N_1178,N_1141,N_1134);
or U1179 (N_1179,N_1149,N_1133);
nand U1180 (N_1180,N_1134,N_1112);
or U1181 (N_1181,N_1103,N_1140);
nand U1182 (N_1182,N_1129,N_1112);
or U1183 (N_1183,N_1138,N_1122);
nand U1184 (N_1184,N_1104,N_1123);
nor U1185 (N_1185,N_1119,N_1120);
nor U1186 (N_1186,N_1117,N_1106);
nand U1187 (N_1187,N_1146,N_1129);
nand U1188 (N_1188,N_1132,N_1110);
and U1189 (N_1189,N_1120,N_1141);
and U1190 (N_1190,N_1105,N_1141);
or U1191 (N_1191,N_1132,N_1131);
nor U1192 (N_1192,N_1115,N_1123);
nor U1193 (N_1193,N_1118,N_1129);
or U1194 (N_1194,N_1118,N_1122);
or U1195 (N_1195,N_1117,N_1136);
nand U1196 (N_1196,N_1145,N_1107);
or U1197 (N_1197,N_1134,N_1108);
nand U1198 (N_1198,N_1100,N_1109);
xor U1199 (N_1199,N_1148,N_1102);
nor U1200 (N_1200,N_1195,N_1177);
and U1201 (N_1201,N_1151,N_1161);
and U1202 (N_1202,N_1196,N_1156);
and U1203 (N_1203,N_1194,N_1160);
or U1204 (N_1204,N_1184,N_1178);
or U1205 (N_1205,N_1166,N_1163);
and U1206 (N_1206,N_1183,N_1192);
and U1207 (N_1207,N_1182,N_1159);
and U1208 (N_1208,N_1165,N_1172);
nor U1209 (N_1209,N_1181,N_1197);
nor U1210 (N_1210,N_1168,N_1162);
or U1211 (N_1211,N_1153,N_1170);
nor U1212 (N_1212,N_1175,N_1169);
nand U1213 (N_1213,N_1167,N_1164);
nor U1214 (N_1214,N_1188,N_1193);
or U1215 (N_1215,N_1173,N_1186);
and U1216 (N_1216,N_1191,N_1199);
nand U1217 (N_1217,N_1180,N_1179);
or U1218 (N_1218,N_1185,N_1155);
xor U1219 (N_1219,N_1171,N_1157);
xor U1220 (N_1220,N_1189,N_1190);
and U1221 (N_1221,N_1154,N_1150);
or U1222 (N_1222,N_1187,N_1152);
xor U1223 (N_1223,N_1174,N_1176);
or U1224 (N_1224,N_1198,N_1158);
nand U1225 (N_1225,N_1167,N_1163);
nor U1226 (N_1226,N_1181,N_1166);
nand U1227 (N_1227,N_1159,N_1176);
and U1228 (N_1228,N_1188,N_1186);
nand U1229 (N_1229,N_1167,N_1150);
or U1230 (N_1230,N_1170,N_1182);
nor U1231 (N_1231,N_1192,N_1152);
or U1232 (N_1232,N_1183,N_1157);
nor U1233 (N_1233,N_1172,N_1191);
nor U1234 (N_1234,N_1194,N_1154);
nor U1235 (N_1235,N_1165,N_1193);
nor U1236 (N_1236,N_1175,N_1181);
nand U1237 (N_1237,N_1157,N_1150);
nor U1238 (N_1238,N_1173,N_1172);
xor U1239 (N_1239,N_1171,N_1160);
and U1240 (N_1240,N_1168,N_1155);
or U1241 (N_1241,N_1189,N_1199);
or U1242 (N_1242,N_1151,N_1189);
and U1243 (N_1243,N_1167,N_1174);
and U1244 (N_1244,N_1176,N_1163);
nand U1245 (N_1245,N_1161,N_1195);
or U1246 (N_1246,N_1196,N_1194);
or U1247 (N_1247,N_1180,N_1165);
nand U1248 (N_1248,N_1194,N_1197);
or U1249 (N_1249,N_1187,N_1181);
and U1250 (N_1250,N_1204,N_1206);
nor U1251 (N_1251,N_1207,N_1249);
or U1252 (N_1252,N_1224,N_1246);
nand U1253 (N_1253,N_1210,N_1247);
nor U1254 (N_1254,N_1211,N_1244);
nor U1255 (N_1255,N_1245,N_1235);
or U1256 (N_1256,N_1232,N_1201);
or U1257 (N_1257,N_1203,N_1200);
nand U1258 (N_1258,N_1225,N_1236);
and U1259 (N_1259,N_1222,N_1228);
and U1260 (N_1260,N_1234,N_1216);
nand U1261 (N_1261,N_1214,N_1227);
or U1262 (N_1262,N_1248,N_1229);
nand U1263 (N_1263,N_1217,N_1213);
nand U1264 (N_1264,N_1243,N_1215);
nor U1265 (N_1265,N_1239,N_1220);
nor U1266 (N_1266,N_1231,N_1219);
nand U1267 (N_1267,N_1223,N_1221);
nor U1268 (N_1268,N_1208,N_1230);
nor U1269 (N_1269,N_1209,N_1233);
and U1270 (N_1270,N_1205,N_1241);
or U1271 (N_1271,N_1242,N_1226);
nand U1272 (N_1272,N_1240,N_1218);
nor U1273 (N_1273,N_1202,N_1238);
nand U1274 (N_1274,N_1212,N_1237);
nor U1275 (N_1275,N_1235,N_1247);
or U1276 (N_1276,N_1211,N_1245);
nand U1277 (N_1277,N_1230,N_1202);
or U1278 (N_1278,N_1219,N_1200);
nor U1279 (N_1279,N_1244,N_1241);
nor U1280 (N_1280,N_1215,N_1202);
nand U1281 (N_1281,N_1234,N_1242);
and U1282 (N_1282,N_1224,N_1215);
or U1283 (N_1283,N_1248,N_1208);
nand U1284 (N_1284,N_1211,N_1200);
nor U1285 (N_1285,N_1212,N_1228);
and U1286 (N_1286,N_1212,N_1244);
and U1287 (N_1287,N_1237,N_1214);
and U1288 (N_1288,N_1213,N_1215);
nand U1289 (N_1289,N_1216,N_1215);
nor U1290 (N_1290,N_1204,N_1228);
nand U1291 (N_1291,N_1209,N_1211);
or U1292 (N_1292,N_1236,N_1207);
and U1293 (N_1293,N_1204,N_1222);
and U1294 (N_1294,N_1217,N_1204);
nor U1295 (N_1295,N_1202,N_1233);
and U1296 (N_1296,N_1218,N_1238);
xor U1297 (N_1297,N_1210,N_1237);
nor U1298 (N_1298,N_1249,N_1219);
nand U1299 (N_1299,N_1217,N_1239);
nand U1300 (N_1300,N_1288,N_1279);
or U1301 (N_1301,N_1262,N_1271);
xor U1302 (N_1302,N_1261,N_1292);
nor U1303 (N_1303,N_1289,N_1250);
nor U1304 (N_1304,N_1270,N_1268);
xnor U1305 (N_1305,N_1266,N_1283);
nor U1306 (N_1306,N_1278,N_1298);
xnor U1307 (N_1307,N_1251,N_1256);
nor U1308 (N_1308,N_1282,N_1272);
and U1309 (N_1309,N_1296,N_1265);
nand U1310 (N_1310,N_1258,N_1269);
nand U1311 (N_1311,N_1264,N_1252);
or U1312 (N_1312,N_1285,N_1267);
nand U1313 (N_1313,N_1275,N_1260);
nor U1314 (N_1314,N_1253,N_1294);
nand U1315 (N_1315,N_1255,N_1286);
and U1316 (N_1316,N_1297,N_1273);
nor U1317 (N_1317,N_1254,N_1290);
nor U1318 (N_1318,N_1299,N_1263);
nand U1319 (N_1319,N_1280,N_1276);
or U1320 (N_1320,N_1257,N_1291);
and U1321 (N_1321,N_1274,N_1277);
and U1322 (N_1322,N_1284,N_1259);
nor U1323 (N_1323,N_1295,N_1287);
and U1324 (N_1324,N_1293,N_1281);
nor U1325 (N_1325,N_1253,N_1281);
nand U1326 (N_1326,N_1276,N_1253);
nor U1327 (N_1327,N_1266,N_1272);
xnor U1328 (N_1328,N_1270,N_1254);
or U1329 (N_1329,N_1270,N_1278);
or U1330 (N_1330,N_1273,N_1250);
or U1331 (N_1331,N_1283,N_1290);
nor U1332 (N_1332,N_1287,N_1257);
nor U1333 (N_1333,N_1252,N_1296);
and U1334 (N_1334,N_1273,N_1262);
nor U1335 (N_1335,N_1281,N_1280);
nand U1336 (N_1336,N_1269,N_1279);
or U1337 (N_1337,N_1275,N_1298);
nand U1338 (N_1338,N_1267,N_1286);
nor U1339 (N_1339,N_1260,N_1273);
and U1340 (N_1340,N_1296,N_1272);
or U1341 (N_1341,N_1277,N_1288);
or U1342 (N_1342,N_1250,N_1280);
and U1343 (N_1343,N_1261,N_1287);
or U1344 (N_1344,N_1273,N_1263);
nand U1345 (N_1345,N_1290,N_1255);
nand U1346 (N_1346,N_1251,N_1275);
and U1347 (N_1347,N_1266,N_1263);
nand U1348 (N_1348,N_1298,N_1272);
and U1349 (N_1349,N_1270,N_1277);
nor U1350 (N_1350,N_1300,N_1318);
and U1351 (N_1351,N_1335,N_1326);
nand U1352 (N_1352,N_1325,N_1310);
nand U1353 (N_1353,N_1338,N_1308);
or U1354 (N_1354,N_1327,N_1343);
nor U1355 (N_1355,N_1322,N_1301);
or U1356 (N_1356,N_1336,N_1305);
or U1357 (N_1357,N_1345,N_1323);
or U1358 (N_1358,N_1304,N_1348);
nor U1359 (N_1359,N_1328,N_1332);
xnor U1360 (N_1360,N_1317,N_1319);
or U1361 (N_1361,N_1333,N_1315);
or U1362 (N_1362,N_1330,N_1346);
nor U1363 (N_1363,N_1320,N_1339);
nand U1364 (N_1364,N_1321,N_1331);
and U1365 (N_1365,N_1342,N_1347);
nor U1366 (N_1366,N_1313,N_1302);
nor U1367 (N_1367,N_1337,N_1312);
nor U1368 (N_1368,N_1344,N_1306);
nand U1369 (N_1369,N_1311,N_1309);
nor U1370 (N_1370,N_1324,N_1329);
nor U1371 (N_1371,N_1334,N_1314);
nor U1372 (N_1372,N_1307,N_1340);
nor U1373 (N_1373,N_1316,N_1349);
nand U1374 (N_1374,N_1303,N_1341);
or U1375 (N_1375,N_1336,N_1327);
nor U1376 (N_1376,N_1348,N_1316);
nor U1377 (N_1377,N_1321,N_1340);
and U1378 (N_1378,N_1329,N_1348);
nand U1379 (N_1379,N_1329,N_1326);
nor U1380 (N_1380,N_1317,N_1300);
or U1381 (N_1381,N_1313,N_1344);
nand U1382 (N_1382,N_1338,N_1344);
xnor U1383 (N_1383,N_1308,N_1318);
nor U1384 (N_1384,N_1339,N_1325);
nor U1385 (N_1385,N_1335,N_1318);
nor U1386 (N_1386,N_1305,N_1326);
and U1387 (N_1387,N_1302,N_1340);
and U1388 (N_1388,N_1336,N_1319);
nand U1389 (N_1389,N_1304,N_1339);
and U1390 (N_1390,N_1346,N_1322);
nand U1391 (N_1391,N_1327,N_1341);
xnor U1392 (N_1392,N_1346,N_1320);
nand U1393 (N_1393,N_1330,N_1342);
nand U1394 (N_1394,N_1328,N_1344);
and U1395 (N_1395,N_1349,N_1325);
nand U1396 (N_1396,N_1333,N_1305);
and U1397 (N_1397,N_1326,N_1331);
and U1398 (N_1398,N_1311,N_1349);
nand U1399 (N_1399,N_1313,N_1334);
nand U1400 (N_1400,N_1391,N_1350);
xor U1401 (N_1401,N_1359,N_1371);
xor U1402 (N_1402,N_1372,N_1392);
or U1403 (N_1403,N_1356,N_1379);
or U1404 (N_1404,N_1377,N_1374);
nand U1405 (N_1405,N_1362,N_1390);
nor U1406 (N_1406,N_1389,N_1367);
xor U1407 (N_1407,N_1394,N_1360);
nand U1408 (N_1408,N_1355,N_1366);
nor U1409 (N_1409,N_1363,N_1393);
and U1410 (N_1410,N_1375,N_1381);
and U1411 (N_1411,N_1357,N_1397);
or U1412 (N_1412,N_1354,N_1370);
xor U1413 (N_1413,N_1369,N_1368);
and U1414 (N_1414,N_1386,N_1388);
nand U1415 (N_1415,N_1382,N_1376);
nor U1416 (N_1416,N_1358,N_1387);
and U1417 (N_1417,N_1373,N_1399);
or U1418 (N_1418,N_1361,N_1364);
nor U1419 (N_1419,N_1380,N_1352);
or U1420 (N_1420,N_1365,N_1384);
nor U1421 (N_1421,N_1383,N_1378);
and U1422 (N_1422,N_1396,N_1395);
nor U1423 (N_1423,N_1353,N_1398);
and U1424 (N_1424,N_1385,N_1351);
nor U1425 (N_1425,N_1355,N_1394);
and U1426 (N_1426,N_1397,N_1398);
or U1427 (N_1427,N_1399,N_1359);
and U1428 (N_1428,N_1352,N_1364);
nand U1429 (N_1429,N_1375,N_1393);
nand U1430 (N_1430,N_1383,N_1354);
or U1431 (N_1431,N_1389,N_1397);
and U1432 (N_1432,N_1373,N_1360);
nand U1433 (N_1433,N_1359,N_1353);
and U1434 (N_1434,N_1367,N_1363);
nand U1435 (N_1435,N_1356,N_1359);
nand U1436 (N_1436,N_1385,N_1393);
nand U1437 (N_1437,N_1379,N_1372);
and U1438 (N_1438,N_1358,N_1388);
or U1439 (N_1439,N_1377,N_1372);
or U1440 (N_1440,N_1359,N_1382);
and U1441 (N_1441,N_1383,N_1372);
and U1442 (N_1442,N_1390,N_1359);
nand U1443 (N_1443,N_1375,N_1362);
or U1444 (N_1444,N_1367,N_1376);
or U1445 (N_1445,N_1396,N_1367);
or U1446 (N_1446,N_1380,N_1353);
nor U1447 (N_1447,N_1385,N_1350);
nand U1448 (N_1448,N_1375,N_1353);
xor U1449 (N_1449,N_1397,N_1375);
and U1450 (N_1450,N_1448,N_1423);
and U1451 (N_1451,N_1444,N_1446);
or U1452 (N_1452,N_1427,N_1414);
nor U1453 (N_1453,N_1402,N_1431);
nor U1454 (N_1454,N_1426,N_1418);
nor U1455 (N_1455,N_1403,N_1442);
nand U1456 (N_1456,N_1412,N_1428);
nor U1457 (N_1457,N_1413,N_1409);
and U1458 (N_1458,N_1439,N_1416);
or U1459 (N_1459,N_1449,N_1435);
nand U1460 (N_1460,N_1445,N_1407);
xor U1461 (N_1461,N_1400,N_1419);
and U1462 (N_1462,N_1417,N_1415);
or U1463 (N_1463,N_1406,N_1422);
and U1464 (N_1464,N_1438,N_1410);
nand U1465 (N_1465,N_1434,N_1429);
nand U1466 (N_1466,N_1436,N_1437);
or U1467 (N_1467,N_1405,N_1404);
nor U1468 (N_1468,N_1447,N_1443);
nand U1469 (N_1469,N_1408,N_1420);
nand U1470 (N_1470,N_1433,N_1425);
nand U1471 (N_1471,N_1401,N_1411);
or U1472 (N_1472,N_1441,N_1421);
or U1473 (N_1473,N_1440,N_1430);
and U1474 (N_1474,N_1424,N_1432);
xnor U1475 (N_1475,N_1432,N_1423);
or U1476 (N_1476,N_1428,N_1424);
nor U1477 (N_1477,N_1416,N_1426);
or U1478 (N_1478,N_1440,N_1412);
or U1479 (N_1479,N_1406,N_1444);
and U1480 (N_1480,N_1431,N_1429);
or U1481 (N_1481,N_1426,N_1435);
nor U1482 (N_1482,N_1445,N_1415);
and U1483 (N_1483,N_1437,N_1422);
and U1484 (N_1484,N_1410,N_1417);
xor U1485 (N_1485,N_1445,N_1431);
or U1486 (N_1486,N_1443,N_1401);
nor U1487 (N_1487,N_1410,N_1420);
and U1488 (N_1488,N_1447,N_1434);
and U1489 (N_1489,N_1426,N_1429);
nand U1490 (N_1490,N_1405,N_1401);
nand U1491 (N_1491,N_1447,N_1420);
nand U1492 (N_1492,N_1433,N_1403);
xnor U1493 (N_1493,N_1406,N_1439);
nand U1494 (N_1494,N_1405,N_1439);
nand U1495 (N_1495,N_1421,N_1418);
xor U1496 (N_1496,N_1411,N_1436);
nand U1497 (N_1497,N_1440,N_1446);
nand U1498 (N_1498,N_1435,N_1443);
and U1499 (N_1499,N_1407,N_1403);
nor U1500 (N_1500,N_1473,N_1456);
nor U1501 (N_1501,N_1488,N_1499);
xor U1502 (N_1502,N_1450,N_1472);
nand U1503 (N_1503,N_1458,N_1462);
and U1504 (N_1504,N_1477,N_1465);
nor U1505 (N_1505,N_1481,N_1490);
nand U1506 (N_1506,N_1461,N_1491);
nor U1507 (N_1507,N_1463,N_1489);
or U1508 (N_1508,N_1471,N_1467);
and U1509 (N_1509,N_1482,N_1480);
nor U1510 (N_1510,N_1484,N_1495);
and U1511 (N_1511,N_1493,N_1498);
nand U1512 (N_1512,N_1464,N_1468);
and U1513 (N_1513,N_1454,N_1451);
and U1514 (N_1514,N_1497,N_1452);
nor U1515 (N_1515,N_1453,N_1496);
and U1516 (N_1516,N_1470,N_1486);
or U1517 (N_1517,N_1487,N_1457);
nand U1518 (N_1518,N_1455,N_1474);
or U1519 (N_1519,N_1479,N_1492);
and U1520 (N_1520,N_1459,N_1460);
nand U1521 (N_1521,N_1478,N_1476);
or U1522 (N_1522,N_1475,N_1469);
nor U1523 (N_1523,N_1485,N_1494);
and U1524 (N_1524,N_1466,N_1483);
nand U1525 (N_1525,N_1469,N_1499);
nand U1526 (N_1526,N_1453,N_1473);
nand U1527 (N_1527,N_1489,N_1487);
or U1528 (N_1528,N_1454,N_1458);
and U1529 (N_1529,N_1499,N_1494);
nand U1530 (N_1530,N_1460,N_1484);
nand U1531 (N_1531,N_1493,N_1491);
and U1532 (N_1532,N_1455,N_1499);
nor U1533 (N_1533,N_1490,N_1470);
or U1534 (N_1534,N_1481,N_1455);
nand U1535 (N_1535,N_1477,N_1480);
xnor U1536 (N_1536,N_1453,N_1493);
nand U1537 (N_1537,N_1451,N_1452);
and U1538 (N_1538,N_1454,N_1493);
and U1539 (N_1539,N_1473,N_1484);
nand U1540 (N_1540,N_1451,N_1466);
and U1541 (N_1541,N_1459,N_1471);
and U1542 (N_1542,N_1495,N_1464);
or U1543 (N_1543,N_1452,N_1492);
nand U1544 (N_1544,N_1460,N_1498);
nand U1545 (N_1545,N_1465,N_1460);
or U1546 (N_1546,N_1466,N_1464);
or U1547 (N_1547,N_1459,N_1467);
xnor U1548 (N_1548,N_1498,N_1495);
nand U1549 (N_1549,N_1486,N_1484);
or U1550 (N_1550,N_1526,N_1502);
or U1551 (N_1551,N_1548,N_1542);
and U1552 (N_1552,N_1543,N_1529);
or U1553 (N_1553,N_1532,N_1538);
and U1554 (N_1554,N_1534,N_1531);
and U1555 (N_1555,N_1528,N_1517);
nor U1556 (N_1556,N_1509,N_1525);
xnor U1557 (N_1557,N_1540,N_1516);
xor U1558 (N_1558,N_1505,N_1547);
nand U1559 (N_1559,N_1510,N_1535);
and U1560 (N_1560,N_1507,N_1515);
nor U1561 (N_1561,N_1511,N_1527);
nand U1562 (N_1562,N_1539,N_1503);
nand U1563 (N_1563,N_1523,N_1508);
nand U1564 (N_1564,N_1545,N_1520);
nand U1565 (N_1565,N_1546,N_1519);
and U1566 (N_1566,N_1512,N_1518);
nor U1567 (N_1567,N_1501,N_1536);
nor U1568 (N_1568,N_1549,N_1521);
nor U1569 (N_1569,N_1522,N_1524);
xnor U1570 (N_1570,N_1506,N_1544);
and U1571 (N_1571,N_1541,N_1533);
or U1572 (N_1572,N_1513,N_1514);
and U1573 (N_1573,N_1537,N_1500);
and U1574 (N_1574,N_1504,N_1530);
nor U1575 (N_1575,N_1530,N_1521);
nand U1576 (N_1576,N_1534,N_1547);
or U1577 (N_1577,N_1521,N_1539);
and U1578 (N_1578,N_1543,N_1542);
xor U1579 (N_1579,N_1537,N_1501);
xor U1580 (N_1580,N_1513,N_1505);
and U1581 (N_1581,N_1549,N_1518);
and U1582 (N_1582,N_1541,N_1510);
nand U1583 (N_1583,N_1505,N_1532);
nor U1584 (N_1584,N_1511,N_1516);
nor U1585 (N_1585,N_1535,N_1509);
nand U1586 (N_1586,N_1512,N_1528);
nor U1587 (N_1587,N_1501,N_1519);
nand U1588 (N_1588,N_1544,N_1501);
nand U1589 (N_1589,N_1532,N_1543);
nor U1590 (N_1590,N_1534,N_1503);
nand U1591 (N_1591,N_1524,N_1511);
or U1592 (N_1592,N_1515,N_1543);
xor U1593 (N_1593,N_1546,N_1544);
and U1594 (N_1594,N_1547,N_1520);
or U1595 (N_1595,N_1504,N_1545);
nor U1596 (N_1596,N_1535,N_1522);
nor U1597 (N_1597,N_1507,N_1510);
nand U1598 (N_1598,N_1514,N_1537);
nand U1599 (N_1599,N_1505,N_1509);
or U1600 (N_1600,N_1575,N_1554);
and U1601 (N_1601,N_1571,N_1569);
nand U1602 (N_1602,N_1551,N_1559);
or U1603 (N_1603,N_1588,N_1589);
nor U1604 (N_1604,N_1592,N_1553);
nand U1605 (N_1605,N_1579,N_1598);
nor U1606 (N_1606,N_1555,N_1597);
or U1607 (N_1607,N_1593,N_1576);
nor U1608 (N_1608,N_1584,N_1590);
nor U1609 (N_1609,N_1582,N_1585);
and U1610 (N_1610,N_1570,N_1552);
nor U1611 (N_1611,N_1566,N_1568);
or U1612 (N_1612,N_1564,N_1558);
nor U1613 (N_1613,N_1595,N_1596);
and U1614 (N_1614,N_1587,N_1565);
nor U1615 (N_1615,N_1561,N_1583);
or U1616 (N_1616,N_1581,N_1580);
or U1617 (N_1617,N_1573,N_1599);
nor U1618 (N_1618,N_1556,N_1586);
nor U1619 (N_1619,N_1577,N_1550);
and U1620 (N_1620,N_1591,N_1557);
nor U1621 (N_1621,N_1560,N_1572);
and U1622 (N_1622,N_1574,N_1578);
or U1623 (N_1623,N_1562,N_1567);
nor U1624 (N_1624,N_1563,N_1594);
or U1625 (N_1625,N_1578,N_1567);
or U1626 (N_1626,N_1585,N_1557);
nor U1627 (N_1627,N_1573,N_1591);
or U1628 (N_1628,N_1582,N_1551);
nor U1629 (N_1629,N_1582,N_1565);
or U1630 (N_1630,N_1566,N_1562);
or U1631 (N_1631,N_1583,N_1580);
or U1632 (N_1632,N_1598,N_1592);
nor U1633 (N_1633,N_1585,N_1553);
or U1634 (N_1634,N_1562,N_1561);
or U1635 (N_1635,N_1568,N_1586);
and U1636 (N_1636,N_1559,N_1584);
and U1637 (N_1637,N_1568,N_1578);
and U1638 (N_1638,N_1593,N_1560);
and U1639 (N_1639,N_1596,N_1597);
or U1640 (N_1640,N_1581,N_1575);
or U1641 (N_1641,N_1596,N_1585);
and U1642 (N_1642,N_1561,N_1557);
nand U1643 (N_1643,N_1562,N_1589);
nor U1644 (N_1644,N_1594,N_1564);
or U1645 (N_1645,N_1580,N_1587);
and U1646 (N_1646,N_1594,N_1565);
and U1647 (N_1647,N_1584,N_1575);
nor U1648 (N_1648,N_1554,N_1567);
or U1649 (N_1649,N_1575,N_1550);
xor U1650 (N_1650,N_1630,N_1624);
nand U1651 (N_1651,N_1632,N_1641);
nand U1652 (N_1652,N_1629,N_1604);
or U1653 (N_1653,N_1649,N_1609);
nor U1654 (N_1654,N_1648,N_1611);
nand U1655 (N_1655,N_1610,N_1612);
xor U1656 (N_1656,N_1634,N_1608);
nor U1657 (N_1657,N_1619,N_1635);
and U1658 (N_1658,N_1623,N_1617);
or U1659 (N_1659,N_1640,N_1605);
nor U1660 (N_1660,N_1603,N_1636);
xnor U1661 (N_1661,N_1642,N_1647);
or U1662 (N_1662,N_1620,N_1613);
or U1663 (N_1663,N_1644,N_1614);
and U1664 (N_1664,N_1646,N_1622);
nand U1665 (N_1665,N_1621,N_1639);
nand U1666 (N_1666,N_1600,N_1615);
xnor U1667 (N_1667,N_1607,N_1643);
and U1668 (N_1668,N_1618,N_1645);
and U1669 (N_1669,N_1631,N_1616);
nor U1670 (N_1670,N_1626,N_1625);
or U1671 (N_1671,N_1638,N_1637);
nand U1672 (N_1672,N_1628,N_1602);
xor U1673 (N_1673,N_1601,N_1627);
and U1674 (N_1674,N_1606,N_1633);
or U1675 (N_1675,N_1623,N_1603);
nor U1676 (N_1676,N_1629,N_1615);
and U1677 (N_1677,N_1611,N_1635);
nand U1678 (N_1678,N_1640,N_1607);
or U1679 (N_1679,N_1626,N_1629);
or U1680 (N_1680,N_1600,N_1633);
nor U1681 (N_1681,N_1623,N_1631);
nand U1682 (N_1682,N_1616,N_1623);
or U1683 (N_1683,N_1612,N_1633);
nor U1684 (N_1684,N_1619,N_1640);
and U1685 (N_1685,N_1605,N_1639);
nor U1686 (N_1686,N_1605,N_1611);
xnor U1687 (N_1687,N_1630,N_1647);
nor U1688 (N_1688,N_1602,N_1627);
and U1689 (N_1689,N_1624,N_1643);
and U1690 (N_1690,N_1622,N_1635);
xnor U1691 (N_1691,N_1639,N_1631);
nor U1692 (N_1692,N_1627,N_1616);
nor U1693 (N_1693,N_1610,N_1628);
and U1694 (N_1694,N_1641,N_1607);
or U1695 (N_1695,N_1617,N_1619);
nor U1696 (N_1696,N_1613,N_1642);
or U1697 (N_1697,N_1606,N_1649);
xor U1698 (N_1698,N_1635,N_1648);
nor U1699 (N_1699,N_1617,N_1601);
or U1700 (N_1700,N_1693,N_1685);
nor U1701 (N_1701,N_1669,N_1658);
or U1702 (N_1702,N_1652,N_1675);
nand U1703 (N_1703,N_1666,N_1691);
xor U1704 (N_1704,N_1663,N_1662);
nand U1705 (N_1705,N_1697,N_1683);
xor U1706 (N_1706,N_1690,N_1676);
nor U1707 (N_1707,N_1654,N_1672);
nor U1708 (N_1708,N_1692,N_1664);
nand U1709 (N_1709,N_1679,N_1670);
or U1710 (N_1710,N_1695,N_1650);
xor U1711 (N_1711,N_1660,N_1671);
and U1712 (N_1712,N_1680,N_1681);
or U1713 (N_1713,N_1696,N_1661);
or U1714 (N_1714,N_1688,N_1655);
and U1715 (N_1715,N_1659,N_1699);
and U1716 (N_1716,N_1698,N_1656);
nor U1717 (N_1717,N_1684,N_1694);
nor U1718 (N_1718,N_1689,N_1668);
nor U1719 (N_1719,N_1665,N_1653);
nand U1720 (N_1720,N_1687,N_1657);
nor U1721 (N_1721,N_1674,N_1673);
nand U1722 (N_1722,N_1678,N_1682);
or U1723 (N_1723,N_1667,N_1677);
nand U1724 (N_1724,N_1686,N_1651);
and U1725 (N_1725,N_1699,N_1669);
or U1726 (N_1726,N_1654,N_1656);
xnor U1727 (N_1727,N_1653,N_1695);
nand U1728 (N_1728,N_1662,N_1657);
xnor U1729 (N_1729,N_1665,N_1656);
xor U1730 (N_1730,N_1651,N_1653);
and U1731 (N_1731,N_1671,N_1697);
or U1732 (N_1732,N_1688,N_1698);
and U1733 (N_1733,N_1662,N_1658);
and U1734 (N_1734,N_1680,N_1689);
nor U1735 (N_1735,N_1665,N_1691);
xnor U1736 (N_1736,N_1689,N_1678);
nor U1737 (N_1737,N_1670,N_1666);
nand U1738 (N_1738,N_1691,N_1651);
nand U1739 (N_1739,N_1651,N_1696);
and U1740 (N_1740,N_1669,N_1681);
and U1741 (N_1741,N_1693,N_1683);
nand U1742 (N_1742,N_1679,N_1693);
or U1743 (N_1743,N_1688,N_1653);
nor U1744 (N_1744,N_1652,N_1698);
nor U1745 (N_1745,N_1650,N_1682);
and U1746 (N_1746,N_1695,N_1680);
and U1747 (N_1747,N_1669,N_1653);
nand U1748 (N_1748,N_1661,N_1655);
nor U1749 (N_1749,N_1666,N_1699);
nor U1750 (N_1750,N_1734,N_1725);
or U1751 (N_1751,N_1715,N_1738);
and U1752 (N_1752,N_1728,N_1726);
nor U1753 (N_1753,N_1710,N_1729);
or U1754 (N_1754,N_1741,N_1749);
and U1755 (N_1755,N_1713,N_1724);
or U1756 (N_1756,N_1737,N_1742);
nor U1757 (N_1757,N_1736,N_1743);
nand U1758 (N_1758,N_1746,N_1744);
or U1759 (N_1759,N_1714,N_1727);
nand U1760 (N_1760,N_1709,N_1700);
and U1761 (N_1761,N_1748,N_1733);
xor U1762 (N_1762,N_1718,N_1723);
nand U1763 (N_1763,N_1717,N_1716);
xor U1764 (N_1764,N_1706,N_1739);
or U1765 (N_1765,N_1730,N_1722);
nor U1766 (N_1766,N_1719,N_1721);
nand U1767 (N_1767,N_1720,N_1707);
and U1768 (N_1768,N_1704,N_1711);
or U1769 (N_1769,N_1705,N_1701);
nor U1770 (N_1770,N_1740,N_1745);
nor U1771 (N_1771,N_1732,N_1702);
and U1772 (N_1772,N_1747,N_1731);
and U1773 (N_1773,N_1712,N_1703);
nand U1774 (N_1774,N_1735,N_1708);
nand U1775 (N_1775,N_1745,N_1729);
xnor U1776 (N_1776,N_1711,N_1730);
nand U1777 (N_1777,N_1709,N_1701);
nor U1778 (N_1778,N_1748,N_1707);
nand U1779 (N_1779,N_1712,N_1727);
nand U1780 (N_1780,N_1746,N_1731);
nand U1781 (N_1781,N_1722,N_1717);
or U1782 (N_1782,N_1723,N_1728);
xnor U1783 (N_1783,N_1735,N_1737);
and U1784 (N_1784,N_1728,N_1708);
nor U1785 (N_1785,N_1720,N_1725);
and U1786 (N_1786,N_1719,N_1714);
nor U1787 (N_1787,N_1736,N_1720);
nand U1788 (N_1788,N_1716,N_1742);
or U1789 (N_1789,N_1700,N_1727);
xnor U1790 (N_1790,N_1721,N_1706);
xor U1791 (N_1791,N_1728,N_1701);
and U1792 (N_1792,N_1721,N_1741);
nor U1793 (N_1793,N_1707,N_1729);
nor U1794 (N_1794,N_1731,N_1725);
nor U1795 (N_1795,N_1700,N_1734);
nor U1796 (N_1796,N_1715,N_1705);
nand U1797 (N_1797,N_1722,N_1741);
nor U1798 (N_1798,N_1705,N_1736);
nand U1799 (N_1799,N_1724,N_1737);
nor U1800 (N_1800,N_1797,N_1751);
xor U1801 (N_1801,N_1786,N_1774);
nand U1802 (N_1802,N_1761,N_1788);
and U1803 (N_1803,N_1771,N_1793);
nor U1804 (N_1804,N_1759,N_1791);
and U1805 (N_1805,N_1770,N_1796);
and U1806 (N_1806,N_1752,N_1792);
nor U1807 (N_1807,N_1795,N_1750);
nand U1808 (N_1808,N_1782,N_1783);
or U1809 (N_1809,N_1779,N_1756);
xor U1810 (N_1810,N_1785,N_1789);
and U1811 (N_1811,N_1798,N_1772);
nor U1812 (N_1812,N_1764,N_1794);
nor U1813 (N_1813,N_1754,N_1758);
nor U1814 (N_1814,N_1781,N_1753);
nand U1815 (N_1815,N_1769,N_1757);
xor U1816 (N_1816,N_1767,N_1799);
nand U1817 (N_1817,N_1762,N_1787);
nor U1818 (N_1818,N_1784,N_1776);
and U1819 (N_1819,N_1760,N_1778);
and U1820 (N_1820,N_1790,N_1755);
and U1821 (N_1821,N_1780,N_1766);
nor U1822 (N_1822,N_1777,N_1765);
nor U1823 (N_1823,N_1763,N_1775);
or U1824 (N_1824,N_1773,N_1768);
nor U1825 (N_1825,N_1792,N_1758);
and U1826 (N_1826,N_1781,N_1785);
nor U1827 (N_1827,N_1753,N_1770);
nor U1828 (N_1828,N_1783,N_1797);
and U1829 (N_1829,N_1758,N_1790);
nor U1830 (N_1830,N_1797,N_1755);
xnor U1831 (N_1831,N_1787,N_1792);
xnor U1832 (N_1832,N_1787,N_1764);
or U1833 (N_1833,N_1761,N_1786);
xnor U1834 (N_1834,N_1751,N_1777);
nand U1835 (N_1835,N_1781,N_1762);
nor U1836 (N_1836,N_1780,N_1759);
nand U1837 (N_1837,N_1769,N_1798);
and U1838 (N_1838,N_1773,N_1793);
and U1839 (N_1839,N_1764,N_1768);
nor U1840 (N_1840,N_1796,N_1779);
and U1841 (N_1841,N_1785,N_1787);
and U1842 (N_1842,N_1798,N_1751);
nor U1843 (N_1843,N_1796,N_1787);
nor U1844 (N_1844,N_1781,N_1769);
nand U1845 (N_1845,N_1752,N_1761);
nand U1846 (N_1846,N_1760,N_1754);
nand U1847 (N_1847,N_1767,N_1758);
and U1848 (N_1848,N_1773,N_1791);
and U1849 (N_1849,N_1756,N_1757);
or U1850 (N_1850,N_1812,N_1828);
xnor U1851 (N_1851,N_1831,N_1835);
and U1852 (N_1852,N_1849,N_1829);
or U1853 (N_1853,N_1816,N_1817);
and U1854 (N_1854,N_1800,N_1810);
and U1855 (N_1855,N_1842,N_1801);
nand U1856 (N_1856,N_1809,N_1834);
nand U1857 (N_1857,N_1820,N_1848);
or U1858 (N_1858,N_1802,N_1805);
or U1859 (N_1859,N_1811,N_1838);
or U1860 (N_1860,N_1815,N_1823);
or U1861 (N_1861,N_1804,N_1819);
and U1862 (N_1862,N_1843,N_1808);
nor U1863 (N_1863,N_1825,N_1827);
nor U1864 (N_1864,N_1844,N_1830);
or U1865 (N_1865,N_1833,N_1814);
nand U1866 (N_1866,N_1841,N_1837);
nand U1867 (N_1867,N_1806,N_1822);
xnor U1868 (N_1868,N_1824,N_1832);
nand U1869 (N_1869,N_1807,N_1818);
or U1870 (N_1870,N_1803,N_1839);
nand U1871 (N_1871,N_1826,N_1813);
or U1872 (N_1872,N_1845,N_1840);
and U1873 (N_1873,N_1847,N_1846);
nand U1874 (N_1874,N_1836,N_1821);
nand U1875 (N_1875,N_1821,N_1830);
or U1876 (N_1876,N_1839,N_1824);
or U1877 (N_1877,N_1838,N_1800);
or U1878 (N_1878,N_1816,N_1849);
or U1879 (N_1879,N_1836,N_1813);
and U1880 (N_1880,N_1845,N_1819);
nand U1881 (N_1881,N_1819,N_1841);
and U1882 (N_1882,N_1813,N_1844);
nor U1883 (N_1883,N_1800,N_1831);
nor U1884 (N_1884,N_1820,N_1837);
nand U1885 (N_1885,N_1808,N_1815);
and U1886 (N_1886,N_1832,N_1810);
xnor U1887 (N_1887,N_1826,N_1827);
nor U1888 (N_1888,N_1816,N_1839);
and U1889 (N_1889,N_1801,N_1831);
and U1890 (N_1890,N_1840,N_1827);
and U1891 (N_1891,N_1839,N_1831);
nand U1892 (N_1892,N_1807,N_1842);
xor U1893 (N_1893,N_1810,N_1812);
or U1894 (N_1894,N_1823,N_1811);
nand U1895 (N_1895,N_1842,N_1848);
and U1896 (N_1896,N_1810,N_1842);
nor U1897 (N_1897,N_1815,N_1831);
or U1898 (N_1898,N_1807,N_1836);
and U1899 (N_1899,N_1818,N_1849);
nor U1900 (N_1900,N_1870,N_1861);
nor U1901 (N_1901,N_1869,N_1853);
nor U1902 (N_1902,N_1876,N_1859);
nand U1903 (N_1903,N_1889,N_1854);
nor U1904 (N_1904,N_1890,N_1899);
nor U1905 (N_1905,N_1893,N_1865);
or U1906 (N_1906,N_1872,N_1866);
nand U1907 (N_1907,N_1886,N_1898);
nand U1908 (N_1908,N_1851,N_1863);
xnor U1909 (N_1909,N_1855,N_1852);
and U1910 (N_1910,N_1874,N_1882);
or U1911 (N_1911,N_1891,N_1856);
nand U1912 (N_1912,N_1885,N_1879);
or U1913 (N_1913,N_1896,N_1873);
or U1914 (N_1914,N_1883,N_1871);
nor U1915 (N_1915,N_1868,N_1887);
nor U1916 (N_1916,N_1867,N_1877);
nor U1917 (N_1917,N_1880,N_1895);
nand U1918 (N_1918,N_1858,N_1875);
nand U1919 (N_1919,N_1892,N_1897);
nor U1920 (N_1920,N_1860,N_1888);
or U1921 (N_1921,N_1884,N_1864);
or U1922 (N_1922,N_1862,N_1894);
nor U1923 (N_1923,N_1850,N_1878);
or U1924 (N_1924,N_1857,N_1881);
nand U1925 (N_1925,N_1856,N_1864);
and U1926 (N_1926,N_1895,N_1881);
xnor U1927 (N_1927,N_1883,N_1886);
and U1928 (N_1928,N_1878,N_1875);
nor U1929 (N_1929,N_1896,N_1861);
or U1930 (N_1930,N_1893,N_1871);
or U1931 (N_1931,N_1888,N_1871);
or U1932 (N_1932,N_1852,N_1871);
xnor U1933 (N_1933,N_1853,N_1896);
and U1934 (N_1934,N_1887,N_1870);
and U1935 (N_1935,N_1866,N_1896);
and U1936 (N_1936,N_1883,N_1876);
nor U1937 (N_1937,N_1886,N_1885);
nand U1938 (N_1938,N_1893,N_1877);
xnor U1939 (N_1939,N_1865,N_1850);
xor U1940 (N_1940,N_1854,N_1893);
nand U1941 (N_1941,N_1875,N_1887);
nand U1942 (N_1942,N_1858,N_1869);
or U1943 (N_1943,N_1880,N_1890);
nor U1944 (N_1944,N_1860,N_1850);
nor U1945 (N_1945,N_1874,N_1877);
nor U1946 (N_1946,N_1889,N_1899);
nor U1947 (N_1947,N_1885,N_1863);
nor U1948 (N_1948,N_1874,N_1853);
and U1949 (N_1949,N_1858,N_1886);
xnor U1950 (N_1950,N_1905,N_1916);
or U1951 (N_1951,N_1939,N_1920);
and U1952 (N_1952,N_1922,N_1906);
or U1953 (N_1953,N_1943,N_1923);
nand U1954 (N_1954,N_1907,N_1928);
xnor U1955 (N_1955,N_1919,N_1942);
xor U1956 (N_1956,N_1938,N_1918);
or U1957 (N_1957,N_1902,N_1940);
xnor U1958 (N_1958,N_1949,N_1930);
nand U1959 (N_1959,N_1913,N_1908);
and U1960 (N_1960,N_1910,N_1909);
nand U1961 (N_1961,N_1925,N_1926);
nor U1962 (N_1962,N_1911,N_1921);
xor U1963 (N_1963,N_1946,N_1947);
or U1964 (N_1964,N_1932,N_1924);
nand U1965 (N_1965,N_1900,N_1929);
nor U1966 (N_1966,N_1904,N_1948);
and U1967 (N_1967,N_1927,N_1903);
or U1968 (N_1968,N_1933,N_1937);
nor U1969 (N_1969,N_1912,N_1917);
nor U1970 (N_1970,N_1914,N_1944);
nand U1971 (N_1971,N_1936,N_1941);
and U1972 (N_1972,N_1945,N_1935);
or U1973 (N_1973,N_1901,N_1915);
xor U1974 (N_1974,N_1931,N_1934);
and U1975 (N_1975,N_1944,N_1943);
or U1976 (N_1976,N_1901,N_1921);
or U1977 (N_1977,N_1903,N_1924);
or U1978 (N_1978,N_1939,N_1933);
nor U1979 (N_1979,N_1911,N_1925);
xor U1980 (N_1980,N_1939,N_1907);
nor U1981 (N_1981,N_1916,N_1902);
nand U1982 (N_1982,N_1909,N_1948);
xor U1983 (N_1983,N_1908,N_1937);
nand U1984 (N_1984,N_1945,N_1902);
xnor U1985 (N_1985,N_1931,N_1946);
nand U1986 (N_1986,N_1936,N_1947);
nor U1987 (N_1987,N_1913,N_1937);
or U1988 (N_1988,N_1920,N_1934);
xor U1989 (N_1989,N_1915,N_1949);
and U1990 (N_1990,N_1932,N_1915);
nor U1991 (N_1991,N_1934,N_1938);
nand U1992 (N_1992,N_1936,N_1906);
nand U1993 (N_1993,N_1927,N_1923);
nor U1994 (N_1994,N_1932,N_1909);
and U1995 (N_1995,N_1922,N_1946);
or U1996 (N_1996,N_1906,N_1932);
and U1997 (N_1997,N_1935,N_1941);
and U1998 (N_1998,N_1909,N_1935);
or U1999 (N_1999,N_1924,N_1945);
nand U2000 (N_2000,N_1976,N_1977);
nand U2001 (N_2001,N_1984,N_1954);
or U2002 (N_2002,N_1974,N_1951);
nor U2003 (N_2003,N_1997,N_1986);
nor U2004 (N_2004,N_1964,N_1967);
nor U2005 (N_2005,N_1961,N_1953);
and U2006 (N_2006,N_1998,N_1989);
nand U2007 (N_2007,N_1970,N_1996);
or U2008 (N_2008,N_1994,N_1992);
and U2009 (N_2009,N_1980,N_1962);
and U2010 (N_2010,N_1972,N_1993);
xnor U2011 (N_2011,N_1958,N_1968);
nand U2012 (N_2012,N_1969,N_1965);
nor U2013 (N_2013,N_1983,N_1975);
and U2014 (N_2014,N_1950,N_1990);
xnor U2015 (N_2015,N_1971,N_1959);
nand U2016 (N_2016,N_1956,N_1966);
and U2017 (N_2017,N_1999,N_1991);
nand U2018 (N_2018,N_1979,N_1963);
or U2019 (N_2019,N_1985,N_1988);
nor U2020 (N_2020,N_1957,N_1978);
nor U2021 (N_2021,N_1960,N_1955);
nor U2022 (N_2022,N_1995,N_1987);
or U2023 (N_2023,N_1973,N_1982);
and U2024 (N_2024,N_1952,N_1981);
nand U2025 (N_2025,N_1985,N_1982);
nor U2026 (N_2026,N_1982,N_1954);
xor U2027 (N_2027,N_1950,N_1968);
and U2028 (N_2028,N_1997,N_1965);
and U2029 (N_2029,N_1974,N_1995);
and U2030 (N_2030,N_1993,N_1994);
or U2031 (N_2031,N_1997,N_1992);
nand U2032 (N_2032,N_1989,N_1986);
xor U2033 (N_2033,N_1978,N_1956);
and U2034 (N_2034,N_1957,N_1989);
or U2035 (N_2035,N_1961,N_1979);
xor U2036 (N_2036,N_1970,N_1997);
nor U2037 (N_2037,N_1980,N_1959);
nor U2038 (N_2038,N_1998,N_1999);
xor U2039 (N_2039,N_1978,N_1955);
or U2040 (N_2040,N_1974,N_1955);
nand U2041 (N_2041,N_1955,N_1994);
or U2042 (N_2042,N_1965,N_1970);
nand U2043 (N_2043,N_1961,N_1994);
nand U2044 (N_2044,N_1995,N_1956);
xor U2045 (N_2045,N_1958,N_1960);
nor U2046 (N_2046,N_1975,N_1950);
xor U2047 (N_2047,N_1970,N_1951);
or U2048 (N_2048,N_1970,N_1992);
and U2049 (N_2049,N_1965,N_1952);
or U2050 (N_2050,N_2028,N_2026);
and U2051 (N_2051,N_2049,N_2044);
nand U2052 (N_2052,N_2027,N_2045);
or U2053 (N_2053,N_2022,N_2043);
or U2054 (N_2054,N_2015,N_2004);
and U2055 (N_2055,N_2031,N_2037);
and U2056 (N_2056,N_2020,N_2033);
nand U2057 (N_2057,N_2032,N_2041);
nand U2058 (N_2058,N_2019,N_2014);
nand U2059 (N_2059,N_2011,N_2042);
or U2060 (N_2060,N_2047,N_2023);
nor U2061 (N_2061,N_2000,N_2006);
and U2062 (N_2062,N_2008,N_2017);
and U2063 (N_2063,N_2039,N_2002);
nor U2064 (N_2064,N_2010,N_2035);
and U2065 (N_2065,N_2007,N_2034);
nor U2066 (N_2066,N_2013,N_2003);
nand U2067 (N_2067,N_2040,N_2009);
xnor U2068 (N_2068,N_2029,N_2036);
nand U2069 (N_2069,N_2012,N_2005);
nand U2070 (N_2070,N_2021,N_2024);
or U2071 (N_2071,N_2046,N_2016);
and U2072 (N_2072,N_2001,N_2030);
nor U2073 (N_2073,N_2048,N_2038);
and U2074 (N_2074,N_2018,N_2025);
or U2075 (N_2075,N_2048,N_2043);
nand U2076 (N_2076,N_2003,N_2035);
or U2077 (N_2077,N_2027,N_2042);
nand U2078 (N_2078,N_2014,N_2024);
or U2079 (N_2079,N_2009,N_2002);
and U2080 (N_2080,N_2001,N_2020);
nor U2081 (N_2081,N_2022,N_2039);
or U2082 (N_2082,N_2016,N_2023);
or U2083 (N_2083,N_2037,N_2011);
nand U2084 (N_2084,N_2001,N_2033);
nor U2085 (N_2085,N_2003,N_2008);
nor U2086 (N_2086,N_2049,N_2035);
and U2087 (N_2087,N_2018,N_2002);
nand U2088 (N_2088,N_2038,N_2008);
nor U2089 (N_2089,N_2043,N_2008);
and U2090 (N_2090,N_2046,N_2003);
xnor U2091 (N_2091,N_2014,N_2048);
xnor U2092 (N_2092,N_2024,N_2040);
and U2093 (N_2093,N_2046,N_2001);
xnor U2094 (N_2094,N_2007,N_2026);
and U2095 (N_2095,N_2042,N_2020);
nand U2096 (N_2096,N_2048,N_2030);
nor U2097 (N_2097,N_2018,N_2027);
nand U2098 (N_2098,N_2000,N_2013);
or U2099 (N_2099,N_2009,N_2029);
and U2100 (N_2100,N_2097,N_2071);
nand U2101 (N_2101,N_2063,N_2096);
and U2102 (N_2102,N_2087,N_2051);
and U2103 (N_2103,N_2088,N_2072);
nor U2104 (N_2104,N_2074,N_2075);
xnor U2105 (N_2105,N_2069,N_2089);
or U2106 (N_2106,N_2094,N_2076);
nand U2107 (N_2107,N_2077,N_2064);
or U2108 (N_2108,N_2084,N_2073);
or U2109 (N_2109,N_2099,N_2055);
nor U2110 (N_2110,N_2093,N_2095);
nand U2111 (N_2111,N_2066,N_2068);
or U2112 (N_2112,N_2078,N_2059);
and U2113 (N_2113,N_2054,N_2086);
and U2114 (N_2114,N_2053,N_2060);
nand U2115 (N_2115,N_2091,N_2079);
nand U2116 (N_2116,N_2062,N_2090);
and U2117 (N_2117,N_2052,N_2082);
and U2118 (N_2118,N_2083,N_2050);
or U2119 (N_2119,N_2065,N_2056);
and U2120 (N_2120,N_2081,N_2080);
and U2121 (N_2121,N_2058,N_2061);
xor U2122 (N_2122,N_2098,N_2092);
nor U2123 (N_2123,N_2057,N_2067);
or U2124 (N_2124,N_2085,N_2070);
nor U2125 (N_2125,N_2053,N_2074);
nand U2126 (N_2126,N_2074,N_2073);
nor U2127 (N_2127,N_2071,N_2056);
or U2128 (N_2128,N_2068,N_2095);
and U2129 (N_2129,N_2096,N_2092);
nand U2130 (N_2130,N_2077,N_2076);
nor U2131 (N_2131,N_2055,N_2072);
nor U2132 (N_2132,N_2050,N_2077);
and U2133 (N_2133,N_2061,N_2069);
nand U2134 (N_2134,N_2063,N_2072);
and U2135 (N_2135,N_2080,N_2066);
and U2136 (N_2136,N_2086,N_2071);
and U2137 (N_2137,N_2068,N_2077);
or U2138 (N_2138,N_2069,N_2098);
nand U2139 (N_2139,N_2097,N_2050);
nand U2140 (N_2140,N_2064,N_2071);
xnor U2141 (N_2141,N_2070,N_2090);
nand U2142 (N_2142,N_2070,N_2066);
and U2143 (N_2143,N_2052,N_2089);
and U2144 (N_2144,N_2064,N_2059);
and U2145 (N_2145,N_2091,N_2097);
and U2146 (N_2146,N_2088,N_2084);
and U2147 (N_2147,N_2055,N_2070);
nand U2148 (N_2148,N_2073,N_2088);
nor U2149 (N_2149,N_2060,N_2062);
or U2150 (N_2150,N_2108,N_2120);
or U2151 (N_2151,N_2137,N_2135);
nor U2152 (N_2152,N_2114,N_2115);
nand U2153 (N_2153,N_2144,N_2147);
nand U2154 (N_2154,N_2111,N_2128);
nor U2155 (N_2155,N_2103,N_2126);
and U2156 (N_2156,N_2107,N_2101);
or U2157 (N_2157,N_2139,N_2142);
nor U2158 (N_2158,N_2117,N_2146);
xor U2159 (N_2159,N_2118,N_2116);
xor U2160 (N_2160,N_2112,N_2140);
nand U2161 (N_2161,N_2105,N_2121);
and U2162 (N_2162,N_2129,N_2136);
nand U2163 (N_2163,N_2109,N_2134);
nand U2164 (N_2164,N_2100,N_2102);
nand U2165 (N_2165,N_2104,N_2130);
nand U2166 (N_2166,N_2141,N_2125);
and U2167 (N_2167,N_2143,N_2124);
nand U2168 (N_2168,N_2110,N_2127);
and U2169 (N_2169,N_2149,N_2145);
or U2170 (N_2170,N_2113,N_2148);
and U2171 (N_2171,N_2138,N_2119);
or U2172 (N_2172,N_2131,N_2132);
or U2173 (N_2173,N_2106,N_2122);
and U2174 (N_2174,N_2123,N_2133);
and U2175 (N_2175,N_2136,N_2147);
and U2176 (N_2176,N_2141,N_2112);
xor U2177 (N_2177,N_2109,N_2126);
and U2178 (N_2178,N_2146,N_2104);
nand U2179 (N_2179,N_2131,N_2114);
xor U2180 (N_2180,N_2148,N_2128);
nand U2181 (N_2181,N_2131,N_2125);
or U2182 (N_2182,N_2139,N_2116);
or U2183 (N_2183,N_2141,N_2105);
nand U2184 (N_2184,N_2149,N_2125);
or U2185 (N_2185,N_2148,N_2116);
and U2186 (N_2186,N_2115,N_2120);
xor U2187 (N_2187,N_2113,N_2111);
and U2188 (N_2188,N_2149,N_2143);
nand U2189 (N_2189,N_2139,N_2149);
nand U2190 (N_2190,N_2125,N_2105);
nor U2191 (N_2191,N_2113,N_2123);
nor U2192 (N_2192,N_2139,N_2105);
nor U2193 (N_2193,N_2104,N_2143);
nor U2194 (N_2194,N_2117,N_2129);
nor U2195 (N_2195,N_2149,N_2107);
nor U2196 (N_2196,N_2133,N_2139);
or U2197 (N_2197,N_2148,N_2139);
or U2198 (N_2198,N_2144,N_2103);
nand U2199 (N_2199,N_2132,N_2144);
xnor U2200 (N_2200,N_2186,N_2176);
nand U2201 (N_2201,N_2195,N_2166);
and U2202 (N_2202,N_2153,N_2151);
xor U2203 (N_2203,N_2190,N_2185);
and U2204 (N_2204,N_2173,N_2160);
or U2205 (N_2205,N_2158,N_2187);
and U2206 (N_2206,N_2175,N_2199);
nand U2207 (N_2207,N_2150,N_2194);
or U2208 (N_2208,N_2164,N_2197);
nor U2209 (N_2209,N_2172,N_2170);
and U2210 (N_2210,N_2184,N_2189);
and U2211 (N_2211,N_2168,N_2163);
nor U2212 (N_2212,N_2152,N_2161);
nor U2213 (N_2213,N_2183,N_2159);
or U2214 (N_2214,N_2180,N_2196);
or U2215 (N_2215,N_2182,N_2157);
nor U2216 (N_2216,N_2171,N_2167);
and U2217 (N_2217,N_2162,N_2156);
nor U2218 (N_2218,N_2188,N_2154);
or U2219 (N_2219,N_2165,N_2179);
nand U2220 (N_2220,N_2177,N_2198);
and U2221 (N_2221,N_2192,N_2155);
nor U2222 (N_2222,N_2193,N_2181);
or U2223 (N_2223,N_2191,N_2169);
and U2224 (N_2224,N_2178,N_2174);
and U2225 (N_2225,N_2157,N_2165);
nor U2226 (N_2226,N_2199,N_2182);
nand U2227 (N_2227,N_2172,N_2186);
xnor U2228 (N_2228,N_2158,N_2169);
xnor U2229 (N_2229,N_2176,N_2167);
and U2230 (N_2230,N_2175,N_2188);
nand U2231 (N_2231,N_2164,N_2176);
or U2232 (N_2232,N_2190,N_2196);
and U2233 (N_2233,N_2156,N_2179);
and U2234 (N_2234,N_2170,N_2160);
or U2235 (N_2235,N_2158,N_2183);
or U2236 (N_2236,N_2159,N_2170);
nor U2237 (N_2237,N_2168,N_2156);
nor U2238 (N_2238,N_2150,N_2192);
xor U2239 (N_2239,N_2181,N_2160);
xnor U2240 (N_2240,N_2170,N_2192);
nand U2241 (N_2241,N_2196,N_2173);
or U2242 (N_2242,N_2180,N_2194);
nand U2243 (N_2243,N_2197,N_2198);
xnor U2244 (N_2244,N_2186,N_2158);
nor U2245 (N_2245,N_2168,N_2150);
or U2246 (N_2246,N_2152,N_2171);
nand U2247 (N_2247,N_2181,N_2192);
nor U2248 (N_2248,N_2170,N_2169);
nand U2249 (N_2249,N_2162,N_2182);
or U2250 (N_2250,N_2243,N_2247);
nor U2251 (N_2251,N_2249,N_2221);
and U2252 (N_2252,N_2201,N_2244);
and U2253 (N_2253,N_2208,N_2219);
and U2254 (N_2254,N_2225,N_2202);
or U2255 (N_2255,N_2206,N_2241);
and U2256 (N_2256,N_2212,N_2238);
nand U2257 (N_2257,N_2224,N_2245);
and U2258 (N_2258,N_2205,N_2216);
or U2259 (N_2259,N_2236,N_2204);
nor U2260 (N_2260,N_2207,N_2242);
and U2261 (N_2261,N_2234,N_2226);
nand U2262 (N_2262,N_2230,N_2227);
or U2263 (N_2263,N_2213,N_2203);
or U2264 (N_2264,N_2210,N_2217);
or U2265 (N_2265,N_2218,N_2233);
nor U2266 (N_2266,N_2246,N_2223);
and U2267 (N_2267,N_2231,N_2214);
or U2268 (N_2268,N_2211,N_2200);
or U2269 (N_2269,N_2209,N_2215);
or U2270 (N_2270,N_2235,N_2222);
nor U2271 (N_2271,N_2239,N_2228);
and U2272 (N_2272,N_2240,N_2232);
or U2273 (N_2273,N_2229,N_2248);
nor U2274 (N_2274,N_2237,N_2220);
nand U2275 (N_2275,N_2217,N_2230);
and U2276 (N_2276,N_2212,N_2236);
xnor U2277 (N_2277,N_2246,N_2228);
xor U2278 (N_2278,N_2216,N_2227);
nor U2279 (N_2279,N_2205,N_2232);
and U2280 (N_2280,N_2241,N_2201);
nor U2281 (N_2281,N_2241,N_2248);
nand U2282 (N_2282,N_2245,N_2244);
nand U2283 (N_2283,N_2210,N_2220);
nand U2284 (N_2284,N_2221,N_2204);
xnor U2285 (N_2285,N_2230,N_2206);
nand U2286 (N_2286,N_2215,N_2248);
and U2287 (N_2287,N_2205,N_2214);
or U2288 (N_2288,N_2236,N_2220);
nand U2289 (N_2289,N_2232,N_2248);
or U2290 (N_2290,N_2249,N_2233);
nor U2291 (N_2291,N_2232,N_2211);
nand U2292 (N_2292,N_2225,N_2236);
nand U2293 (N_2293,N_2225,N_2246);
nand U2294 (N_2294,N_2225,N_2230);
or U2295 (N_2295,N_2207,N_2204);
nand U2296 (N_2296,N_2221,N_2243);
nand U2297 (N_2297,N_2216,N_2219);
xnor U2298 (N_2298,N_2218,N_2207);
or U2299 (N_2299,N_2203,N_2220);
and U2300 (N_2300,N_2295,N_2258);
nor U2301 (N_2301,N_2262,N_2252);
and U2302 (N_2302,N_2280,N_2255);
nand U2303 (N_2303,N_2267,N_2287);
xor U2304 (N_2304,N_2270,N_2291);
and U2305 (N_2305,N_2286,N_2275);
nand U2306 (N_2306,N_2296,N_2288);
nor U2307 (N_2307,N_2250,N_2294);
nand U2308 (N_2308,N_2274,N_2271);
nand U2309 (N_2309,N_2261,N_2273);
nand U2310 (N_2310,N_2268,N_2251);
nor U2311 (N_2311,N_2297,N_2254);
nand U2312 (N_2312,N_2263,N_2260);
nand U2313 (N_2313,N_2285,N_2299);
nand U2314 (N_2314,N_2278,N_2266);
nand U2315 (N_2315,N_2282,N_2292);
and U2316 (N_2316,N_2277,N_2264);
and U2317 (N_2317,N_2256,N_2298);
or U2318 (N_2318,N_2259,N_2289);
nand U2319 (N_2319,N_2265,N_2283);
and U2320 (N_2320,N_2269,N_2276);
xnor U2321 (N_2321,N_2279,N_2257);
nor U2322 (N_2322,N_2290,N_2284);
and U2323 (N_2323,N_2293,N_2272);
nand U2324 (N_2324,N_2281,N_2253);
and U2325 (N_2325,N_2266,N_2250);
xnor U2326 (N_2326,N_2279,N_2269);
nand U2327 (N_2327,N_2272,N_2286);
or U2328 (N_2328,N_2280,N_2262);
or U2329 (N_2329,N_2270,N_2279);
nor U2330 (N_2330,N_2271,N_2269);
nor U2331 (N_2331,N_2270,N_2285);
or U2332 (N_2332,N_2277,N_2269);
and U2333 (N_2333,N_2292,N_2259);
nor U2334 (N_2334,N_2282,N_2262);
nand U2335 (N_2335,N_2272,N_2291);
or U2336 (N_2336,N_2278,N_2253);
or U2337 (N_2337,N_2298,N_2254);
nand U2338 (N_2338,N_2289,N_2260);
xnor U2339 (N_2339,N_2257,N_2273);
and U2340 (N_2340,N_2278,N_2290);
and U2341 (N_2341,N_2297,N_2256);
and U2342 (N_2342,N_2285,N_2277);
nor U2343 (N_2343,N_2266,N_2256);
or U2344 (N_2344,N_2276,N_2258);
and U2345 (N_2345,N_2267,N_2288);
nor U2346 (N_2346,N_2278,N_2271);
or U2347 (N_2347,N_2274,N_2262);
and U2348 (N_2348,N_2271,N_2268);
nand U2349 (N_2349,N_2286,N_2263);
nor U2350 (N_2350,N_2310,N_2319);
or U2351 (N_2351,N_2324,N_2302);
and U2352 (N_2352,N_2343,N_2316);
nor U2353 (N_2353,N_2336,N_2347);
or U2354 (N_2354,N_2329,N_2333);
nand U2355 (N_2355,N_2304,N_2300);
nand U2356 (N_2356,N_2345,N_2317);
or U2357 (N_2357,N_2301,N_2348);
nand U2358 (N_2358,N_2313,N_2327);
nor U2359 (N_2359,N_2323,N_2339);
nand U2360 (N_2360,N_2306,N_2330);
nand U2361 (N_2361,N_2307,N_2312);
or U2362 (N_2362,N_2337,N_2308);
nand U2363 (N_2363,N_2309,N_2303);
and U2364 (N_2364,N_2318,N_2346);
and U2365 (N_2365,N_2325,N_2322);
and U2366 (N_2366,N_2315,N_2314);
or U2367 (N_2367,N_2338,N_2334);
or U2368 (N_2368,N_2320,N_2326);
and U2369 (N_2369,N_2335,N_2331);
and U2370 (N_2370,N_2328,N_2349);
and U2371 (N_2371,N_2340,N_2305);
nor U2372 (N_2372,N_2311,N_2332);
and U2373 (N_2373,N_2342,N_2321);
nand U2374 (N_2374,N_2344,N_2341);
and U2375 (N_2375,N_2314,N_2305);
and U2376 (N_2376,N_2346,N_2307);
and U2377 (N_2377,N_2335,N_2326);
nand U2378 (N_2378,N_2307,N_2341);
and U2379 (N_2379,N_2341,N_2308);
or U2380 (N_2380,N_2315,N_2301);
xor U2381 (N_2381,N_2305,N_2342);
or U2382 (N_2382,N_2346,N_2335);
xor U2383 (N_2383,N_2335,N_2311);
nand U2384 (N_2384,N_2303,N_2343);
nor U2385 (N_2385,N_2342,N_2337);
and U2386 (N_2386,N_2326,N_2314);
and U2387 (N_2387,N_2322,N_2308);
nor U2388 (N_2388,N_2304,N_2317);
nor U2389 (N_2389,N_2300,N_2306);
nand U2390 (N_2390,N_2327,N_2333);
nor U2391 (N_2391,N_2336,N_2334);
nand U2392 (N_2392,N_2309,N_2315);
and U2393 (N_2393,N_2326,N_2344);
nand U2394 (N_2394,N_2306,N_2333);
xnor U2395 (N_2395,N_2344,N_2304);
or U2396 (N_2396,N_2319,N_2326);
or U2397 (N_2397,N_2322,N_2340);
or U2398 (N_2398,N_2346,N_2328);
xor U2399 (N_2399,N_2322,N_2311);
and U2400 (N_2400,N_2394,N_2383);
nand U2401 (N_2401,N_2354,N_2364);
and U2402 (N_2402,N_2372,N_2356);
nand U2403 (N_2403,N_2393,N_2382);
or U2404 (N_2404,N_2353,N_2385);
xor U2405 (N_2405,N_2380,N_2370);
or U2406 (N_2406,N_2389,N_2392);
xnor U2407 (N_2407,N_2352,N_2398);
nand U2408 (N_2408,N_2390,N_2366);
nor U2409 (N_2409,N_2360,N_2362);
or U2410 (N_2410,N_2367,N_2384);
nor U2411 (N_2411,N_2388,N_2395);
and U2412 (N_2412,N_2358,N_2386);
nand U2413 (N_2413,N_2377,N_2361);
and U2414 (N_2414,N_2368,N_2379);
nand U2415 (N_2415,N_2397,N_2399);
xnor U2416 (N_2416,N_2387,N_2351);
nand U2417 (N_2417,N_2371,N_2350);
or U2418 (N_2418,N_2381,N_2376);
nand U2419 (N_2419,N_2373,N_2355);
nand U2420 (N_2420,N_2378,N_2375);
or U2421 (N_2421,N_2365,N_2359);
nor U2422 (N_2422,N_2363,N_2396);
xnor U2423 (N_2423,N_2369,N_2391);
or U2424 (N_2424,N_2357,N_2374);
or U2425 (N_2425,N_2392,N_2365);
nor U2426 (N_2426,N_2378,N_2395);
nor U2427 (N_2427,N_2389,N_2397);
or U2428 (N_2428,N_2365,N_2397);
nand U2429 (N_2429,N_2353,N_2386);
and U2430 (N_2430,N_2381,N_2358);
nand U2431 (N_2431,N_2387,N_2398);
nand U2432 (N_2432,N_2383,N_2390);
and U2433 (N_2433,N_2359,N_2350);
nor U2434 (N_2434,N_2359,N_2354);
nand U2435 (N_2435,N_2351,N_2377);
or U2436 (N_2436,N_2358,N_2361);
nand U2437 (N_2437,N_2377,N_2398);
and U2438 (N_2438,N_2352,N_2399);
or U2439 (N_2439,N_2352,N_2383);
and U2440 (N_2440,N_2378,N_2376);
nor U2441 (N_2441,N_2397,N_2378);
or U2442 (N_2442,N_2389,N_2391);
and U2443 (N_2443,N_2367,N_2377);
or U2444 (N_2444,N_2362,N_2361);
nor U2445 (N_2445,N_2373,N_2385);
and U2446 (N_2446,N_2351,N_2378);
and U2447 (N_2447,N_2362,N_2381);
nor U2448 (N_2448,N_2364,N_2392);
and U2449 (N_2449,N_2355,N_2397);
nor U2450 (N_2450,N_2418,N_2402);
and U2451 (N_2451,N_2419,N_2400);
nor U2452 (N_2452,N_2435,N_2426);
or U2453 (N_2453,N_2440,N_2442);
nor U2454 (N_2454,N_2445,N_2408);
nor U2455 (N_2455,N_2414,N_2449);
nor U2456 (N_2456,N_2444,N_2403);
nor U2457 (N_2457,N_2431,N_2446);
and U2458 (N_2458,N_2406,N_2429);
nand U2459 (N_2459,N_2427,N_2411);
nand U2460 (N_2460,N_2439,N_2422);
nand U2461 (N_2461,N_2447,N_2430);
xnor U2462 (N_2462,N_2415,N_2434);
and U2463 (N_2463,N_2416,N_2433);
or U2464 (N_2464,N_2441,N_2413);
nor U2465 (N_2465,N_2405,N_2437);
xor U2466 (N_2466,N_2407,N_2409);
and U2467 (N_2467,N_2412,N_2423);
xor U2468 (N_2468,N_2428,N_2410);
nor U2469 (N_2469,N_2448,N_2424);
nor U2470 (N_2470,N_2417,N_2401);
or U2471 (N_2471,N_2432,N_2438);
and U2472 (N_2472,N_2421,N_2443);
nand U2473 (N_2473,N_2436,N_2425);
or U2474 (N_2474,N_2404,N_2420);
nand U2475 (N_2475,N_2406,N_2443);
nor U2476 (N_2476,N_2440,N_2436);
xor U2477 (N_2477,N_2433,N_2435);
nand U2478 (N_2478,N_2410,N_2433);
and U2479 (N_2479,N_2433,N_2446);
or U2480 (N_2480,N_2417,N_2427);
or U2481 (N_2481,N_2430,N_2407);
and U2482 (N_2482,N_2445,N_2440);
nor U2483 (N_2483,N_2404,N_2434);
and U2484 (N_2484,N_2449,N_2424);
and U2485 (N_2485,N_2410,N_2435);
or U2486 (N_2486,N_2438,N_2435);
or U2487 (N_2487,N_2410,N_2447);
xnor U2488 (N_2488,N_2446,N_2449);
nand U2489 (N_2489,N_2443,N_2426);
and U2490 (N_2490,N_2408,N_2417);
or U2491 (N_2491,N_2437,N_2442);
nor U2492 (N_2492,N_2425,N_2405);
nand U2493 (N_2493,N_2405,N_2432);
xor U2494 (N_2494,N_2409,N_2449);
or U2495 (N_2495,N_2421,N_2406);
nand U2496 (N_2496,N_2406,N_2400);
or U2497 (N_2497,N_2422,N_2428);
nand U2498 (N_2498,N_2447,N_2412);
nor U2499 (N_2499,N_2411,N_2438);
and U2500 (N_2500,N_2486,N_2471);
nor U2501 (N_2501,N_2463,N_2498);
or U2502 (N_2502,N_2473,N_2472);
and U2503 (N_2503,N_2462,N_2455);
nor U2504 (N_2504,N_2450,N_2457);
nand U2505 (N_2505,N_2496,N_2451);
nor U2506 (N_2506,N_2465,N_2468);
or U2507 (N_2507,N_2477,N_2460);
and U2508 (N_2508,N_2485,N_2474);
and U2509 (N_2509,N_2492,N_2481);
nor U2510 (N_2510,N_2453,N_2464);
nor U2511 (N_2511,N_2478,N_2452);
nor U2512 (N_2512,N_2475,N_2497);
and U2513 (N_2513,N_2470,N_2479);
or U2514 (N_2514,N_2458,N_2484);
xor U2515 (N_2515,N_2480,N_2490);
or U2516 (N_2516,N_2454,N_2483);
and U2517 (N_2517,N_2467,N_2487);
or U2518 (N_2518,N_2456,N_2499);
or U2519 (N_2519,N_2459,N_2493);
nand U2520 (N_2520,N_2466,N_2488);
xnor U2521 (N_2521,N_2461,N_2469);
or U2522 (N_2522,N_2495,N_2482);
nor U2523 (N_2523,N_2489,N_2494);
nor U2524 (N_2524,N_2476,N_2491);
and U2525 (N_2525,N_2478,N_2477);
and U2526 (N_2526,N_2452,N_2455);
nand U2527 (N_2527,N_2473,N_2474);
nor U2528 (N_2528,N_2473,N_2493);
nand U2529 (N_2529,N_2452,N_2473);
and U2530 (N_2530,N_2470,N_2481);
nor U2531 (N_2531,N_2480,N_2476);
nand U2532 (N_2532,N_2450,N_2459);
xnor U2533 (N_2533,N_2462,N_2495);
and U2534 (N_2534,N_2457,N_2495);
nor U2535 (N_2535,N_2492,N_2487);
nor U2536 (N_2536,N_2478,N_2495);
or U2537 (N_2537,N_2465,N_2494);
or U2538 (N_2538,N_2469,N_2459);
or U2539 (N_2539,N_2476,N_2489);
and U2540 (N_2540,N_2490,N_2486);
or U2541 (N_2541,N_2479,N_2487);
or U2542 (N_2542,N_2453,N_2459);
or U2543 (N_2543,N_2492,N_2455);
xnor U2544 (N_2544,N_2464,N_2473);
and U2545 (N_2545,N_2487,N_2478);
xor U2546 (N_2546,N_2485,N_2484);
nand U2547 (N_2547,N_2488,N_2493);
nand U2548 (N_2548,N_2483,N_2459);
nor U2549 (N_2549,N_2478,N_2472);
or U2550 (N_2550,N_2540,N_2547);
nor U2551 (N_2551,N_2517,N_2533);
and U2552 (N_2552,N_2509,N_2506);
or U2553 (N_2553,N_2516,N_2548);
or U2554 (N_2554,N_2546,N_2528);
nor U2555 (N_2555,N_2500,N_2519);
nand U2556 (N_2556,N_2527,N_2523);
nor U2557 (N_2557,N_2542,N_2545);
nand U2558 (N_2558,N_2525,N_2539);
and U2559 (N_2559,N_2504,N_2502);
or U2560 (N_2560,N_2510,N_2524);
nor U2561 (N_2561,N_2530,N_2536);
and U2562 (N_2562,N_2515,N_2529);
nand U2563 (N_2563,N_2543,N_2513);
nor U2564 (N_2564,N_2549,N_2501);
and U2565 (N_2565,N_2520,N_2503);
xor U2566 (N_2566,N_2508,N_2531);
and U2567 (N_2567,N_2507,N_2537);
nor U2568 (N_2568,N_2521,N_2512);
xnor U2569 (N_2569,N_2522,N_2514);
nand U2570 (N_2570,N_2544,N_2538);
and U2571 (N_2571,N_2534,N_2535);
nand U2572 (N_2572,N_2532,N_2511);
nand U2573 (N_2573,N_2518,N_2526);
nand U2574 (N_2574,N_2505,N_2541);
nand U2575 (N_2575,N_2532,N_2507);
nand U2576 (N_2576,N_2510,N_2531);
or U2577 (N_2577,N_2548,N_2530);
nand U2578 (N_2578,N_2518,N_2535);
and U2579 (N_2579,N_2515,N_2523);
and U2580 (N_2580,N_2526,N_2530);
and U2581 (N_2581,N_2528,N_2505);
or U2582 (N_2582,N_2523,N_2518);
nor U2583 (N_2583,N_2539,N_2531);
nand U2584 (N_2584,N_2536,N_2539);
xor U2585 (N_2585,N_2529,N_2533);
and U2586 (N_2586,N_2515,N_2535);
nand U2587 (N_2587,N_2548,N_2542);
nor U2588 (N_2588,N_2500,N_2534);
xor U2589 (N_2589,N_2502,N_2542);
and U2590 (N_2590,N_2538,N_2530);
and U2591 (N_2591,N_2506,N_2511);
or U2592 (N_2592,N_2515,N_2541);
nand U2593 (N_2593,N_2502,N_2539);
nor U2594 (N_2594,N_2522,N_2501);
nand U2595 (N_2595,N_2510,N_2502);
xnor U2596 (N_2596,N_2506,N_2528);
xor U2597 (N_2597,N_2546,N_2511);
nand U2598 (N_2598,N_2518,N_2515);
and U2599 (N_2599,N_2508,N_2518);
nand U2600 (N_2600,N_2592,N_2593);
nand U2601 (N_2601,N_2558,N_2594);
nor U2602 (N_2602,N_2553,N_2557);
or U2603 (N_2603,N_2582,N_2555);
nor U2604 (N_2604,N_2571,N_2570);
nand U2605 (N_2605,N_2573,N_2581);
nand U2606 (N_2606,N_2598,N_2597);
nor U2607 (N_2607,N_2551,N_2595);
or U2608 (N_2608,N_2561,N_2572);
nor U2609 (N_2609,N_2585,N_2559);
nand U2610 (N_2610,N_2591,N_2563);
or U2611 (N_2611,N_2584,N_2596);
nand U2612 (N_2612,N_2589,N_2568);
and U2613 (N_2613,N_2586,N_2554);
or U2614 (N_2614,N_2560,N_2580);
and U2615 (N_2615,N_2587,N_2566);
nor U2616 (N_2616,N_2588,N_2583);
xor U2617 (N_2617,N_2556,N_2599);
or U2618 (N_2618,N_2577,N_2567);
nor U2619 (N_2619,N_2590,N_2575);
or U2620 (N_2620,N_2578,N_2550);
xnor U2621 (N_2621,N_2579,N_2562);
and U2622 (N_2622,N_2565,N_2564);
nand U2623 (N_2623,N_2552,N_2569);
nand U2624 (N_2624,N_2576,N_2574);
or U2625 (N_2625,N_2585,N_2569);
or U2626 (N_2626,N_2591,N_2561);
nor U2627 (N_2627,N_2574,N_2593);
nand U2628 (N_2628,N_2573,N_2568);
nand U2629 (N_2629,N_2591,N_2577);
xnor U2630 (N_2630,N_2569,N_2557);
xor U2631 (N_2631,N_2586,N_2580);
and U2632 (N_2632,N_2561,N_2589);
nand U2633 (N_2633,N_2590,N_2591);
or U2634 (N_2634,N_2557,N_2578);
nand U2635 (N_2635,N_2580,N_2571);
and U2636 (N_2636,N_2574,N_2591);
nor U2637 (N_2637,N_2584,N_2568);
or U2638 (N_2638,N_2570,N_2562);
or U2639 (N_2639,N_2570,N_2555);
or U2640 (N_2640,N_2550,N_2563);
and U2641 (N_2641,N_2597,N_2596);
nand U2642 (N_2642,N_2577,N_2580);
nor U2643 (N_2643,N_2575,N_2580);
or U2644 (N_2644,N_2571,N_2593);
or U2645 (N_2645,N_2567,N_2556);
nand U2646 (N_2646,N_2590,N_2568);
or U2647 (N_2647,N_2596,N_2592);
and U2648 (N_2648,N_2578,N_2567);
or U2649 (N_2649,N_2573,N_2572);
or U2650 (N_2650,N_2647,N_2615);
xnor U2651 (N_2651,N_2624,N_2607);
or U2652 (N_2652,N_2612,N_2622);
and U2653 (N_2653,N_2630,N_2645);
nand U2654 (N_2654,N_2603,N_2601);
or U2655 (N_2655,N_2641,N_2649);
nor U2656 (N_2656,N_2637,N_2643);
nand U2657 (N_2657,N_2626,N_2602);
or U2658 (N_2658,N_2605,N_2617);
nor U2659 (N_2659,N_2631,N_2638);
nor U2660 (N_2660,N_2633,N_2610);
and U2661 (N_2661,N_2616,N_2648);
nand U2662 (N_2662,N_2639,N_2609);
nor U2663 (N_2663,N_2635,N_2642);
nor U2664 (N_2664,N_2627,N_2618);
or U2665 (N_2665,N_2606,N_2625);
nor U2666 (N_2666,N_2608,N_2614);
or U2667 (N_2667,N_2621,N_2619);
and U2668 (N_2668,N_2646,N_2620);
xor U2669 (N_2669,N_2604,N_2613);
or U2670 (N_2670,N_2629,N_2600);
and U2671 (N_2671,N_2636,N_2634);
or U2672 (N_2672,N_2623,N_2611);
nor U2673 (N_2673,N_2644,N_2628);
and U2674 (N_2674,N_2632,N_2640);
and U2675 (N_2675,N_2601,N_2622);
nand U2676 (N_2676,N_2619,N_2628);
nand U2677 (N_2677,N_2636,N_2638);
and U2678 (N_2678,N_2616,N_2613);
nand U2679 (N_2679,N_2626,N_2615);
nand U2680 (N_2680,N_2610,N_2645);
xnor U2681 (N_2681,N_2633,N_2627);
and U2682 (N_2682,N_2644,N_2648);
nand U2683 (N_2683,N_2619,N_2633);
nand U2684 (N_2684,N_2632,N_2643);
nand U2685 (N_2685,N_2606,N_2617);
and U2686 (N_2686,N_2622,N_2605);
nor U2687 (N_2687,N_2644,N_2604);
nand U2688 (N_2688,N_2645,N_2616);
and U2689 (N_2689,N_2632,N_2644);
nor U2690 (N_2690,N_2600,N_2645);
and U2691 (N_2691,N_2634,N_2622);
nand U2692 (N_2692,N_2630,N_2640);
nand U2693 (N_2693,N_2637,N_2615);
and U2694 (N_2694,N_2639,N_2617);
nor U2695 (N_2695,N_2634,N_2610);
or U2696 (N_2696,N_2623,N_2636);
or U2697 (N_2697,N_2626,N_2634);
or U2698 (N_2698,N_2648,N_2619);
and U2699 (N_2699,N_2625,N_2607);
nand U2700 (N_2700,N_2667,N_2688);
or U2701 (N_2701,N_2650,N_2691);
xor U2702 (N_2702,N_2656,N_2659);
nor U2703 (N_2703,N_2697,N_2664);
nor U2704 (N_2704,N_2696,N_2679);
and U2705 (N_2705,N_2660,N_2694);
or U2706 (N_2706,N_2680,N_2665);
nor U2707 (N_2707,N_2678,N_2689);
and U2708 (N_2708,N_2686,N_2658);
nand U2709 (N_2709,N_2666,N_2693);
nand U2710 (N_2710,N_2655,N_2699);
or U2711 (N_2711,N_2692,N_2681);
and U2712 (N_2712,N_2651,N_2683);
xnor U2713 (N_2713,N_2661,N_2698);
or U2714 (N_2714,N_2695,N_2673);
xnor U2715 (N_2715,N_2663,N_2657);
nand U2716 (N_2716,N_2671,N_2672);
and U2717 (N_2717,N_2669,N_2662);
or U2718 (N_2718,N_2654,N_2668);
nand U2719 (N_2719,N_2687,N_2682);
and U2720 (N_2720,N_2684,N_2675);
xor U2721 (N_2721,N_2670,N_2674);
or U2722 (N_2722,N_2677,N_2676);
or U2723 (N_2723,N_2685,N_2690);
nand U2724 (N_2724,N_2653,N_2652);
or U2725 (N_2725,N_2660,N_2670);
and U2726 (N_2726,N_2674,N_2694);
xnor U2727 (N_2727,N_2695,N_2681);
or U2728 (N_2728,N_2685,N_2669);
and U2729 (N_2729,N_2652,N_2691);
nand U2730 (N_2730,N_2688,N_2689);
and U2731 (N_2731,N_2654,N_2662);
nor U2732 (N_2732,N_2662,N_2678);
nor U2733 (N_2733,N_2661,N_2665);
nor U2734 (N_2734,N_2697,N_2654);
or U2735 (N_2735,N_2689,N_2672);
nor U2736 (N_2736,N_2662,N_2660);
nand U2737 (N_2737,N_2661,N_2654);
xor U2738 (N_2738,N_2691,N_2676);
nor U2739 (N_2739,N_2657,N_2653);
nand U2740 (N_2740,N_2684,N_2686);
nor U2741 (N_2741,N_2662,N_2650);
or U2742 (N_2742,N_2678,N_2687);
nor U2743 (N_2743,N_2675,N_2662);
or U2744 (N_2744,N_2667,N_2653);
nand U2745 (N_2745,N_2694,N_2653);
or U2746 (N_2746,N_2660,N_2680);
nor U2747 (N_2747,N_2681,N_2698);
or U2748 (N_2748,N_2697,N_2677);
nor U2749 (N_2749,N_2698,N_2663);
nand U2750 (N_2750,N_2730,N_2722);
nand U2751 (N_2751,N_2742,N_2728);
or U2752 (N_2752,N_2734,N_2741);
or U2753 (N_2753,N_2713,N_2708);
and U2754 (N_2754,N_2743,N_2738);
nand U2755 (N_2755,N_2737,N_2716);
or U2756 (N_2756,N_2702,N_2749);
and U2757 (N_2757,N_2706,N_2707);
nor U2758 (N_2758,N_2703,N_2748);
xor U2759 (N_2759,N_2725,N_2735);
and U2760 (N_2760,N_2726,N_2731);
or U2761 (N_2761,N_2744,N_2732);
and U2762 (N_2762,N_2746,N_2739);
or U2763 (N_2763,N_2714,N_2704);
nand U2764 (N_2764,N_2724,N_2740);
or U2765 (N_2765,N_2719,N_2717);
and U2766 (N_2766,N_2715,N_2723);
nor U2767 (N_2767,N_2701,N_2711);
and U2768 (N_2768,N_2720,N_2721);
or U2769 (N_2769,N_2705,N_2709);
nor U2770 (N_2770,N_2718,N_2729);
xor U2771 (N_2771,N_2747,N_2712);
nor U2772 (N_2772,N_2700,N_2736);
xnor U2773 (N_2773,N_2733,N_2710);
nor U2774 (N_2774,N_2745,N_2727);
nor U2775 (N_2775,N_2708,N_2721);
nor U2776 (N_2776,N_2743,N_2713);
nor U2777 (N_2777,N_2718,N_2728);
and U2778 (N_2778,N_2737,N_2723);
and U2779 (N_2779,N_2726,N_2721);
nand U2780 (N_2780,N_2732,N_2709);
or U2781 (N_2781,N_2705,N_2727);
nor U2782 (N_2782,N_2714,N_2735);
nand U2783 (N_2783,N_2703,N_2741);
nor U2784 (N_2784,N_2738,N_2725);
and U2785 (N_2785,N_2701,N_2726);
and U2786 (N_2786,N_2740,N_2701);
or U2787 (N_2787,N_2719,N_2721);
and U2788 (N_2788,N_2742,N_2730);
nand U2789 (N_2789,N_2744,N_2719);
nor U2790 (N_2790,N_2727,N_2714);
and U2791 (N_2791,N_2736,N_2728);
and U2792 (N_2792,N_2733,N_2715);
nand U2793 (N_2793,N_2733,N_2707);
nand U2794 (N_2794,N_2737,N_2707);
nor U2795 (N_2795,N_2736,N_2742);
or U2796 (N_2796,N_2725,N_2730);
and U2797 (N_2797,N_2706,N_2701);
or U2798 (N_2798,N_2700,N_2747);
or U2799 (N_2799,N_2732,N_2721);
nor U2800 (N_2800,N_2799,N_2779);
or U2801 (N_2801,N_2788,N_2774);
or U2802 (N_2802,N_2798,N_2791);
nand U2803 (N_2803,N_2793,N_2760);
nor U2804 (N_2804,N_2750,N_2766);
and U2805 (N_2805,N_2768,N_2780);
and U2806 (N_2806,N_2759,N_2755);
or U2807 (N_2807,N_2795,N_2758);
nand U2808 (N_2808,N_2762,N_2751);
or U2809 (N_2809,N_2773,N_2790);
or U2810 (N_2810,N_2778,N_2781);
nand U2811 (N_2811,N_2777,N_2783);
xor U2812 (N_2812,N_2789,N_2792);
nor U2813 (N_2813,N_2782,N_2752);
xnor U2814 (N_2814,N_2765,N_2796);
nor U2815 (N_2815,N_2785,N_2775);
xnor U2816 (N_2816,N_2786,N_2770);
xor U2817 (N_2817,N_2784,N_2772);
and U2818 (N_2818,N_2771,N_2754);
and U2819 (N_2819,N_2767,N_2787);
nor U2820 (N_2820,N_2756,N_2753);
nor U2821 (N_2821,N_2797,N_2764);
nor U2822 (N_2822,N_2763,N_2794);
and U2823 (N_2823,N_2757,N_2761);
or U2824 (N_2824,N_2776,N_2769);
and U2825 (N_2825,N_2752,N_2767);
and U2826 (N_2826,N_2752,N_2769);
and U2827 (N_2827,N_2776,N_2785);
nand U2828 (N_2828,N_2754,N_2759);
and U2829 (N_2829,N_2765,N_2767);
xnor U2830 (N_2830,N_2785,N_2798);
nor U2831 (N_2831,N_2767,N_2753);
or U2832 (N_2832,N_2772,N_2754);
xor U2833 (N_2833,N_2789,N_2791);
xor U2834 (N_2834,N_2795,N_2793);
and U2835 (N_2835,N_2780,N_2750);
and U2836 (N_2836,N_2796,N_2786);
nand U2837 (N_2837,N_2793,N_2763);
nor U2838 (N_2838,N_2767,N_2793);
nor U2839 (N_2839,N_2751,N_2774);
or U2840 (N_2840,N_2774,N_2786);
nand U2841 (N_2841,N_2775,N_2771);
and U2842 (N_2842,N_2792,N_2797);
xnor U2843 (N_2843,N_2795,N_2785);
or U2844 (N_2844,N_2775,N_2774);
nand U2845 (N_2845,N_2786,N_2762);
nand U2846 (N_2846,N_2757,N_2799);
nand U2847 (N_2847,N_2779,N_2764);
nor U2848 (N_2848,N_2787,N_2753);
and U2849 (N_2849,N_2778,N_2786);
nand U2850 (N_2850,N_2810,N_2811);
nand U2851 (N_2851,N_2816,N_2821);
or U2852 (N_2852,N_2819,N_2831);
and U2853 (N_2853,N_2833,N_2820);
or U2854 (N_2854,N_2823,N_2803);
nor U2855 (N_2855,N_2838,N_2801);
nor U2856 (N_2856,N_2836,N_2818);
or U2857 (N_2857,N_2802,N_2849);
nor U2858 (N_2858,N_2835,N_2812);
nand U2859 (N_2859,N_2817,N_2805);
and U2860 (N_2860,N_2824,N_2845);
nand U2861 (N_2861,N_2830,N_2846);
nand U2862 (N_2862,N_2815,N_2829);
nor U2863 (N_2863,N_2800,N_2848);
or U2864 (N_2864,N_2809,N_2837);
nor U2865 (N_2865,N_2844,N_2826);
nor U2866 (N_2866,N_2808,N_2822);
and U2867 (N_2867,N_2839,N_2841);
nor U2868 (N_2868,N_2840,N_2807);
xnor U2869 (N_2869,N_2825,N_2843);
nor U2870 (N_2870,N_2814,N_2828);
or U2871 (N_2871,N_2847,N_2827);
xor U2872 (N_2872,N_2813,N_2842);
and U2873 (N_2873,N_2804,N_2834);
nand U2874 (N_2874,N_2806,N_2832);
or U2875 (N_2875,N_2803,N_2800);
nand U2876 (N_2876,N_2802,N_2806);
nand U2877 (N_2877,N_2816,N_2842);
nand U2878 (N_2878,N_2807,N_2819);
nor U2879 (N_2879,N_2820,N_2814);
xor U2880 (N_2880,N_2816,N_2832);
nand U2881 (N_2881,N_2807,N_2844);
nand U2882 (N_2882,N_2823,N_2846);
nor U2883 (N_2883,N_2835,N_2807);
nor U2884 (N_2884,N_2808,N_2801);
nand U2885 (N_2885,N_2814,N_2819);
nand U2886 (N_2886,N_2841,N_2815);
nor U2887 (N_2887,N_2819,N_2832);
and U2888 (N_2888,N_2833,N_2815);
nor U2889 (N_2889,N_2836,N_2846);
nor U2890 (N_2890,N_2840,N_2811);
nor U2891 (N_2891,N_2845,N_2800);
xnor U2892 (N_2892,N_2836,N_2845);
or U2893 (N_2893,N_2801,N_2841);
nand U2894 (N_2894,N_2821,N_2827);
and U2895 (N_2895,N_2800,N_2849);
or U2896 (N_2896,N_2813,N_2801);
or U2897 (N_2897,N_2816,N_2822);
xnor U2898 (N_2898,N_2802,N_2801);
and U2899 (N_2899,N_2804,N_2807);
nor U2900 (N_2900,N_2863,N_2894);
or U2901 (N_2901,N_2872,N_2855);
nor U2902 (N_2902,N_2893,N_2852);
or U2903 (N_2903,N_2876,N_2895);
xnor U2904 (N_2904,N_2862,N_2864);
and U2905 (N_2905,N_2897,N_2881);
and U2906 (N_2906,N_2880,N_2853);
nand U2907 (N_2907,N_2851,N_2857);
nor U2908 (N_2908,N_2882,N_2885);
and U2909 (N_2909,N_2890,N_2892);
nand U2910 (N_2910,N_2854,N_2883);
or U2911 (N_2911,N_2859,N_2875);
or U2912 (N_2912,N_2856,N_2896);
or U2913 (N_2913,N_2887,N_2871);
and U2914 (N_2914,N_2858,N_2899);
nor U2915 (N_2915,N_2886,N_2874);
nand U2916 (N_2916,N_2866,N_2868);
nand U2917 (N_2917,N_2891,N_2869);
nand U2918 (N_2918,N_2867,N_2861);
and U2919 (N_2919,N_2878,N_2884);
and U2920 (N_2920,N_2850,N_2879);
nor U2921 (N_2921,N_2865,N_2889);
and U2922 (N_2922,N_2873,N_2888);
xnor U2923 (N_2923,N_2898,N_2860);
nand U2924 (N_2924,N_2877,N_2870);
or U2925 (N_2925,N_2896,N_2851);
xnor U2926 (N_2926,N_2889,N_2857);
nand U2927 (N_2927,N_2871,N_2864);
or U2928 (N_2928,N_2854,N_2853);
nand U2929 (N_2929,N_2874,N_2854);
and U2930 (N_2930,N_2872,N_2886);
or U2931 (N_2931,N_2881,N_2894);
and U2932 (N_2932,N_2899,N_2884);
nand U2933 (N_2933,N_2861,N_2881);
or U2934 (N_2934,N_2858,N_2891);
nor U2935 (N_2935,N_2898,N_2862);
or U2936 (N_2936,N_2893,N_2860);
and U2937 (N_2937,N_2870,N_2865);
and U2938 (N_2938,N_2880,N_2897);
or U2939 (N_2939,N_2892,N_2861);
nand U2940 (N_2940,N_2859,N_2894);
nand U2941 (N_2941,N_2858,N_2887);
nand U2942 (N_2942,N_2897,N_2873);
nor U2943 (N_2943,N_2859,N_2854);
or U2944 (N_2944,N_2865,N_2858);
nand U2945 (N_2945,N_2850,N_2854);
nor U2946 (N_2946,N_2894,N_2891);
and U2947 (N_2947,N_2857,N_2855);
nand U2948 (N_2948,N_2870,N_2851);
nand U2949 (N_2949,N_2882,N_2857);
and U2950 (N_2950,N_2949,N_2931);
and U2951 (N_2951,N_2947,N_2911);
nor U2952 (N_2952,N_2934,N_2904);
or U2953 (N_2953,N_2940,N_2939);
nor U2954 (N_2954,N_2943,N_2928);
nor U2955 (N_2955,N_2945,N_2908);
nor U2956 (N_2956,N_2900,N_2913);
nor U2957 (N_2957,N_2935,N_2941);
or U2958 (N_2958,N_2917,N_2910);
nor U2959 (N_2959,N_2902,N_2912);
xor U2960 (N_2960,N_2905,N_2901);
nor U2961 (N_2961,N_2937,N_2942);
nand U2962 (N_2962,N_2948,N_2933);
nand U2963 (N_2963,N_2938,N_2946);
and U2964 (N_2964,N_2944,N_2927);
nor U2965 (N_2965,N_2932,N_2921);
or U2966 (N_2966,N_2918,N_2936);
and U2967 (N_2967,N_2926,N_2919);
and U2968 (N_2968,N_2909,N_2906);
nor U2969 (N_2969,N_2903,N_2929);
nand U2970 (N_2970,N_2916,N_2915);
or U2971 (N_2971,N_2920,N_2922);
nor U2972 (N_2972,N_2907,N_2923);
nand U2973 (N_2973,N_2924,N_2930);
nor U2974 (N_2974,N_2914,N_2925);
nor U2975 (N_2975,N_2900,N_2940);
nand U2976 (N_2976,N_2912,N_2900);
nand U2977 (N_2977,N_2938,N_2908);
xor U2978 (N_2978,N_2901,N_2903);
or U2979 (N_2979,N_2907,N_2900);
xor U2980 (N_2980,N_2949,N_2916);
and U2981 (N_2981,N_2948,N_2932);
and U2982 (N_2982,N_2909,N_2947);
xnor U2983 (N_2983,N_2930,N_2948);
and U2984 (N_2984,N_2932,N_2910);
or U2985 (N_2985,N_2940,N_2947);
nand U2986 (N_2986,N_2913,N_2907);
nor U2987 (N_2987,N_2928,N_2916);
nand U2988 (N_2988,N_2922,N_2936);
nor U2989 (N_2989,N_2932,N_2935);
or U2990 (N_2990,N_2932,N_2909);
nand U2991 (N_2991,N_2948,N_2946);
nor U2992 (N_2992,N_2909,N_2937);
and U2993 (N_2993,N_2903,N_2927);
nand U2994 (N_2994,N_2943,N_2931);
xor U2995 (N_2995,N_2907,N_2924);
nand U2996 (N_2996,N_2930,N_2927);
nor U2997 (N_2997,N_2926,N_2900);
nor U2998 (N_2998,N_2915,N_2918);
nand U2999 (N_2999,N_2923,N_2924);
nand UO_0 (O_0,N_2988,N_2979);
or UO_1 (O_1,N_2994,N_2968);
nand UO_2 (O_2,N_2996,N_2954);
and UO_3 (O_3,N_2974,N_2973);
and UO_4 (O_4,N_2986,N_2984);
and UO_5 (O_5,N_2990,N_2961);
nor UO_6 (O_6,N_2971,N_2951);
and UO_7 (O_7,N_2956,N_2965);
nand UO_8 (O_8,N_2959,N_2982);
nor UO_9 (O_9,N_2983,N_2963);
nand UO_10 (O_10,N_2952,N_2972);
or UO_11 (O_11,N_2970,N_2975);
nand UO_12 (O_12,N_2950,N_2999);
nand UO_13 (O_13,N_2992,N_2967);
nand UO_14 (O_14,N_2955,N_2981);
and UO_15 (O_15,N_2969,N_2993);
nand UO_16 (O_16,N_2997,N_2957);
nor UO_17 (O_17,N_2962,N_2995);
or UO_18 (O_18,N_2958,N_2998);
and UO_19 (O_19,N_2953,N_2985);
and UO_20 (O_20,N_2989,N_2964);
and UO_21 (O_21,N_2987,N_2960);
or UO_22 (O_22,N_2978,N_2980);
nand UO_23 (O_23,N_2976,N_2991);
and UO_24 (O_24,N_2966,N_2977);
and UO_25 (O_25,N_2973,N_2958);
nor UO_26 (O_26,N_2980,N_2970);
nor UO_27 (O_27,N_2973,N_2950);
nor UO_28 (O_28,N_2997,N_2983);
and UO_29 (O_29,N_2966,N_2965);
and UO_30 (O_30,N_2997,N_2987);
nand UO_31 (O_31,N_2960,N_2984);
or UO_32 (O_32,N_2976,N_2962);
xor UO_33 (O_33,N_2977,N_2968);
or UO_34 (O_34,N_2969,N_2981);
nand UO_35 (O_35,N_2981,N_2958);
xor UO_36 (O_36,N_2967,N_2955);
nor UO_37 (O_37,N_2952,N_2962);
or UO_38 (O_38,N_2997,N_2974);
or UO_39 (O_39,N_2999,N_2988);
nand UO_40 (O_40,N_2955,N_2959);
and UO_41 (O_41,N_2992,N_2956);
nor UO_42 (O_42,N_2981,N_2968);
nor UO_43 (O_43,N_2954,N_2965);
or UO_44 (O_44,N_2957,N_2952);
nor UO_45 (O_45,N_2991,N_2960);
nor UO_46 (O_46,N_2977,N_2970);
and UO_47 (O_47,N_2997,N_2961);
and UO_48 (O_48,N_2977,N_2974);
nor UO_49 (O_49,N_2991,N_2985);
or UO_50 (O_50,N_2963,N_2967);
and UO_51 (O_51,N_2967,N_2991);
nand UO_52 (O_52,N_2963,N_2975);
nor UO_53 (O_53,N_2968,N_2952);
or UO_54 (O_54,N_2979,N_2998);
or UO_55 (O_55,N_2985,N_2978);
nor UO_56 (O_56,N_2967,N_2972);
and UO_57 (O_57,N_2965,N_2989);
and UO_58 (O_58,N_2956,N_2988);
nor UO_59 (O_59,N_2994,N_2955);
and UO_60 (O_60,N_2978,N_2953);
xor UO_61 (O_61,N_2982,N_2995);
nor UO_62 (O_62,N_2979,N_2959);
xor UO_63 (O_63,N_2999,N_2951);
xor UO_64 (O_64,N_2969,N_2952);
and UO_65 (O_65,N_2966,N_2964);
or UO_66 (O_66,N_2965,N_2978);
nand UO_67 (O_67,N_2960,N_2979);
nor UO_68 (O_68,N_2958,N_2995);
nand UO_69 (O_69,N_2953,N_2974);
nor UO_70 (O_70,N_2952,N_2963);
nor UO_71 (O_71,N_2988,N_2987);
xnor UO_72 (O_72,N_2993,N_2984);
nand UO_73 (O_73,N_2980,N_2963);
nor UO_74 (O_74,N_2998,N_2997);
nand UO_75 (O_75,N_2990,N_2974);
or UO_76 (O_76,N_2991,N_2984);
nand UO_77 (O_77,N_2983,N_2956);
or UO_78 (O_78,N_2990,N_2992);
and UO_79 (O_79,N_2963,N_2955);
nand UO_80 (O_80,N_2983,N_2984);
nor UO_81 (O_81,N_2993,N_2957);
and UO_82 (O_82,N_2955,N_2998);
or UO_83 (O_83,N_2998,N_2956);
or UO_84 (O_84,N_2988,N_2984);
and UO_85 (O_85,N_2995,N_2979);
nand UO_86 (O_86,N_2994,N_2952);
nand UO_87 (O_87,N_2969,N_2990);
or UO_88 (O_88,N_2965,N_2993);
nor UO_89 (O_89,N_2998,N_2982);
or UO_90 (O_90,N_2997,N_2955);
nand UO_91 (O_91,N_2984,N_2970);
nor UO_92 (O_92,N_2964,N_2980);
nand UO_93 (O_93,N_2964,N_2984);
nor UO_94 (O_94,N_2965,N_2992);
and UO_95 (O_95,N_2980,N_2979);
nand UO_96 (O_96,N_2965,N_2999);
nor UO_97 (O_97,N_2967,N_2952);
xor UO_98 (O_98,N_2954,N_2991);
or UO_99 (O_99,N_2994,N_2973);
or UO_100 (O_100,N_2984,N_2974);
nand UO_101 (O_101,N_2991,N_2972);
xnor UO_102 (O_102,N_2985,N_2968);
xnor UO_103 (O_103,N_2995,N_2988);
xor UO_104 (O_104,N_2974,N_2999);
or UO_105 (O_105,N_2987,N_2980);
nor UO_106 (O_106,N_2962,N_2985);
xor UO_107 (O_107,N_2990,N_2987);
or UO_108 (O_108,N_2991,N_2953);
nor UO_109 (O_109,N_2999,N_2967);
or UO_110 (O_110,N_2982,N_2955);
nand UO_111 (O_111,N_2981,N_2967);
or UO_112 (O_112,N_2991,N_2993);
and UO_113 (O_113,N_2992,N_2959);
or UO_114 (O_114,N_2974,N_2964);
nor UO_115 (O_115,N_2976,N_2975);
or UO_116 (O_116,N_2964,N_2995);
nand UO_117 (O_117,N_2957,N_2985);
nand UO_118 (O_118,N_2989,N_2950);
nand UO_119 (O_119,N_2966,N_2951);
nand UO_120 (O_120,N_2966,N_2959);
and UO_121 (O_121,N_2968,N_2953);
nor UO_122 (O_122,N_2973,N_2964);
and UO_123 (O_123,N_2985,N_2993);
nor UO_124 (O_124,N_2987,N_2974);
xor UO_125 (O_125,N_2978,N_2988);
and UO_126 (O_126,N_2951,N_2964);
xor UO_127 (O_127,N_2961,N_2999);
or UO_128 (O_128,N_2977,N_2999);
xnor UO_129 (O_129,N_2971,N_2969);
and UO_130 (O_130,N_2991,N_2983);
nor UO_131 (O_131,N_2970,N_2999);
nor UO_132 (O_132,N_2974,N_2956);
and UO_133 (O_133,N_2964,N_2987);
nor UO_134 (O_134,N_2997,N_2956);
nor UO_135 (O_135,N_2964,N_2953);
nand UO_136 (O_136,N_2961,N_2998);
or UO_137 (O_137,N_2960,N_2972);
or UO_138 (O_138,N_2970,N_2963);
nand UO_139 (O_139,N_2970,N_2972);
nor UO_140 (O_140,N_2992,N_2981);
xnor UO_141 (O_141,N_2993,N_2960);
xor UO_142 (O_142,N_2979,N_2963);
nand UO_143 (O_143,N_2992,N_2982);
xnor UO_144 (O_144,N_2988,N_2980);
or UO_145 (O_145,N_2958,N_2974);
and UO_146 (O_146,N_2951,N_2990);
or UO_147 (O_147,N_2987,N_2975);
and UO_148 (O_148,N_2975,N_2981);
or UO_149 (O_149,N_2996,N_2957);
xnor UO_150 (O_150,N_2967,N_2969);
and UO_151 (O_151,N_2961,N_2995);
and UO_152 (O_152,N_2990,N_2972);
nand UO_153 (O_153,N_2979,N_2987);
or UO_154 (O_154,N_2979,N_2984);
nand UO_155 (O_155,N_2983,N_2968);
xor UO_156 (O_156,N_2965,N_2977);
and UO_157 (O_157,N_2968,N_2950);
and UO_158 (O_158,N_2971,N_2991);
and UO_159 (O_159,N_2955,N_2988);
and UO_160 (O_160,N_2999,N_2998);
nor UO_161 (O_161,N_2958,N_2960);
nand UO_162 (O_162,N_2956,N_2952);
or UO_163 (O_163,N_2977,N_2990);
nor UO_164 (O_164,N_2950,N_2982);
nand UO_165 (O_165,N_2969,N_2974);
or UO_166 (O_166,N_2954,N_2952);
nor UO_167 (O_167,N_2970,N_2973);
nor UO_168 (O_168,N_2995,N_2999);
and UO_169 (O_169,N_2994,N_2964);
or UO_170 (O_170,N_2980,N_2973);
nand UO_171 (O_171,N_2992,N_2977);
or UO_172 (O_172,N_2996,N_2993);
nor UO_173 (O_173,N_2986,N_2998);
nand UO_174 (O_174,N_2951,N_2956);
nor UO_175 (O_175,N_2952,N_2978);
xor UO_176 (O_176,N_2959,N_2981);
nor UO_177 (O_177,N_2999,N_2981);
or UO_178 (O_178,N_2968,N_2992);
or UO_179 (O_179,N_2966,N_2954);
nand UO_180 (O_180,N_2950,N_2993);
nor UO_181 (O_181,N_2994,N_2975);
nor UO_182 (O_182,N_2984,N_2972);
and UO_183 (O_183,N_2988,N_2966);
nand UO_184 (O_184,N_2950,N_2985);
nor UO_185 (O_185,N_2965,N_2972);
nand UO_186 (O_186,N_2952,N_2974);
nor UO_187 (O_187,N_2957,N_2966);
and UO_188 (O_188,N_2983,N_2975);
nand UO_189 (O_189,N_2996,N_2951);
or UO_190 (O_190,N_2979,N_2969);
and UO_191 (O_191,N_2989,N_2968);
or UO_192 (O_192,N_2984,N_2968);
nand UO_193 (O_193,N_2973,N_2969);
xor UO_194 (O_194,N_2958,N_2996);
nand UO_195 (O_195,N_2976,N_2968);
and UO_196 (O_196,N_2952,N_2996);
or UO_197 (O_197,N_2958,N_2969);
nand UO_198 (O_198,N_2966,N_2967);
or UO_199 (O_199,N_2959,N_2976);
or UO_200 (O_200,N_2959,N_2950);
nor UO_201 (O_201,N_2963,N_2951);
xor UO_202 (O_202,N_2969,N_2987);
xor UO_203 (O_203,N_2999,N_2997);
nor UO_204 (O_204,N_2985,N_2958);
and UO_205 (O_205,N_2961,N_2971);
nand UO_206 (O_206,N_2953,N_2956);
nand UO_207 (O_207,N_2979,N_2994);
nor UO_208 (O_208,N_2992,N_2951);
and UO_209 (O_209,N_2964,N_2957);
and UO_210 (O_210,N_2962,N_2977);
or UO_211 (O_211,N_2970,N_2991);
and UO_212 (O_212,N_2957,N_2954);
or UO_213 (O_213,N_2977,N_2967);
nor UO_214 (O_214,N_2957,N_2960);
xor UO_215 (O_215,N_2965,N_2953);
nor UO_216 (O_216,N_2983,N_2952);
or UO_217 (O_217,N_2971,N_2955);
and UO_218 (O_218,N_2987,N_2971);
nor UO_219 (O_219,N_2957,N_2999);
and UO_220 (O_220,N_2963,N_2973);
and UO_221 (O_221,N_2997,N_2995);
nand UO_222 (O_222,N_2976,N_2978);
xnor UO_223 (O_223,N_2972,N_2992);
nand UO_224 (O_224,N_2979,N_2975);
nand UO_225 (O_225,N_2982,N_2951);
nor UO_226 (O_226,N_2977,N_2985);
nor UO_227 (O_227,N_2985,N_2996);
nand UO_228 (O_228,N_2966,N_2998);
nor UO_229 (O_229,N_2964,N_2986);
and UO_230 (O_230,N_2951,N_2954);
nor UO_231 (O_231,N_2999,N_2980);
nor UO_232 (O_232,N_2979,N_2952);
and UO_233 (O_233,N_2972,N_2974);
nor UO_234 (O_234,N_2971,N_2967);
nor UO_235 (O_235,N_2993,N_2968);
and UO_236 (O_236,N_2965,N_2969);
or UO_237 (O_237,N_2956,N_2981);
xor UO_238 (O_238,N_2972,N_2971);
nor UO_239 (O_239,N_2951,N_2962);
and UO_240 (O_240,N_2997,N_2991);
and UO_241 (O_241,N_2970,N_2950);
or UO_242 (O_242,N_2996,N_2962);
nand UO_243 (O_243,N_2985,N_2994);
nor UO_244 (O_244,N_2982,N_2972);
or UO_245 (O_245,N_2989,N_2982);
and UO_246 (O_246,N_2988,N_2997);
nand UO_247 (O_247,N_2980,N_2958);
xor UO_248 (O_248,N_2959,N_2987);
or UO_249 (O_249,N_2998,N_2989);
or UO_250 (O_250,N_2962,N_2993);
nand UO_251 (O_251,N_2995,N_2998);
xor UO_252 (O_252,N_2978,N_2983);
xor UO_253 (O_253,N_2996,N_2955);
nand UO_254 (O_254,N_2958,N_2994);
xnor UO_255 (O_255,N_2971,N_2989);
nand UO_256 (O_256,N_2950,N_2951);
nand UO_257 (O_257,N_2991,N_2986);
or UO_258 (O_258,N_2969,N_2956);
nor UO_259 (O_259,N_2960,N_2956);
nor UO_260 (O_260,N_2952,N_2964);
nor UO_261 (O_261,N_2990,N_2954);
nor UO_262 (O_262,N_2967,N_2951);
nor UO_263 (O_263,N_2994,N_2962);
nor UO_264 (O_264,N_2976,N_2996);
nor UO_265 (O_265,N_2953,N_2990);
nand UO_266 (O_266,N_2953,N_2950);
and UO_267 (O_267,N_2976,N_2950);
or UO_268 (O_268,N_2994,N_2983);
and UO_269 (O_269,N_2977,N_2959);
or UO_270 (O_270,N_2964,N_2961);
nand UO_271 (O_271,N_2972,N_2975);
nor UO_272 (O_272,N_2984,N_2994);
and UO_273 (O_273,N_2997,N_2985);
nor UO_274 (O_274,N_2992,N_2955);
nor UO_275 (O_275,N_2984,N_2976);
or UO_276 (O_276,N_2982,N_2961);
nor UO_277 (O_277,N_2984,N_2969);
nor UO_278 (O_278,N_2960,N_2953);
nand UO_279 (O_279,N_2985,N_2984);
xor UO_280 (O_280,N_2978,N_2962);
and UO_281 (O_281,N_2976,N_2998);
or UO_282 (O_282,N_2953,N_2984);
or UO_283 (O_283,N_2954,N_2989);
nand UO_284 (O_284,N_2962,N_2988);
nor UO_285 (O_285,N_2961,N_2984);
nand UO_286 (O_286,N_2978,N_2971);
nor UO_287 (O_287,N_2997,N_2963);
or UO_288 (O_288,N_2969,N_2964);
nor UO_289 (O_289,N_2959,N_2958);
nand UO_290 (O_290,N_2981,N_2982);
and UO_291 (O_291,N_2955,N_2950);
or UO_292 (O_292,N_2987,N_2998);
xor UO_293 (O_293,N_2965,N_2962);
xor UO_294 (O_294,N_2998,N_2980);
and UO_295 (O_295,N_2969,N_2966);
or UO_296 (O_296,N_2999,N_2971);
nor UO_297 (O_297,N_2987,N_2989);
and UO_298 (O_298,N_2979,N_2981);
xnor UO_299 (O_299,N_2982,N_2986);
nor UO_300 (O_300,N_2988,N_2977);
or UO_301 (O_301,N_2971,N_2962);
nor UO_302 (O_302,N_2978,N_2979);
nor UO_303 (O_303,N_2971,N_2964);
and UO_304 (O_304,N_2975,N_2980);
xor UO_305 (O_305,N_2979,N_2976);
nand UO_306 (O_306,N_2984,N_2973);
nor UO_307 (O_307,N_2999,N_2984);
and UO_308 (O_308,N_2980,N_2991);
and UO_309 (O_309,N_2992,N_2969);
nor UO_310 (O_310,N_2992,N_2962);
or UO_311 (O_311,N_2971,N_2965);
nor UO_312 (O_312,N_2956,N_2955);
nand UO_313 (O_313,N_2991,N_2965);
or UO_314 (O_314,N_2981,N_2978);
nand UO_315 (O_315,N_2992,N_2995);
nand UO_316 (O_316,N_2979,N_2958);
nor UO_317 (O_317,N_2996,N_2984);
nand UO_318 (O_318,N_2976,N_2973);
nor UO_319 (O_319,N_2990,N_2978);
nor UO_320 (O_320,N_2983,N_2988);
xnor UO_321 (O_321,N_2971,N_2954);
nand UO_322 (O_322,N_2996,N_2970);
or UO_323 (O_323,N_2979,N_2950);
nand UO_324 (O_324,N_2990,N_2968);
or UO_325 (O_325,N_2975,N_2959);
and UO_326 (O_326,N_2951,N_2974);
nor UO_327 (O_327,N_2991,N_2950);
nand UO_328 (O_328,N_2989,N_2992);
and UO_329 (O_329,N_2963,N_2954);
nor UO_330 (O_330,N_2978,N_2986);
nand UO_331 (O_331,N_2955,N_2991);
nor UO_332 (O_332,N_2958,N_2991);
and UO_333 (O_333,N_2988,N_2994);
nor UO_334 (O_334,N_2972,N_2987);
or UO_335 (O_335,N_2957,N_2970);
and UO_336 (O_336,N_2973,N_2967);
nand UO_337 (O_337,N_2974,N_2981);
nand UO_338 (O_338,N_2959,N_2996);
and UO_339 (O_339,N_2982,N_2988);
or UO_340 (O_340,N_2963,N_2991);
xor UO_341 (O_341,N_2986,N_2959);
and UO_342 (O_342,N_2976,N_2997);
and UO_343 (O_343,N_2990,N_2956);
or UO_344 (O_344,N_2978,N_2961);
or UO_345 (O_345,N_2990,N_2985);
nand UO_346 (O_346,N_2950,N_2965);
or UO_347 (O_347,N_2965,N_2986);
and UO_348 (O_348,N_2974,N_2965);
nor UO_349 (O_349,N_2981,N_2987);
nor UO_350 (O_350,N_2975,N_2989);
or UO_351 (O_351,N_2997,N_2953);
nand UO_352 (O_352,N_2969,N_2985);
nor UO_353 (O_353,N_2996,N_2997);
xor UO_354 (O_354,N_2966,N_2952);
nor UO_355 (O_355,N_2977,N_2976);
nor UO_356 (O_356,N_2950,N_2963);
or UO_357 (O_357,N_2957,N_2986);
and UO_358 (O_358,N_2955,N_2977);
nor UO_359 (O_359,N_2971,N_2986);
xnor UO_360 (O_360,N_2971,N_2966);
and UO_361 (O_361,N_2996,N_2961);
nand UO_362 (O_362,N_2959,N_2999);
nor UO_363 (O_363,N_2974,N_2967);
and UO_364 (O_364,N_2950,N_2952);
nor UO_365 (O_365,N_2999,N_2985);
nor UO_366 (O_366,N_2991,N_2979);
and UO_367 (O_367,N_2954,N_2987);
and UO_368 (O_368,N_2983,N_2969);
or UO_369 (O_369,N_2966,N_2984);
or UO_370 (O_370,N_2991,N_2989);
or UO_371 (O_371,N_2966,N_2953);
xnor UO_372 (O_372,N_2983,N_2989);
nor UO_373 (O_373,N_2998,N_2996);
nand UO_374 (O_374,N_2996,N_2974);
xor UO_375 (O_375,N_2983,N_2993);
and UO_376 (O_376,N_2951,N_2961);
and UO_377 (O_377,N_2990,N_2988);
nand UO_378 (O_378,N_2971,N_2970);
nor UO_379 (O_379,N_2988,N_2965);
and UO_380 (O_380,N_2986,N_2955);
or UO_381 (O_381,N_2989,N_2974);
or UO_382 (O_382,N_2974,N_2961);
or UO_383 (O_383,N_2960,N_2997);
nand UO_384 (O_384,N_2985,N_2956);
or UO_385 (O_385,N_2970,N_2983);
xor UO_386 (O_386,N_2994,N_2966);
xor UO_387 (O_387,N_2959,N_2974);
and UO_388 (O_388,N_2968,N_2966);
or UO_389 (O_389,N_2959,N_2964);
nand UO_390 (O_390,N_2965,N_2970);
nand UO_391 (O_391,N_2982,N_2962);
nand UO_392 (O_392,N_2995,N_2994);
nand UO_393 (O_393,N_2957,N_2981);
nand UO_394 (O_394,N_2956,N_2970);
nor UO_395 (O_395,N_2988,N_2992);
nand UO_396 (O_396,N_2973,N_2987);
nand UO_397 (O_397,N_2959,N_2971);
and UO_398 (O_398,N_2989,N_2985);
or UO_399 (O_399,N_2963,N_2992);
nand UO_400 (O_400,N_2958,N_2984);
and UO_401 (O_401,N_2987,N_2978);
and UO_402 (O_402,N_2951,N_2989);
and UO_403 (O_403,N_2963,N_2957);
and UO_404 (O_404,N_2961,N_2994);
or UO_405 (O_405,N_2954,N_2970);
nand UO_406 (O_406,N_2986,N_2974);
nand UO_407 (O_407,N_2993,N_2955);
nand UO_408 (O_408,N_2950,N_2986);
or UO_409 (O_409,N_2974,N_2979);
nor UO_410 (O_410,N_2992,N_2953);
and UO_411 (O_411,N_2980,N_2953);
nand UO_412 (O_412,N_2977,N_2953);
nor UO_413 (O_413,N_2988,N_2958);
or UO_414 (O_414,N_2986,N_2966);
and UO_415 (O_415,N_2973,N_2975);
or UO_416 (O_416,N_2988,N_2973);
or UO_417 (O_417,N_2974,N_2993);
or UO_418 (O_418,N_2963,N_2958);
or UO_419 (O_419,N_2978,N_2982);
nor UO_420 (O_420,N_2984,N_2954);
and UO_421 (O_421,N_2951,N_2985);
and UO_422 (O_422,N_2979,N_2964);
xor UO_423 (O_423,N_2996,N_2994);
or UO_424 (O_424,N_2977,N_2981);
nor UO_425 (O_425,N_2960,N_2994);
or UO_426 (O_426,N_2953,N_2969);
and UO_427 (O_427,N_2954,N_2968);
nor UO_428 (O_428,N_2991,N_2998);
nand UO_429 (O_429,N_2996,N_2953);
nand UO_430 (O_430,N_2993,N_2981);
and UO_431 (O_431,N_2997,N_2952);
xnor UO_432 (O_432,N_2981,N_2986);
or UO_433 (O_433,N_2984,N_2989);
and UO_434 (O_434,N_2966,N_2963);
and UO_435 (O_435,N_2994,N_2954);
nand UO_436 (O_436,N_2962,N_2950);
and UO_437 (O_437,N_2952,N_2985);
and UO_438 (O_438,N_2961,N_2992);
nor UO_439 (O_439,N_2997,N_2994);
xnor UO_440 (O_440,N_2979,N_2957);
and UO_441 (O_441,N_2950,N_2969);
nor UO_442 (O_442,N_2965,N_2990);
nor UO_443 (O_443,N_2998,N_2970);
xor UO_444 (O_444,N_2996,N_2991);
nand UO_445 (O_445,N_2998,N_2957);
nor UO_446 (O_446,N_2974,N_2968);
or UO_447 (O_447,N_2973,N_2972);
or UO_448 (O_448,N_2952,N_2992);
or UO_449 (O_449,N_2968,N_2951);
or UO_450 (O_450,N_2977,N_2980);
nand UO_451 (O_451,N_2957,N_2974);
nor UO_452 (O_452,N_2953,N_2961);
nand UO_453 (O_453,N_2991,N_2987);
nor UO_454 (O_454,N_2961,N_2968);
and UO_455 (O_455,N_2994,N_2972);
and UO_456 (O_456,N_2965,N_2982);
and UO_457 (O_457,N_2961,N_2960);
nand UO_458 (O_458,N_2976,N_2961);
xnor UO_459 (O_459,N_2953,N_2979);
nand UO_460 (O_460,N_2970,N_2976);
nor UO_461 (O_461,N_2992,N_2966);
nor UO_462 (O_462,N_2994,N_2992);
and UO_463 (O_463,N_2968,N_2969);
and UO_464 (O_464,N_2990,N_2983);
nand UO_465 (O_465,N_2986,N_2973);
nand UO_466 (O_466,N_2969,N_2977);
nand UO_467 (O_467,N_2991,N_2968);
or UO_468 (O_468,N_2993,N_2997);
or UO_469 (O_469,N_2979,N_2961);
nor UO_470 (O_470,N_2961,N_2987);
nor UO_471 (O_471,N_2996,N_2981);
and UO_472 (O_472,N_2987,N_2970);
and UO_473 (O_473,N_2994,N_2987);
xnor UO_474 (O_474,N_2965,N_2979);
nand UO_475 (O_475,N_2997,N_2973);
or UO_476 (O_476,N_2959,N_2983);
or UO_477 (O_477,N_2964,N_2993);
or UO_478 (O_478,N_2969,N_2955);
nand UO_479 (O_479,N_2987,N_2962);
nor UO_480 (O_480,N_2966,N_2991);
nand UO_481 (O_481,N_2960,N_2976);
nand UO_482 (O_482,N_2976,N_2995);
and UO_483 (O_483,N_2976,N_2966);
nor UO_484 (O_484,N_2975,N_2964);
xnor UO_485 (O_485,N_2980,N_2995);
nand UO_486 (O_486,N_2977,N_2951);
nand UO_487 (O_487,N_2970,N_2982);
or UO_488 (O_488,N_2968,N_2957);
nand UO_489 (O_489,N_2969,N_2976);
xor UO_490 (O_490,N_2966,N_2974);
nand UO_491 (O_491,N_2966,N_2995);
nor UO_492 (O_492,N_2993,N_2951);
and UO_493 (O_493,N_2999,N_2983);
nor UO_494 (O_494,N_2956,N_2976);
nand UO_495 (O_495,N_2962,N_2989);
and UO_496 (O_496,N_2955,N_2985);
nand UO_497 (O_497,N_2984,N_2957);
and UO_498 (O_498,N_2991,N_2990);
or UO_499 (O_499,N_2989,N_2993);
endmodule