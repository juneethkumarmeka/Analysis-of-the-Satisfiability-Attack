module basic_1000_10000_1500_2_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5001,N_5002,N_5003,N_5005,N_5006,N_5007,N_5009,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5019,N_5021,N_5022,N_5023,N_5025,N_5026,N_5027,N_5031,N_5033,N_5034,N_5035,N_5036,N_5037,N_5042,N_5043,N_5049,N_5051,N_5053,N_5054,N_5055,N_5059,N_5060,N_5062,N_5063,N_5065,N_5068,N_5069,N_5070,N_5071,N_5074,N_5075,N_5076,N_5078,N_5079,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5096,N_5097,N_5098,N_5104,N_5105,N_5106,N_5110,N_5112,N_5113,N_5114,N_5115,N_5117,N_5118,N_5121,N_5122,N_5124,N_5125,N_5126,N_5127,N_5129,N_5130,N_5131,N_5132,N_5137,N_5138,N_5142,N_5144,N_5145,N_5149,N_5151,N_5154,N_5155,N_5156,N_5158,N_5159,N_5160,N_5162,N_5163,N_5164,N_5167,N_5168,N_5169,N_5171,N_5172,N_5174,N_5175,N_5182,N_5186,N_5188,N_5191,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5204,N_5206,N_5209,N_5210,N_5211,N_5212,N_5214,N_5215,N_5216,N_5218,N_5220,N_5221,N_5222,N_5226,N_5227,N_5229,N_5230,N_5231,N_5233,N_5234,N_5235,N_5236,N_5239,N_5240,N_5242,N_5245,N_5247,N_5252,N_5253,N_5254,N_5255,N_5256,N_5258,N_5259,N_5261,N_5262,N_5263,N_5264,N_5266,N_5267,N_5268,N_5271,N_5272,N_5273,N_5277,N_5279,N_5280,N_5283,N_5285,N_5286,N_5289,N_5291,N_5292,N_5295,N_5297,N_5298,N_5300,N_5301,N_5302,N_5303,N_5305,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5317,N_5318,N_5321,N_5323,N_5324,N_5325,N_5326,N_5328,N_5329,N_5330,N_5332,N_5333,N_5334,N_5335,N_5337,N_5338,N_5339,N_5340,N_5341,N_5343,N_5345,N_5347,N_5348,N_5349,N_5351,N_5352,N_5354,N_5355,N_5356,N_5358,N_5360,N_5364,N_5367,N_5369,N_5374,N_5376,N_5377,N_5380,N_5381,N_5383,N_5385,N_5387,N_5388,N_5390,N_5391,N_5393,N_5394,N_5396,N_5397,N_5398,N_5399,N_5400,N_5402,N_5403,N_5404,N_5406,N_5410,N_5411,N_5413,N_5414,N_5415,N_5421,N_5426,N_5427,N_5431,N_5432,N_5443,N_5444,N_5445,N_5447,N_5448,N_5449,N_5450,N_5452,N_5453,N_5454,N_5455,N_5459,N_5460,N_5462,N_5463,N_5466,N_5470,N_5471,N_5472,N_5473,N_5477,N_5483,N_5486,N_5491,N_5493,N_5495,N_5496,N_5498,N_5499,N_5501,N_5502,N_5504,N_5506,N_5507,N_5509,N_5510,N_5515,N_5516,N_5522,N_5524,N_5525,N_5527,N_5528,N_5529,N_5530,N_5532,N_5533,N_5534,N_5535,N_5536,N_5538,N_5542,N_5544,N_5546,N_5547,N_5549,N_5550,N_5551,N_5553,N_5554,N_5555,N_5556,N_5557,N_5559,N_5561,N_5562,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5575,N_5576,N_5577,N_5579,N_5580,N_5581,N_5583,N_5585,N_5586,N_5587,N_5588,N_5590,N_5591,N_5593,N_5595,N_5598,N_5599,N_5601,N_5602,N_5603,N_5605,N_5606,N_5607,N_5609,N_5610,N_5611,N_5616,N_5617,N_5618,N_5622,N_5623,N_5624,N_5625,N_5627,N_5628,N_5633,N_5635,N_5636,N_5637,N_5639,N_5640,N_5648,N_5649,N_5650,N_5652,N_5657,N_5658,N_5660,N_5661,N_5662,N_5664,N_5665,N_5666,N_5667,N_5671,N_5672,N_5673,N_5675,N_5676,N_5678,N_5682,N_5684,N_5685,N_5686,N_5687,N_5689,N_5690,N_5691,N_5694,N_5696,N_5697,N_5698,N_5700,N_5701,N_5702,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5714,N_5715,N_5716,N_5720,N_5721,N_5723,N_5725,N_5726,N_5727,N_5728,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5737,N_5740,N_5743,N_5745,N_5747,N_5748,N_5749,N_5750,N_5752,N_5755,N_5758,N_5760,N_5761,N_5762,N_5763,N_5764,N_5766,N_5767,N_5768,N_5771,N_5773,N_5774,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5785,N_5788,N_5789,N_5791,N_5792,N_5793,N_5794,N_5795,N_5797,N_5800,N_5801,N_5802,N_5804,N_5806,N_5809,N_5812,N_5814,N_5815,N_5816,N_5818,N_5819,N_5823,N_5825,N_5829,N_5832,N_5833,N_5834,N_5835,N_5836,N_5839,N_5840,N_5842,N_5844,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5858,N_5859,N_5860,N_5861,N_5863,N_5864,N_5867,N_5868,N_5869,N_5870,N_5872,N_5874,N_5875,N_5876,N_5877,N_5879,N_5880,N_5881,N_5883,N_5885,N_5886,N_5888,N_5890,N_5891,N_5892,N_5898,N_5899,N_5900,N_5903,N_5904,N_5905,N_5907,N_5909,N_5910,N_5911,N_5915,N_5918,N_5919,N_5922,N_5925,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5940,N_5941,N_5942,N_5945,N_5947,N_5948,N_5949,N_5950,N_5951,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5960,N_5961,N_5962,N_5963,N_5966,N_5967,N_5968,N_5969,N_5970,N_5974,N_5975,N_5978,N_5980,N_5983,N_5985,N_5987,N_5988,N_5989,N_5991,N_5992,N_5993,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6002,N_6003,N_6004,N_6006,N_6011,N_6012,N_6013,N_6014,N_6015,N_6017,N_6020,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6031,N_6034,N_6036,N_6039,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6050,N_6051,N_6052,N_6053,N_6054,N_6056,N_6058,N_6059,N_6060,N_6064,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6075,N_6076,N_6077,N_6078,N_6079,N_6081,N_6082,N_6083,N_6084,N_6085,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6104,N_6105,N_6106,N_6109,N_6110,N_6111,N_6115,N_6116,N_6117,N_6118,N_6122,N_6124,N_6125,N_6127,N_6128,N_6131,N_6133,N_6136,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6146,N_6147,N_6148,N_6150,N_6152,N_6154,N_6155,N_6156,N_6157,N_6158,N_6160,N_6161,N_6166,N_6167,N_6168,N_6169,N_6172,N_6175,N_6176,N_6177,N_6178,N_6180,N_6181,N_6183,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6204,N_6208,N_6209,N_6210,N_6211,N_6213,N_6214,N_6216,N_6217,N_6218,N_6220,N_6224,N_6225,N_6227,N_6228,N_6231,N_6233,N_6235,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6249,N_6251,N_6253,N_6254,N_6255,N_6257,N_6258,N_6260,N_6261,N_6263,N_6265,N_6269,N_6270,N_6271,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6281,N_6282,N_6283,N_6285,N_6287,N_6288,N_6289,N_6291,N_6293,N_6294,N_6296,N_6297,N_6298,N_6299,N_6300,N_6304,N_6305,N_6306,N_6308,N_6309,N_6311,N_6314,N_6315,N_6316,N_6317,N_6319,N_6320,N_6321,N_6323,N_6324,N_6325,N_6327,N_6328,N_6329,N_6330,N_6334,N_6335,N_6338,N_6339,N_6340,N_6341,N_6344,N_6346,N_6348,N_6351,N_6353,N_6355,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6373,N_6374,N_6375,N_6377,N_6378,N_6379,N_6384,N_6385,N_6386,N_6388,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6405,N_6407,N_6409,N_6410,N_6411,N_6412,N_6415,N_6416,N_6422,N_6424,N_6426,N_6427,N_6428,N_6429,N_6430,N_6432,N_6434,N_6435,N_6436,N_6440,N_6441,N_6444,N_6447,N_6449,N_6451,N_6452,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6462,N_6463,N_6465,N_6467,N_6469,N_6470,N_6471,N_6472,N_6473,N_6477,N_6479,N_6480,N_6482,N_6483,N_6484,N_6487,N_6489,N_6490,N_6493,N_6496,N_6499,N_6501,N_6503,N_6505,N_6506,N_6509,N_6512,N_6514,N_6515,N_6516,N_6519,N_6520,N_6521,N_6523,N_6524,N_6525,N_6526,N_6528,N_6531,N_6532,N_6533,N_6534,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6551,N_6553,N_6554,N_6556,N_6557,N_6559,N_6560,N_6561,N_6563,N_6565,N_6566,N_6567,N_6569,N_6570,N_6572,N_6574,N_6575,N_6577,N_6578,N_6579,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6590,N_6594,N_6596,N_6597,N_6598,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6621,N_6623,N_6625,N_6626,N_6629,N_6630,N_6635,N_6636,N_6638,N_6639,N_6640,N_6643,N_6644,N_6648,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6660,N_6661,N_6662,N_6664,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6673,N_6674,N_6676,N_6678,N_6679,N_6681,N_6682,N_6683,N_6684,N_6685,N_6689,N_6690,N_6692,N_6694,N_6695,N_6696,N_6698,N_6699,N_6701,N_6703,N_6704,N_6705,N_6710,N_6711,N_6712,N_6713,N_6715,N_6716,N_6717,N_6721,N_6722,N_6727,N_6729,N_6730,N_6732,N_6733,N_6735,N_6739,N_6740,N_6742,N_6743,N_6744,N_6746,N_6749,N_6751,N_6752,N_6753,N_6755,N_6757,N_6759,N_6763,N_6764,N_6765,N_6766,N_6768,N_6769,N_6771,N_6772,N_6775,N_6776,N_6777,N_6779,N_6781,N_6783,N_6784,N_6786,N_6787,N_6788,N_6789,N_6790,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6800,N_6801,N_6803,N_6806,N_6807,N_6809,N_6810,N_6812,N_6813,N_6814,N_6815,N_6816,N_6819,N_6821,N_6822,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6832,N_6833,N_6838,N_6840,N_6841,N_6843,N_6847,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6867,N_6868,N_6870,N_6874,N_6876,N_6881,N_6882,N_6884,N_6887,N_6888,N_6889,N_6890,N_6899,N_6900,N_6901,N_6904,N_6905,N_6907,N_6908,N_6909,N_6916,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6929,N_6930,N_6931,N_6933,N_6934,N_6935,N_6938,N_6939,N_6942,N_6943,N_6944,N_6946,N_6949,N_6952,N_6954,N_6958,N_6961,N_6964,N_6968,N_6969,N_6971,N_6972,N_6978,N_6979,N_6980,N_6982,N_6983,N_6985,N_6986,N_6989,N_6990,N_6991,N_6992,N_6996,N_6997,N_6998,N_6999,N_7000,N_7003,N_7004,N_7007,N_7008,N_7009,N_7011,N_7012,N_7013,N_7014,N_7016,N_7017,N_7018,N_7020,N_7021,N_7022,N_7027,N_7028,N_7029,N_7031,N_7032,N_7034,N_7036,N_7037,N_7038,N_7039,N_7040,N_7043,N_7044,N_7046,N_7048,N_7049,N_7050,N_7052,N_7053,N_7054,N_7055,N_7056,N_7058,N_7062,N_7065,N_7068,N_7069,N_7070,N_7072,N_7073,N_7075,N_7076,N_7077,N_7078,N_7082,N_7083,N_7084,N_7085,N_7087,N_7089,N_7090,N_7093,N_7094,N_7095,N_7097,N_7098,N_7099,N_7100,N_7102,N_7103,N_7104,N_7107,N_7108,N_7111,N_7113,N_7114,N_7117,N_7118,N_7121,N_7122,N_7123,N_7127,N_7130,N_7131,N_7135,N_7136,N_7137,N_7142,N_7145,N_7146,N_7147,N_7148,N_7149,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7160,N_7162,N_7163,N_7164,N_7165,N_7166,N_7168,N_7169,N_7171,N_7172,N_7174,N_7176,N_7179,N_7180,N_7181,N_7183,N_7185,N_7186,N_7187,N_7188,N_7191,N_7192,N_7195,N_7196,N_7197,N_7198,N_7199,N_7201,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7225,N_7226,N_7227,N_7228,N_7230,N_7233,N_7234,N_7235,N_7236,N_7238,N_7239,N_7240,N_7241,N_7243,N_7245,N_7248,N_7249,N_7251,N_7252,N_7259,N_7260,N_7261,N_7262,N_7264,N_7266,N_7269,N_7270,N_7273,N_7276,N_7280,N_7281,N_7282,N_7283,N_7285,N_7286,N_7289,N_7290,N_7295,N_7301,N_7303,N_7304,N_7305,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7316,N_7317,N_7321,N_7323,N_7324,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7336,N_7338,N_7339,N_7342,N_7344,N_7345,N_7346,N_7348,N_7349,N_7352,N_7353,N_7354,N_7357,N_7358,N_7359,N_7360,N_7361,N_7363,N_7364,N_7365,N_7366,N_7368,N_7369,N_7370,N_7371,N_7372,N_7374,N_7375,N_7376,N_7377,N_7379,N_7380,N_7383,N_7384,N_7386,N_7389,N_7390,N_7395,N_7397,N_7398,N_7399,N_7401,N_7403,N_7404,N_7406,N_7407,N_7408,N_7409,N_7412,N_7413,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7424,N_7425,N_7426,N_7427,N_7428,N_7431,N_7433,N_7434,N_7435,N_7436,N_7437,N_7439,N_7441,N_7442,N_7443,N_7445,N_7446,N_7447,N_7448,N_7452,N_7453,N_7454,N_7455,N_7457,N_7460,N_7461,N_7462,N_7463,N_7465,N_7467,N_7468,N_7469,N_7470,N_7472,N_7474,N_7475,N_7476,N_7478,N_7480,N_7482,N_7483,N_7484,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7494,N_7495,N_7497,N_7500,N_7501,N_7502,N_7503,N_7505,N_7508,N_7510,N_7511,N_7513,N_7514,N_7515,N_7516,N_7517,N_7522,N_7523,N_7524,N_7526,N_7527,N_7528,N_7529,N_7533,N_7535,N_7536,N_7537,N_7538,N_7540,N_7544,N_7545,N_7546,N_7547,N_7548,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7558,N_7559,N_7562,N_7565,N_7566,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7585,N_7589,N_7590,N_7591,N_7594,N_7595,N_7596,N_7597,N_7598,N_7601,N_7602,N_7603,N_7605,N_7606,N_7607,N_7611,N_7612,N_7613,N_7615,N_7618,N_7620,N_7621,N_7622,N_7623,N_7624,N_7628,N_7629,N_7631,N_7634,N_7635,N_7640,N_7641,N_7643,N_7646,N_7647,N_7648,N_7649,N_7650,N_7653,N_7654,N_7659,N_7660,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7669,N_7670,N_7672,N_7673,N_7674,N_7675,N_7676,N_7680,N_7681,N_7682,N_7683,N_7685,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7698,N_7699,N_7701,N_7704,N_7705,N_7706,N_7707,N_7708,N_7711,N_7715,N_7716,N_7717,N_7719,N_7721,N_7722,N_7725,N_7729,N_7730,N_7732,N_7734,N_7737,N_7738,N_7739,N_7740,N_7741,N_7745,N_7746,N_7747,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7756,N_7758,N_7759,N_7760,N_7762,N_7763,N_7769,N_7770,N_7771,N_7773,N_7774,N_7775,N_7777,N_7780,N_7782,N_7784,N_7786,N_7787,N_7788,N_7789,N_7791,N_7792,N_7794,N_7795,N_7797,N_7799,N_7800,N_7802,N_7805,N_7806,N_7810,N_7812,N_7813,N_7814,N_7815,N_7816,N_7818,N_7819,N_7820,N_7824,N_7825,N_7826,N_7831,N_7832,N_7833,N_7834,N_7836,N_7837,N_7838,N_7839,N_7840,N_7843,N_7845,N_7846,N_7847,N_7849,N_7852,N_7855,N_7856,N_7857,N_7860,N_7861,N_7862,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7884,N_7885,N_7886,N_7887,N_7888,N_7890,N_7894,N_7896,N_7898,N_7900,N_7901,N_7903,N_7904,N_7908,N_7909,N_7910,N_7911,N_7913,N_7914,N_7917,N_7918,N_7920,N_7921,N_7922,N_7923,N_7925,N_7926,N_7927,N_7928,N_7931,N_7932,N_7933,N_7935,N_7936,N_7939,N_7941,N_7942,N_7943,N_7945,N_7946,N_7947,N_7949,N_7950,N_7952,N_7953,N_7956,N_7957,N_7960,N_7962,N_7963,N_7965,N_7966,N_7968,N_7969,N_7972,N_7973,N_7974,N_7975,N_7976,N_7979,N_7981,N_7982,N_7983,N_7984,N_7987,N_7988,N_7989,N_7992,N_7997,N_7999,N_8001,N_8004,N_8005,N_8012,N_8014,N_8015,N_8016,N_8017,N_8019,N_8020,N_8022,N_8023,N_8024,N_8027,N_8030,N_8035,N_8037,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8049,N_8051,N_8058,N_8062,N_8064,N_8065,N_8068,N_8070,N_8071,N_8074,N_8076,N_8078,N_8079,N_8081,N_8082,N_8084,N_8086,N_8087,N_8088,N_8091,N_8093,N_8094,N_8099,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8110,N_8111,N_8114,N_8116,N_8119,N_8122,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8133,N_8134,N_8135,N_8139,N_8140,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8159,N_8160,N_8161,N_8163,N_8166,N_8168,N_8172,N_8173,N_8175,N_8176,N_8177,N_8181,N_8183,N_8186,N_8189,N_8190,N_8192,N_8193,N_8196,N_8199,N_8200,N_8203,N_8204,N_8205,N_8206,N_8208,N_8210,N_8212,N_8213,N_8214,N_8216,N_8217,N_8219,N_8220,N_8226,N_8227,N_8228,N_8229,N_8230,N_8232,N_8233,N_8234,N_8235,N_8236,N_8239,N_8241,N_8242,N_8243,N_8247,N_8248,N_8249,N_8251,N_8255,N_8256,N_8258,N_8259,N_8260,N_8262,N_8263,N_8264,N_8265,N_8266,N_8269,N_8272,N_8274,N_8275,N_8276,N_8279,N_8282,N_8284,N_8285,N_8286,N_8288,N_8292,N_8301,N_8303,N_8304,N_8306,N_8307,N_8308,N_8309,N_8310,N_8312,N_8314,N_8316,N_8317,N_8318,N_8320,N_8321,N_8324,N_8326,N_8327,N_8329,N_8330,N_8331,N_8333,N_8334,N_8335,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8349,N_8352,N_8353,N_8354,N_8356,N_8359,N_8361,N_8366,N_8368,N_8370,N_8371,N_8372,N_8375,N_8380,N_8382,N_8383,N_8386,N_8387,N_8388,N_8390,N_8400,N_8401,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8411,N_8416,N_8417,N_8419,N_8420,N_8422,N_8423,N_8424,N_8426,N_8428,N_8430,N_8432,N_8433,N_8436,N_8437,N_8439,N_8441,N_8444,N_8446,N_8448,N_8450,N_8451,N_8452,N_8455,N_8457,N_8461,N_8462,N_8463,N_8466,N_8468,N_8469,N_8471,N_8474,N_8475,N_8477,N_8478,N_8481,N_8485,N_8486,N_8487,N_8488,N_8489,N_8492,N_8493,N_8494,N_8495,N_8500,N_8502,N_8503,N_8504,N_8507,N_8508,N_8510,N_8511,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8528,N_8530,N_8531,N_8532,N_8533,N_8535,N_8537,N_8539,N_8540,N_8541,N_8542,N_8543,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8555,N_8556,N_8559,N_8560,N_8561,N_8563,N_8566,N_8567,N_8568,N_8570,N_8571,N_8572,N_8574,N_8575,N_8579,N_8580,N_8581,N_8582,N_8584,N_8586,N_8587,N_8588,N_8589,N_8590,N_8592,N_8595,N_8597,N_8603,N_8606,N_8608,N_8610,N_8611,N_8614,N_8615,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8625,N_8626,N_8627,N_8632,N_8633,N_8634,N_8635,N_8639,N_8640,N_8641,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8650,N_8652,N_8655,N_8657,N_8658,N_8659,N_8660,N_8662,N_8665,N_8666,N_8668,N_8669,N_8670,N_8672,N_8674,N_8676,N_8677,N_8678,N_8680,N_8681,N_8682,N_8684,N_8685,N_8686,N_8687,N_8688,N_8690,N_8691,N_8692,N_8694,N_8695,N_8698,N_8701,N_8702,N_8703,N_8704,N_8705,N_8707,N_8708,N_8710,N_8711,N_8713,N_8714,N_8716,N_8719,N_8720,N_8721,N_8724,N_8725,N_8726,N_8729,N_8731,N_8732,N_8733,N_8737,N_8738,N_8739,N_8742,N_8743,N_8744,N_8745,N_8746,N_8748,N_8749,N_8750,N_8755,N_8756,N_8758,N_8759,N_8760,N_8761,N_8762,N_8764,N_8765,N_8768,N_8769,N_8771,N_8772,N_8773,N_8775,N_8777,N_8778,N_8779,N_8780,N_8782,N_8783,N_8784,N_8785,N_8787,N_8790,N_8794,N_8795,N_8796,N_8797,N_8799,N_8800,N_8801,N_8802,N_8803,N_8806,N_8807,N_8809,N_8810,N_8811,N_8815,N_8816,N_8819,N_8821,N_8823,N_8824,N_8825,N_8826,N_8827,N_8829,N_8831,N_8833,N_8834,N_8837,N_8839,N_8841,N_8843,N_8846,N_8847,N_8848,N_8849,N_8850,N_8854,N_8855,N_8857,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8866,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8880,N_8884,N_8885,N_8886,N_8887,N_8888,N_8891,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8903,N_8904,N_8905,N_8907,N_8910,N_8912,N_8913,N_8915,N_8917,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8931,N_8932,N_8933,N_8934,N_8936,N_8939,N_8941,N_8942,N_8945,N_8947,N_8950,N_8951,N_8953,N_8957,N_8958,N_8962,N_8967,N_8971,N_8973,N_8975,N_8976,N_8978,N_8979,N_8980,N_8981,N_8982,N_8986,N_8987,N_8989,N_8992,N_8993,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9007,N_9009,N_9010,N_9011,N_9012,N_9014,N_9015,N_9016,N_9017,N_9019,N_9024,N_9025,N_9029,N_9032,N_9033,N_9035,N_9036,N_9037,N_9042,N_9046,N_9047,N_9048,N_9050,N_9051,N_9053,N_9055,N_9056,N_9058,N_9059,N_9061,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9070,N_9071,N_9073,N_9075,N_9077,N_9078,N_9079,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9089,N_9091,N_9093,N_9095,N_9096,N_9099,N_9104,N_9105,N_9106,N_9107,N_9108,N_9111,N_9112,N_9113,N_9114,N_9116,N_9117,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9134,N_9136,N_9137,N_9138,N_9140,N_9142,N_9145,N_9146,N_9149,N_9150,N_9152,N_9153,N_9154,N_9155,N_9157,N_9162,N_9163,N_9165,N_9169,N_9170,N_9174,N_9175,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9191,N_9192,N_9193,N_9194,N_9196,N_9197,N_9198,N_9199,N_9202,N_9206,N_9207,N_9209,N_9210,N_9212,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9221,N_9222,N_9227,N_9228,N_9229,N_9230,N_9233,N_9236,N_9239,N_9240,N_9243,N_9244,N_9245,N_9246,N_9247,N_9251,N_9256,N_9257,N_9258,N_9261,N_9262,N_9265,N_9266,N_9267,N_9268,N_9270,N_9272,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9282,N_9283,N_9284,N_9285,N_9286,N_9288,N_9289,N_9290,N_9292,N_9294,N_9296,N_9298,N_9299,N_9301,N_9302,N_9304,N_9307,N_9308,N_9309,N_9310,N_9312,N_9313,N_9314,N_9316,N_9318,N_9319,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9330,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9340,N_9341,N_9342,N_9343,N_9346,N_9348,N_9349,N_9355,N_9356,N_9358,N_9361,N_9362,N_9364,N_9369,N_9373,N_9374,N_9376,N_9386,N_9387,N_9388,N_9390,N_9391,N_9392,N_9395,N_9396,N_9397,N_9400,N_9402,N_9403,N_9404,N_9406,N_9408,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9419,N_9420,N_9422,N_9423,N_9424,N_9425,N_9427,N_9429,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9438,N_9440,N_9448,N_9449,N_9451,N_9452,N_9453,N_9454,N_9455,N_9457,N_9458,N_9460,N_9463,N_9468,N_9470,N_9471,N_9472,N_9475,N_9476,N_9477,N_9478,N_9480,N_9482,N_9483,N_9485,N_9489,N_9492,N_9493,N_9495,N_9496,N_9497,N_9499,N_9503,N_9506,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9516,N_9518,N_9519,N_9523,N_9524,N_9525,N_9529,N_9530,N_9531,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9540,N_9541,N_9542,N_9544,N_9545,N_9546,N_9550,N_9551,N_9552,N_9553,N_9556,N_9557,N_9559,N_9560,N_9562,N_9563,N_9564,N_9567,N_9571,N_9574,N_9577,N_9579,N_9580,N_9581,N_9584,N_9587,N_9589,N_9591,N_9592,N_9594,N_9595,N_9597,N_9599,N_9600,N_9601,N_9602,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9612,N_9616,N_9617,N_9619,N_9620,N_9621,N_9622,N_9623,N_9625,N_9626,N_9627,N_9630,N_9633,N_9634,N_9635,N_9637,N_9640,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9651,N_9653,N_9654,N_9655,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9667,N_9668,N_9669,N_9674,N_9675,N_9676,N_9679,N_9680,N_9681,N_9684,N_9687,N_9688,N_9689,N_9690,N_9691,N_9693,N_9696,N_9697,N_9698,N_9702,N_9703,N_9705,N_9708,N_9709,N_9710,N_9711,N_9713,N_9714,N_9716,N_9717,N_9720,N_9722,N_9723,N_9725,N_9726,N_9727,N_9728,N_9733,N_9734,N_9735,N_9736,N_9737,N_9739,N_9740,N_9741,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9751,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9762,N_9764,N_9765,N_9766,N_9768,N_9769,N_9770,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9781,N_9782,N_9785,N_9786,N_9789,N_9791,N_9792,N_9793,N_9795,N_9796,N_9797,N_9798,N_9799,N_9801,N_9803,N_9804,N_9805,N_9806,N_9808,N_9809,N_9811,N_9812,N_9813,N_9815,N_9816,N_9817,N_9818,N_9820,N_9821,N_9823,N_9826,N_9828,N_9829,N_9830,N_9832,N_9833,N_9836,N_9841,N_9842,N_9843,N_9844,N_9846,N_9848,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9864,N_9869,N_9871,N_9874,N_9875,N_9876,N_9878,N_9880,N_9881,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9892,N_9893,N_9894,N_9896,N_9897,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9911,N_9912,N_9913,N_9914,N_9915,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9924,N_9925,N_9927,N_9930,N_9931,N_9935,N_9938,N_9939,N_9940,N_9943,N_9944,N_9946,N_9947,N_9948,N_9949,N_9950,N_9952,N_9953,N_9955,N_9956,N_9957,N_9960,N_9964,N_9965,N_9966,N_9969,N_9970,N_9972,N_9974,N_9975,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9984,N_9985,N_9986,N_9989,N_9991,N_9992,N_9993,N_9995,N_9996,N_9997,N_9999;
or U0 (N_0,In_233,In_497);
or U1 (N_1,In_267,In_942);
or U2 (N_2,In_637,In_59);
or U3 (N_3,In_683,In_677);
xnor U4 (N_4,In_384,In_748);
nor U5 (N_5,In_588,In_853);
nand U6 (N_6,In_951,In_899);
or U7 (N_7,In_916,In_232);
nand U8 (N_8,In_591,In_430);
nand U9 (N_9,In_4,In_70);
nor U10 (N_10,In_937,In_204);
xnor U11 (N_11,In_858,In_728);
and U12 (N_12,In_504,In_646);
nand U13 (N_13,In_699,In_872);
and U14 (N_14,In_451,In_411);
nand U15 (N_15,In_444,In_630);
nand U16 (N_16,In_344,In_999);
and U17 (N_17,In_27,In_634);
nor U18 (N_18,In_163,In_84);
or U19 (N_19,In_322,In_211);
nor U20 (N_20,In_626,In_765);
or U21 (N_21,In_182,In_517);
and U22 (N_22,In_289,In_323);
and U23 (N_23,In_548,In_834);
nor U24 (N_24,In_889,In_96);
nand U25 (N_25,In_394,In_854);
or U26 (N_26,In_208,In_724);
nor U27 (N_27,In_442,In_439);
and U28 (N_28,In_127,In_892);
nand U29 (N_29,In_791,In_968);
nor U30 (N_30,In_374,In_906);
nor U31 (N_31,In_828,In_111);
nor U32 (N_32,In_249,In_429);
nor U33 (N_33,In_882,In_901);
nor U34 (N_34,In_353,In_237);
nor U35 (N_35,In_918,In_513);
or U36 (N_36,In_19,In_216);
nand U37 (N_37,In_514,In_152);
nand U38 (N_38,In_939,In_109);
or U39 (N_39,In_376,In_848);
nand U40 (N_40,In_799,In_814);
xnor U41 (N_41,In_707,In_930);
or U42 (N_42,In_986,In_871);
or U43 (N_43,In_43,In_469);
xnor U44 (N_44,In_101,In_191);
or U45 (N_45,In_841,In_678);
nand U46 (N_46,In_18,In_553);
nor U47 (N_47,In_31,In_800);
or U48 (N_48,In_99,In_961);
and U49 (N_49,In_483,In_518);
or U50 (N_50,In_623,In_744);
nor U51 (N_51,In_658,In_29);
and U52 (N_52,In_402,In_365);
or U53 (N_53,In_957,In_761);
or U54 (N_54,In_958,In_845);
nand U55 (N_55,In_425,In_572);
nand U56 (N_56,In_946,In_562);
nand U57 (N_57,In_994,In_22);
nor U58 (N_58,In_352,In_87);
xor U59 (N_59,In_717,In_740);
and U60 (N_60,In_253,In_114);
nand U61 (N_61,In_285,In_488);
xor U62 (N_62,In_149,In_381);
nand U63 (N_63,In_5,In_38);
nand U64 (N_64,In_137,In_252);
xnor U65 (N_65,In_122,In_94);
or U66 (N_66,In_822,In_909);
nor U67 (N_67,In_341,In_783);
nand U68 (N_68,In_293,In_62);
or U69 (N_69,In_960,In_118);
nor U70 (N_70,In_276,In_15);
nand U71 (N_71,In_105,In_516);
nor U72 (N_72,In_46,In_346);
nor U73 (N_73,In_56,In_780);
nand U74 (N_74,In_522,In_415);
nor U75 (N_75,In_556,In_511);
and U76 (N_76,In_966,In_3);
xnor U77 (N_77,In_829,In_325);
and U78 (N_78,In_866,In_505);
and U79 (N_79,In_527,In_512);
nor U80 (N_80,In_320,In_856);
nor U81 (N_81,In_218,In_804);
or U82 (N_82,In_407,In_921);
nor U83 (N_83,In_794,In_715);
or U84 (N_84,In_400,In_492);
nor U85 (N_85,In_142,In_300);
nor U86 (N_86,In_337,In_652);
nor U87 (N_87,In_977,In_455);
nand U88 (N_88,In_161,In_378);
xor U89 (N_89,In_190,In_819);
or U90 (N_90,In_143,In_368);
and U91 (N_91,In_36,In_107);
and U92 (N_92,In_850,In_536);
nand U93 (N_93,In_825,In_543);
nand U94 (N_94,In_885,In_690);
and U95 (N_95,In_335,In_45);
xnor U96 (N_96,In_119,In_836);
or U97 (N_97,In_91,In_176);
xnor U98 (N_98,In_979,In_656);
or U99 (N_99,In_21,In_302);
nand U100 (N_100,In_154,In_597);
nor U101 (N_101,In_818,In_414);
nand U102 (N_102,In_840,In_682);
and U103 (N_103,In_813,In_399);
or U104 (N_104,In_980,In_196);
or U105 (N_105,In_236,In_771);
nor U106 (N_106,In_371,In_277);
nor U107 (N_107,In_25,In_531);
nand U108 (N_108,In_729,In_259);
nor U109 (N_109,In_478,In_558);
or U110 (N_110,In_116,In_348);
and U111 (N_111,In_164,In_338);
or U112 (N_112,In_132,In_759);
nor U113 (N_113,In_427,In_826);
nand U114 (N_114,In_723,In_925);
nand U115 (N_115,In_460,In_601);
nand U116 (N_116,In_489,In_621);
or U117 (N_117,In_653,In_857);
or U118 (N_118,In_491,In_767);
and U119 (N_119,In_534,In_576);
and U120 (N_120,In_446,In_355);
nor U121 (N_121,In_681,In_648);
xnor U122 (N_122,In_185,In_875);
nand U123 (N_123,In_148,In_228);
or U124 (N_124,In_490,In_903);
or U125 (N_125,In_862,In_789);
nand U126 (N_126,In_612,In_12);
and U127 (N_127,In_162,In_452);
nor U128 (N_128,In_719,In_265);
and U129 (N_129,In_959,In_608);
nor U130 (N_130,In_817,In_766);
nor U131 (N_131,In_778,In_736);
nand U132 (N_132,In_902,In_806);
and U133 (N_133,In_777,In_784);
nand U134 (N_134,In_71,In_312);
nor U135 (N_135,In_987,In_287);
nor U136 (N_136,In_238,In_565);
or U137 (N_137,In_832,In_217);
nor U138 (N_138,In_650,In_340);
and U139 (N_139,In_474,In_847);
nand U140 (N_140,In_508,In_611);
or U141 (N_141,In_546,In_952);
nor U142 (N_142,In_718,In_37);
nand U143 (N_143,In_750,In_581);
and U144 (N_144,In_879,In_403);
or U145 (N_145,In_223,In_754);
and U146 (N_146,In_8,In_192);
nand U147 (N_147,In_10,In_870);
or U148 (N_148,In_580,In_863);
nand U149 (N_149,In_891,In_125);
and U150 (N_150,In_391,In_904);
or U151 (N_151,In_711,In_470);
xnor U152 (N_152,In_502,In_245);
or U153 (N_153,In_423,In_13);
xor U154 (N_154,In_709,In_257);
nand U155 (N_155,In_573,In_471);
nor U156 (N_156,In_934,In_227);
or U157 (N_157,In_173,In_108);
or U158 (N_158,In_129,In_998);
and U159 (N_159,In_532,In_336);
nor U160 (N_160,In_643,In_795);
nor U161 (N_161,In_200,In_398);
or U162 (N_162,In_619,In_792);
and U163 (N_163,In_640,In_53);
and U164 (N_164,In_575,In_453);
and U165 (N_165,In_35,In_821);
or U166 (N_166,In_121,In_803);
and U167 (N_167,In_938,In_589);
nand U168 (N_168,In_753,In_698);
nand U169 (N_169,In_663,In_738);
xor U170 (N_170,In_254,In_30);
and U171 (N_171,In_625,In_297);
nor U172 (N_172,In_975,In_450);
or U173 (N_173,In_291,In_385);
nand U174 (N_174,In_897,In_389);
nor U175 (N_175,In_90,In_243);
and U176 (N_176,In_797,In_660);
nor U177 (N_177,In_641,In_842);
nor U178 (N_178,In_367,In_742);
or U179 (N_179,In_867,In_569);
or U180 (N_180,In_387,In_97);
xor U181 (N_181,In_131,In_726);
or U182 (N_182,In_635,In_790);
nand U183 (N_183,In_628,In_417);
xnor U184 (N_184,In_786,In_808);
or U185 (N_185,In_95,In_295);
or U186 (N_186,In_544,In_144);
nor U187 (N_187,In_883,In_503);
nand U188 (N_188,In_234,In_486);
nand U189 (N_189,In_275,In_473);
xor U190 (N_190,In_331,In_616);
xnor U191 (N_191,In_333,In_855);
nor U192 (N_192,In_272,In_128);
nand U193 (N_193,In_466,In_298);
xnor U194 (N_194,In_940,In_482);
and U195 (N_195,In_28,In_454);
nor U196 (N_196,In_55,In_746);
or U197 (N_197,In_271,In_815);
nand U198 (N_198,In_869,In_342);
xor U199 (N_199,In_535,In_993);
nor U200 (N_200,In_20,In_706);
nand U201 (N_201,In_278,In_997);
nand U202 (N_202,In_345,In_755);
and U203 (N_203,In_306,In_927);
nor U204 (N_204,In_213,In_447);
nand U205 (N_205,In_199,In_226);
and U206 (N_206,In_397,In_457);
nor U207 (N_207,In_170,In_865);
nor U208 (N_208,In_135,In_315);
xnor U209 (N_209,In_123,In_476);
or U210 (N_210,In_620,In_689);
or U211 (N_211,In_448,In_554);
nand U212 (N_212,In_802,In_622);
nand U213 (N_213,In_24,In_837);
or U214 (N_214,In_721,In_432);
nand U215 (N_215,In_11,In_433);
and U216 (N_216,In_89,In_773);
nand U217 (N_217,In_67,In_354);
nand U218 (N_218,In_919,In_500);
xnor U219 (N_219,In_0,In_487);
nand U220 (N_220,In_263,In_421);
and U221 (N_221,In_555,In_372);
or U222 (N_222,In_393,In_509);
nand U223 (N_223,In_47,In_379);
nor U224 (N_224,In_989,In_214);
and U225 (N_225,In_893,In_846);
and U226 (N_226,In_48,In_413);
and U227 (N_227,In_545,In_664);
or U228 (N_228,In_976,In_382);
xor U229 (N_229,In_79,In_110);
and U230 (N_230,In_568,In_657);
or U231 (N_231,In_26,In_395);
nand U232 (N_232,In_592,In_66);
or U233 (N_233,In_283,In_933);
and U234 (N_234,In_936,In_896);
nand U235 (N_235,In_359,In_582);
nor U236 (N_236,In_409,In_964);
and U237 (N_237,In_552,In_313);
or U238 (N_238,In_201,In_849);
or U239 (N_239,In_538,In_990);
nand U240 (N_240,In_932,In_41);
nor U241 (N_241,In_907,In_205);
or U242 (N_242,In_324,In_260);
or U243 (N_243,In_134,In_603);
nand U244 (N_244,In_262,In_58);
or U245 (N_245,In_184,In_456);
or U246 (N_246,In_186,In_969);
xor U247 (N_247,In_230,In_499);
xnor U248 (N_248,In_563,In_120);
nand U249 (N_249,In_593,In_714);
nor U250 (N_250,In_730,In_973);
nand U251 (N_251,In_189,In_244);
nand U252 (N_252,In_316,In_188);
and U253 (N_253,In_14,In_688);
or U254 (N_254,In_624,In_947);
or U255 (N_255,In_364,In_443);
nand U256 (N_256,In_811,In_310);
or U257 (N_257,In_844,In_687);
nand U258 (N_258,In_670,In_496);
xor U259 (N_259,In_655,In_733);
or U260 (N_260,In_60,In_584);
nor U261 (N_261,In_225,In_136);
nand U262 (N_262,In_422,In_126);
nor U263 (N_263,In_595,In_284);
and U264 (N_264,In_988,In_326);
and U265 (N_265,In_661,In_756);
xor U266 (N_266,In_361,In_805);
or U267 (N_267,In_197,In_63);
nor U268 (N_268,In_177,In_317);
nand U269 (N_269,In_629,In_525);
or U270 (N_270,In_329,In_133);
nor U271 (N_271,In_281,In_370);
nand U272 (N_272,In_945,In_984);
and U273 (N_273,In_768,In_93);
nor U274 (N_274,In_542,In_350);
or U275 (N_275,In_524,In_319);
or U276 (N_276,In_145,In_65);
and U277 (N_277,In_944,In_294);
nor U278 (N_278,In_156,In_712);
nand U279 (N_279,In_100,In_760);
or U280 (N_280,In_550,In_72);
nor U281 (N_281,In_716,In_831);
and U282 (N_282,In_181,In_17);
and U283 (N_283,In_878,In_528);
or U284 (N_284,In_465,In_735);
or U285 (N_285,In_138,In_519);
nand U286 (N_286,In_533,In_985);
xor U287 (N_287,In_436,In_559);
or U288 (N_288,In_801,In_438);
or U289 (N_289,In_820,In_510);
and U290 (N_290,In_665,In_739);
or U291 (N_291,In_720,In_861);
nor U292 (N_292,In_461,In_713);
or U293 (N_293,In_299,In_375);
or U294 (N_294,In_467,In_179);
nand U295 (N_295,In_599,In_810);
or U296 (N_296,In_130,In_437);
or U297 (N_297,In_369,In_685);
nand U298 (N_298,In_732,In_540);
nand U299 (N_299,In_587,In_406);
or U300 (N_300,In_80,In_917);
xor U301 (N_301,In_741,In_153);
or U302 (N_302,In_693,In_649);
or U303 (N_303,In_363,In_146);
nor U304 (N_304,In_737,In_775);
nor U305 (N_305,In_905,In_113);
nand U306 (N_306,In_73,In_250);
and U307 (N_307,In_241,In_541);
or U308 (N_308,In_602,In_662);
nand U309 (N_309,In_900,In_373);
nand U310 (N_310,In_914,In_751);
nor U311 (N_311,In_701,In_967);
nand U312 (N_312,In_557,In_703);
or U313 (N_313,In_675,In_991);
or U314 (N_314,In_282,In_594);
xor U315 (N_315,In_954,In_224);
and U316 (N_316,In_539,In_112);
xor U317 (N_317,In_155,In_928);
or U318 (N_318,In_671,In_64);
and U319 (N_319,In_210,In_212);
or U320 (N_320,In_632,In_408);
nand U321 (N_321,In_290,In_42);
and U322 (N_322,In_308,In_416);
nor U323 (N_323,In_209,In_674);
or U324 (N_324,In_974,In_982);
nor U325 (N_325,In_104,In_686);
nand U326 (N_326,In_852,In_659);
nor U327 (N_327,In_231,In_668);
or U328 (N_328,In_195,In_51);
nand U329 (N_329,In_859,In_75);
and U330 (N_330,In_357,In_304);
and U331 (N_331,In_561,In_972);
nor U332 (N_332,In_388,In_647);
nand U333 (N_333,In_877,In_157);
and U334 (N_334,In_307,In_248);
or U335 (N_335,In_950,In_33);
and U336 (N_336,In_349,In_923);
nor U337 (N_337,In_955,In_610);
or U338 (N_338,In_705,In_910);
and U339 (N_339,In_251,In_410);
nor U340 (N_340,In_695,In_40);
or U341 (N_341,In_6,In_931);
nand U342 (N_342,In_358,In_32);
or U343 (N_343,In_420,In_633);
and U344 (N_344,In_963,In_258);
nand U345 (N_345,In_229,In_604);
or U346 (N_346,In_949,In_360);
nand U347 (N_347,In_645,In_288);
and U348 (N_348,In_788,In_605);
nand U349 (N_349,In_1,In_762);
nand U350 (N_350,In_876,In_279);
or U351 (N_351,In_710,In_956);
nor U352 (N_352,In_507,In_669);
nand U353 (N_353,In_160,In_679);
or U354 (N_354,In_970,In_757);
nand U355 (N_355,In_202,In_183);
nor U356 (N_356,In_428,In_484);
nand U357 (N_357,In_330,In_567);
and U358 (N_358,In_725,In_412);
nand U359 (N_359,In_667,In_34);
and U360 (N_360,In_431,In_139);
and U361 (N_361,In_579,In_779);
or U362 (N_362,In_607,In_390);
nand U363 (N_363,In_798,In_419);
nor U364 (N_364,In_631,In_274);
nor U365 (N_365,In_600,In_311);
or U366 (N_366,In_380,In_493);
nor U367 (N_367,In_39,In_680);
nor U368 (N_368,In_194,In_140);
nor U369 (N_369,In_613,In_61);
and U370 (N_370,In_995,In_401);
nand U371 (N_371,In_948,In_943);
nor U372 (N_372,In_49,In_747);
or U373 (N_373,In_318,In_115);
nand U374 (N_374,In_560,In_743);
nand U375 (N_375,In_684,In_85);
and U376 (N_376,In_468,In_911);
nand U377 (N_377,In_240,In_426);
nor U378 (N_378,In_158,In_920);
or U379 (N_379,In_764,In_888);
nor U380 (N_380,In_570,In_16);
nand U381 (N_381,In_141,In_694);
and U382 (N_382,In_435,In_702);
or U383 (N_383,In_103,In_328);
and U384 (N_384,In_356,In_774);
and U385 (N_385,In_464,In_971);
or U386 (N_386,In_636,In_585);
and U387 (N_387,In_796,In_255);
and U388 (N_388,In_639,In_981);
or U389 (N_389,In_642,In_292);
nand U390 (N_390,In_651,In_941);
or U391 (N_391,In_835,In_377);
and U392 (N_392,In_449,In_459);
nand U393 (N_393,In_666,In_586);
xnor U394 (N_394,In_734,In_102);
and U395 (N_395,In_458,In_480);
or U396 (N_396,In_77,In_722);
nand U397 (N_397,In_424,In_445);
nand U398 (N_398,In_700,In_884);
or U399 (N_399,In_691,In_785);
nand U400 (N_400,In_965,In_463);
and U401 (N_401,In_88,In_405);
and U402 (N_402,In_83,In_547);
and U403 (N_403,In_763,In_770);
or U404 (N_404,In_221,In_485);
and U405 (N_405,In_74,In_807);
nand U406 (N_406,In_574,In_498);
nor U407 (N_407,In_261,In_566);
and U408 (N_408,In_273,In_860);
and U409 (N_409,In_246,In_50);
nor U410 (N_410,In_617,In_305);
xor U411 (N_411,In_873,In_78);
nand U412 (N_412,In_479,In_752);
nand U413 (N_413,In_321,In_598);
nand U414 (N_414,In_838,In_551);
or U415 (N_415,In_913,In_571);
nor U416 (N_416,In_696,In_440);
or U417 (N_417,In_172,In_915);
nor U418 (N_418,In_81,In_150);
nor U419 (N_419,In_206,In_147);
xnor U420 (N_420,In_477,In_929);
nand U421 (N_421,In_269,In_175);
and U422 (N_422,In_881,In_166);
or U423 (N_423,In_69,In_57);
nand U424 (N_424,In_7,In_124);
nor U425 (N_425,In_247,In_992);
and U426 (N_426,In_23,In_169);
nor U427 (N_427,In_441,In_781);
and U428 (N_428,In_782,In_264);
nand U429 (N_429,In_583,In_731);
and U430 (N_430,In_2,In_880);
nor U431 (N_431,In_638,In_745);
or U432 (N_432,In_286,In_615);
nand U433 (N_433,In_314,In_614);
and U434 (N_434,In_922,In_874);
nand U435 (N_435,In_596,In_833);
or U436 (N_436,In_577,In_830);
xnor U437 (N_437,In_268,In_339);
nor U438 (N_438,In_220,In_222);
or U439 (N_439,In_654,In_362);
nand U440 (N_440,In_898,In_851);
nand U441 (N_441,In_462,In_886);
and U442 (N_442,In_697,In_926);
nand U443 (N_443,In_996,In_704);
or U444 (N_444,In_890,In_787);
or U445 (N_445,In_506,In_270);
or U446 (N_446,In_351,In_912);
and U447 (N_447,In_526,In_827);
or U448 (N_448,In_296,In_168);
nand U449 (N_449,In_676,In_606);
xnor U450 (N_450,In_256,In_908);
or U451 (N_451,In_418,In_327);
and U452 (N_452,In_332,In_198);
nand U453 (N_453,In_520,In_868);
and U454 (N_454,In_537,In_303);
nand U455 (N_455,In_749,In_117);
and U456 (N_456,In_521,In_174);
or U457 (N_457,In_86,In_864);
nor U458 (N_458,In_280,In_215);
nor U459 (N_459,In_266,In_962);
nand U460 (N_460,In_301,In_590);
and U461 (N_461,In_242,In_727);
and U462 (N_462,In_180,In_52);
nand U463 (N_463,In_673,In_809);
or U464 (N_464,In_165,In_812);
or U465 (N_465,In_495,In_549);
nor U466 (N_466,In_235,In_207);
xnor U467 (N_467,In_203,In_396);
nand U468 (N_468,In_9,In_159);
xor U469 (N_469,In_167,In_515);
nor U470 (N_470,In_894,In_758);
nor U471 (N_471,In_627,In_178);
or U472 (N_472,In_935,In_772);
or U473 (N_473,In_816,In_392);
or U474 (N_474,In_54,In_776);
or U475 (N_475,In_219,In_309);
nand U476 (N_476,In_404,In_708);
nor U477 (N_477,In_347,In_978);
nor U478 (N_478,In_334,In_386);
or U479 (N_479,In_924,In_472);
and U480 (N_480,In_895,In_983);
and U481 (N_481,In_823,In_106);
nor U482 (N_482,In_793,In_475);
or U483 (N_483,In_383,In_530);
nor U484 (N_484,In_171,In_366);
nand U485 (N_485,In_523,In_839);
and U486 (N_486,In_98,In_76);
and U487 (N_487,In_692,In_644);
xnor U488 (N_488,In_82,In_481);
and U489 (N_489,In_824,In_92);
nand U490 (N_490,In_887,In_44);
xnor U491 (N_491,In_578,In_843);
xor U492 (N_492,In_343,In_193);
xnor U493 (N_493,In_564,In_187);
nor U494 (N_494,In_239,In_501);
nor U495 (N_495,In_529,In_151);
nor U496 (N_496,In_494,In_769);
or U497 (N_497,In_672,In_953);
and U498 (N_498,In_618,In_434);
nand U499 (N_499,In_609,In_68);
nand U500 (N_500,In_560,In_277);
nor U501 (N_501,In_629,In_850);
or U502 (N_502,In_905,In_108);
or U503 (N_503,In_51,In_143);
nand U504 (N_504,In_741,In_249);
nor U505 (N_505,In_34,In_262);
and U506 (N_506,In_714,In_162);
or U507 (N_507,In_582,In_62);
nor U508 (N_508,In_858,In_493);
or U509 (N_509,In_913,In_770);
and U510 (N_510,In_432,In_175);
nand U511 (N_511,In_58,In_814);
nor U512 (N_512,In_676,In_478);
and U513 (N_513,In_495,In_785);
nand U514 (N_514,In_967,In_679);
nand U515 (N_515,In_223,In_319);
nor U516 (N_516,In_399,In_240);
nand U517 (N_517,In_550,In_748);
and U518 (N_518,In_577,In_50);
nand U519 (N_519,In_799,In_69);
or U520 (N_520,In_502,In_401);
nand U521 (N_521,In_975,In_638);
xor U522 (N_522,In_978,In_291);
nor U523 (N_523,In_851,In_226);
nand U524 (N_524,In_920,In_303);
xor U525 (N_525,In_417,In_158);
and U526 (N_526,In_186,In_582);
nand U527 (N_527,In_650,In_456);
nand U528 (N_528,In_268,In_411);
nor U529 (N_529,In_492,In_554);
nand U530 (N_530,In_557,In_517);
or U531 (N_531,In_105,In_252);
nor U532 (N_532,In_227,In_756);
nor U533 (N_533,In_266,In_745);
nand U534 (N_534,In_779,In_641);
nand U535 (N_535,In_387,In_213);
and U536 (N_536,In_678,In_52);
nand U537 (N_537,In_622,In_565);
or U538 (N_538,In_264,In_309);
nor U539 (N_539,In_667,In_851);
nor U540 (N_540,In_711,In_638);
nand U541 (N_541,In_5,In_6);
and U542 (N_542,In_611,In_433);
or U543 (N_543,In_743,In_285);
or U544 (N_544,In_737,In_969);
nor U545 (N_545,In_655,In_918);
or U546 (N_546,In_799,In_786);
nor U547 (N_547,In_674,In_447);
and U548 (N_548,In_739,In_362);
or U549 (N_549,In_923,In_957);
or U550 (N_550,In_702,In_590);
nor U551 (N_551,In_266,In_270);
and U552 (N_552,In_849,In_155);
nor U553 (N_553,In_185,In_239);
and U554 (N_554,In_980,In_937);
xor U555 (N_555,In_578,In_182);
or U556 (N_556,In_191,In_666);
or U557 (N_557,In_950,In_184);
nor U558 (N_558,In_180,In_369);
or U559 (N_559,In_47,In_213);
and U560 (N_560,In_631,In_115);
nand U561 (N_561,In_827,In_501);
or U562 (N_562,In_610,In_483);
or U563 (N_563,In_70,In_179);
nand U564 (N_564,In_213,In_991);
or U565 (N_565,In_451,In_428);
nand U566 (N_566,In_997,In_701);
or U567 (N_567,In_14,In_39);
and U568 (N_568,In_369,In_392);
and U569 (N_569,In_321,In_902);
or U570 (N_570,In_730,In_822);
and U571 (N_571,In_79,In_198);
or U572 (N_572,In_869,In_518);
nand U573 (N_573,In_575,In_497);
nor U574 (N_574,In_237,In_723);
nand U575 (N_575,In_713,In_551);
or U576 (N_576,In_37,In_398);
xor U577 (N_577,In_460,In_182);
nand U578 (N_578,In_117,In_232);
nand U579 (N_579,In_71,In_804);
and U580 (N_580,In_582,In_787);
nor U581 (N_581,In_953,In_876);
nor U582 (N_582,In_463,In_731);
nand U583 (N_583,In_580,In_143);
or U584 (N_584,In_214,In_927);
and U585 (N_585,In_161,In_372);
or U586 (N_586,In_459,In_75);
nand U587 (N_587,In_164,In_576);
nor U588 (N_588,In_932,In_955);
xnor U589 (N_589,In_553,In_489);
nor U590 (N_590,In_491,In_574);
and U591 (N_591,In_264,In_709);
xnor U592 (N_592,In_113,In_50);
nand U593 (N_593,In_786,In_258);
nand U594 (N_594,In_389,In_237);
nand U595 (N_595,In_624,In_558);
or U596 (N_596,In_192,In_401);
and U597 (N_597,In_73,In_206);
xor U598 (N_598,In_998,In_46);
nor U599 (N_599,In_759,In_705);
and U600 (N_600,In_225,In_901);
and U601 (N_601,In_656,In_458);
xor U602 (N_602,In_231,In_136);
or U603 (N_603,In_847,In_253);
nand U604 (N_604,In_184,In_820);
nand U605 (N_605,In_392,In_400);
nand U606 (N_606,In_189,In_450);
nor U607 (N_607,In_148,In_668);
nand U608 (N_608,In_782,In_856);
and U609 (N_609,In_451,In_57);
nand U610 (N_610,In_644,In_475);
nor U611 (N_611,In_244,In_768);
or U612 (N_612,In_820,In_241);
or U613 (N_613,In_24,In_928);
nor U614 (N_614,In_311,In_255);
nand U615 (N_615,In_54,In_583);
and U616 (N_616,In_97,In_85);
nor U617 (N_617,In_291,In_713);
and U618 (N_618,In_545,In_930);
nand U619 (N_619,In_380,In_973);
xor U620 (N_620,In_562,In_481);
nor U621 (N_621,In_213,In_801);
nor U622 (N_622,In_988,In_835);
xnor U623 (N_623,In_161,In_819);
nand U624 (N_624,In_782,In_515);
or U625 (N_625,In_620,In_406);
and U626 (N_626,In_631,In_794);
xor U627 (N_627,In_78,In_878);
nor U628 (N_628,In_2,In_428);
nand U629 (N_629,In_277,In_236);
nor U630 (N_630,In_488,In_311);
and U631 (N_631,In_30,In_318);
xnor U632 (N_632,In_937,In_108);
and U633 (N_633,In_806,In_605);
nand U634 (N_634,In_922,In_148);
nand U635 (N_635,In_965,In_592);
and U636 (N_636,In_493,In_12);
nor U637 (N_637,In_292,In_310);
nor U638 (N_638,In_382,In_219);
and U639 (N_639,In_529,In_866);
nor U640 (N_640,In_611,In_786);
and U641 (N_641,In_392,In_308);
nor U642 (N_642,In_979,In_417);
nor U643 (N_643,In_584,In_306);
or U644 (N_644,In_490,In_266);
nor U645 (N_645,In_40,In_172);
xor U646 (N_646,In_375,In_31);
or U647 (N_647,In_972,In_823);
or U648 (N_648,In_259,In_439);
nor U649 (N_649,In_437,In_358);
and U650 (N_650,In_81,In_382);
or U651 (N_651,In_868,In_144);
nor U652 (N_652,In_956,In_929);
nor U653 (N_653,In_173,In_739);
nor U654 (N_654,In_580,In_135);
or U655 (N_655,In_185,In_85);
or U656 (N_656,In_654,In_128);
nand U657 (N_657,In_48,In_15);
nand U658 (N_658,In_552,In_419);
nand U659 (N_659,In_390,In_394);
xor U660 (N_660,In_975,In_973);
nand U661 (N_661,In_151,In_877);
xor U662 (N_662,In_968,In_508);
xor U663 (N_663,In_630,In_923);
nand U664 (N_664,In_621,In_210);
or U665 (N_665,In_725,In_99);
or U666 (N_666,In_130,In_65);
nor U667 (N_667,In_439,In_224);
nor U668 (N_668,In_851,In_204);
nor U669 (N_669,In_573,In_197);
nand U670 (N_670,In_603,In_5);
nor U671 (N_671,In_785,In_478);
nor U672 (N_672,In_495,In_239);
nand U673 (N_673,In_713,In_322);
xnor U674 (N_674,In_636,In_567);
nor U675 (N_675,In_772,In_185);
and U676 (N_676,In_386,In_65);
or U677 (N_677,In_158,In_485);
xnor U678 (N_678,In_288,In_196);
nor U679 (N_679,In_824,In_227);
nand U680 (N_680,In_997,In_509);
nand U681 (N_681,In_990,In_466);
nor U682 (N_682,In_668,In_31);
or U683 (N_683,In_534,In_395);
nand U684 (N_684,In_599,In_367);
and U685 (N_685,In_936,In_406);
and U686 (N_686,In_327,In_607);
or U687 (N_687,In_152,In_764);
nor U688 (N_688,In_634,In_922);
and U689 (N_689,In_332,In_897);
and U690 (N_690,In_316,In_931);
and U691 (N_691,In_643,In_76);
nor U692 (N_692,In_50,In_82);
nand U693 (N_693,In_2,In_27);
or U694 (N_694,In_479,In_124);
nor U695 (N_695,In_90,In_884);
nand U696 (N_696,In_870,In_539);
xnor U697 (N_697,In_655,In_159);
or U698 (N_698,In_945,In_675);
or U699 (N_699,In_658,In_875);
nor U700 (N_700,In_885,In_80);
and U701 (N_701,In_633,In_43);
nand U702 (N_702,In_525,In_739);
xnor U703 (N_703,In_930,In_876);
and U704 (N_704,In_709,In_659);
nor U705 (N_705,In_659,In_749);
or U706 (N_706,In_340,In_331);
or U707 (N_707,In_696,In_557);
or U708 (N_708,In_977,In_118);
or U709 (N_709,In_781,In_584);
and U710 (N_710,In_667,In_739);
and U711 (N_711,In_533,In_359);
and U712 (N_712,In_423,In_88);
nor U713 (N_713,In_833,In_471);
nor U714 (N_714,In_450,In_200);
or U715 (N_715,In_235,In_150);
nand U716 (N_716,In_491,In_404);
nand U717 (N_717,In_309,In_74);
or U718 (N_718,In_919,In_65);
and U719 (N_719,In_697,In_281);
or U720 (N_720,In_319,In_230);
nand U721 (N_721,In_831,In_607);
nand U722 (N_722,In_41,In_832);
and U723 (N_723,In_877,In_655);
nand U724 (N_724,In_360,In_36);
nand U725 (N_725,In_822,In_811);
nand U726 (N_726,In_676,In_746);
nand U727 (N_727,In_270,In_913);
and U728 (N_728,In_806,In_416);
nor U729 (N_729,In_878,In_834);
xor U730 (N_730,In_205,In_254);
nand U731 (N_731,In_874,In_128);
nor U732 (N_732,In_264,In_878);
and U733 (N_733,In_886,In_961);
nand U734 (N_734,In_287,In_901);
nand U735 (N_735,In_759,In_500);
or U736 (N_736,In_55,In_569);
and U737 (N_737,In_829,In_165);
nand U738 (N_738,In_819,In_330);
or U739 (N_739,In_682,In_638);
nor U740 (N_740,In_192,In_753);
and U741 (N_741,In_46,In_485);
and U742 (N_742,In_802,In_226);
and U743 (N_743,In_957,In_455);
or U744 (N_744,In_658,In_353);
or U745 (N_745,In_110,In_505);
or U746 (N_746,In_824,In_823);
nand U747 (N_747,In_797,In_852);
or U748 (N_748,In_545,In_122);
nor U749 (N_749,In_150,In_44);
nor U750 (N_750,In_995,In_486);
nand U751 (N_751,In_683,In_398);
nor U752 (N_752,In_762,In_951);
nand U753 (N_753,In_397,In_496);
nand U754 (N_754,In_786,In_52);
xnor U755 (N_755,In_46,In_297);
and U756 (N_756,In_172,In_820);
or U757 (N_757,In_421,In_338);
or U758 (N_758,In_963,In_309);
nor U759 (N_759,In_567,In_54);
or U760 (N_760,In_962,In_576);
nor U761 (N_761,In_314,In_340);
nand U762 (N_762,In_331,In_263);
nor U763 (N_763,In_243,In_177);
and U764 (N_764,In_91,In_971);
or U765 (N_765,In_447,In_925);
nand U766 (N_766,In_796,In_451);
nor U767 (N_767,In_562,In_477);
and U768 (N_768,In_196,In_331);
or U769 (N_769,In_746,In_23);
and U770 (N_770,In_417,In_217);
or U771 (N_771,In_325,In_833);
and U772 (N_772,In_635,In_453);
nand U773 (N_773,In_782,In_409);
or U774 (N_774,In_632,In_805);
xor U775 (N_775,In_924,In_812);
nor U776 (N_776,In_63,In_984);
and U777 (N_777,In_359,In_78);
nand U778 (N_778,In_788,In_870);
and U779 (N_779,In_427,In_396);
nor U780 (N_780,In_228,In_973);
or U781 (N_781,In_356,In_763);
nand U782 (N_782,In_270,In_373);
nand U783 (N_783,In_306,In_883);
xor U784 (N_784,In_794,In_321);
or U785 (N_785,In_992,In_491);
and U786 (N_786,In_259,In_472);
nor U787 (N_787,In_508,In_679);
xnor U788 (N_788,In_936,In_634);
nand U789 (N_789,In_428,In_610);
nor U790 (N_790,In_233,In_550);
nor U791 (N_791,In_828,In_497);
and U792 (N_792,In_240,In_577);
nand U793 (N_793,In_622,In_964);
and U794 (N_794,In_391,In_93);
nand U795 (N_795,In_755,In_415);
nand U796 (N_796,In_529,In_667);
xnor U797 (N_797,In_204,In_323);
xor U798 (N_798,In_783,In_242);
nand U799 (N_799,In_16,In_975);
and U800 (N_800,In_561,In_930);
xnor U801 (N_801,In_251,In_348);
nand U802 (N_802,In_710,In_698);
or U803 (N_803,In_229,In_871);
nor U804 (N_804,In_997,In_955);
nor U805 (N_805,In_447,In_145);
nor U806 (N_806,In_837,In_998);
nand U807 (N_807,In_538,In_770);
or U808 (N_808,In_757,In_928);
and U809 (N_809,In_563,In_825);
and U810 (N_810,In_66,In_297);
and U811 (N_811,In_349,In_880);
nor U812 (N_812,In_224,In_164);
or U813 (N_813,In_573,In_831);
nand U814 (N_814,In_11,In_720);
nand U815 (N_815,In_328,In_139);
nand U816 (N_816,In_805,In_785);
and U817 (N_817,In_352,In_152);
and U818 (N_818,In_774,In_159);
or U819 (N_819,In_850,In_945);
nor U820 (N_820,In_949,In_52);
xor U821 (N_821,In_899,In_602);
nand U822 (N_822,In_162,In_113);
xor U823 (N_823,In_2,In_434);
and U824 (N_824,In_890,In_18);
nor U825 (N_825,In_51,In_172);
or U826 (N_826,In_31,In_426);
nand U827 (N_827,In_956,In_774);
nor U828 (N_828,In_976,In_361);
xnor U829 (N_829,In_103,In_284);
nor U830 (N_830,In_630,In_794);
nor U831 (N_831,In_564,In_907);
or U832 (N_832,In_929,In_50);
or U833 (N_833,In_971,In_252);
or U834 (N_834,In_413,In_786);
nor U835 (N_835,In_861,In_287);
and U836 (N_836,In_586,In_383);
nor U837 (N_837,In_910,In_515);
xor U838 (N_838,In_244,In_41);
and U839 (N_839,In_237,In_278);
and U840 (N_840,In_359,In_119);
xnor U841 (N_841,In_532,In_234);
xor U842 (N_842,In_712,In_286);
nand U843 (N_843,In_180,In_216);
nand U844 (N_844,In_0,In_32);
or U845 (N_845,In_837,In_801);
and U846 (N_846,In_811,In_96);
nor U847 (N_847,In_50,In_582);
or U848 (N_848,In_291,In_398);
nand U849 (N_849,In_158,In_748);
nor U850 (N_850,In_992,In_967);
nor U851 (N_851,In_618,In_225);
or U852 (N_852,In_892,In_830);
nand U853 (N_853,In_919,In_468);
xnor U854 (N_854,In_973,In_830);
xnor U855 (N_855,In_582,In_774);
and U856 (N_856,In_147,In_280);
nor U857 (N_857,In_854,In_406);
nand U858 (N_858,In_240,In_985);
nand U859 (N_859,In_858,In_519);
and U860 (N_860,In_62,In_249);
nor U861 (N_861,In_588,In_667);
and U862 (N_862,In_648,In_564);
or U863 (N_863,In_702,In_823);
nor U864 (N_864,In_735,In_846);
and U865 (N_865,In_820,In_803);
nand U866 (N_866,In_724,In_34);
or U867 (N_867,In_404,In_617);
nand U868 (N_868,In_799,In_519);
nor U869 (N_869,In_336,In_157);
nor U870 (N_870,In_495,In_849);
and U871 (N_871,In_316,In_58);
nor U872 (N_872,In_573,In_375);
or U873 (N_873,In_226,In_447);
nand U874 (N_874,In_819,In_995);
and U875 (N_875,In_25,In_491);
nand U876 (N_876,In_305,In_69);
nor U877 (N_877,In_885,In_937);
and U878 (N_878,In_515,In_537);
nor U879 (N_879,In_799,In_40);
xor U880 (N_880,In_400,In_516);
and U881 (N_881,In_291,In_645);
xnor U882 (N_882,In_389,In_241);
or U883 (N_883,In_186,In_21);
xnor U884 (N_884,In_682,In_750);
nand U885 (N_885,In_210,In_879);
nor U886 (N_886,In_710,In_943);
nand U887 (N_887,In_454,In_823);
nor U888 (N_888,In_268,In_439);
or U889 (N_889,In_309,In_162);
and U890 (N_890,In_538,In_54);
or U891 (N_891,In_807,In_166);
or U892 (N_892,In_723,In_942);
nor U893 (N_893,In_613,In_345);
nand U894 (N_894,In_891,In_463);
or U895 (N_895,In_806,In_479);
nor U896 (N_896,In_859,In_421);
or U897 (N_897,In_109,In_56);
nor U898 (N_898,In_906,In_621);
and U899 (N_899,In_619,In_4);
or U900 (N_900,In_498,In_47);
xnor U901 (N_901,In_784,In_616);
and U902 (N_902,In_278,In_569);
and U903 (N_903,In_276,In_849);
xor U904 (N_904,In_600,In_308);
nor U905 (N_905,In_494,In_554);
and U906 (N_906,In_507,In_788);
and U907 (N_907,In_47,In_788);
nand U908 (N_908,In_468,In_931);
nand U909 (N_909,In_587,In_804);
nor U910 (N_910,In_876,In_218);
nor U911 (N_911,In_798,In_45);
or U912 (N_912,In_919,In_23);
and U913 (N_913,In_152,In_908);
nand U914 (N_914,In_919,In_715);
nor U915 (N_915,In_68,In_334);
xor U916 (N_916,In_722,In_464);
nand U917 (N_917,In_220,In_966);
nand U918 (N_918,In_216,In_33);
nand U919 (N_919,In_489,In_508);
nand U920 (N_920,In_970,In_295);
or U921 (N_921,In_429,In_553);
or U922 (N_922,In_826,In_713);
nand U923 (N_923,In_368,In_22);
and U924 (N_924,In_802,In_463);
nand U925 (N_925,In_657,In_830);
nand U926 (N_926,In_244,In_746);
xor U927 (N_927,In_717,In_542);
nor U928 (N_928,In_851,In_506);
or U929 (N_929,In_631,In_560);
nand U930 (N_930,In_134,In_941);
or U931 (N_931,In_492,In_685);
nor U932 (N_932,In_435,In_511);
and U933 (N_933,In_680,In_827);
nand U934 (N_934,In_750,In_861);
or U935 (N_935,In_703,In_615);
nor U936 (N_936,In_512,In_974);
or U937 (N_937,In_281,In_407);
and U938 (N_938,In_263,In_289);
or U939 (N_939,In_8,In_183);
nand U940 (N_940,In_308,In_808);
nand U941 (N_941,In_10,In_464);
nor U942 (N_942,In_88,In_279);
nand U943 (N_943,In_322,In_657);
or U944 (N_944,In_615,In_591);
nand U945 (N_945,In_463,In_113);
nand U946 (N_946,In_298,In_203);
nand U947 (N_947,In_470,In_697);
and U948 (N_948,In_44,In_658);
nand U949 (N_949,In_741,In_447);
xor U950 (N_950,In_426,In_194);
nand U951 (N_951,In_269,In_527);
xor U952 (N_952,In_606,In_623);
nor U953 (N_953,In_5,In_998);
nand U954 (N_954,In_336,In_201);
nand U955 (N_955,In_119,In_978);
nand U956 (N_956,In_271,In_594);
nor U957 (N_957,In_466,In_495);
or U958 (N_958,In_263,In_181);
xnor U959 (N_959,In_703,In_465);
and U960 (N_960,In_280,In_284);
and U961 (N_961,In_345,In_21);
or U962 (N_962,In_439,In_222);
nand U963 (N_963,In_91,In_28);
nor U964 (N_964,In_343,In_565);
and U965 (N_965,In_837,In_423);
nand U966 (N_966,In_608,In_328);
and U967 (N_967,In_912,In_867);
nand U968 (N_968,In_607,In_175);
and U969 (N_969,In_552,In_615);
nand U970 (N_970,In_756,In_521);
nand U971 (N_971,In_133,In_459);
and U972 (N_972,In_75,In_328);
nor U973 (N_973,In_767,In_927);
or U974 (N_974,In_988,In_246);
nand U975 (N_975,In_393,In_810);
or U976 (N_976,In_727,In_651);
or U977 (N_977,In_489,In_780);
or U978 (N_978,In_124,In_155);
and U979 (N_979,In_142,In_564);
xor U980 (N_980,In_744,In_526);
nor U981 (N_981,In_248,In_162);
and U982 (N_982,In_492,In_717);
nor U983 (N_983,In_254,In_884);
nor U984 (N_984,In_234,In_209);
nand U985 (N_985,In_898,In_401);
nor U986 (N_986,In_706,In_532);
and U987 (N_987,In_273,In_225);
and U988 (N_988,In_372,In_988);
xor U989 (N_989,In_49,In_874);
nand U990 (N_990,In_381,In_289);
and U991 (N_991,In_631,In_145);
xor U992 (N_992,In_962,In_95);
nor U993 (N_993,In_187,In_927);
nand U994 (N_994,In_899,In_353);
and U995 (N_995,In_278,In_575);
xor U996 (N_996,In_176,In_253);
nor U997 (N_997,In_688,In_85);
nand U998 (N_998,In_713,In_346);
nand U999 (N_999,In_192,In_73);
and U1000 (N_1000,In_97,In_613);
or U1001 (N_1001,In_723,In_181);
or U1002 (N_1002,In_918,In_92);
or U1003 (N_1003,In_621,In_289);
and U1004 (N_1004,In_267,In_596);
nand U1005 (N_1005,In_24,In_637);
nand U1006 (N_1006,In_767,In_26);
nand U1007 (N_1007,In_89,In_445);
nand U1008 (N_1008,In_383,In_336);
and U1009 (N_1009,In_479,In_260);
nor U1010 (N_1010,In_961,In_68);
or U1011 (N_1011,In_543,In_688);
nor U1012 (N_1012,In_390,In_540);
nand U1013 (N_1013,In_805,In_142);
nor U1014 (N_1014,In_536,In_144);
nand U1015 (N_1015,In_287,In_648);
or U1016 (N_1016,In_538,In_497);
and U1017 (N_1017,In_185,In_41);
and U1018 (N_1018,In_627,In_923);
xnor U1019 (N_1019,In_45,In_553);
and U1020 (N_1020,In_815,In_372);
or U1021 (N_1021,In_12,In_42);
nand U1022 (N_1022,In_879,In_721);
and U1023 (N_1023,In_186,In_792);
nand U1024 (N_1024,In_225,In_32);
and U1025 (N_1025,In_869,In_937);
and U1026 (N_1026,In_242,In_380);
nand U1027 (N_1027,In_589,In_20);
or U1028 (N_1028,In_876,In_236);
or U1029 (N_1029,In_605,In_306);
nor U1030 (N_1030,In_139,In_184);
nand U1031 (N_1031,In_267,In_910);
and U1032 (N_1032,In_452,In_416);
nor U1033 (N_1033,In_254,In_646);
nor U1034 (N_1034,In_738,In_276);
nor U1035 (N_1035,In_233,In_572);
nand U1036 (N_1036,In_34,In_18);
nor U1037 (N_1037,In_380,In_538);
nand U1038 (N_1038,In_638,In_29);
nor U1039 (N_1039,In_268,In_735);
nand U1040 (N_1040,In_0,In_914);
or U1041 (N_1041,In_84,In_845);
xor U1042 (N_1042,In_537,In_572);
xor U1043 (N_1043,In_986,In_624);
nor U1044 (N_1044,In_675,In_312);
or U1045 (N_1045,In_560,In_445);
nor U1046 (N_1046,In_123,In_937);
nor U1047 (N_1047,In_884,In_671);
nor U1048 (N_1048,In_28,In_394);
nand U1049 (N_1049,In_507,In_773);
xnor U1050 (N_1050,In_807,In_385);
and U1051 (N_1051,In_89,In_495);
nand U1052 (N_1052,In_186,In_307);
and U1053 (N_1053,In_998,In_806);
and U1054 (N_1054,In_987,In_610);
nor U1055 (N_1055,In_974,In_361);
and U1056 (N_1056,In_680,In_498);
xnor U1057 (N_1057,In_369,In_820);
nor U1058 (N_1058,In_172,In_338);
or U1059 (N_1059,In_74,In_34);
or U1060 (N_1060,In_707,In_651);
nor U1061 (N_1061,In_754,In_653);
and U1062 (N_1062,In_680,In_850);
and U1063 (N_1063,In_636,In_714);
nand U1064 (N_1064,In_639,In_180);
or U1065 (N_1065,In_667,In_454);
nor U1066 (N_1066,In_366,In_435);
and U1067 (N_1067,In_706,In_770);
or U1068 (N_1068,In_428,In_914);
nand U1069 (N_1069,In_539,In_44);
nand U1070 (N_1070,In_72,In_12);
and U1071 (N_1071,In_260,In_420);
nor U1072 (N_1072,In_442,In_298);
and U1073 (N_1073,In_733,In_55);
nand U1074 (N_1074,In_723,In_626);
or U1075 (N_1075,In_472,In_744);
or U1076 (N_1076,In_557,In_199);
or U1077 (N_1077,In_464,In_538);
or U1078 (N_1078,In_58,In_592);
xor U1079 (N_1079,In_39,In_85);
and U1080 (N_1080,In_395,In_802);
or U1081 (N_1081,In_24,In_55);
nand U1082 (N_1082,In_492,In_166);
and U1083 (N_1083,In_829,In_121);
and U1084 (N_1084,In_240,In_305);
nand U1085 (N_1085,In_772,In_800);
and U1086 (N_1086,In_185,In_790);
and U1087 (N_1087,In_122,In_386);
or U1088 (N_1088,In_899,In_264);
nor U1089 (N_1089,In_71,In_915);
xor U1090 (N_1090,In_429,In_557);
nor U1091 (N_1091,In_508,In_854);
xor U1092 (N_1092,In_639,In_785);
or U1093 (N_1093,In_55,In_189);
nor U1094 (N_1094,In_947,In_602);
or U1095 (N_1095,In_796,In_163);
nor U1096 (N_1096,In_379,In_574);
or U1097 (N_1097,In_510,In_993);
or U1098 (N_1098,In_931,In_269);
nor U1099 (N_1099,In_899,In_755);
nand U1100 (N_1100,In_240,In_96);
nand U1101 (N_1101,In_16,In_712);
nor U1102 (N_1102,In_543,In_545);
and U1103 (N_1103,In_652,In_983);
nand U1104 (N_1104,In_663,In_261);
nor U1105 (N_1105,In_378,In_784);
and U1106 (N_1106,In_239,In_895);
nor U1107 (N_1107,In_83,In_610);
or U1108 (N_1108,In_84,In_59);
or U1109 (N_1109,In_555,In_463);
nor U1110 (N_1110,In_360,In_397);
and U1111 (N_1111,In_137,In_585);
or U1112 (N_1112,In_730,In_65);
and U1113 (N_1113,In_9,In_106);
nor U1114 (N_1114,In_407,In_489);
nor U1115 (N_1115,In_930,In_640);
nand U1116 (N_1116,In_641,In_91);
or U1117 (N_1117,In_269,In_288);
and U1118 (N_1118,In_436,In_81);
and U1119 (N_1119,In_663,In_997);
and U1120 (N_1120,In_34,In_677);
nand U1121 (N_1121,In_91,In_800);
xnor U1122 (N_1122,In_62,In_521);
or U1123 (N_1123,In_678,In_128);
or U1124 (N_1124,In_197,In_832);
or U1125 (N_1125,In_951,In_222);
nor U1126 (N_1126,In_644,In_417);
and U1127 (N_1127,In_606,In_759);
nor U1128 (N_1128,In_792,In_266);
nand U1129 (N_1129,In_851,In_807);
and U1130 (N_1130,In_945,In_883);
or U1131 (N_1131,In_808,In_53);
nand U1132 (N_1132,In_448,In_195);
nand U1133 (N_1133,In_264,In_317);
and U1134 (N_1134,In_66,In_548);
nand U1135 (N_1135,In_539,In_743);
xnor U1136 (N_1136,In_985,In_816);
nor U1137 (N_1137,In_703,In_322);
nand U1138 (N_1138,In_793,In_444);
nor U1139 (N_1139,In_807,In_632);
nand U1140 (N_1140,In_96,In_391);
or U1141 (N_1141,In_539,In_0);
and U1142 (N_1142,In_497,In_837);
nor U1143 (N_1143,In_427,In_730);
xor U1144 (N_1144,In_207,In_716);
nor U1145 (N_1145,In_271,In_485);
and U1146 (N_1146,In_248,In_759);
nor U1147 (N_1147,In_556,In_836);
and U1148 (N_1148,In_284,In_110);
nor U1149 (N_1149,In_862,In_944);
nor U1150 (N_1150,In_269,In_137);
and U1151 (N_1151,In_899,In_297);
xor U1152 (N_1152,In_76,In_990);
nor U1153 (N_1153,In_949,In_925);
nor U1154 (N_1154,In_964,In_700);
and U1155 (N_1155,In_326,In_714);
nand U1156 (N_1156,In_275,In_494);
nand U1157 (N_1157,In_100,In_797);
nor U1158 (N_1158,In_934,In_97);
nand U1159 (N_1159,In_189,In_921);
and U1160 (N_1160,In_792,In_4);
xor U1161 (N_1161,In_286,In_885);
and U1162 (N_1162,In_100,In_30);
nor U1163 (N_1163,In_101,In_273);
xor U1164 (N_1164,In_385,In_684);
or U1165 (N_1165,In_743,In_417);
or U1166 (N_1166,In_630,In_643);
or U1167 (N_1167,In_233,In_863);
nand U1168 (N_1168,In_741,In_580);
xor U1169 (N_1169,In_498,In_70);
and U1170 (N_1170,In_447,In_913);
xor U1171 (N_1171,In_304,In_132);
or U1172 (N_1172,In_848,In_318);
xor U1173 (N_1173,In_139,In_478);
nor U1174 (N_1174,In_264,In_302);
and U1175 (N_1175,In_35,In_771);
or U1176 (N_1176,In_534,In_333);
and U1177 (N_1177,In_769,In_601);
nor U1178 (N_1178,In_452,In_586);
and U1179 (N_1179,In_86,In_731);
or U1180 (N_1180,In_504,In_719);
and U1181 (N_1181,In_809,In_942);
xnor U1182 (N_1182,In_779,In_105);
nor U1183 (N_1183,In_585,In_560);
and U1184 (N_1184,In_479,In_400);
or U1185 (N_1185,In_328,In_962);
or U1186 (N_1186,In_120,In_568);
or U1187 (N_1187,In_103,In_106);
nand U1188 (N_1188,In_15,In_478);
nor U1189 (N_1189,In_406,In_316);
nand U1190 (N_1190,In_810,In_425);
or U1191 (N_1191,In_525,In_636);
or U1192 (N_1192,In_438,In_215);
nand U1193 (N_1193,In_134,In_640);
and U1194 (N_1194,In_425,In_189);
xnor U1195 (N_1195,In_159,In_816);
nand U1196 (N_1196,In_173,In_396);
nand U1197 (N_1197,In_363,In_938);
nor U1198 (N_1198,In_289,In_815);
nand U1199 (N_1199,In_646,In_947);
nand U1200 (N_1200,In_527,In_557);
nor U1201 (N_1201,In_558,In_726);
xor U1202 (N_1202,In_171,In_428);
xor U1203 (N_1203,In_307,In_135);
or U1204 (N_1204,In_608,In_225);
and U1205 (N_1205,In_181,In_217);
and U1206 (N_1206,In_713,In_770);
xnor U1207 (N_1207,In_324,In_441);
nand U1208 (N_1208,In_158,In_701);
nand U1209 (N_1209,In_3,In_642);
or U1210 (N_1210,In_757,In_406);
nor U1211 (N_1211,In_746,In_255);
nor U1212 (N_1212,In_190,In_319);
nand U1213 (N_1213,In_227,In_868);
nor U1214 (N_1214,In_711,In_389);
and U1215 (N_1215,In_130,In_790);
or U1216 (N_1216,In_698,In_464);
nand U1217 (N_1217,In_144,In_190);
and U1218 (N_1218,In_946,In_828);
nor U1219 (N_1219,In_305,In_64);
or U1220 (N_1220,In_312,In_278);
nand U1221 (N_1221,In_819,In_328);
nor U1222 (N_1222,In_944,In_291);
or U1223 (N_1223,In_152,In_533);
or U1224 (N_1224,In_443,In_699);
or U1225 (N_1225,In_134,In_550);
nand U1226 (N_1226,In_416,In_629);
nor U1227 (N_1227,In_376,In_730);
or U1228 (N_1228,In_990,In_748);
and U1229 (N_1229,In_679,In_826);
nor U1230 (N_1230,In_120,In_518);
nand U1231 (N_1231,In_452,In_108);
xor U1232 (N_1232,In_817,In_714);
xnor U1233 (N_1233,In_648,In_15);
or U1234 (N_1234,In_64,In_670);
or U1235 (N_1235,In_859,In_42);
xor U1236 (N_1236,In_977,In_755);
or U1237 (N_1237,In_653,In_805);
nand U1238 (N_1238,In_86,In_650);
or U1239 (N_1239,In_395,In_967);
nand U1240 (N_1240,In_20,In_833);
xor U1241 (N_1241,In_118,In_979);
nor U1242 (N_1242,In_869,In_579);
and U1243 (N_1243,In_300,In_973);
or U1244 (N_1244,In_489,In_173);
xor U1245 (N_1245,In_720,In_410);
nor U1246 (N_1246,In_1,In_915);
nand U1247 (N_1247,In_277,In_846);
nand U1248 (N_1248,In_509,In_434);
xnor U1249 (N_1249,In_487,In_827);
and U1250 (N_1250,In_862,In_767);
or U1251 (N_1251,In_184,In_438);
xnor U1252 (N_1252,In_886,In_278);
nand U1253 (N_1253,In_209,In_991);
and U1254 (N_1254,In_901,In_314);
nand U1255 (N_1255,In_657,In_246);
or U1256 (N_1256,In_876,In_934);
and U1257 (N_1257,In_75,In_853);
nand U1258 (N_1258,In_913,In_29);
or U1259 (N_1259,In_526,In_606);
and U1260 (N_1260,In_763,In_430);
or U1261 (N_1261,In_740,In_252);
nand U1262 (N_1262,In_796,In_11);
or U1263 (N_1263,In_516,In_197);
and U1264 (N_1264,In_88,In_651);
and U1265 (N_1265,In_310,In_122);
and U1266 (N_1266,In_182,In_478);
or U1267 (N_1267,In_761,In_114);
or U1268 (N_1268,In_954,In_226);
and U1269 (N_1269,In_197,In_939);
nand U1270 (N_1270,In_689,In_60);
and U1271 (N_1271,In_763,In_891);
xnor U1272 (N_1272,In_510,In_963);
xnor U1273 (N_1273,In_508,In_58);
or U1274 (N_1274,In_23,In_373);
or U1275 (N_1275,In_606,In_28);
or U1276 (N_1276,In_758,In_12);
nand U1277 (N_1277,In_793,In_570);
and U1278 (N_1278,In_948,In_17);
or U1279 (N_1279,In_372,In_810);
nand U1280 (N_1280,In_221,In_785);
or U1281 (N_1281,In_339,In_886);
or U1282 (N_1282,In_256,In_451);
and U1283 (N_1283,In_766,In_454);
nor U1284 (N_1284,In_282,In_771);
or U1285 (N_1285,In_401,In_34);
nand U1286 (N_1286,In_281,In_686);
and U1287 (N_1287,In_90,In_704);
xor U1288 (N_1288,In_157,In_105);
nand U1289 (N_1289,In_374,In_940);
or U1290 (N_1290,In_5,In_379);
nor U1291 (N_1291,In_601,In_107);
and U1292 (N_1292,In_90,In_954);
and U1293 (N_1293,In_771,In_113);
and U1294 (N_1294,In_587,In_141);
and U1295 (N_1295,In_496,In_825);
and U1296 (N_1296,In_299,In_922);
nor U1297 (N_1297,In_337,In_827);
or U1298 (N_1298,In_773,In_566);
nand U1299 (N_1299,In_871,In_18);
nor U1300 (N_1300,In_912,In_132);
or U1301 (N_1301,In_941,In_234);
nand U1302 (N_1302,In_100,In_142);
nor U1303 (N_1303,In_916,In_574);
and U1304 (N_1304,In_341,In_204);
nor U1305 (N_1305,In_347,In_395);
nor U1306 (N_1306,In_260,In_704);
and U1307 (N_1307,In_397,In_680);
nand U1308 (N_1308,In_908,In_391);
nand U1309 (N_1309,In_624,In_627);
and U1310 (N_1310,In_60,In_653);
xnor U1311 (N_1311,In_484,In_149);
nand U1312 (N_1312,In_269,In_909);
and U1313 (N_1313,In_703,In_340);
xor U1314 (N_1314,In_810,In_715);
or U1315 (N_1315,In_255,In_680);
nor U1316 (N_1316,In_613,In_947);
xor U1317 (N_1317,In_103,In_835);
and U1318 (N_1318,In_951,In_393);
or U1319 (N_1319,In_487,In_943);
or U1320 (N_1320,In_883,In_676);
xor U1321 (N_1321,In_703,In_445);
and U1322 (N_1322,In_276,In_339);
and U1323 (N_1323,In_661,In_55);
xnor U1324 (N_1324,In_196,In_0);
nor U1325 (N_1325,In_950,In_51);
nand U1326 (N_1326,In_242,In_188);
nor U1327 (N_1327,In_291,In_265);
nand U1328 (N_1328,In_0,In_913);
and U1329 (N_1329,In_554,In_15);
nand U1330 (N_1330,In_272,In_402);
nand U1331 (N_1331,In_712,In_208);
nand U1332 (N_1332,In_986,In_816);
nor U1333 (N_1333,In_102,In_350);
and U1334 (N_1334,In_210,In_432);
and U1335 (N_1335,In_93,In_650);
nor U1336 (N_1336,In_673,In_362);
nor U1337 (N_1337,In_321,In_901);
nor U1338 (N_1338,In_909,In_52);
nand U1339 (N_1339,In_274,In_757);
xor U1340 (N_1340,In_331,In_458);
or U1341 (N_1341,In_542,In_123);
nor U1342 (N_1342,In_214,In_905);
nor U1343 (N_1343,In_183,In_694);
nor U1344 (N_1344,In_840,In_10);
or U1345 (N_1345,In_782,In_275);
xnor U1346 (N_1346,In_168,In_366);
nand U1347 (N_1347,In_955,In_767);
nand U1348 (N_1348,In_367,In_48);
or U1349 (N_1349,In_674,In_206);
xor U1350 (N_1350,In_444,In_45);
nand U1351 (N_1351,In_759,In_801);
nand U1352 (N_1352,In_523,In_767);
nand U1353 (N_1353,In_217,In_468);
nor U1354 (N_1354,In_95,In_994);
nand U1355 (N_1355,In_828,In_746);
and U1356 (N_1356,In_646,In_897);
or U1357 (N_1357,In_878,In_365);
and U1358 (N_1358,In_338,In_835);
nand U1359 (N_1359,In_818,In_34);
nand U1360 (N_1360,In_802,In_814);
and U1361 (N_1361,In_678,In_463);
nand U1362 (N_1362,In_688,In_483);
nor U1363 (N_1363,In_344,In_548);
or U1364 (N_1364,In_45,In_816);
xor U1365 (N_1365,In_216,In_349);
and U1366 (N_1366,In_232,In_503);
nand U1367 (N_1367,In_7,In_449);
nand U1368 (N_1368,In_719,In_449);
nand U1369 (N_1369,In_826,In_291);
and U1370 (N_1370,In_102,In_865);
nand U1371 (N_1371,In_406,In_315);
and U1372 (N_1372,In_610,In_244);
and U1373 (N_1373,In_877,In_35);
and U1374 (N_1374,In_181,In_615);
nand U1375 (N_1375,In_195,In_391);
nand U1376 (N_1376,In_859,In_177);
nand U1377 (N_1377,In_597,In_710);
nor U1378 (N_1378,In_666,In_437);
nand U1379 (N_1379,In_6,In_712);
or U1380 (N_1380,In_55,In_424);
or U1381 (N_1381,In_125,In_61);
and U1382 (N_1382,In_102,In_124);
or U1383 (N_1383,In_935,In_947);
and U1384 (N_1384,In_439,In_897);
nor U1385 (N_1385,In_530,In_51);
or U1386 (N_1386,In_656,In_915);
and U1387 (N_1387,In_850,In_1);
nand U1388 (N_1388,In_147,In_799);
nor U1389 (N_1389,In_684,In_772);
and U1390 (N_1390,In_125,In_228);
and U1391 (N_1391,In_187,In_157);
nor U1392 (N_1392,In_452,In_672);
nor U1393 (N_1393,In_922,In_633);
nand U1394 (N_1394,In_345,In_32);
or U1395 (N_1395,In_539,In_631);
nor U1396 (N_1396,In_89,In_388);
and U1397 (N_1397,In_226,In_744);
and U1398 (N_1398,In_416,In_389);
nand U1399 (N_1399,In_332,In_670);
nor U1400 (N_1400,In_278,In_974);
or U1401 (N_1401,In_648,In_384);
nand U1402 (N_1402,In_809,In_266);
nor U1403 (N_1403,In_539,In_292);
or U1404 (N_1404,In_488,In_525);
nor U1405 (N_1405,In_348,In_14);
nand U1406 (N_1406,In_905,In_765);
and U1407 (N_1407,In_76,In_157);
nand U1408 (N_1408,In_856,In_2);
or U1409 (N_1409,In_475,In_226);
or U1410 (N_1410,In_629,In_274);
and U1411 (N_1411,In_608,In_579);
nor U1412 (N_1412,In_782,In_757);
nor U1413 (N_1413,In_151,In_491);
nand U1414 (N_1414,In_654,In_392);
and U1415 (N_1415,In_534,In_28);
or U1416 (N_1416,In_453,In_924);
or U1417 (N_1417,In_374,In_91);
nor U1418 (N_1418,In_447,In_413);
or U1419 (N_1419,In_526,In_208);
nor U1420 (N_1420,In_846,In_32);
nor U1421 (N_1421,In_624,In_669);
nand U1422 (N_1422,In_273,In_128);
nand U1423 (N_1423,In_160,In_565);
or U1424 (N_1424,In_470,In_641);
and U1425 (N_1425,In_495,In_457);
nor U1426 (N_1426,In_382,In_362);
nand U1427 (N_1427,In_149,In_885);
nor U1428 (N_1428,In_94,In_878);
xnor U1429 (N_1429,In_815,In_662);
or U1430 (N_1430,In_203,In_911);
nor U1431 (N_1431,In_709,In_945);
and U1432 (N_1432,In_947,In_434);
xnor U1433 (N_1433,In_99,In_231);
and U1434 (N_1434,In_265,In_310);
xnor U1435 (N_1435,In_179,In_141);
and U1436 (N_1436,In_556,In_8);
nand U1437 (N_1437,In_928,In_269);
xor U1438 (N_1438,In_747,In_96);
or U1439 (N_1439,In_0,In_974);
xor U1440 (N_1440,In_325,In_632);
and U1441 (N_1441,In_716,In_914);
nand U1442 (N_1442,In_898,In_676);
and U1443 (N_1443,In_423,In_853);
or U1444 (N_1444,In_847,In_610);
or U1445 (N_1445,In_227,In_443);
or U1446 (N_1446,In_977,In_401);
and U1447 (N_1447,In_394,In_622);
and U1448 (N_1448,In_343,In_279);
xor U1449 (N_1449,In_169,In_125);
or U1450 (N_1450,In_438,In_641);
nor U1451 (N_1451,In_965,In_709);
nor U1452 (N_1452,In_238,In_262);
or U1453 (N_1453,In_496,In_411);
nor U1454 (N_1454,In_899,In_835);
or U1455 (N_1455,In_759,In_388);
and U1456 (N_1456,In_106,In_568);
or U1457 (N_1457,In_407,In_446);
nand U1458 (N_1458,In_558,In_481);
or U1459 (N_1459,In_873,In_663);
nor U1460 (N_1460,In_759,In_154);
nor U1461 (N_1461,In_563,In_393);
nand U1462 (N_1462,In_61,In_272);
nand U1463 (N_1463,In_433,In_467);
and U1464 (N_1464,In_111,In_574);
xnor U1465 (N_1465,In_788,In_927);
or U1466 (N_1466,In_259,In_96);
nor U1467 (N_1467,In_451,In_74);
nor U1468 (N_1468,In_496,In_850);
nor U1469 (N_1469,In_308,In_36);
xor U1470 (N_1470,In_458,In_312);
nor U1471 (N_1471,In_520,In_896);
or U1472 (N_1472,In_968,In_42);
or U1473 (N_1473,In_142,In_579);
nor U1474 (N_1474,In_689,In_755);
or U1475 (N_1475,In_49,In_205);
nor U1476 (N_1476,In_369,In_909);
nand U1477 (N_1477,In_865,In_257);
nand U1478 (N_1478,In_415,In_590);
or U1479 (N_1479,In_54,In_173);
nand U1480 (N_1480,In_991,In_99);
or U1481 (N_1481,In_189,In_790);
or U1482 (N_1482,In_557,In_491);
and U1483 (N_1483,In_902,In_993);
or U1484 (N_1484,In_60,In_148);
or U1485 (N_1485,In_902,In_800);
nand U1486 (N_1486,In_197,In_17);
or U1487 (N_1487,In_329,In_471);
or U1488 (N_1488,In_278,In_251);
nor U1489 (N_1489,In_887,In_538);
or U1490 (N_1490,In_955,In_361);
nor U1491 (N_1491,In_313,In_888);
and U1492 (N_1492,In_123,In_825);
nor U1493 (N_1493,In_888,In_333);
nor U1494 (N_1494,In_430,In_323);
xor U1495 (N_1495,In_534,In_241);
xor U1496 (N_1496,In_350,In_373);
xor U1497 (N_1497,In_632,In_922);
or U1498 (N_1498,In_812,In_895);
and U1499 (N_1499,In_798,In_611);
xor U1500 (N_1500,In_680,In_282);
nand U1501 (N_1501,In_25,In_224);
and U1502 (N_1502,In_746,In_437);
nor U1503 (N_1503,In_55,In_419);
nor U1504 (N_1504,In_877,In_768);
xor U1505 (N_1505,In_66,In_27);
nand U1506 (N_1506,In_284,In_207);
and U1507 (N_1507,In_161,In_604);
or U1508 (N_1508,In_614,In_305);
nor U1509 (N_1509,In_232,In_641);
and U1510 (N_1510,In_420,In_190);
or U1511 (N_1511,In_117,In_313);
or U1512 (N_1512,In_623,In_537);
nand U1513 (N_1513,In_610,In_308);
nor U1514 (N_1514,In_730,In_103);
or U1515 (N_1515,In_134,In_898);
and U1516 (N_1516,In_422,In_343);
nand U1517 (N_1517,In_774,In_194);
xor U1518 (N_1518,In_333,In_413);
nor U1519 (N_1519,In_29,In_992);
xor U1520 (N_1520,In_199,In_760);
and U1521 (N_1521,In_966,In_101);
and U1522 (N_1522,In_873,In_86);
xnor U1523 (N_1523,In_73,In_557);
and U1524 (N_1524,In_918,In_246);
xnor U1525 (N_1525,In_785,In_193);
or U1526 (N_1526,In_352,In_627);
nand U1527 (N_1527,In_160,In_264);
and U1528 (N_1528,In_241,In_846);
or U1529 (N_1529,In_798,In_138);
and U1530 (N_1530,In_360,In_530);
nor U1531 (N_1531,In_268,In_893);
or U1532 (N_1532,In_537,In_654);
and U1533 (N_1533,In_569,In_938);
and U1534 (N_1534,In_995,In_533);
and U1535 (N_1535,In_367,In_105);
nor U1536 (N_1536,In_630,In_828);
and U1537 (N_1537,In_74,In_696);
nor U1538 (N_1538,In_224,In_129);
xor U1539 (N_1539,In_969,In_613);
nand U1540 (N_1540,In_855,In_981);
or U1541 (N_1541,In_596,In_372);
nand U1542 (N_1542,In_104,In_512);
nor U1543 (N_1543,In_148,In_414);
or U1544 (N_1544,In_138,In_402);
nor U1545 (N_1545,In_976,In_464);
nor U1546 (N_1546,In_724,In_695);
nand U1547 (N_1547,In_616,In_122);
xnor U1548 (N_1548,In_794,In_896);
nand U1549 (N_1549,In_480,In_847);
nor U1550 (N_1550,In_334,In_70);
nand U1551 (N_1551,In_397,In_846);
nor U1552 (N_1552,In_19,In_353);
and U1553 (N_1553,In_225,In_932);
and U1554 (N_1554,In_44,In_987);
nand U1555 (N_1555,In_692,In_345);
nor U1556 (N_1556,In_671,In_388);
nand U1557 (N_1557,In_65,In_33);
nand U1558 (N_1558,In_781,In_855);
and U1559 (N_1559,In_370,In_99);
nor U1560 (N_1560,In_773,In_453);
nor U1561 (N_1561,In_151,In_952);
or U1562 (N_1562,In_813,In_869);
nor U1563 (N_1563,In_285,In_424);
and U1564 (N_1564,In_861,In_369);
nor U1565 (N_1565,In_537,In_803);
nor U1566 (N_1566,In_203,In_508);
nor U1567 (N_1567,In_562,In_811);
nor U1568 (N_1568,In_173,In_603);
nand U1569 (N_1569,In_955,In_979);
or U1570 (N_1570,In_652,In_767);
nor U1571 (N_1571,In_241,In_897);
and U1572 (N_1572,In_419,In_876);
and U1573 (N_1573,In_298,In_212);
and U1574 (N_1574,In_741,In_782);
nor U1575 (N_1575,In_632,In_186);
and U1576 (N_1576,In_389,In_403);
nand U1577 (N_1577,In_780,In_830);
and U1578 (N_1578,In_775,In_1);
nand U1579 (N_1579,In_327,In_48);
nand U1580 (N_1580,In_71,In_475);
nand U1581 (N_1581,In_354,In_246);
and U1582 (N_1582,In_261,In_708);
nand U1583 (N_1583,In_58,In_441);
and U1584 (N_1584,In_59,In_862);
or U1585 (N_1585,In_887,In_442);
nor U1586 (N_1586,In_661,In_5);
or U1587 (N_1587,In_211,In_731);
or U1588 (N_1588,In_858,In_267);
and U1589 (N_1589,In_982,In_374);
and U1590 (N_1590,In_665,In_440);
nand U1591 (N_1591,In_522,In_729);
xor U1592 (N_1592,In_636,In_274);
nor U1593 (N_1593,In_150,In_12);
and U1594 (N_1594,In_296,In_598);
and U1595 (N_1595,In_689,In_962);
and U1596 (N_1596,In_224,In_525);
nor U1597 (N_1597,In_216,In_974);
xnor U1598 (N_1598,In_63,In_811);
and U1599 (N_1599,In_938,In_50);
and U1600 (N_1600,In_83,In_756);
and U1601 (N_1601,In_949,In_616);
nor U1602 (N_1602,In_601,In_152);
nor U1603 (N_1603,In_651,In_20);
or U1604 (N_1604,In_721,In_584);
or U1605 (N_1605,In_634,In_919);
nor U1606 (N_1606,In_523,In_618);
nor U1607 (N_1607,In_497,In_900);
and U1608 (N_1608,In_562,In_845);
and U1609 (N_1609,In_240,In_40);
nand U1610 (N_1610,In_782,In_138);
and U1611 (N_1611,In_396,In_373);
xor U1612 (N_1612,In_616,In_759);
and U1613 (N_1613,In_623,In_174);
nand U1614 (N_1614,In_870,In_938);
or U1615 (N_1615,In_486,In_616);
nand U1616 (N_1616,In_201,In_643);
nand U1617 (N_1617,In_565,In_661);
and U1618 (N_1618,In_104,In_384);
or U1619 (N_1619,In_350,In_764);
nand U1620 (N_1620,In_581,In_678);
nand U1621 (N_1621,In_218,In_293);
xnor U1622 (N_1622,In_947,In_440);
nand U1623 (N_1623,In_755,In_64);
nand U1624 (N_1624,In_137,In_85);
and U1625 (N_1625,In_882,In_793);
nor U1626 (N_1626,In_523,In_755);
and U1627 (N_1627,In_382,In_962);
nor U1628 (N_1628,In_370,In_253);
or U1629 (N_1629,In_471,In_118);
or U1630 (N_1630,In_500,In_595);
nor U1631 (N_1631,In_704,In_360);
nand U1632 (N_1632,In_460,In_818);
nand U1633 (N_1633,In_850,In_871);
nor U1634 (N_1634,In_867,In_303);
or U1635 (N_1635,In_916,In_395);
nand U1636 (N_1636,In_297,In_788);
nor U1637 (N_1637,In_483,In_290);
nand U1638 (N_1638,In_770,In_985);
and U1639 (N_1639,In_27,In_180);
nand U1640 (N_1640,In_814,In_95);
xnor U1641 (N_1641,In_251,In_434);
nor U1642 (N_1642,In_762,In_67);
xor U1643 (N_1643,In_886,In_170);
nor U1644 (N_1644,In_754,In_642);
nor U1645 (N_1645,In_971,In_885);
and U1646 (N_1646,In_815,In_993);
nor U1647 (N_1647,In_804,In_303);
nor U1648 (N_1648,In_532,In_887);
xor U1649 (N_1649,In_751,In_823);
nor U1650 (N_1650,In_533,In_552);
or U1651 (N_1651,In_715,In_809);
and U1652 (N_1652,In_549,In_127);
nand U1653 (N_1653,In_284,In_590);
or U1654 (N_1654,In_728,In_64);
nand U1655 (N_1655,In_168,In_119);
or U1656 (N_1656,In_554,In_784);
nor U1657 (N_1657,In_391,In_203);
and U1658 (N_1658,In_43,In_307);
nor U1659 (N_1659,In_71,In_84);
nand U1660 (N_1660,In_15,In_964);
and U1661 (N_1661,In_488,In_0);
and U1662 (N_1662,In_338,In_459);
nand U1663 (N_1663,In_176,In_354);
and U1664 (N_1664,In_462,In_704);
or U1665 (N_1665,In_426,In_801);
nand U1666 (N_1666,In_984,In_869);
nor U1667 (N_1667,In_862,In_62);
nor U1668 (N_1668,In_341,In_241);
and U1669 (N_1669,In_104,In_172);
nand U1670 (N_1670,In_589,In_353);
nand U1671 (N_1671,In_734,In_373);
nor U1672 (N_1672,In_795,In_184);
nand U1673 (N_1673,In_820,In_335);
nor U1674 (N_1674,In_829,In_24);
nand U1675 (N_1675,In_623,In_675);
or U1676 (N_1676,In_836,In_981);
nand U1677 (N_1677,In_656,In_775);
nand U1678 (N_1678,In_749,In_241);
and U1679 (N_1679,In_796,In_331);
nand U1680 (N_1680,In_162,In_355);
nand U1681 (N_1681,In_259,In_177);
and U1682 (N_1682,In_460,In_102);
or U1683 (N_1683,In_748,In_365);
nor U1684 (N_1684,In_362,In_913);
or U1685 (N_1685,In_876,In_686);
nor U1686 (N_1686,In_561,In_563);
and U1687 (N_1687,In_927,In_211);
nor U1688 (N_1688,In_473,In_246);
nor U1689 (N_1689,In_955,In_301);
and U1690 (N_1690,In_325,In_501);
xnor U1691 (N_1691,In_223,In_742);
or U1692 (N_1692,In_932,In_630);
nor U1693 (N_1693,In_286,In_976);
nand U1694 (N_1694,In_672,In_851);
or U1695 (N_1695,In_351,In_222);
and U1696 (N_1696,In_909,In_854);
or U1697 (N_1697,In_397,In_141);
nand U1698 (N_1698,In_676,In_35);
and U1699 (N_1699,In_58,In_756);
nand U1700 (N_1700,In_112,In_1);
or U1701 (N_1701,In_463,In_632);
or U1702 (N_1702,In_380,In_393);
nor U1703 (N_1703,In_833,In_401);
and U1704 (N_1704,In_201,In_420);
nor U1705 (N_1705,In_593,In_658);
or U1706 (N_1706,In_512,In_738);
nor U1707 (N_1707,In_23,In_503);
nor U1708 (N_1708,In_49,In_942);
and U1709 (N_1709,In_66,In_3);
nor U1710 (N_1710,In_809,In_842);
xor U1711 (N_1711,In_565,In_801);
nor U1712 (N_1712,In_904,In_154);
nand U1713 (N_1713,In_680,In_371);
nand U1714 (N_1714,In_913,In_574);
xnor U1715 (N_1715,In_319,In_871);
nand U1716 (N_1716,In_423,In_943);
nor U1717 (N_1717,In_259,In_463);
and U1718 (N_1718,In_338,In_672);
and U1719 (N_1719,In_232,In_988);
and U1720 (N_1720,In_519,In_536);
and U1721 (N_1721,In_135,In_153);
and U1722 (N_1722,In_526,In_728);
and U1723 (N_1723,In_616,In_8);
nand U1724 (N_1724,In_356,In_290);
nand U1725 (N_1725,In_106,In_500);
and U1726 (N_1726,In_967,In_953);
or U1727 (N_1727,In_849,In_718);
xnor U1728 (N_1728,In_83,In_261);
and U1729 (N_1729,In_137,In_911);
and U1730 (N_1730,In_880,In_394);
nand U1731 (N_1731,In_366,In_313);
nand U1732 (N_1732,In_859,In_104);
or U1733 (N_1733,In_338,In_365);
xor U1734 (N_1734,In_186,In_174);
nand U1735 (N_1735,In_801,In_805);
nand U1736 (N_1736,In_651,In_990);
nor U1737 (N_1737,In_97,In_96);
xor U1738 (N_1738,In_407,In_266);
nor U1739 (N_1739,In_888,In_913);
or U1740 (N_1740,In_215,In_476);
or U1741 (N_1741,In_383,In_872);
nand U1742 (N_1742,In_970,In_202);
or U1743 (N_1743,In_890,In_671);
xor U1744 (N_1744,In_439,In_336);
nor U1745 (N_1745,In_671,In_78);
or U1746 (N_1746,In_86,In_868);
or U1747 (N_1747,In_303,In_411);
or U1748 (N_1748,In_683,In_968);
and U1749 (N_1749,In_670,In_675);
or U1750 (N_1750,In_405,In_447);
nand U1751 (N_1751,In_875,In_524);
and U1752 (N_1752,In_881,In_465);
nand U1753 (N_1753,In_858,In_113);
nand U1754 (N_1754,In_898,In_155);
or U1755 (N_1755,In_328,In_843);
nand U1756 (N_1756,In_142,In_791);
or U1757 (N_1757,In_682,In_296);
xnor U1758 (N_1758,In_804,In_417);
nand U1759 (N_1759,In_667,In_122);
xor U1760 (N_1760,In_98,In_126);
nand U1761 (N_1761,In_816,In_204);
nand U1762 (N_1762,In_1,In_947);
nor U1763 (N_1763,In_496,In_833);
xnor U1764 (N_1764,In_938,In_700);
or U1765 (N_1765,In_47,In_408);
and U1766 (N_1766,In_677,In_330);
and U1767 (N_1767,In_455,In_701);
nand U1768 (N_1768,In_19,In_21);
or U1769 (N_1769,In_166,In_71);
xor U1770 (N_1770,In_655,In_24);
nor U1771 (N_1771,In_924,In_161);
or U1772 (N_1772,In_433,In_774);
nor U1773 (N_1773,In_303,In_313);
nor U1774 (N_1774,In_299,In_84);
or U1775 (N_1775,In_830,In_938);
or U1776 (N_1776,In_975,In_750);
nand U1777 (N_1777,In_103,In_155);
and U1778 (N_1778,In_67,In_547);
nand U1779 (N_1779,In_288,In_496);
xnor U1780 (N_1780,In_98,In_722);
nand U1781 (N_1781,In_277,In_757);
and U1782 (N_1782,In_142,In_888);
xor U1783 (N_1783,In_925,In_814);
and U1784 (N_1784,In_435,In_82);
nand U1785 (N_1785,In_58,In_711);
nand U1786 (N_1786,In_708,In_267);
and U1787 (N_1787,In_418,In_153);
and U1788 (N_1788,In_186,In_258);
and U1789 (N_1789,In_436,In_590);
or U1790 (N_1790,In_485,In_586);
nor U1791 (N_1791,In_192,In_741);
nand U1792 (N_1792,In_527,In_699);
nand U1793 (N_1793,In_609,In_349);
nand U1794 (N_1794,In_161,In_151);
and U1795 (N_1795,In_819,In_174);
nor U1796 (N_1796,In_911,In_412);
nor U1797 (N_1797,In_819,In_225);
xor U1798 (N_1798,In_119,In_83);
or U1799 (N_1799,In_896,In_426);
or U1800 (N_1800,In_898,In_713);
nor U1801 (N_1801,In_621,In_412);
nand U1802 (N_1802,In_114,In_919);
nand U1803 (N_1803,In_239,In_823);
nor U1804 (N_1804,In_895,In_39);
or U1805 (N_1805,In_610,In_950);
or U1806 (N_1806,In_981,In_450);
nor U1807 (N_1807,In_132,In_32);
xor U1808 (N_1808,In_605,In_73);
nor U1809 (N_1809,In_209,In_819);
or U1810 (N_1810,In_838,In_258);
and U1811 (N_1811,In_632,In_534);
nor U1812 (N_1812,In_208,In_119);
xor U1813 (N_1813,In_57,In_285);
nand U1814 (N_1814,In_611,In_361);
and U1815 (N_1815,In_468,In_941);
and U1816 (N_1816,In_983,In_670);
nor U1817 (N_1817,In_510,In_595);
xor U1818 (N_1818,In_725,In_900);
nand U1819 (N_1819,In_134,In_568);
nand U1820 (N_1820,In_684,In_493);
nor U1821 (N_1821,In_61,In_793);
xor U1822 (N_1822,In_433,In_636);
nand U1823 (N_1823,In_589,In_342);
nor U1824 (N_1824,In_486,In_460);
nor U1825 (N_1825,In_901,In_227);
nor U1826 (N_1826,In_519,In_771);
and U1827 (N_1827,In_720,In_799);
nor U1828 (N_1828,In_742,In_631);
nand U1829 (N_1829,In_593,In_111);
or U1830 (N_1830,In_550,In_100);
xnor U1831 (N_1831,In_372,In_197);
nor U1832 (N_1832,In_121,In_45);
nor U1833 (N_1833,In_407,In_305);
nor U1834 (N_1834,In_378,In_28);
or U1835 (N_1835,In_259,In_765);
or U1836 (N_1836,In_134,In_366);
or U1837 (N_1837,In_569,In_527);
nand U1838 (N_1838,In_943,In_799);
nand U1839 (N_1839,In_557,In_255);
nor U1840 (N_1840,In_51,In_191);
xnor U1841 (N_1841,In_521,In_624);
and U1842 (N_1842,In_642,In_821);
nand U1843 (N_1843,In_902,In_605);
nand U1844 (N_1844,In_629,In_99);
xor U1845 (N_1845,In_402,In_14);
nand U1846 (N_1846,In_310,In_838);
nand U1847 (N_1847,In_465,In_407);
and U1848 (N_1848,In_500,In_959);
nand U1849 (N_1849,In_195,In_487);
or U1850 (N_1850,In_507,In_15);
nand U1851 (N_1851,In_817,In_533);
nand U1852 (N_1852,In_293,In_161);
and U1853 (N_1853,In_116,In_434);
or U1854 (N_1854,In_664,In_61);
and U1855 (N_1855,In_574,In_586);
nand U1856 (N_1856,In_351,In_24);
and U1857 (N_1857,In_732,In_753);
nand U1858 (N_1858,In_475,In_461);
nor U1859 (N_1859,In_619,In_60);
and U1860 (N_1860,In_650,In_731);
nand U1861 (N_1861,In_264,In_675);
nand U1862 (N_1862,In_389,In_131);
and U1863 (N_1863,In_847,In_741);
and U1864 (N_1864,In_848,In_328);
nor U1865 (N_1865,In_120,In_679);
nor U1866 (N_1866,In_875,In_527);
and U1867 (N_1867,In_373,In_879);
or U1868 (N_1868,In_121,In_142);
and U1869 (N_1869,In_820,In_399);
nand U1870 (N_1870,In_96,In_717);
or U1871 (N_1871,In_859,In_785);
nand U1872 (N_1872,In_13,In_249);
or U1873 (N_1873,In_206,In_342);
nand U1874 (N_1874,In_454,In_774);
nor U1875 (N_1875,In_644,In_168);
nor U1876 (N_1876,In_350,In_11);
or U1877 (N_1877,In_219,In_627);
and U1878 (N_1878,In_871,In_661);
and U1879 (N_1879,In_166,In_458);
or U1880 (N_1880,In_919,In_15);
nand U1881 (N_1881,In_790,In_533);
nand U1882 (N_1882,In_254,In_428);
nor U1883 (N_1883,In_560,In_243);
or U1884 (N_1884,In_306,In_369);
nor U1885 (N_1885,In_838,In_864);
nand U1886 (N_1886,In_150,In_785);
and U1887 (N_1887,In_670,In_885);
and U1888 (N_1888,In_696,In_352);
nand U1889 (N_1889,In_302,In_565);
nand U1890 (N_1890,In_526,In_959);
or U1891 (N_1891,In_868,In_148);
nor U1892 (N_1892,In_552,In_584);
or U1893 (N_1893,In_315,In_858);
nor U1894 (N_1894,In_135,In_383);
xor U1895 (N_1895,In_900,In_580);
or U1896 (N_1896,In_349,In_70);
and U1897 (N_1897,In_406,In_796);
or U1898 (N_1898,In_598,In_42);
nor U1899 (N_1899,In_82,In_901);
or U1900 (N_1900,In_141,In_222);
xnor U1901 (N_1901,In_232,In_479);
and U1902 (N_1902,In_187,In_413);
nand U1903 (N_1903,In_377,In_613);
and U1904 (N_1904,In_954,In_250);
or U1905 (N_1905,In_677,In_476);
xnor U1906 (N_1906,In_335,In_654);
and U1907 (N_1907,In_644,In_688);
and U1908 (N_1908,In_634,In_573);
nand U1909 (N_1909,In_121,In_725);
and U1910 (N_1910,In_900,In_714);
nor U1911 (N_1911,In_330,In_903);
and U1912 (N_1912,In_489,In_917);
xnor U1913 (N_1913,In_0,In_173);
or U1914 (N_1914,In_79,In_668);
xnor U1915 (N_1915,In_250,In_699);
nor U1916 (N_1916,In_149,In_241);
xnor U1917 (N_1917,In_887,In_915);
nor U1918 (N_1918,In_487,In_244);
and U1919 (N_1919,In_739,In_294);
and U1920 (N_1920,In_855,In_786);
nand U1921 (N_1921,In_738,In_735);
or U1922 (N_1922,In_794,In_24);
xnor U1923 (N_1923,In_39,In_899);
or U1924 (N_1924,In_680,In_720);
or U1925 (N_1925,In_952,In_979);
xor U1926 (N_1926,In_952,In_499);
and U1927 (N_1927,In_313,In_44);
nand U1928 (N_1928,In_381,In_617);
or U1929 (N_1929,In_133,In_931);
or U1930 (N_1930,In_702,In_114);
nand U1931 (N_1931,In_762,In_209);
nand U1932 (N_1932,In_78,In_421);
or U1933 (N_1933,In_807,In_109);
xor U1934 (N_1934,In_183,In_764);
or U1935 (N_1935,In_620,In_218);
xor U1936 (N_1936,In_437,In_947);
xor U1937 (N_1937,In_151,In_340);
nor U1938 (N_1938,In_659,In_154);
and U1939 (N_1939,In_168,In_972);
or U1940 (N_1940,In_48,In_387);
and U1941 (N_1941,In_131,In_101);
or U1942 (N_1942,In_199,In_491);
and U1943 (N_1943,In_226,In_588);
and U1944 (N_1944,In_781,In_344);
and U1945 (N_1945,In_519,In_706);
and U1946 (N_1946,In_400,In_384);
nor U1947 (N_1947,In_944,In_958);
and U1948 (N_1948,In_202,In_725);
nand U1949 (N_1949,In_231,In_880);
and U1950 (N_1950,In_222,In_11);
nor U1951 (N_1951,In_180,In_964);
and U1952 (N_1952,In_173,In_38);
nor U1953 (N_1953,In_386,In_51);
and U1954 (N_1954,In_560,In_703);
xor U1955 (N_1955,In_468,In_314);
xor U1956 (N_1956,In_101,In_644);
nand U1957 (N_1957,In_214,In_547);
nor U1958 (N_1958,In_859,In_327);
nor U1959 (N_1959,In_240,In_596);
nand U1960 (N_1960,In_50,In_541);
nor U1961 (N_1961,In_102,In_851);
and U1962 (N_1962,In_408,In_433);
or U1963 (N_1963,In_345,In_175);
nor U1964 (N_1964,In_330,In_348);
or U1965 (N_1965,In_110,In_946);
nor U1966 (N_1966,In_421,In_613);
nor U1967 (N_1967,In_577,In_540);
or U1968 (N_1968,In_1,In_869);
or U1969 (N_1969,In_931,In_65);
or U1970 (N_1970,In_448,In_273);
nand U1971 (N_1971,In_324,In_106);
nand U1972 (N_1972,In_250,In_345);
nor U1973 (N_1973,In_585,In_55);
and U1974 (N_1974,In_907,In_385);
xor U1975 (N_1975,In_844,In_976);
nand U1976 (N_1976,In_935,In_277);
or U1977 (N_1977,In_802,In_984);
or U1978 (N_1978,In_330,In_742);
or U1979 (N_1979,In_742,In_63);
or U1980 (N_1980,In_219,In_631);
nand U1981 (N_1981,In_996,In_528);
xnor U1982 (N_1982,In_979,In_792);
nor U1983 (N_1983,In_275,In_247);
and U1984 (N_1984,In_802,In_865);
nor U1985 (N_1985,In_318,In_269);
nor U1986 (N_1986,In_826,In_18);
or U1987 (N_1987,In_664,In_509);
nor U1988 (N_1988,In_272,In_329);
nand U1989 (N_1989,In_351,In_414);
nand U1990 (N_1990,In_578,In_849);
and U1991 (N_1991,In_966,In_553);
nor U1992 (N_1992,In_754,In_132);
nor U1993 (N_1993,In_16,In_376);
or U1994 (N_1994,In_904,In_883);
nor U1995 (N_1995,In_73,In_722);
or U1996 (N_1996,In_47,In_765);
xnor U1997 (N_1997,In_739,In_298);
nand U1998 (N_1998,In_879,In_104);
xnor U1999 (N_1999,In_693,In_82);
or U2000 (N_2000,In_105,In_233);
or U2001 (N_2001,In_124,In_891);
xor U2002 (N_2002,In_384,In_596);
nand U2003 (N_2003,In_625,In_266);
nand U2004 (N_2004,In_914,In_121);
nand U2005 (N_2005,In_191,In_450);
nand U2006 (N_2006,In_220,In_457);
nor U2007 (N_2007,In_23,In_708);
and U2008 (N_2008,In_288,In_271);
nor U2009 (N_2009,In_807,In_608);
or U2010 (N_2010,In_269,In_487);
and U2011 (N_2011,In_566,In_93);
nand U2012 (N_2012,In_655,In_208);
and U2013 (N_2013,In_771,In_96);
and U2014 (N_2014,In_302,In_718);
or U2015 (N_2015,In_909,In_244);
xnor U2016 (N_2016,In_99,In_564);
or U2017 (N_2017,In_751,In_463);
and U2018 (N_2018,In_269,In_759);
nand U2019 (N_2019,In_778,In_917);
nor U2020 (N_2020,In_372,In_931);
nor U2021 (N_2021,In_966,In_193);
and U2022 (N_2022,In_759,In_341);
or U2023 (N_2023,In_597,In_587);
or U2024 (N_2024,In_807,In_652);
xnor U2025 (N_2025,In_182,In_705);
and U2026 (N_2026,In_673,In_103);
xnor U2027 (N_2027,In_408,In_710);
or U2028 (N_2028,In_254,In_880);
or U2029 (N_2029,In_38,In_46);
or U2030 (N_2030,In_633,In_338);
or U2031 (N_2031,In_266,In_734);
nand U2032 (N_2032,In_759,In_795);
xnor U2033 (N_2033,In_28,In_717);
nand U2034 (N_2034,In_1,In_271);
nand U2035 (N_2035,In_85,In_393);
and U2036 (N_2036,In_881,In_764);
and U2037 (N_2037,In_353,In_572);
nor U2038 (N_2038,In_337,In_873);
and U2039 (N_2039,In_697,In_768);
and U2040 (N_2040,In_428,In_46);
and U2041 (N_2041,In_281,In_924);
or U2042 (N_2042,In_846,In_547);
nor U2043 (N_2043,In_532,In_653);
and U2044 (N_2044,In_536,In_914);
and U2045 (N_2045,In_847,In_941);
nand U2046 (N_2046,In_354,In_623);
nor U2047 (N_2047,In_358,In_796);
nor U2048 (N_2048,In_2,In_511);
nor U2049 (N_2049,In_19,In_306);
or U2050 (N_2050,In_559,In_817);
and U2051 (N_2051,In_475,In_922);
nor U2052 (N_2052,In_162,In_874);
nor U2053 (N_2053,In_54,In_405);
nand U2054 (N_2054,In_966,In_628);
nand U2055 (N_2055,In_127,In_512);
nor U2056 (N_2056,In_30,In_617);
and U2057 (N_2057,In_134,In_309);
xnor U2058 (N_2058,In_370,In_859);
nand U2059 (N_2059,In_215,In_620);
xor U2060 (N_2060,In_275,In_479);
and U2061 (N_2061,In_465,In_921);
nor U2062 (N_2062,In_450,In_245);
nand U2063 (N_2063,In_720,In_269);
and U2064 (N_2064,In_435,In_732);
nand U2065 (N_2065,In_865,In_28);
or U2066 (N_2066,In_42,In_585);
nor U2067 (N_2067,In_550,In_187);
nor U2068 (N_2068,In_389,In_658);
xnor U2069 (N_2069,In_570,In_765);
nor U2070 (N_2070,In_189,In_46);
nand U2071 (N_2071,In_277,In_807);
and U2072 (N_2072,In_136,In_151);
and U2073 (N_2073,In_670,In_758);
nor U2074 (N_2074,In_228,In_831);
nor U2075 (N_2075,In_336,In_998);
or U2076 (N_2076,In_375,In_277);
xnor U2077 (N_2077,In_15,In_828);
and U2078 (N_2078,In_736,In_670);
nor U2079 (N_2079,In_13,In_229);
and U2080 (N_2080,In_740,In_638);
nor U2081 (N_2081,In_831,In_320);
and U2082 (N_2082,In_766,In_744);
nand U2083 (N_2083,In_439,In_851);
and U2084 (N_2084,In_833,In_662);
nor U2085 (N_2085,In_248,In_715);
nand U2086 (N_2086,In_639,In_320);
and U2087 (N_2087,In_507,In_683);
nand U2088 (N_2088,In_505,In_271);
nor U2089 (N_2089,In_838,In_401);
nor U2090 (N_2090,In_43,In_457);
nor U2091 (N_2091,In_562,In_309);
nand U2092 (N_2092,In_188,In_584);
nor U2093 (N_2093,In_711,In_944);
and U2094 (N_2094,In_648,In_645);
and U2095 (N_2095,In_654,In_137);
and U2096 (N_2096,In_286,In_284);
xor U2097 (N_2097,In_199,In_79);
or U2098 (N_2098,In_667,In_622);
nand U2099 (N_2099,In_252,In_656);
and U2100 (N_2100,In_980,In_244);
nand U2101 (N_2101,In_400,In_956);
nor U2102 (N_2102,In_755,In_668);
and U2103 (N_2103,In_146,In_739);
nor U2104 (N_2104,In_484,In_758);
nor U2105 (N_2105,In_749,In_435);
and U2106 (N_2106,In_775,In_772);
nand U2107 (N_2107,In_456,In_830);
nand U2108 (N_2108,In_593,In_989);
nand U2109 (N_2109,In_986,In_804);
nand U2110 (N_2110,In_173,In_394);
xor U2111 (N_2111,In_533,In_39);
nand U2112 (N_2112,In_763,In_164);
nand U2113 (N_2113,In_67,In_446);
nor U2114 (N_2114,In_101,In_690);
and U2115 (N_2115,In_997,In_537);
nor U2116 (N_2116,In_376,In_398);
nand U2117 (N_2117,In_347,In_728);
nand U2118 (N_2118,In_836,In_204);
xor U2119 (N_2119,In_797,In_480);
nand U2120 (N_2120,In_383,In_313);
or U2121 (N_2121,In_199,In_91);
xnor U2122 (N_2122,In_811,In_323);
and U2123 (N_2123,In_485,In_634);
and U2124 (N_2124,In_45,In_7);
xnor U2125 (N_2125,In_290,In_672);
nor U2126 (N_2126,In_226,In_700);
or U2127 (N_2127,In_788,In_533);
or U2128 (N_2128,In_851,In_922);
nand U2129 (N_2129,In_862,In_714);
nand U2130 (N_2130,In_72,In_240);
nor U2131 (N_2131,In_742,In_951);
and U2132 (N_2132,In_663,In_752);
nor U2133 (N_2133,In_591,In_509);
nand U2134 (N_2134,In_947,In_615);
nand U2135 (N_2135,In_368,In_255);
nor U2136 (N_2136,In_311,In_857);
and U2137 (N_2137,In_172,In_605);
xor U2138 (N_2138,In_893,In_363);
nor U2139 (N_2139,In_614,In_66);
nor U2140 (N_2140,In_455,In_481);
and U2141 (N_2141,In_350,In_452);
and U2142 (N_2142,In_766,In_931);
and U2143 (N_2143,In_626,In_122);
nor U2144 (N_2144,In_65,In_848);
and U2145 (N_2145,In_4,In_526);
and U2146 (N_2146,In_573,In_972);
and U2147 (N_2147,In_46,In_474);
nor U2148 (N_2148,In_451,In_839);
and U2149 (N_2149,In_698,In_437);
or U2150 (N_2150,In_624,In_751);
or U2151 (N_2151,In_220,In_465);
or U2152 (N_2152,In_853,In_805);
and U2153 (N_2153,In_264,In_985);
or U2154 (N_2154,In_868,In_130);
nand U2155 (N_2155,In_550,In_96);
nor U2156 (N_2156,In_738,In_822);
nand U2157 (N_2157,In_246,In_506);
nand U2158 (N_2158,In_864,In_570);
nor U2159 (N_2159,In_157,In_738);
nor U2160 (N_2160,In_342,In_527);
xor U2161 (N_2161,In_281,In_42);
and U2162 (N_2162,In_17,In_33);
nor U2163 (N_2163,In_620,In_500);
and U2164 (N_2164,In_811,In_994);
nor U2165 (N_2165,In_68,In_680);
nor U2166 (N_2166,In_584,In_428);
nor U2167 (N_2167,In_34,In_651);
nor U2168 (N_2168,In_579,In_240);
nor U2169 (N_2169,In_470,In_737);
or U2170 (N_2170,In_315,In_162);
nor U2171 (N_2171,In_93,In_953);
xnor U2172 (N_2172,In_867,In_207);
xor U2173 (N_2173,In_965,In_270);
and U2174 (N_2174,In_841,In_183);
nor U2175 (N_2175,In_757,In_193);
nor U2176 (N_2176,In_241,In_606);
and U2177 (N_2177,In_184,In_664);
and U2178 (N_2178,In_78,In_377);
xnor U2179 (N_2179,In_897,In_428);
or U2180 (N_2180,In_581,In_711);
or U2181 (N_2181,In_533,In_558);
nor U2182 (N_2182,In_648,In_934);
and U2183 (N_2183,In_409,In_437);
nor U2184 (N_2184,In_207,In_809);
nor U2185 (N_2185,In_640,In_414);
or U2186 (N_2186,In_366,In_608);
nor U2187 (N_2187,In_624,In_612);
or U2188 (N_2188,In_385,In_496);
and U2189 (N_2189,In_863,In_521);
nand U2190 (N_2190,In_904,In_334);
or U2191 (N_2191,In_560,In_456);
or U2192 (N_2192,In_10,In_724);
xor U2193 (N_2193,In_928,In_590);
or U2194 (N_2194,In_697,In_251);
and U2195 (N_2195,In_393,In_768);
and U2196 (N_2196,In_555,In_331);
and U2197 (N_2197,In_810,In_24);
nand U2198 (N_2198,In_612,In_403);
and U2199 (N_2199,In_690,In_692);
nor U2200 (N_2200,In_415,In_679);
nand U2201 (N_2201,In_944,In_802);
nand U2202 (N_2202,In_421,In_271);
or U2203 (N_2203,In_588,In_643);
nor U2204 (N_2204,In_267,In_2);
xor U2205 (N_2205,In_842,In_450);
nor U2206 (N_2206,In_568,In_71);
nand U2207 (N_2207,In_702,In_643);
nor U2208 (N_2208,In_870,In_221);
nand U2209 (N_2209,In_924,In_465);
and U2210 (N_2210,In_528,In_947);
nand U2211 (N_2211,In_306,In_960);
nand U2212 (N_2212,In_615,In_982);
nor U2213 (N_2213,In_112,In_255);
or U2214 (N_2214,In_664,In_972);
and U2215 (N_2215,In_701,In_99);
nor U2216 (N_2216,In_479,In_405);
nor U2217 (N_2217,In_360,In_930);
nand U2218 (N_2218,In_282,In_621);
nor U2219 (N_2219,In_425,In_981);
nand U2220 (N_2220,In_480,In_771);
nand U2221 (N_2221,In_499,In_600);
nor U2222 (N_2222,In_845,In_192);
nand U2223 (N_2223,In_296,In_185);
nor U2224 (N_2224,In_760,In_132);
and U2225 (N_2225,In_736,In_593);
xnor U2226 (N_2226,In_785,In_809);
and U2227 (N_2227,In_938,In_930);
or U2228 (N_2228,In_77,In_100);
and U2229 (N_2229,In_25,In_953);
or U2230 (N_2230,In_981,In_242);
or U2231 (N_2231,In_111,In_743);
and U2232 (N_2232,In_682,In_329);
nor U2233 (N_2233,In_108,In_253);
and U2234 (N_2234,In_411,In_554);
and U2235 (N_2235,In_868,In_914);
or U2236 (N_2236,In_66,In_6);
or U2237 (N_2237,In_254,In_599);
or U2238 (N_2238,In_175,In_511);
or U2239 (N_2239,In_293,In_683);
nor U2240 (N_2240,In_645,In_47);
xnor U2241 (N_2241,In_804,In_203);
and U2242 (N_2242,In_835,In_724);
and U2243 (N_2243,In_230,In_271);
nor U2244 (N_2244,In_96,In_272);
and U2245 (N_2245,In_783,In_202);
or U2246 (N_2246,In_669,In_66);
xor U2247 (N_2247,In_281,In_450);
and U2248 (N_2248,In_5,In_425);
xor U2249 (N_2249,In_607,In_279);
and U2250 (N_2250,In_657,In_641);
or U2251 (N_2251,In_63,In_925);
nand U2252 (N_2252,In_526,In_942);
and U2253 (N_2253,In_774,In_42);
or U2254 (N_2254,In_3,In_533);
and U2255 (N_2255,In_562,In_68);
and U2256 (N_2256,In_658,In_196);
or U2257 (N_2257,In_807,In_273);
or U2258 (N_2258,In_348,In_938);
or U2259 (N_2259,In_904,In_803);
nand U2260 (N_2260,In_800,In_507);
nand U2261 (N_2261,In_111,In_252);
or U2262 (N_2262,In_18,In_953);
and U2263 (N_2263,In_959,In_425);
or U2264 (N_2264,In_714,In_201);
or U2265 (N_2265,In_518,In_832);
and U2266 (N_2266,In_629,In_348);
or U2267 (N_2267,In_861,In_174);
nor U2268 (N_2268,In_774,In_997);
or U2269 (N_2269,In_648,In_172);
or U2270 (N_2270,In_529,In_459);
nor U2271 (N_2271,In_129,In_511);
or U2272 (N_2272,In_349,In_86);
and U2273 (N_2273,In_818,In_79);
nor U2274 (N_2274,In_327,In_172);
nor U2275 (N_2275,In_994,In_588);
nor U2276 (N_2276,In_250,In_725);
nor U2277 (N_2277,In_52,In_634);
nor U2278 (N_2278,In_525,In_465);
or U2279 (N_2279,In_856,In_72);
and U2280 (N_2280,In_159,In_772);
nand U2281 (N_2281,In_489,In_270);
nand U2282 (N_2282,In_358,In_800);
and U2283 (N_2283,In_424,In_416);
or U2284 (N_2284,In_305,In_161);
and U2285 (N_2285,In_820,In_47);
nand U2286 (N_2286,In_754,In_900);
xnor U2287 (N_2287,In_497,In_960);
and U2288 (N_2288,In_859,In_581);
or U2289 (N_2289,In_481,In_130);
or U2290 (N_2290,In_927,In_265);
xor U2291 (N_2291,In_919,In_815);
nand U2292 (N_2292,In_457,In_566);
xnor U2293 (N_2293,In_905,In_914);
or U2294 (N_2294,In_577,In_381);
or U2295 (N_2295,In_148,In_955);
nor U2296 (N_2296,In_729,In_647);
nand U2297 (N_2297,In_626,In_3);
nand U2298 (N_2298,In_822,In_763);
and U2299 (N_2299,In_957,In_711);
or U2300 (N_2300,In_432,In_462);
or U2301 (N_2301,In_242,In_112);
nand U2302 (N_2302,In_938,In_996);
nor U2303 (N_2303,In_858,In_407);
and U2304 (N_2304,In_795,In_189);
nand U2305 (N_2305,In_4,In_810);
or U2306 (N_2306,In_405,In_717);
and U2307 (N_2307,In_784,In_92);
or U2308 (N_2308,In_864,In_361);
and U2309 (N_2309,In_971,In_281);
xor U2310 (N_2310,In_854,In_587);
xor U2311 (N_2311,In_768,In_563);
and U2312 (N_2312,In_34,In_329);
nand U2313 (N_2313,In_374,In_795);
nand U2314 (N_2314,In_977,In_774);
or U2315 (N_2315,In_490,In_841);
xnor U2316 (N_2316,In_391,In_978);
nand U2317 (N_2317,In_737,In_688);
and U2318 (N_2318,In_954,In_590);
nand U2319 (N_2319,In_673,In_889);
and U2320 (N_2320,In_304,In_784);
nand U2321 (N_2321,In_379,In_383);
and U2322 (N_2322,In_916,In_477);
and U2323 (N_2323,In_791,In_772);
nand U2324 (N_2324,In_738,In_981);
nand U2325 (N_2325,In_295,In_436);
xnor U2326 (N_2326,In_94,In_174);
and U2327 (N_2327,In_529,In_750);
or U2328 (N_2328,In_41,In_762);
nand U2329 (N_2329,In_213,In_688);
or U2330 (N_2330,In_970,In_849);
nor U2331 (N_2331,In_987,In_240);
nor U2332 (N_2332,In_738,In_971);
and U2333 (N_2333,In_401,In_592);
and U2334 (N_2334,In_224,In_905);
nor U2335 (N_2335,In_116,In_569);
or U2336 (N_2336,In_755,In_710);
and U2337 (N_2337,In_232,In_364);
or U2338 (N_2338,In_741,In_518);
xnor U2339 (N_2339,In_659,In_520);
nand U2340 (N_2340,In_765,In_103);
nand U2341 (N_2341,In_731,In_286);
nor U2342 (N_2342,In_200,In_628);
or U2343 (N_2343,In_377,In_184);
or U2344 (N_2344,In_221,In_709);
nor U2345 (N_2345,In_251,In_235);
nand U2346 (N_2346,In_908,In_71);
nand U2347 (N_2347,In_731,In_11);
or U2348 (N_2348,In_659,In_741);
or U2349 (N_2349,In_67,In_5);
nor U2350 (N_2350,In_109,In_998);
nor U2351 (N_2351,In_964,In_937);
or U2352 (N_2352,In_678,In_227);
and U2353 (N_2353,In_270,In_683);
and U2354 (N_2354,In_353,In_799);
nand U2355 (N_2355,In_656,In_38);
nor U2356 (N_2356,In_918,In_144);
nand U2357 (N_2357,In_874,In_484);
or U2358 (N_2358,In_50,In_492);
and U2359 (N_2359,In_838,In_752);
and U2360 (N_2360,In_22,In_723);
or U2361 (N_2361,In_720,In_63);
and U2362 (N_2362,In_463,In_274);
or U2363 (N_2363,In_814,In_83);
or U2364 (N_2364,In_834,In_189);
or U2365 (N_2365,In_950,In_209);
or U2366 (N_2366,In_178,In_214);
and U2367 (N_2367,In_125,In_411);
nor U2368 (N_2368,In_608,In_995);
nand U2369 (N_2369,In_449,In_536);
nand U2370 (N_2370,In_524,In_127);
nor U2371 (N_2371,In_129,In_855);
or U2372 (N_2372,In_211,In_186);
nand U2373 (N_2373,In_795,In_23);
or U2374 (N_2374,In_874,In_714);
nor U2375 (N_2375,In_578,In_567);
nor U2376 (N_2376,In_63,In_240);
nor U2377 (N_2377,In_465,In_385);
nor U2378 (N_2378,In_486,In_324);
and U2379 (N_2379,In_699,In_120);
nor U2380 (N_2380,In_871,In_704);
nor U2381 (N_2381,In_72,In_413);
and U2382 (N_2382,In_420,In_475);
or U2383 (N_2383,In_171,In_294);
nor U2384 (N_2384,In_15,In_524);
and U2385 (N_2385,In_877,In_741);
nand U2386 (N_2386,In_144,In_466);
and U2387 (N_2387,In_29,In_34);
and U2388 (N_2388,In_624,In_611);
or U2389 (N_2389,In_990,In_151);
or U2390 (N_2390,In_975,In_3);
and U2391 (N_2391,In_882,In_653);
nand U2392 (N_2392,In_201,In_1);
and U2393 (N_2393,In_421,In_13);
and U2394 (N_2394,In_878,In_988);
or U2395 (N_2395,In_27,In_480);
xor U2396 (N_2396,In_534,In_482);
or U2397 (N_2397,In_475,In_353);
and U2398 (N_2398,In_546,In_987);
nand U2399 (N_2399,In_815,In_610);
or U2400 (N_2400,In_233,In_313);
nand U2401 (N_2401,In_595,In_75);
nand U2402 (N_2402,In_70,In_234);
xnor U2403 (N_2403,In_225,In_7);
nand U2404 (N_2404,In_999,In_390);
nor U2405 (N_2405,In_565,In_840);
nand U2406 (N_2406,In_40,In_768);
nor U2407 (N_2407,In_330,In_421);
nor U2408 (N_2408,In_584,In_123);
xor U2409 (N_2409,In_579,In_372);
nand U2410 (N_2410,In_612,In_40);
nand U2411 (N_2411,In_879,In_609);
nand U2412 (N_2412,In_76,In_698);
nand U2413 (N_2413,In_81,In_877);
and U2414 (N_2414,In_909,In_749);
nand U2415 (N_2415,In_581,In_843);
nand U2416 (N_2416,In_0,In_843);
or U2417 (N_2417,In_982,In_541);
nand U2418 (N_2418,In_331,In_912);
and U2419 (N_2419,In_602,In_476);
or U2420 (N_2420,In_289,In_519);
nor U2421 (N_2421,In_466,In_496);
nor U2422 (N_2422,In_409,In_183);
xnor U2423 (N_2423,In_711,In_50);
nand U2424 (N_2424,In_401,In_603);
or U2425 (N_2425,In_551,In_471);
nand U2426 (N_2426,In_640,In_62);
and U2427 (N_2427,In_580,In_481);
or U2428 (N_2428,In_264,In_516);
nor U2429 (N_2429,In_494,In_762);
xor U2430 (N_2430,In_482,In_945);
nor U2431 (N_2431,In_605,In_760);
nor U2432 (N_2432,In_622,In_8);
and U2433 (N_2433,In_323,In_74);
or U2434 (N_2434,In_407,In_651);
nor U2435 (N_2435,In_832,In_163);
nand U2436 (N_2436,In_45,In_657);
nand U2437 (N_2437,In_724,In_760);
and U2438 (N_2438,In_157,In_200);
or U2439 (N_2439,In_429,In_438);
xnor U2440 (N_2440,In_539,In_92);
or U2441 (N_2441,In_870,In_112);
and U2442 (N_2442,In_868,In_374);
and U2443 (N_2443,In_140,In_959);
and U2444 (N_2444,In_728,In_918);
xnor U2445 (N_2445,In_689,In_2);
and U2446 (N_2446,In_188,In_314);
nor U2447 (N_2447,In_324,In_537);
or U2448 (N_2448,In_895,In_568);
or U2449 (N_2449,In_903,In_788);
nor U2450 (N_2450,In_392,In_689);
and U2451 (N_2451,In_87,In_881);
or U2452 (N_2452,In_967,In_831);
and U2453 (N_2453,In_946,In_993);
and U2454 (N_2454,In_711,In_180);
nor U2455 (N_2455,In_442,In_969);
and U2456 (N_2456,In_13,In_763);
nand U2457 (N_2457,In_929,In_299);
or U2458 (N_2458,In_819,In_77);
xnor U2459 (N_2459,In_669,In_743);
xnor U2460 (N_2460,In_882,In_241);
nand U2461 (N_2461,In_66,In_487);
or U2462 (N_2462,In_251,In_273);
nor U2463 (N_2463,In_632,In_804);
xnor U2464 (N_2464,In_513,In_867);
or U2465 (N_2465,In_598,In_130);
xor U2466 (N_2466,In_662,In_823);
nor U2467 (N_2467,In_828,In_495);
nand U2468 (N_2468,In_873,In_749);
and U2469 (N_2469,In_278,In_657);
xnor U2470 (N_2470,In_34,In_365);
nand U2471 (N_2471,In_577,In_134);
nor U2472 (N_2472,In_810,In_660);
nor U2473 (N_2473,In_140,In_916);
and U2474 (N_2474,In_471,In_488);
nand U2475 (N_2475,In_311,In_333);
and U2476 (N_2476,In_939,In_415);
nand U2477 (N_2477,In_545,In_987);
nor U2478 (N_2478,In_714,In_247);
and U2479 (N_2479,In_580,In_785);
nor U2480 (N_2480,In_30,In_871);
nor U2481 (N_2481,In_447,In_770);
xnor U2482 (N_2482,In_495,In_121);
nand U2483 (N_2483,In_491,In_244);
and U2484 (N_2484,In_23,In_495);
nor U2485 (N_2485,In_395,In_96);
nor U2486 (N_2486,In_955,In_906);
xnor U2487 (N_2487,In_525,In_620);
and U2488 (N_2488,In_749,In_677);
and U2489 (N_2489,In_935,In_777);
nand U2490 (N_2490,In_558,In_148);
or U2491 (N_2491,In_730,In_978);
and U2492 (N_2492,In_213,In_7);
or U2493 (N_2493,In_613,In_784);
and U2494 (N_2494,In_660,In_450);
and U2495 (N_2495,In_873,In_557);
nand U2496 (N_2496,In_690,In_527);
or U2497 (N_2497,In_543,In_734);
nand U2498 (N_2498,In_656,In_512);
and U2499 (N_2499,In_280,In_159);
and U2500 (N_2500,In_562,In_510);
and U2501 (N_2501,In_834,In_659);
nor U2502 (N_2502,In_496,In_359);
nand U2503 (N_2503,In_244,In_52);
or U2504 (N_2504,In_315,In_62);
or U2505 (N_2505,In_619,In_380);
nor U2506 (N_2506,In_267,In_367);
nand U2507 (N_2507,In_77,In_230);
or U2508 (N_2508,In_694,In_596);
or U2509 (N_2509,In_627,In_9);
and U2510 (N_2510,In_21,In_872);
or U2511 (N_2511,In_826,In_148);
or U2512 (N_2512,In_51,In_196);
or U2513 (N_2513,In_334,In_262);
or U2514 (N_2514,In_398,In_151);
and U2515 (N_2515,In_983,In_158);
and U2516 (N_2516,In_189,In_118);
or U2517 (N_2517,In_649,In_661);
and U2518 (N_2518,In_18,In_152);
nor U2519 (N_2519,In_971,In_179);
nand U2520 (N_2520,In_591,In_816);
xnor U2521 (N_2521,In_708,In_695);
nand U2522 (N_2522,In_758,In_271);
or U2523 (N_2523,In_693,In_820);
or U2524 (N_2524,In_711,In_993);
nand U2525 (N_2525,In_243,In_353);
nand U2526 (N_2526,In_853,In_625);
or U2527 (N_2527,In_239,In_863);
nor U2528 (N_2528,In_356,In_842);
and U2529 (N_2529,In_996,In_76);
and U2530 (N_2530,In_442,In_22);
or U2531 (N_2531,In_458,In_450);
or U2532 (N_2532,In_817,In_814);
nand U2533 (N_2533,In_366,In_427);
nor U2534 (N_2534,In_361,In_861);
or U2535 (N_2535,In_775,In_13);
or U2536 (N_2536,In_297,In_426);
xnor U2537 (N_2537,In_663,In_194);
xor U2538 (N_2538,In_523,In_43);
and U2539 (N_2539,In_534,In_855);
and U2540 (N_2540,In_858,In_759);
nand U2541 (N_2541,In_641,In_753);
nor U2542 (N_2542,In_644,In_125);
xor U2543 (N_2543,In_743,In_408);
or U2544 (N_2544,In_771,In_847);
or U2545 (N_2545,In_959,In_536);
nor U2546 (N_2546,In_605,In_689);
or U2547 (N_2547,In_287,In_919);
or U2548 (N_2548,In_585,In_0);
or U2549 (N_2549,In_57,In_48);
nor U2550 (N_2550,In_21,In_377);
nor U2551 (N_2551,In_898,In_288);
or U2552 (N_2552,In_180,In_830);
xor U2553 (N_2553,In_510,In_234);
and U2554 (N_2554,In_842,In_858);
nand U2555 (N_2555,In_203,In_334);
and U2556 (N_2556,In_129,In_656);
or U2557 (N_2557,In_343,In_993);
xor U2558 (N_2558,In_820,In_173);
nand U2559 (N_2559,In_762,In_557);
nor U2560 (N_2560,In_996,In_881);
or U2561 (N_2561,In_840,In_784);
and U2562 (N_2562,In_474,In_430);
nand U2563 (N_2563,In_127,In_870);
nand U2564 (N_2564,In_637,In_411);
xor U2565 (N_2565,In_769,In_11);
nor U2566 (N_2566,In_138,In_808);
and U2567 (N_2567,In_909,In_175);
nor U2568 (N_2568,In_565,In_986);
xnor U2569 (N_2569,In_396,In_215);
or U2570 (N_2570,In_133,In_705);
nor U2571 (N_2571,In_207,In_765);
nand U2572 (N_2572,In_563,In_599);
nor U2573 (N_2573,In_827,In_199);
xnor U2574 (N_2574,In_487,In_310);
nand U2575 (N_2575,In_818,In_7);
nor U2576 (N_2576,In_357,In_330);
or U2577 (N_2577,In_286,In_376);
or U2578 (N_2578,In_450,In_583);
or U2579 (N_2579,In_60,In_62);
nand U2580 (N_2580,In_485,In_24);
and U2581 (N_2581,In_479,In_461);
or U2582 (N_2582,In_808,In_481);
nand U2583 (N_2583,In_806,In_197);
nor U2584 (N_2584,In_801,In_702);
nand U2585 (N_2585,In_937,In_295);
nor U2586 (N_2586,In_526,In_104);
or U2587 (N_2587,In_101,In_24);
xnor U2588 (N_2588,In_174,In_70);
and U2589 (N_2589,In_113,In_602);
and U2590 (N_2590,In_850,In_446);
or U2591 (N_2591,In_830,In_208);
nor U2592 (N_2592,In_230,In_273);
or U2593 (N_2593,In_674,In_965);
nor U2594 (N_2594,In_212,In_441);
or U2595 (N_2595,In_500,In_190);
and U2596 (N_2596,In_228,In_825);
nand U2597 (N_2597,In_943,In_92);
and U2598 (N_2598,In_178,In_456);
or U2599 (N_2599,In_516,In_368);
nor U2600 (N_2600,In_407,In_212);
nand U2601 (N_2601,In_52,In_288);
nor U2602 (N_2602,In_157,In_996);
and U2603 (N_2603,In_52,In_243);
and U2604 (N_2604,In_784,In_229);
xnor U2605 (N_2605,In_33,In_82);
or U2606 (N_2606,In_810,In_957);
nor U2607 (N_2607,In_175,In_719);
and U2608 (N_2608,In_597,In_697);
or U2609 (N_2609,In_88,In_761);
and U2610 (N_2610,In_392,In_202);
nand U2611 (N_2611,In_24,In_496);
and U2612 (N_2612,In_408,In_817);
xnor U2613 (N_2613,In_633,In_221);
nor U2614 (N_2614,In_749,In_621);
or U2615 (N_2615,In_257,In_645);
and U2616 (N_2616,In_114,In_836);
xor U2617 (N_2617,In_192,In_174);
xor U2618 (N_2618,In_62,In_590);
nand U2619 (N_2619,In_65,In_912);
or U2620 (N_2620,In_221,In_327);
or U2621 (N_2621,In_416,In_955);
nand U2622 (N_2622,In_277,In_52);
and U2623 (N_2623,In_548,In_306);
and U2624 (N_2624,In_804,In_988);
and U2625 (N_2625,In_64,In_602);
nand U2626 (N_2626,In_889,In_777);
or U2627 (N_2627,In_832,In_705);
or U2628 (N_2628,In_866,In_794);
nor U2629 (N_2629,In_876,In_499);
and U2630 (N_2630,In_191,In_260);
nand U2631 (N_2631,In_235,In_816);
nor U2632 (N_2632,In_538,In_939);
and U2633 (N_2633,In_989,In_707);
nand U2634 (N_2634,In_437,In_99);
and U2635 (N_2635,In_148,In_41);
nor U2636 (N_2636,In_809,In_74);
xor U2637 (N_2637,In_549,In_130);
nand U2638 (N_2638,In_353,In_126);
nand U2639 (N_2639,In_876,In_83);
nand U2640 (N_2640,In_935,In_821);
nand U2641 (N_2641,In_555,In_746);
nor U2642 (N_2642,In_230,In_996);
and U2643 (N_2643,In_918,In_183);
nand U2644 (N_2644,In_326,In_803);
nor U2645 (N_2645,In_808,In_830);
or U2646 (N_2646,In_377,In_693);
and U2647 (N_2647,In_539,In_215);
nand U2648 (N_2648,In_21,In_896);
and U2649 (N_2649,In_155,In_987);
nand U2650 (N_2650,In_371,In_366);
nor U2651 (N_2651,In_42,In_467);
and U2652 (N_2652,In_761,In_635);
or U2653 (N_2653,In_331,In_725);
nor U2654 (N_2654,In_121,In_979);
nand U2655 (N_2655,In_335,In_187);
nor U2656 (N_2656,In_92,In_364);
and U2657 (N_2657,In_252,In_563);
nor U2658 (N_2658,In_56,In_201);
and U2659 (N_2659,In_706,In_699);
and U2660 (N_2660,In_374,In_607);
and U2661 (N_2661,In_329,In_650);
or U2662 (N_2662,In_232,In_634);
nand U2663 (N_2663,In_40,In_777);
or U2664 (N_2664,In_238,In_597);
nand U2665 (N_2665,In_459,In_677);
and U2666 (N_2666,In_348,In_81);
nor U2667 (N_2667,In_238,In_293);
and U2668 (N_2668,In_671,In_663);
nand U2669 (N_2669,In_128,In_327);
nand U2670 (N_2670,In_557,In_413);
nor U2671 (N_2671,In_912,In_70);
or U2672 (N_2672,In_18,In_476);
nand U2673 (N_2673,In_299,In_493);
xor U2674 (N_2674,In_928,In_399);
and U2675 (N_2675,In_699,In_538);
or U2676 (N_2676,In_491,In_18);
nand U2677 (N_2677,In_619,In_137);
nand U2678 (N_2678,In_202,In_279);
and U2679 (N_2679,In_328,In_900);
nand U2680 (N_2680,In_22,In_968);
nor U2681 (N_2681,In_681,In_269);
nand U2682 (N_2682,In_181,In_854);
xor U2683 (N_2683,In_462,In_105);
and U2684 (N_2684,In_442,In_869);
and U2685 (N_2685,In_398,In_604);
nor U2686 (N_2686,In_46,In_809);
or U2687 (N_2687,In_378,In_87);
and U2688 (N_2688,In_958,In_754);
nor U2689 (N_2689,In_539,In_577);
nor U2690 (N_2690,In_290,In_9);
nor U2691 (N_2691,In_205,In_281);
nor U2692 (N_2692,In_256,In_249);
xnor U2693 (N_2693,In_17,In_170);
nor U2694 (N_2694,In_893,In_520);
nand U2695 (N_2695,In_928,In_333);
or U2696 (N_2696,In_824,In_323);
and U2697 (N_2697,In_709,In_861);
nor U2698 (N_2698,In_639,In_268);
and U2699 (N_2699,In_682,In_239);
and U2700 (N_2700,In_115,In_715);
and U2701 (N_2701,In_78,In_729);
nor U2702 (N_2702,In_720,In_705);
nand U2703 (N_2703,In_833,In_605);
nand U2704 (N_2704,In_112,In_317);
and U2705 (N_2705,In_84,In_199);
xor U2706 (N_2706,In_884,In_944);
and U2707 (N_2707,In_920,In_183);
nor U2708 (N_2708,In_239,In_726);
or U2709 (N_2709,In_489,In_195);
and U2710 (N_2710,In_547,In_787);
nand U2711 (N_2711,In_382,In_302);
nand U2712 (N_2712,In_355,In_139);
nand U2713 (N_2713,In_64,In_685);
or U2714 (N_2714,In_829,In_450);
and U2715 (N_2715,In_717,In_905);
nor U2716 (N_2716,In_9,In_336);
and U2717 (N_2717,In_800,In_175);
or U2718 (N_2718,In_626,In_539);
and U2719 (N_2719,In_860,In_834);
and U2720 (N_2720,In_771,In_453);
nor U2721 (N_2721,In_841,In_739);
xor U2722 (N_2722,In_726,In_135);
nand U2723 (N_2723,In_775,In_833);
nand U2724 (N_2724,In_194,In_595);
or U2725 (N_2725,In_639,In_171);
nand U2726 (N_2726,In_186,In_31);
nand U2727 (N_2727,In_509,In_552);
nor U2728 (N_2728,In_168,In_621);
nor U2729 (N_2729,In_118,In_734);
nor U2730 (N_2730,In_262,In_791);
xor U2731 (N_2731,In_333,In_788);
or U2732 (N_2732,In_861,In_260);
and U2733 (N_2733,In_931,In_222);
or U2734 (N_2734,In_302,In_206);
or U2735 (N_2735,In_121,In_286);
nand U2736 (N_2736,In_6,In_184);
nand U2737 (N_2737,In_797,In_216);
nor U2738 (N_2738,In_831,In_538);
or U2739 (N_2739,In_229,In_397);
nand U2740 (N_2740,In_372,In_275);
or U2741 (N_2741,In_645,In_157);
and U2742 (N_2742,In_890,In_328);
and U2743 (N_2743,In_606,In_499);
and U2744 (N_2744,In_1,In_580);
nor U2745 (N_2745,In_571,In_60);
nand U2746 (N_2746,In_95,In_505);
or U2747 (N_2747,In_826,In_9);
nor U2748 (N_2748,In_250,In_458);
nand U2749 (N_2749,In_564,In_454);
and U2750 (N_2750,In_254,In_947);
or U2751 (N_2751,In_410,In_159);
or U2752 (N_2752,In_385,In_234);
and U2753 (N_2753,In_825,In_247);
or U2754 (N_2754,In_550,In_687);
nor U2755 (N_2755,In_41,In_865);
nand U2756 (N_2756,In_320,In_292);
and U2757 (N_2757,In_886,In_512);
nand U2758 (N_2758,In_665,In_103);
nor U2759 (N_2759,In_488,In_159);
and U2760 (N_2760,In_61,In_989);
xnor U2761 (N_2761,In_869,In_899);
xor U2762 (N_2762,In_493,In_601);
or U2763 (N_2763,In_764,In_542);
or U2764 (N_2764,In_35,In_893);
xnor U2765 (N_2765,In_979,In_727);
or U2766 (N_2766,In_533,In_560);
nor U2767 (N_2767,In_597,In_900);
nor U2768 (N_2768,In_360,In_4);
and U2769 (N_2769,In_678,In_370);
or U2770 (N_2770,In_208,In_922);
nor U2771 (N_2771,In_42,In_825);
or U2772 (N_2772,In_376,In_731);
and U2773 (N_2773,In_206,In_388);
nand U2774 (N_2774,In_747,In_587);
or U2775 (N_2775,In_567,In_580);
nor U2776 (N_2776,In_642,In_598);
nand U2777 (N_2777,In_671,In_390);
nor U2778 (N_2778,In_652,In_826);
or U2779 (N_2779,In_36,In_92);
or U2780 (N_2780,In_61,In_307);
nand U2781 (N_2781,In_544,In_893);
or U2782 (N_2782,In_468,In_706);
nand U2783 (N_2783,In_331,In_861);
or U2784 (N_2784,In_250,In_363);
nand U2785 (N_2785,In_217,In_768);
and U2786 (N_2786,In_237,In_752);
nand U2787 (N_2787,In_747,In_258);
nand U2788 (N_2788,In_666,In_918);
or U2789 (N_2789,In_322,In_276);
xor U2790 (N_2790,In_358,In_491);
or U2791 (N_2791,In_909,In_326);
and U2792 (N_2792,In_464,In_380);
nor U2793 (N_2793,In_301,In_821);
or U2794 (N_2794,In_514,In_862);
nor U2795 (N_2795,In_545,In_785);
nor U2796 (N_2796,In_334,In_623);
or U2797 (N_2797,In_376,In_830);
nand U2798 (N_2798,In_570,In_921);
nand U2799 (N_2799,In_45,In_501);
or U2800 (N_2800,In_206,In_923);
nor U2801 (N_2801,In_883,In_46);
or U2802 (N_2802,In_443,In_373);
nor U2803 (N_2803,In_596,In_153);
nand U2804 (N_2804,In_55,In_114);
nand U2805 (N_2805,In_968,In_211);
nand U2806 (N_2806,In_812,In_886);
nand U2807 (N_2807,In_862,In_230);
nand U2808 (N_2808,In_570,In_744);
or U2809 (N_2809,In_272,In_472);
or U2810 (N_2810,In_312,In_252);
and U2811 (N_2811,In_113,In_869);
nor U2812 (N_2812,In_4,In_262);
nor U2813 (N_2813,In_500,In_875);
nand U2814 (N_2814,In_668,In_441);
and U2815 (N_2815,In_245,In_966);
nand U2816 (N_2816,In_254,In_391);
nor U2817 (N_2817,In_529,In_558);
and U2818 (N_2818,In_697,In_667);
or U2819 (N_2819,In_722,In_900);
nor U2820 (N_2820,In_366,In_96);
or U2821 (N_2821,In_14,In_133);
nor U2822 (N_2822,In_412,In_227);
nor U2823 (N_2823,In_2,In_207);
and U2824 (N_2824,In_453,In_416);
nand U2825 (N_2825,In_532,In_485);
and U2826 (N_2826,In_173,In_991);
nand U2827 (N_2827,In_216,In_711);
and U2828 (N_2828,In_188,In_722);
nor U2829 (N_2829,In_537,In_562);
and U2830 (N_2830,In_494,In_460);
nand U2831 (N_2831,In_728,In_795);
xnor U2832 (N_2832,In_539,In_329);
and U2833 (N_2833,In_528,In_218);
and U2834 (N_2834,In_74,In_904);
and U2835 (N_2835,In_787,In_488);
xor U2836 (N_2836,In_330,In_485);
and U2837 (N_2837,In_161,In_488);
nand U2838 (N_2838,In_964,In_629);
nor U2839 (N_2839,In_867,In_455);
nand U2840 (N_2840,In_362,In_88);
and U2841 (N_2841,In_76,In_207);
or U2842 (N_2842,In_708,In_723);
or U2843 (N_2843,In_178,In_799);
or U2844 (N_2844,In_946,In_866);
nand U2845 (N_2845,In_210,In_178);
or U2846 (N_2846,In_536,In_405);
or U2847 (N_2847,In_222,In_606);
and U2848 (N_2848,In_34,In_514);
and U2849 (N_2849,In_292,In_607);
xnor U2850 (N_2850,In_962,In_527);
and U2851 (N_2851,In_310,In_494);
or U2852 (N_2852,In_537,In_971);
or U2853 (N_2853,In_674,In_111);
or U2854 (N_2854,In_457,In_179);
xor U2855 (N_2855,In_730,In_35);
nor U2856 (N_2856,In_350,In_851);
nor U2857 (N_2857,In_11,In_134);
and U2858 (N_2858,In_619,In_547);
nand U2859 (N_2859,In_957,In_616);
and U2860 (N_2860,In_882,In_279);
nand U2861 (N_2861,In_105,In_180);
xnor U2862 (N_2862,In_533,In_200);
and U2863 (N_2863,In_746,In_118);
nor U2864 (N_2864,In_330,In_16);
or U2865 (N_2865,In_746,In_126);
nor U2866 (N_2866,In_200,In_353);
nor U2867 (N_2867,In_633,In_540);
or U2868 (N_2868,In_767,In_40);
nand U2869 (N_2869,In_540,In_629);
nor U2870 (N_2870,In_5,In_26);
nor U2871 (N_2871,In_391,In_442);
xnor U2872 (N_2872,In_26,In_852);
nor U2873 (N_2873,In_748,In_420);
nor U2874 (N_2874,In_400,In_352);
nor U2875 (N_2875,In_133,In_111);
nor U2876 (N_2876,In_70,In_48);
nand U2877 (N_2877,In_272,In_325);
nand U2878 (N_2878,In_832,In_107);
nor U2879 (N_2879,In_771,In_273);
nand U2880 (N_2880,In_150,In_337);
or U2881 (N_2881,In_545,In_134);
nor U2882 (N_2882,In_394,In_713);
and U2883 (N_2883,In_300,In_432);
and U2884 (N_2884,In_257,In_495);
or U2885 (N_2885,In_763,In_502);
nand U2886 (N_2886,In_930,In_19);
nand U2887 (N_2887,In_601,In_567);
nor U2888 (N_2888,In_496,In_30);
nor U2889 (N_2889,In_528,In_687);
nor U2890 (N_2890,In_520,In_487);
nor U2891 (N_2891,In_476,In_721);
nor U2892 (N_2892,In_993,In_737);
nor U2893 (N_2893,In_876,In_577);
xnor U2894 (N_2894,In_671,In_939);
and U2895 (N_2895,In_111,In_969);
nand U2896 (N_2896,In_144,In_847);
or U2897 (N_2897,In_898,In_700);
or U2898 (N_2898,In_490,In_224);
and U2899 (N_2899,In_958,In_218);
xnor U2900 (N_2900,In_297,In_279);
nand U2901 (N_2901,In_111,In_646);
xnor U2902 (N_2902,In_43,In_622);
or U2903 (N_2903,In_214,In_707);
and U2904 (N_2904,In_247,In_744);
xor U2905 (N_2905,In_314,In_125);
nor U2906 (N_2906,In_817,In_583);
or U2907 (N_2907,In_674,In_80);
nor U2908 (N_2908,In_693,In_670);
xor U2909 (N_2909,In_343,In_728);
nand U2910 (N_2910,In_448,In_807);
xor U2911 (N_2911,In_54,In_73);
or U2912 (N_2912,In_559,In_164);
xor U2913 (N_2913,In_953,In_899);
and U2914 (N_2914,In_509,In_172);
xnor U2915 (N_2915,In_522,In_409);
nor U2916 (N_2916,In_779,In_193);
xor U2917 (N_2917,In_943,In_700);
or U2918 (N_2918,In_605,In_256);
nand U2919 (N_2919,In_415,In_986);
or U2920 (N_2920,In_105,In_409);
nor U2921 (N_2921,In_599,In_32);
and U2922 (N_2922,In_398,In_359);
and U2923 (N_2923,In_788,In_277);
nor U2924 (N_2924,In_824,In_828);
nand U2925 (N_2925,In_986,In_615);
xor U2926 (N_2926,In_609,In_396);
nor U2927 (N_2927,In_866,In_80);
nor U2928 (N_2928,In_389,In_641);
or U2929 (N_2929,In_32,In_498);
and U2930 (N_2930,In_650,In_587);
and U2931 (N_2931,In_49,In_896);
nand U2932 (N_2932,In_446,In_124);
or U2933 (N_2933,In_845,In_162);
nand U2934 (N_2934,In_214,In_339);
nand U2935 (N_2935,In_823,In_796);
nand U2936 (N_2936,In_473,In_884);
or U2937 (N_2937,In_903,In_641);
or U2938 (N_2938,In_739,In_345);
or U2939 (N_2939,In_537,In_345);
nor U2940 (N_2940,In_357,In_217);
xor U2941 (N_2941,In_279,In_237);
and U2942 (N_2942,In_863,In_151);
nand U2943 (N_2943,In_474,In_821);
nor U2944 (N_2944,In_751,In_419);
and U2945 (N_2945,In_513,In_741);
nor U2946 (N_2946,In_235,In_862);
and U2947 (N_2947,In_823,In_504);
and U2948 (N_2948,In_632,In_233);
and U2949 (N_2949,In_331,In_473);
or U2950 (N_2950,In_585,In_104);
or U2951 (N_2951,In_530,In_193);
and U2952 (N_2952,In_716,In_338);
and U2953 (N_2953,In_903,In_306);
nor U2954 (N_2954,In_276,In_45);
or U2955 (N_2955,In_27,In_910);
nor U2956 (N_2956,In_583,In_452);
nor U2957 (N_2957,In_512,In_524);
and U2958 (N_2958,In_771,In_247);
or U2959 (N_2959,In_861,In_661);
nand U2960 (N_2960,In_547,In_228);
nand U2961 (N_2961,In_943,In_919);
and U2962 (N_2962,In_64,In_593);
nand U2963 (N_2963,In_994,In_831);
nor U2964 (N_2964,In_487,In_803);
xor U2965 (N_2965,In_485,In_201);
and U2966 (N_2966,In_566,In_809);
nor U2967 (N_2967,In_498,In_908);
or U2968 (N_2968,In_870,In_571);
nand U2969 (N_2969,In_943,In_123);
and U2970 (N_2970,In_174,In_859);
and U2971 (N_2971,In_142,In_272);
and U2972 (N_2972,In_444,In_384);
nand U2973 (N_2973,In_183,In_645);
nor U2974 (N_2974,In_928,In_390);
nor U2975 (N_2975,In_942,In_124);
xor U2976 (N_2976,In_933,In_680);
xnor U2977 (N_2977,In_702,In_489);
nor U2978 (N_2978,In_406,In_764);
xor U2979 (N_2979,In_92,In_194);
or U2980 (N_2980,In_352,In_947);
nand U2981 (N_2981,In_921,In_53);
nand U2982 (N_2982,In_919,In_421);
nor U2983 (N_2983,In_602,In_701);
nor U2984 (N_2984,In_461,In_245);
and U2985 (N_2985,In_211,In_807);
or U2986 (N_2986,In_547,In_902);
or U2987 (N_2987,In_695,In_447);
nor U2988 (N_2988,In_179,In_987);
and U2989 (N_2989,In_934,In_848);
and U2990 (N_2990,In_732,In_129);
xor U2991 (N_2991,In_860,In_757);
or U2992 (N_2992,In_999,In_488);
nor U2993 (N_2993,In_173,In_883);
and U2994 (N_2994,In_775,In_115);
and U2995 (N_2995,In_724,In_799);
xnor U2996 (N_2996,In_257,In_373);
or U2997 (N_2997,In_657,In_983);
nor U2998 (N_2998,In_500,In_539);
nand U2999 (N_2999,In_751,In_63);
and U3000 (N_3000,In_216,In_101);
or U3001 (N_3001,In_884,In_167);
and U3002 (N_3002,In_978,In_991);
nand U3003 (N_3003,In_545,In_333);
nor U3004 (N_3004,In_425,In_720);
xnor U3005 (N_3005,In_45,In_126);
or U3006 (N_3006,In_560,In_861);
nand U3007 (N_3007,In_235,In_937);
nor U3008 (N_3008,In_558,In_658);
nor U3009 (N_3009,In_491,In_363);
nand U3010 (N_3010,In_143,In_92);
or U3011 (N_3011,In_329,In_426);
nor U3012 (N_3012,In_241,In_839);
or U3013 (N_3013,In_808,In_883);
or U3014 (N_3014,In_470,In_869);
or U3015 (N_3015,In_447,In_306);
xor U3016 (N_3016,In_904,In_868);
or U3017 (N_3017,In_968,In_87);
xnor U3018 (N_3018,In_438,In_953);
nor U3019 (N_3019,In_904,In_833);
xor U3020 (N_3020,In_425,In_972);
and U3021 (N_3021,In_260,In_906);
or U3022 (N_3022,In_550,In_357);
nor U3023 (N_3023,In_488,In_456);
nand U3024 (N_3024,In_851,In_997);
nor U3025 (N_3025,In_976,In_657);
or U3026 (N_3026,In_470,In_109);
and U3027 (N_3027,In_313,In_714);
or U3028 (N_3028,In_588,In_491);
or U3029 (N_3029,In_386,In_509);
xnor U3030 (N_3030,In_64,In_349);
or U3031 (N_3031,In_750,In_719);
and U3032 (N_3032,In_363,In_679);
or U3033 (N_3033,In_463,In_168);
xor U3034 (N_3034,In_382,In_34);
nand U3035 (N_3035,In_727,In_568);
xnor U3036 (N_3036,In_21,In_366);
or U3037 (N_3037,In_721,In_80);
nand U3038 (N_3038,In_151,In_150);
xor U3039 (N_3039,In_981,In_734);
nor U3040 (N_3040,In_399,In_520);
nor U3041 (N_3041,In_359,In_155);
xor U3042 (N_3042,In_811,In_382);
nand U3043 (N_3043,In_520,In_170);
nand U3044 (N_3044,In_468,In_161);
and U3045 (N_3045,In_169,In_503);
nand U3046 (N_3046,In_291,In_256);
nor U3047 (N_3047,In_713,In_480);
nor U3048 (N_3048,In_512,In_643);
nor U3049 (N_3049,In_163,In_718);
or U3050 (N_3050,In_171,In_32);
xnor U3051 (N_3051,In_591,In_153);
nand U3052 (N_3052,In_820,In_509);
nor U3053 (N_3053,In_416,In_534);
nor U3054 (N_3054,In_565,In_80);
or U3055 (N_3055,In_689,In_704);
nor U3056 (N_3056,In_411,In_830);
nor U3057 (N_3057,In_821,In_191);
or U3058 (N_3058,In_471,In_315);
or U3059 (N_3059,In_180,In_4);
xor U3060 (N_3060,In_789,In_664);
nand U3061 (N_3061,In_183,In_915);
nand U3062 (N_3062,In_902,In_880);
nor U3063 (N_3063,In_281,In_530);
nand U3064 (N_3064,In_732,In_826);
and U3065 (N_3065,In_302,In_655);
nor U3066 (N_3066,In_36,In_515);
nand U3067 (N_3067,In_365,In_307);
nand U3068 (N_3068,In_342,In_975);
and U3069 (N_3069,In_208,In_916);
nand U3070 (N_3070,In_262,In_678);
xnor U3071 (N_3071,In_551,In_609);
nor U3072 (N_3072,In_547,In_404);
nand U3073 (N_3073,In_887,In_841);
nor U3074 (N_3074,In_122,In_97);
or U3075 (N_3075,In_369,In_856);
or U3076 (N_3076,In_717,In_367);
nand U3077 (N_3077,In_366,In_241);
nand U3078 (N_3078,In_378,In_450);
xnor U3079 (N_3079,In_564,In_182);
and U3080 (N_3080,In_964,In_656);
and U3081 (N_3081,In_333,In_27);
nand U3082 (N_3082,In_3,In_881);
or U3083 (N_3083,In_70,In_753);
nand U3084 (N_3084,In_238,In_477);
nand U3085 (N_3085,In_175,In_836);
and U3086 (N_3086,In_170,In_860);
xnor U3087 (N_3087,In_526,In_69);
xor U3088 (N_3088,In_544,In_602);
or U3089 (N_3089,In_948,In_770);
or U3090 (N_3090,In_75,In_369);
or U3091 (N_3091,In_839,In_87);
nor U3092 (N_3092,In_532,In_54);
or U3093 (N_3093,In_646,In_470);
and U3094 (N_3094,In_488,In_305);
xnor U3095 (N_3095,In_985,In_363);
nor U3096 (N_3096,In_822,In_495);
nor U3097 (N_3097,In_507,In_983);
and U3098 (N_3098,In_563,In_814);
nor U3099 (N_3099,In_30,In_660);
or U3100 (N_3100,In_926,In_97);
or U3101 (N_3101,In_197,In_26);
or U3102 (N_3102,In_704,In_847);
xnor U3103 (N_3103,In_416,In_166);
xnor U3104 (N_3104,In_691,In_796);
and U3105 (N_3105,In_325,In_507);
nand U3106 (N_3106,In_496,In_910);
nand U3107 (N_3107,In_196,In_768);
and U3108 (N_3108,In_748,In_37);
and U3109 (N_3109,In_939,In_173);
xor U3110 (N_3110,In_955,In_529);
nand U3111 (N_3111,In_153,In_26);
nand U3112 (N_3112,In_811,In_857);
or U3113 (N_3113,In_655,In_154);
and U3114 (N_3114,In_284,In_542);
xnor U3115 (N_3115,In_506,In_631);
or U3116 (N_3116,In_260,In_981);
nor U3117 (N_3117,In_770,In_271);
xor U3118 (N_3118,In_585,In_804);
and U3119 (N_3119,In_122,In_312);
nand U3120 (N_3120,In_818,In_732);
and U3121 (N_3121,In_338,In_309);
nand U3122 (N_3122,In_580,In_462);
nand U3123 (N_3123,In_3,In_693);
nor U3124 (N_3124,In_237,In_608);
nand U3125 (N_3125,In_500,In_580);
and U3126 (N_3126,In_959,In_909);
or U3127 (N_3127,In_523,In_310);
nand U3128 (N_3128,In_228,In_315);
nor U3129 (N_3129,In_341,In_961);
or U3130 (N_3130,In_673,In_702);
nor U3131 (N_3131,In_490,In_599);
nand U3132 (N_3132,In_170,In_671);
or U3133 (N_3133,In_320,In_592);
nor U3134 (N_3134,In_37,In_754);
nor U3135 (N_3135,In_275,In_271);
and U3136 (N_3136,In_868,In_911);
nor U3137 (N_3137,In_203,In_744);
nor U3138 (N_3138,In_561,In_421);
nand U3139 (N_3139,In_357,In_615);
or U3140 (N_3140,In_693,In_137);
xor U3141 (N_3141,In_985,In_857);
and U3142 (N_3142,In_686,In_764);
xnor U3143 (N_3143,In_352,In_991);
and U3144 (N_3144,In_999,In_96);
nand U3145 (N_3145,In_385,In_59);
or U3146 (N_3146,In_839,In_454);
xnor U3147 (N_3147,In_543,In_664);
and U3148 (N_3148,In_795,In_304);
xor U3149 (N_3149,In_135,In_198);
or U3150 (N_3150,In_386,In_515);
nor U3151 (N_3151,In_421,In_776);
or U3152 (N_3152,In_262,In_170);
nand U3153 (N_3153,In_329,In_419);
nor U3154 (N_3154,In_728,In_837);
and U3155 (N_3155,In_513,In_169);
and U3156 (N_3156,In_795,In_547);
nand U3157 (N_3157,In_552,In_77);
xnor U3158 (N_3158,In_425,In_275);
nor U3159 (N_3159,In_510,In_241);
nand U3160 (N_3160,In_681,In_243);
xor U3161 (N_3161,In_137,In_678);
nand U3162 (N_3162,In_345,In_520);
and U3163 (N_3163,In_664,In_624);
nor U3164 (N_3164,In_332,In_501);
and U3165 (N_3165,In_478,In_702);
nand U3166 (N_3166,In_884,In_601);
xnor U3167 (N_3167,In_786,In_297);
nand U3168 (N_3168,In_481,In_456);
nand U3169 (N_3169,In_270,In_818);
and U3170 (N_3170,In_97,In_16);
xor U3171 (N_3171,In_456,In_161);
and U3172 (N_3172,In_244,In_613);
nand U3173 (N_3173,In_12,In_169);
nor U3174 (N_3174,In_121,In_707);
and U3175 (N_3175,In_634,In_709);
nor U3176 (N_3176,In_175,In_956);
and U3177 (N_3177,In_838,In_592);
nand U3178 (N_3178,In_307,In_730);
or U3179 (N_3179,In_23,In_796);
and U3180 (N_3180,In_376,In_172);
xnor U3181 (N_3181,In_322,In_263);
xor U3182 (N_3182,In_608,In_334);
or U3183 (N_3183,In_517,In_492);
and U3184 (N_3184,In_740,In_381);
nand U3185 (N_3185,In_924,In_603);
nor U3186 (N_3186,In_165,In_361);
and U3187 (N_3187,In_312,In_107);
nor U3188 (N_3188,In_176,In_503);
or U3189 (N_3189,In_907,In_535);
and U3190 (N_3190,In_443,In_267);
nor U3191 (N_3191,In_835,In_345);
nor U3192 (N_3192,In_845,In_599);
or U3193 (N_3193,In_975,In_555);
or U3194 (N_3194,In_101,In_924);
nor U3195 (N_3195,In_695,In_260);
nor U3196 (N_3196,In_42,In_540);
nor U3197 (N_3197,In_706,In_844);
nor U3198 (N_3198,In_482,In_161);
nand U3199 (N_3199,In_863,In_353);
nand U3200 (N_3200,In_825,In_201);
and U3201 (N_3201,In_506,In_866);
and U3202 (N_3202,In_944,In_922);
and U3203 (N_3203,In_614,In_722);
or U3204 (N_3204,In_139,In_768);
nand U3205 (N_3205,In_104,In_28);
nand U3206 (N_3206,In_459,In_721);
nand U3207 (N_3207,In_462,In_609);
or U3208 (N_3208,In_664,In_420);
nand U3209 (N_3209,In_600,In_154);
or U3210 (N_3210,In_959,In_457);
or U3211 (N_3211,In_995,In_694);
or U3212 (N_3212,In_986,In_421);
nor U3213 (N_3213,In_10,In_599);
nand U3214 (N_3214,In_635,In_647);
and U3215 (N_3215,In_510,In_533);
and U3216 (N_3216,In_264,In_410);
nor U3217 (N_3217,In_192,In_288);
nand U3218 (N_3218,In_417,In_391);
nor U3219 (N_3219,In_39,In_608);
or U3220 (N_3220,In_527,In_172);
nand U3221 (N_3221,In_93,In_848);
and U3222 (N_3222,In_145,In_253);
and U3223 (N_3223,In_484,In_19);
and U3224 (N_3224,In_41,In_885);
or U3225 (N_3225,In_594,In_192);
nor U3226 (N_3226,In_575,In_588);
nand U3227 (N_3227,In_597,In_396);
nor U3228 (N_3228,In_199,In_546);
xor U3229 (N_3229,In_221,In_849);
nand U3230 (N_3230,In_714,In_256);
nand U3231 (N_3231,In_184,In_373);
nor U3232 (N_3232,In_676,In_941);
or U3233 (N_3233,In_484,In_45);
nor U3234 (N_3234,In_407,In_875);
or U3235 (N_3235,In_898,In_28);
nor U3236 (N_3236,In_630,In_360);
and U3237 (N_3237,In_167,In_795);
and U3238 (N_3238,In_52,In_806);
xnor U3239 (N_3239,In_344,In_713);
nand U3240 (N_3240,In_667,In_507);
nand U3241 (N_3241,In_825,In_417);
or U3242 (N_3242,In_549,In_642);
nor U3243 (N_3243,In_30,In_420);
nand U3244 (N_3244,In_968,In_577);
nor U3245 (N_3245,In_752,In_471);
nor U3246 (N_3246,In_526,In_662);
and U3247 (N_3247,In_481,In_782);
and U3248 (N_3248,In_98,In_527);
and U3249 (N_3249,In_712,In_901);
nand U3250 (N_3250,In_666,In_502);
and U3251 (N_3251,In_312,In_371);
nor U3252 (N_3252,In_119,In_650);
and U3253 (N_3253,In_760,In_539);
nor U3254 (N_3254,In_246,In_654);
or U3255 (N_3255,In_174,In_90);
or U3256 (N_3256,In_368,In_229);
xnor U3257 (N_3257,In_71,In_833);
nor U3258 (N_3258,In_243,In_441);
nand U3259 (N_3259,In_237,In_790);
nor U3260 (N_3260,In_674,In_826);
nor U3261 (N_3261,In_974,In_323);
and U3262 (N_3262,In_367,In_467);
xnor U3263 (N_3263,In_562,In_234);
and U3264 (N_3264,In_841,In_271);
nor U3265 (N_3265,In_58,In_539);
nand U3266 (N_3266,In_823,In_117);
or U3267 (N_3267,In_330,In_977);
or U3268 (N_3268,In_381,In_716);
or U3269 (N_3269,In_468,In_513);
and U3270 (N_3270,In_808,In_874);
nor U3271 (N_3271,In_968,In_702);
nand U3272 (N_3272,In_388,In_330);
nand U3273 (N_3273,In_560,In_553);
or U3274 (N_3274,In_912,In_964);
or U3275 (N_3275,In_604,In_367);
or U3276 (N_3276,In_764,In_974);
nand U3277 (N_3277,In_977,In_573);
and U3278 (N_3278,In_362,In_84);
nand U3279 (N_3279,In_757,In_447);
nor U3280 (N_3280,In_590,In_109);
nand U3281 (N_3281,In_2,In_146);
or U3282 (N_3282,In_950,In_249);
or U3283 (N_3283,In_706,In_777);
or U3284 (N_3284,In_915,In_57);
or U3285 (N_3285,In_822,In_977);
nor U3286 (N_3286,In_96,In_288);
nor U3287 (N_3287,In_810,In_981);
nor U3288 (N_3288,In_222,In_663);
or U3289 (N_3289,In_584,In_2);
nor U3290 (N_3290,In_645,In_920);
and U3291 (N_3291,In_852,In_578);
xor U3292 (N_3292,In_8,In_967);
or U3293 (N_3293,In_225,In_544);
nor U3294 (N_3294,In_706,In_331);
or U3295 (N_3295,In_918,In_675);
nor U3296 (N_3296,In_723,In_384);
nand U3297 (N_3297,In_536,In_881);
nor U3298 (N_3298,In_196,In_470);
nand U3299 (N_3299,In_299,In_307);
or U3300 (N_3300,In_639,In_28);
nor U3301 (N_3301,In_566,In_136);
or U3302 (N_3302,In_689,In_742);
and U3303 (N_3303,In_567,In_603);
nor U3304 (N_3304,In_731,In_454);
nor U3305 (N_3305,In_289,In_467);
or U3306 (N_3306,In_368,In_739);
and U3307 (N_3307,In_691,In_734);
or U3308 (N_3308,In_274,In_975);
or U3309 (N_3309,In_508,In_594);
xor U3310 (N_3310,In_239,In_234);
xor U3311 (N_3311,In_518,In_849);
nor U3312 (N_3312,In_44,In_769);
xor U3313 (N_3313,In_601,In_645);
nand U3314 (N_3314,In_270,In_582);
and U3315 (N_3315,In_610,In_821);
and U3316 (N_3316,In_201,In_943);
or U3317 (N_3317,In_930,In_589);
nand U3318 (N_3318,In_809,In_786);
nand U3319 (N_3319,In_393,In_412);
nand U3320 (N_3320,In_526,In_767);
or U3321 (N_3321,In_423,In_284);
or U3322 (N_3322,In_138,In_44);
or U3323 (N_3323,In_221,In_109);
or U3324 (N_3324,In_167,In_158);
and U3325 (N_3325,In_967,In_795);
and U3326 (N_3326,In_525,In_600);
and U3327 (N_3327,In_666,In_172);
nand U3328 (N_3328,In_465,In_865);
and U3329 (N_3329,In_394,In_356);
or U3330 (N_3330,In_127,In_480);
nand U3331 (N_3331,In_258,In_64);
nand U3332 (N_3332,In_751,In_523);
xor U3333 (N_3333,In_585,In_929);
nor U3334 (N_3334,In_490,In_397);
nand U3335 (N_3335,In_704,In_824);
and U3336 (N_3336,In_723,In_80);
and U3337 (N_3337,In_955,In_624);
or U3338 (N_3338,In_94,In_895);
xor U3339 (N_3339,In_359,In_606);
or U3340 (N_3340,In_227,In_261);
nand U3341 (N_3341,In_352,In_477);
and U3342 (N_3342,In_331,In_212);
nor U3343 (N_3343,In_167,In_218);
and U3344 (N_3344,In_148,In_25);
xnor U3345 (N_3345,In_238,In_871);
or U3346 (N_3346,In_766,In_284);
and U3347 (N_3347,In_973,In_301);
nor U3348 (N_3348,In_51,In_308);
nor U3349 (N_3349,In_651,In_581);
nor U3350 (N_3350,In_73,In_151);
nand U3351 (N_3351,In_118,In_627);
or U3352 (N_3352,In_300,In_156);
nand U3353 (N_3353,In_422,In_309);
or U3354 (N_3354,In_928,In_164);
or U3355 (N_3355,In_897,In_805);
nor U3356 (N_3356,In_275,In_227);
or U3357 (N_3357,In_292,In_34);
nand U3358 (N_3358,In_110,In_143);
and U3359 (N_3359,In_479,In_581);
and U3360 (N_3360,In_546,In_55);
nand U3361 (N_3361,In_445,In_927);
or U3362 (N_3362,In_516,In_507);
nand U3363 (N_3363,In_496,In_755);
and U3364 (N_3364,In_342,In_904);
or U3365 (N_3365,In_764,In_463);
or U3366 (N_3366,In_982,In_635);
and U3367 (N_3367,In_265,In_926);
nor U3368 (N_3368,In_194,In_448);
nor U3369 (N_3369,In_903,In_487);
or U3370 (N_3370,In_243,In_493);
or U3371 (N_3371,In_261,In_869);
nand U3372 (N_3372,In_297,In_375);
or U3373 (N_3373,In_179,In_195);
and U3374 (N_3374,In_540,In_789);
or U3375 (N_3375,In_450,In_81);
nor U3376 (N_3376,In_650,In_643);
xnor U3377 (N_3377,In_778,In_240);
or U3378 (N_3378,In_645,In_893);
or U3379 (N_3379,In_294,In_135);
nor U3380 (N_3380,In_762,In_846);
nand U3381 (N_3381,In_101,In_729);
or U3382 (N_3382,In_588,In_642);
or U3383 (N_3383,In_463,In_708);
nand U3384 (N_3384,In_918,In_233);
nand U3385 (N_3385,In_35,In_800);
nor U3386 (N_3386,In_776,In_964);
nand U3387 (N_3387,In_338,In_449);
and U3388 (N_3388,In_668,In_356);
xnor U3389 (N_3389,In_708,In_761);
nand U3390 (N_3390,In_541,In_510);
nor U3391 (N_3391,In_238,In_287);
nor U3392 (N_3392,In_499,In_919);
nand U3393 (N_3393,In_105,In_898);
nand U3394 (N_3394,In_856,In_18);
xor U3395 (N_3395,In_282,In_16);
and U3396 (N_3396,In_708,In_332);
nand U3397 (N_3397,In_445,In_25);
or U3398 (N_3398,In_755,In_85);
nor U3399 (N_3399,In_232,In_223);
or U3400 (N_3400,In_825,In_569);
nor U3401 (N_3401,In_913,In_321);
and U3402 (N_3402,In_360,In_234);
nand U3403 (N_3403,In_935,In_891);
and U3404 (N_3404,In_853,In_526);
nand U3405 (N_3405,In_265,In_443);
or U3406 (N_3406,In_969,In_228);
nor U3407 (N_3407,In_721,In_816);
nand U3408 (N_3408,In_436,In_867);
or U3409 (N_3409,In_994,In_699);
or U3410 (N_3410,In_966,In_760);
and U3411 (N_3411,In_756,In_284);
or U3412 (N_3412,In_111,In_44);
and U3413 (N_3413,In_182,In_399);
nand U3414 (N_3414,In_115,In_206);
and U3415 (N_3415,In_540,In_507);
nand U3416 (N_3416,In_442,In_502);
nor U3417 (N_3417,In_493,In_580);
nor U3418 (N_3418,In_463,In_885);
or U3419 (N_3419,In_580,In_190);
and U3420 (N_3420,In_968,In_328);
nor U3421 (N_3421,In_888,In_244);
nor U3422 (N_3422,In_993,In_55);
nand U3423 (N_3423,In_890,In_52);
and U3424 (N_3424,In_705,In_737);
and U3425 (N_3425,In_923,In_233);
and U3426 (N_3426,In_517,In_52);
or U3427 (N_3427,In_934,In_994);
or U3428 (N_3428,In_900,In_485);
nand U3429 (N_3429,In_516,In_922);
xnor U3430 (N_3430,In_513,In_619);
or U3431 (N_3431,In_28,In_285);
xnor U3432 (N_3432,In_345,In_565);
nand U3433 (N_3433,In_875,In_559);
xor U3434 (N_3434,In_440,In_773);
or U3435 (N_3435,In_598,In_826);
or U3436 (N_3436,In_884,In_196);
nor U3437 (N_3437,In_911,In_849);
or U3438 (N_3438,In_451,In_908);
or U3439 (N_3439,In_554,In_32);
nand U3440 (N_3440,In_238,In_25);
or U3441 (N_3441,In_798,In_194);
nor U3442 (N_3442,In_586,In_564);
or U3443 (N_3443,In_703,In_584);
and U3444 (N_3444,In_189,In_210);
nor U3445 (N_3445,In_213,In_277);
nand U3446 (N_3446,In_798,In_747);
nand U3447 (N_3447,In_354,In_902);
and U3448 (N_3448,In_931,In_466);
nand U3449 (N_3449,In_198,In_963);
nor U3450 (N_3450,In_557,In_302);
nand U3451 (N_3451,In_99,In_942);
nand U3452 (N_3452,In_169,In_615);
xnor U3453 (N_3453,In_824,In_917);
nand U3454 (N_3454,In_815,In_155);
nor U3455 (N_3455,In_620,In_559);
or U3456 (N_3456,In_73,In_314);
and U3457 (N_3457,In_79,In_426);
or U3458 (N_3458,In_528,In_897);
or U3459 (N_3459,In_903,In_230);
and U3460 (N_3460,In_101,In_208);
or U3461 (N_3461,In_948,In_591);
or U3462 (N_3462,In_69,In_219);
nor U3463 (N_3463,In_305,In_424);
nand U3464 (N_3464,In_97,In_54);
xor U3465 (N_3465,In_728,In_621);
xnor U3466 (N_3466,In_944,In_183);
nor U3467 (N_3467,In_418,In_516);
or U3468 (N_3468,In_12,In_786);
or U3469 (N_3469,In_912,In_416);
or U3470 (N_3470,In_194,In_278);
nor U3471 (N_3471,In_627,In_105);
nor U3472 (N_3472,In_571,In_884);
and U3473 (N_3473,In_779,In_885);
and U3474 (N_3474,In_105,In_895);
nand U3475 (N_3475,In_52,In_357);
nor U3476 (N_3476,In_843,In_140);
xor U3477 (N_3477,In_862,In_11);
and U3478 (N_3478,In_917,In_834);
nor U3479 (N_3479,In_223,In_918);
or U3480 (N_3480,In_380,In_454);
xor U3481 (N_3481,In_273,In_472);
nand U3482 (N_3482,In_388,In_747);
or U3483 (N_3483,In_558,In_286);
or U3484 (N_3484,In_22,In_665);
nor U3485 (N_3485,In_824,In_906);
nand U3486 (N_3486,In_864,In_293);
nor U3487 (N_3487,In_540,In_887);
or U3488 (N_3488,In_809,In_111);
and U3489 (N_3489,In_521,In_448);
and U3490 (N_3490,In_658,In_214);
nand U3491 (N_3491,In_542,In_370);
nor U3492 (N_3492,In_449,In_584);
and U3493 (N_3493,In_12,In_619);
or U3494 (N_3494,In_745,In_961);
nor U3495 (N_3495,In_338,In_747);
and U3496 (N_3496,In_929,In_302);
or U3497 (N_3497,In_275,In_70);
nand U3498 (N_3498,In_555,In_8);
xnor U3499 (N_3499,In_459,In_240);
or U3500 (N_3500,In_937,In_794);
or U3501 (N_3501,In_125,In_167);
nor U3502 (N_3502,In_937,In_878);
and U3503 (N_3503,In_613,In_110);
nor U3504 (N_3504,In_50,In_38);
xor U3505 (N_3505,In_944,In_950);
nand U3506 (N_3506,In_838,In_474);
and U3507 (N_3507,In_47,In_540);
xor U3508 (N_3508,In_964,In_446);
and U3509 (N_3509,In_711,In_143);
nand U3510 (N_3510,In_114,In_255);
and U3511 (N_3511,In_453,In_901);
nor U3512 (N_3512,In_767,In_127);
nor U3513 (N_3513,In_434,In_793);
xnor U3514 (N_3514,In_398,In_213);
nand U3515 (N_3515,In_128,In_195);
and U3516 (N_3516,In_83,In_229);
nor U3517 (N_3517,In_534,In_925);
or U3518 (N_3518,In_461,In_644);
and U3519 (N_3519,In_186,In_758);
and U3520 (N_3520,In_267,In_839);
and U3521 (N_3521,In_709,In_745);
or U3522 (N_3522,In_634,In_782);
nand U3523 (N_3523,In_752,In_157);
or U3524 (N_3524,In_602,In_980);
and U3525 (N_3525,In_736,In_381);
and U3526 (N_3526,In_602,In_735);
nand U3527 (N_3527,In_588,In_923);
nor U3528 (N_3528,In_772,In_432);
and U3529 (N_3529,In_698,In_706);
and U3530 (N_3530,In_286,In_902);
and U3531 (N_3531,In_653,In_672);
nand U3532 (N_3532,In_742,In_3);
nor U3533 (N_3533,In_200,In_655);
and U3534 (N_3534,In_493,In_189);
xor U3535 (N_3535,In_287,In_630);
and U3536 (N_3536,In_74,In_513);
nor U3537 (N_3537,In_873,In_318);
and U3538 (N_3538,In_624,In_34);
nand U3539 (N_3539,In_969,In_394);
nor U3540 (N_3540,In_422,In_458);
xnor U3541 (N_3541,In_454,In_109);
xor U3542 (N_3542,In_791,In_703);
nand U3543 (N_3543,In_865,In_369);
nand U3544 (N_3544,In_595,In_253);
and U3545 (N_3545,In_593,In_928);
and U3546 (N_3546,In_535,In_340);
nor U3547 (N_3547,In_902,In_490);
nand U3548 (N_3548,In_3,In_398);
and U3549 (N_3549,In_778,In_174);
and U3550 (N_3550,In_520,In_771);
and U3551 (N_3551,In_640,In_803);
and U3552 (N_3552,In_176,In_191);
or U3553 (N_3553,In_98,In_634);
xnor U3554 (N_3554,In_609,In_634);
or U3555 (N_3555,In_923,In_292);
or U3556 (N_3556,In_554,In_661);
nor U3557 (N_3557,In_853,In_59);
nor U3558 (N_3558,In_150,In_75);
and U3559 (N_3559,In_654,In_693);
and U3560 (N_3560,In_507,In_851);
or U3561 (N_3561,In_368,In_851);
xnor U3562 (N_3562,In_549,In_383);
xnor U3563 (N_3563,In_280,In_416);
nand U3564 (N_3564,In_798,In_205);
and U3565 (N_3565,In_539,In_701);
or U3566 (N_3566,In_266,In_613);
or U3567 (N_3567,In_139,In_922);
xnor U3568 (N_3568,In_196,In_379);
xor U3569 (N_3569,In_444,In_955);
nor U3570 (N_3570,In_305,In_796);
or U3571 (N_3571,In_829,In_304);
xnor U3572 (N_3572,In_362,In_882);
nor U3573 (N_3573,In_53,In_521);
nand U3574 (N_3574,In_85,In_988);
nand U3575 (N_3575,In_359,In_964);
nand U3576 (N_3576,In_757,In_352);
nand U3577 (N_3577,In_20,In_824);
or U3578 (N_3578,In_533,In_175);
nor U3579 (N_3579,In_516,In_521);
nand U3580 (N_3580,In_57,In_213);
nand U3581 (N_3581,In_641,In_245);
nor U3582 (N_3582,In_578,In_654);
nor U3583 (N_3583,In_525,In_307);
nand U3584 (N_3584,In_163,In_286);
nor U3585 (N_3585,In_810,In_329);
or U3586 (N_3586,In_963,In_815);
nand U3587 (N_3587,In_372,In_518);
xnor U3588 (N_3588,In_801,In_933);
and U3589 (N_3589,In_251,In_475);
and U3590 (N_3590,In_539,In_844);
or U3591 (N_3591,In_863,In_957);
and U3592 (N_3592,In_372,In_316);
nand U3593 (N_3593,In_680,In_636);
or U3594 (N_3594,In_388,In_753);
xor U3595 (N_3595,In_97,In_499);
or U3596 (N_3596,In_679,In_58);
xor U3597 (N_3597,In_569,In_330);
or U3598 (N_3598,In_481,In_319);
nor U3599 (N_3599,In_136,In_199);
xnor U3600 (N_3600,In_467,In_892);
and U3601 (N_3601,In_481,In_61);
or U3602 (N_3602,In_144,In_380);
or U3603 (N_3603,In_192,In_750);
or U3604 (N_3604,In_525,In_634);
nor U3605 (N_3605,In_670,In_755);
or U3606 (N_3606,In_747,In_340);
or U3607 (N_3607,In_303,In_512);
nor U3608 (N_3608,In_737,In_783);
or U3609 (N_3609,In_47,In_318);
or U3610 (N_3610,In_428,In_325);
or U3611 (N_3611,In_22,In_532);
xor U3612 (N_3612,In_505,In_103);
and U3613 (N_3613,In_840,In_89);
nand U3614 (N_3614,In_918,In_863);
and U3615 (N_3615,In_466,In_704);
nor U3616 (N_3616,In_267,In_265);
nand U3617 (N_3617,In_968,In_21);
nor U3618 (N_3618,In_446,In_918);
nand U3619 (N_3619,In_954,In_865);
nand U3620 (N_3620,In_12,In_151);
and U3621 (N_3621,In_837,In_455);
xnor U3622 (N_3622,In_759,In_652);
nor U3623 (N_3623,In_12,In_740);
or U3624 (N_3624,In_592,In_379);
nor U3625 (N_3625,In_161,In_78);
nor U3626 (N_3626,In_308,In_407);
and U3627 (N_3627,In_147,In_439);
nor U3628 (N_3628,In_385,In_15);
and U3629 (N_3629,In_432,In_830);
nor U3630 (N_3630,In_475,In_663);
and U3631 (N_3631,In_644,In_99);
nand U3632 (N_3632,In_915,In_17);
and U3633 (N_3633,In_25,In_821);
or U3634 (N_3634,In_782,In_595);
nor U3635 (N_3635,In_470,In_266);
xor U3636 (N_3636,In_879,In_783);
nor U3637 (N_3637,In_934,In_757);
nor U3638 (N_3638,In_99,In_714);
or U3639 (N_3639,In_937,In_614);
nand U3640 (N_3640,In_203,In_859);
nand U3641 (N_3641,In_683,In_672);
and U3642 (N_3642,In_375,In_991);
and U3643 (N_3643,In_74,In_869);
nor U3644 (N_3644,In_335,In_822);
and U3645 (N_3645,In_20,In_448);
nor U3646 (N_3646,In_448,In_994);
nand U3647 (N_3647,In_365,In_399);
and U3648 (N_3648,In_454,In_801);
and U3649 (N_3649,In_789,In_648);
nand U3650 (N_3650,In_338,In_817);
and U3651 (N_3651,In_760,In_501);
nor U3652 (N_3652,In_852,In_617);
xnor U3653 (N_3653,In_466,In_65);
and U3654 (N_3654,In_301,In_803);
and U3655 (N_3655,In_226,In_659);
or U3656 (N_3656,In_158,In_9);
nand U3657 (N_3657,In_311,In_478);
or U3658 (N_3658,In_0,In_331);
or U3659 (N_3659,In_663,In_211);
or U3660 (N_3660,In_236,In_637);
and U3661 (N_3661,In_584,In_824);
nand U3662 (N_3662,In_283,In_890);
and U3663 (N_3663,In_419,In_288);
and U3664 (N_3664,In_357,In_554);
xor U3665 (N_3665,In_796,In_550);
nor U3666 (N_3666,In_987,In_126);
nand U3667 (N_3667,In_413,In_717);
and U3668 (N_3668,In_658,In_150);
nand U3669 (N_3669,In_367,In_544);
nand U3670 (N_3670,In_996,In_665);
nor U3671 (N_3671,In_722,In_116);
nand U3672 (N_3672,In_421,In_597);
and U3673 (N_3673,In_339,In_584);
or U3674 (N_3674,In_804,In_213);
nor U3675 (N_3675,In_79,In_568);
nor U3676 (N_3676,In_584,In_794);
and U3677 (N_3677,In_889,In_940);
nor U3678 (N_3678,In_304,In_908);
or U3679 (N_3679,In_442,In_946);
nand U3680 (N_3680,In_338,In_623);
nand U3681 (N_3681,In_167,In_407);
and U3682 (N_3682,In_15,In_461);
nand U3683 (N_3683,In_4,In_599);
or U3684 (N_3684,In_430,In_948);
or U3685 (N_3685,In_907,In_693);
and U3686 (N_3686,In_890,In_964);
or U3687 (N_3687,In_275,In_404);
or U3688 (N_3688,In_289,In_202);
xnor U3689 (N_3689,In_858,In_909);
nor U3690 (N_3690,In_210,In_418);
and U3691 (N_3691,In_269,In_265);
nor U3692 (N_3692,In_537,In_490);
nand U3693 (N_3693,In_351,In_394);
xnor U3694 (N_3694,In_457,In_276);
nand U3695 (N_3695,In_847,In_38);
xor U3696 (N_3696,In_39,In_911);
nand U3697 (N_3697,In_129,In_314);
nand U3698 (N_3698,In_985,In_811);
nor U3699 (N_3699,In_188,In_97);
or U3700 (N_3700,In_223,In_18);
nor U3701 (N_3701,In_991,In_744);
or U3702 (N_3702,In_202,In_796);
and U3703 (N_3703,In_359,In_26);
nor U3704 (N_3704,In_228,In_107);
nor U3705 (N_3705,In_5,In_296);
nor U3706 (N_3706,In_826,In_526);
and U3707 (N_3707,In_806,In_552);
nand U3708 (N_3708,In_163,In_288);
xor U3709 (N_3709,In_614,In_914);
xor U3710 (N_3710,In_920,In_132);
nor U3711 (N_3711,In_649,In_715);
and U3712 (N_3712,In_605,In_746);
xor U3713 (N_3713,In_988,In_265);
nor U3714 (N_3714,In_212,In_809);
and U3715 (N_3715,In_752,In_858);
and U3716 (N_3716,In_139,In_153);
and U3717 (N_3717,In_158,In_207);
and U3718 (N_3718,In_227,In_626);
or U3719 (N_3719,In_999,In_551);
nor U3720 (N_3720,In_238,In_665);
xnor U3721 (N_3721,In_223,In_790);
or U3722 (N_3722,In_338,In_248);
xor U3723 (N_3723,In_317,In_291);
or U3724 (N_3724,In_404,In_866);
nand U3725 (N_3725,In_898,In_162);
nor U3726 (N_3726,In_1,In_512);
nor U3727 (N_3727,In_479,In_739);
nor U3728 (N_3728,In_473,In_192);
and U3729 (N_3729,In_145,In_944);
xnor U3730 (N_3730,In_165,In_250);
or U3731 (N_3731,In_667,In_183);
or U3732 (N_3732,In_169,In_713);
xor U3733 (N_3733,In_390,In_836);
nor U3734 (N_3734,In_48,In_140);
and U3735 (N_3735,In_600,In_568);
or U3736 (N_3736,In_324,In_113);
and U3737 (N_3737,In_937,In_858);
and U3738 (N_3738,In_12,In_554);
nor U3739 (N_3739,In_669,In_706);
and U3740 (N_3740,In_640,In_329);
xor U3741 (N_3741,In_789,In_790);
nor U3742 (N_3742,In_178,In_269);
and U3743 (N_3743,In_214,In_605);
or U3744 (N_3744,In_651,In_390);
and U3745 (N_3745,In_862,In_804);
and U3746 (N_3746,In_982,In_198);
nor U3747 (N_3747,In_443,In_326);
xnor U3748 (N_3748,In_16,In_906);
nor U3749 (N_3749,In_885,In_390);
nand U3750 (N_3750,In_539,In_919);
nor U3751 (N_3751,In_548,In_112);
and U3752 (N_3752,In_374,In_610);
and U3753 (N_3753,In_322,In_675);
and U3754 (N_3754,In_855,In_641);
and U3755 (N_3755,In_839,In_735);
or U3756 (N_3756,In_364,In_457);
nand U3757 (N_3757,In_163,In_169);
or U3758 (N_3758,In_158,In_638);
or U3759 (N_3759,In_598,In_376);
and U3760 (N_3760,In_125,In_49);
nand U3761 (N_3761,In_277,In_534);
nor U3762 (N_3762,In_305,In_868);
and U3763 (N_3763,In_513,In_446);
nand U3764 (N_3764,In_243,In_160);
or U3765 (N_3765,In_88,In_550);
and U3766 (N_3766,In_768,In_566);
nand U3767 (N_3767,In_295,In_410);
and U3768 (N_3768,In_757,In_695);
or U3769 (N_3769,In_204,In_868);
nand U3770 (N_3770,In_809,In_651);
nor U3771 (N_3771,In_426,In_941);
or U3772 (N_3772,In_603,In_534);
nor U3773 (N_3773,In_279,In_550);
or U3774 (N_3774,In_668,In_871);
and U3775 (N_3775,In_803,In_575);
nand U3776 (N_3776,In_388,In_678);
and U3777 (N_3777,In_211,In_710);
nand U3778 (N_3778,In_221,In_196);
and U3779 (N_3779,In_987,In_325);
nand U3780 (N_3780,In_609,In_578);
nand U3781 (N_3781,In_356,In_419);
and U3782 (N_3782,In_775,In_109);
and U3783 (N_3783,In_238,In_743);
and U3784 (N_3784,In_268,In_13);
xnor U3785 (N_3785,In_560,In_112);
and U3786 (N_3786,In_355,In_704);
xnor U3787 (N_3787,In_437,In_353);
or U3788 (N_3788,In_350,In_718);
and U3789 (N_3789,In_294,In_328);
nor U3790 (N_3790,In_733,In_604);
or U3791 (N_3791,In_44,In_413);
nor U3792 (N_3792,In_51,In_414);
nor U3793 (N_3793,In_807,In_917);
xnor U3794 (N_3794,In_251,In_480);
and U3795 (N_3795,In_240,In_524);
and U3796 (N_3796,In_771,In_148);
nor U3797 (N_3797,In_543,In_883);
nand U3798 (N_3798,In_92,In_287);
nand U3799 (N_3799,In_757,In_776);
or U3800 (N_3800,In_101,In_267);
and U3801 (N_3801,In_887,In_204);
and U3802 (N_3802,In_761,In_558);
and U3803 (N_3803,In_979,In_907);
nand U3804 (N_3804,In_145,In_140);
and U3805 (N_3805,In_153,In_541);
or U3806 (N_3806,In_648,In_97);
nand U3807 (N_3807,In_468,In_701);
xor U3808 (N_3808,In_195,In_533);
or U3809 (N_3809,In_900,In_213);
and U3810 (N_3810,In_632,In_680);
xor U3811 (N_3811,In_743,In_696);
or U3812 (N_3812,In_272,In_432);
and U3813 (N_3813,In_472,In_102);
xor U3814 (N_3814,In_703,In_76);
or U3815 (N_3815,In_371,In_258);
or U3816 (N_3816,In_807,In_176);
nor U3817 (N_3817,In_879,In_374);
nand U3818 (N_3818,In_891,In_642);
or U3819 (N_3819,In_19,In_423);
or U3820 (N_3820,In_616,In_448);
nor U3821 (N_3821,In_898,In_808);
and U3822 (N_3822,In_815,In_478);
nor U3823 (N_3823,In_175,In_261);
or U3824 (N_3824,In_720,In_842);
or U3825 (N_3825,In_679,In_698);
nor U3826 (N_3826,In_399,In_890);
xor U3827 (N_3827,In_998,In_675);
or U3828 (N_3828,In_699,In_755);
nor U3829 (N_3829,In_464,In_306);
nor U3830 (N_3830,In_519,In_740);
and U3831 (N_3831,In_892,In_590);
and U3832 (N_3832,In_436,In_529);
and U3833 (N_3833,In_212,In_203);
nand U3834 (N_3834,In_53,In_518);
or U3835 (N_3835,In_909,In_459);
or U3836 (N_3836,In_231,In_866);
or U3837 (N_3837,In_731,In_751);
or U3838 (N_3838,In_868,In_103);
xor U3839 (N_3839,In_868,In_783);
nor U3840 (N_3840,In_184,In_299);
nor U3841 (N_3841,In_196,In_349);
nand U3842 (N_3842,In_502,In_775);
or U3843 (N_3843,In_942,In_318);
nand U3844 (N_3844,In_649,In_278);
and U3845 (N_3845,In_387,In_618);
nor U3846 (N_3846,In_987,In_206);
and U3847 (N_3847,In_34,In_968);
or U3848 (N_3848,In_431,In_129);
and U3849 (N_3849,In_83,In_177);
nand U3850 (N_3850,In_446,In_172);
and U3851 (N_3851,In_158,In_621);
and U3852 (N_3852,In_151,In_978);
nand U3853 (N_3853,In_891,In_653);
nor U3854 (N_3854,In_546,In_124);
or U3855 (N_3855,In_186,In_356);
or U3856 (N_3856,In_654,In_550);
nor U3857 (N_3857,In_200,In_932);
nand U3858 (N_3858,In_870,In_349);
nor U3859 (N_3859,In_408,In_342);
and U3860 (N_3860,In_248,In_240);
nand U3861 (N_3861,In_230,In_490);
and U3862 (N_3862,In_276,In_775);
nor U3863 (N_3863,In_320,In_848);
nor U3864 (N_3864,In_840,In_27);
nand U3865 (N_3865,In_444,In_613);
and U3866 (N_3866,In_289,In_779);
nand U3867 (N_3867,In_740,In_432);
nand U3868 (N_3868,In_122,In_185);
nor U3869 (N_3869,In_781,In_794);
and U3870 (N_3870,In_218,In_889);
nor U3871 (N_3871,In_128,In_76);
xor U3872 (N_3872,In_947,In_993);
and U3873 (N_3873,In_461,In_712);
and U3874 (N_3874,In_46,In_397);
xnor U3875 (N_3875,In_728,In_57);
nor U3876 (N_3876,In_170,In_798);
nand U3877 (N_3877,In_533,In_302);
and U3878 (N_3878,In_742,In_442);
and U3879 (N_3879,In_308,In_677);
xor U3880 (N_3880,In_962,In_110);
nand U3881 (N_3881,In_325,In_309);
nor U3882 (N_3882,In_323,In_300);
and U3883 (N_3883,In_68,In_220);
nor U3884 (N_3884,In_941,In_830);
and U3885 (N_3885,In_753,In_548);
nand U3886 (N_3886,In_162,In_980);
nor U3887 (N_3887,In_425,In_291);
nor U3888 (N_3888,In_821,In_753);
nor U3889 (N_3889,In_443,In_441);
nand U3890 (N_3890,In_842,In_762);
and U3891 (N_3891,In_421,In_891);
nor U3892 (N_3892,In_936,In_756);
or U3893 (N_3893,In_393,In_836);
or U3894 (N_3894,In_902,In_457);
nor U3895 (N_3895,In_830,In_499);
nor U3896 (N_3896,In_333,In_136);
or U3897 (N_3897,In_871,In_253);
and U3898 (N_3898,In_94,In_526);
nand U3899 (N_3899,In_195,In_939);
nand U3900 (N_3900,In_971,In_408);
and U3901 (N_3901,In_462,In_890);
xnor U3902 (N_3902,In_830,In_968);
or U3903 (N_3903,In_208,In_91);
xor U3904 (N_3904,In_153,In_724);
and U3905 (N_3905,In_805,In_194);
and U3906 (N_3906,In_803,In_625);
nor U3907 (N_3907,In_47,In_195);
xor U3908 (N_3908,In_659,In_12);
xnor U3909 (N_3909,In_194,In_263);
and U3910 (N_3910,In_212,In_837);
nand U3911 (N_3911,In_539,In_752);
nor U3912 (N_3912,In_819,In_681);
and U3913 (N_3913,In_382,In_750);
nor U3914 (N_3914,In_347,In_802);
or U3915 (N_3915,In_568,In_303);
nor U3916 (N_3916,In_637,In_635);
nand U3917 (N_3917,In_990,In_34);
or U3918 (N_3918,In_501,In_785);
xor U3919 (N_3919,In_894,In_779);
nor U3920 (N_3920,In_936,In_261);
xnor U3921 (N_3921,In_491,In_347);
and U3922 (N_3922,In_921,In_261);
or U3923 (N_3923,In_848,In_177);
and U3924 (N_3924,In_52,In_38);
and U3925 (N_3925,In_478,In_221);
nand U3926 (N_3926,In_322,In_986);
and U3927 (N_3927,In_146,In_321);
nor U3928 (N_3928,In_934,In_393);
or U3929 (N_3929,In_485,In_796);
nand U3930 (N_3930,In_411,In_378);
xor U3931 (N_3931,In_529,In_290);
nand U3932 (N_3932,In_256,In_928);
nand U3933 (N_3933,In_653,In_524);
nand U3934 (N_3934,In_389,In_61);
and U3935 (N_3935,In_763,In_12);
and U3936 (N_3936,In_99,In_93);
or U3937 (N_3937,In_215,In_330);
nand U3938 (N_3938,In_959,In_696);
or U3939 (N_3939,In_376,In_601);
nand U3940 (N_3940,In_179,In_451);
xnor U3941 (N_3941,In_129,In_528);
nand U3942 (N_3942,In_860,In_557);
and U3943 (N_3943,In_915,In_907);
or U3944 (N_3944,In_93,In_851);
nand U3945 (N_3945,In_960,In_189);
and U3946 (N_3946,In_110,In_678);
nand U3947 (N_3947,In_585,In_215);
or U3948 (N_3948,In_878,In_586);
xnor U3949 (N_3949,In_786,In_635);
or U3950 (N_3950,In_35,In_927);
and U3951 (N_3951,In_872,In_418);
or U3952 (N_3952,In_463,In_154);
and U3953 (N_3953,In_221,In_414);
nor U3954 (N_3954,In_138,In_559);
or U3955 (N_3955,In_389,In_518);
nand U3956 (N_3956,In_892,In_93);
or U3957 (N_3957,In_503,In_92);
or U3958 (N_3958,In_842,In_990);
or U3959 (N_3959,In_783,In_657);
and U3960 (N_3960,In_848,In_945);
nor U3961 (N_3961,In_596,In_565);
nand U3962 (N_3962,In_344,In_585);
or U3963 (N_3963,In_850,In_638);
and U3964 (N_3964,In_849,In_812);
xor U3965 (N_3965,In_999,In_404);
and U3966 (N_3966,In_45,In_68);
and U3967 (N_3967,In_905,In_787);
or U3968 (N_3968,In_359,In_295);
nand U3969 (N_3969,In_310,In_6);
nor U3970 (N_3970,In_522,In_625);
or U3971 (N_3971,In_704,In_92);
or U3972 (N_3972,In_203,In_65);
nor U3973 (N_3973,In_395,In_95);
nor U3974 (N_3974,In_674,In_285);
or U3975 (N_3975,In_948,In_737);
nand U3976 (N_3976,In_576,In_778);
and U3977 (N_3977,In_81,In_416);
nor U3978 (N_3978,In_287,In_476);
nor U3979 (N_3979,In_584,In_478);
and U3980 (N_3980,In_973,In_807);
and U3981 (N_3981,In_326,In_647);
and U3982 (N_3982,In_299,In_749);
xnor U3983 (N_3983,In_4,In_949);
nor U3984 (N_3984,In_385,In_23);
nand U3985 (N_3985,In_396,In_112);
and U3986 (N_3986,In_787,In_472);
nand U3987 (N_3987,In_54,In_403);
xor U3988 (N_3988,In_169,In_300);
nor U3989 (N_3989,In_108,In_508);
or U3990 (N_3990,In_337,In_561);
nand U3991 (N_3991,In_359,In_319);
xor U3992 (N_3992,In_425,In_28);
nor U3993 (N_3993,In_846,In_977);
nor U3994 (N_3994,In_76,In_15);
or U3995 (N_3995,In_991,In_520);
and U3996 (N_3996,In_715,In_482);
nand U3997 (N_3997,In_773,In_615);
or U3998 (N_3998,In_514,In_301);
and U3999 (N_3999,In_877,In_369);
xor U4000 (N_4000,In_760,In_607);
or U4001 (N_4001,In_994,In_611);
nand U4002 (N_4002,In_410,In_174);
and U4003 (N_4003,In_949,In_939);
nor U4004 (N_4004,In_524,In_902);
and U4005 (N_4005,In_869,In_358);
or U4006 (N_4006,In_970,In_607);
and U4007 (N_4007,In_150,In_974);
and U4008 (N_4008,In_118,In_134);
xnor U4009 (N_4009,In_980,In_638);
and U4010 (N_4010,In_967,In_821);
nor U4011 (N_4011,In_115,In_471);
nor U4012 (N_4012,In_207,In_290);
nor U4013 (N_4013,In_55,In_219);
and U4014 (N_4014,In_865,In_397);
nor U4015 (N_4015,In_463,In_733);
xnor U4016 (N_4016,In_120,In_361);
or U4017 (N_4017,In_90,In_572);
or U4018 (N_4018,In_88,In_571);
and U4019 (N_4019,In_922,In_880);
nand U4020 (N_4020,In_520,In_875);
and U4021 (N_4021,In_287,In_425);
xor U4022 (N_4022,In_504,In_603);
nand U4023 (N_4023,In_978,In_656);
xnor U4024 (N_4024,In_202,In_276);
and U4025 (N_4025,In_704,In_904);
or U4026 (N_4026,In_141,In_473);
nand U4027 (N_4027,In_657,In_337);
or U4028 (N_4028,In_555,In_803);
nand U4029 (N_4029,In_244,In_193);
nand U4030 (N_4030,In_703,In_795);
nand U4031 (N_4031,In_967,In_749);
xor U4032 (N_4032,In_283,In_586);
xor U4033 (N_4033,In_404,In_806);
or U4034 (N_4034,In_369,In_44);
nor U4035 (N_4035,In_731,In_55);
nand U4036 (N_4036,In_972,In_306);
and U4037 (N_4037,In_419,In_388);
nand U4038 (N_4038,In_896,In_507);
nand U4039 (N_4039,In_62,In_768);
nand U4040 (N_4040,In_667,In_781);
or U4041 (N_4041,In_112,In_518);
nand U4042 (N_4042,In_204,In_713);
and U4043 (N_4043,In_502,In_645);
xnor U4044 (N_4044,In_461,In_243);
nor U4045 (N_4045,In_514,In_962);
nand U4046 (N_4046,In_886,In_996);
xnor U4047 (N_4047,In_55,In_880);
nor U4048 (N_4048,In_700,In_7);
nor U4049 (N_4049,In_80,In_680);
and U4050 (N_4050,In_879,In_973);
nand U4051 (N_4051,In_821,In_600);
nor U4052 (N_4052,In_790,In_741);
nand U4053 (N_4053,In_683,In_496);
and U4054 (N_4054,In_726,In_939);
and U4055 (N_4055,In_364,In_999);
or U4056 (N_4056,In_768,In_789);
nor U4057 (N_4057,In_462,In_810);
or U4058 (N_4058,In_289,In_968);
nand U4059 (N_4059,In_255,In_172);
and U4060 (N_4060,In_605,In_288);
xor U4061 (N_4061,In_488,In_424);
and U4062 (N_4062,In_744,In_626);
or U4063 (N_4063,In_110,In_345);
or U4064 (N_4064,In_609,In_988);
or U4065 (N_4065,In_477,In_873);
or U4066 (N_4066,In_293,In_335);
and U4067 (N_4067,In_553,In_695);
or U4068 (N_4068,In_699,In_383);
or U4069 (N_4069,In_652,In_926);
nor U4070 (N_4070,In_354,In_81);
and U4071 (N_4071,In_702,In_739);
or U4072 (N_4072,In_512,In_206);
or U4073 (N_4073,In_448,In_139);
nor U4074 (N_4074,In_823,In_137);
nand U4075 (N_4075,In_773,In_144);
and U4076 (N_4076,In_800,In_201);
nand U4077 (N_4077,In_176,In_121);
and U4078 (N_4078,In_907,In_186);
nand U4079 (N_4079,In_434,In_5);
nand U4080 (N_4080,In_191,In_373);
xor U4081 (N_4081,In_64,In_89);
xnor U4082 (N_4082,In_455,In_727);
and U4083 (N_4083,In_908,In_24);
nor U4084 (N_4084,In_392,In_691);
or U4085 (N_4085,In_287,In_32);
nand U4086 (N_4086,In_120,In_716);
or U4087 (N_4087,In_101,In_768);
nor U4088 (N_4088,In_816,In_920);
or U4089 (N_4089,In_69,In_833);
nand U4090 (N_4090,In_617,In_165);
nand U4091 (N_4091,In_547,In_529);
nor U4092 (N_4092,In_575,In_60);
and U4093 (N_4093,In_886,In_136);
nand U4094 (N_4094,In_984,In_405);
nor U4095 (N_4095,In_245,In_144);
or U4096 (N_4096,In_694,In_199);
nor U4097 (N_4097,In_662,In_612);
nor U4098 (N_4098,In_541,In_930);
nand U4099 (N_4099,In_137,In_27);
and U4100 (N_4100,In_291,In_372);
nor U4101 (N_4101,In_479,In_36);
and U4102 (N_4102,In_223,In_970);
and U4103 (N_4103,In_393,In_587);
nand U4104 (N_4104,In_131,In_887);
or U4105 (N_4105,In_172,In_808);
and U4106 (N_4106,In_287,In_121);
or U4107 (N_4107,In_388,In_737);
or U4108 (N_4108,In_365,In_384);
xnor U4109 (N_4109,In_785,In_821);
nor U4110 (N_4110,In_497,In_913);
xor U4111 (N_4111,In_370,In_857);
or U4112 (N_4112,In_977,In_253);
nor U4113 (N_4113,In_614,In_328);
or U4114 (N_4114,In_896,In_325);
nor U4115 (N_4115,In_375,In_742);
nor U4116 (N_4116,In_853,In_603);
xnor U4117 (N_4117,In_592,In_164);
or U4118 (N_4118,In_984,In_950);
nor U4119 (N_4119,In_172,In_659);
xor U4120 (N_4120,In_17,In_196);
or U4121 (N_4121,In_753,In_338);
nand U4122 (N_4122,In_872,In_219);
or U4123 (N_4123,In_101,In_506);
or U4124 (N_4124,In_665,In_982);
nor U4125 (N_4125,In_4,In_9);
or U4126 (N_4126,In_519,In_390);
or U4127 (N_4127,In_291,In_174);
nor U4128 (N_4128,In_354,In_824);
or U4129 (N_4129,In_188,In_442);
nand U4130 (N_4130,In_984,In_339);
or U4131 (N_4131,In_739,In_534);
nand U4132 (N_4132,In_258,In_939);
or U4133 (N_4133,In_883,In_214);
or U4134 (N_4134,In_149,In_681);
or U4135 (N_4135,In_379,In_384);
and U4136 (N_4136,In_262,In_353);
xnor U4137 (N_4137,In_15,In_768);
and U4138 (N_4138,In_997,In_378);
xnor U4139 (N_4139,In_626,In_886);
or U4140 (N_4140,In_643,In_946);
and U4141 (N_4141,In_957,In_26);
nor U4142 (N_4142,In_526,In_24);
nor U4143 (N_4143,In_311,In_934);
nor U4144 (N_4144,In_669,In_191);
or U4145 (N_4145,In_728,In_453);
and U4146 (N_4146,In_764,In_352);
nor U4147 (N_4147,In_33,In_328);
and U4148 (N_4148,In_33,In_566);
xor U4149 (N_4149,In_944,In_349);
or U4150 (N_4150,In_522,In_367);
and U4151 (N_4151,In_730,In_872);
nor U4152 (N_4152,In_119,In_127);
xnor U4153 (N_4153,In_317,In_183);
and U4154 (N_4154,In_921,In_372);
nor U4155 (N_4155,In_816,In_39);
nor U4156 (N_4156,In_804,In_123);
nand U4157 (N_4157,In_806,In_250);
and U4158 (N_4158,In_725,In_839);
nor U4159 (N_4159,In_310,In_424);
nor U4160 (N_4160,In_288,In_216);
nor U4161 (N_4161,In_930,In_721);
nand U4162 (N_4162,In_925,In_181);
or U4163 (N_4163,In_884,In_640);
nand U4164 (N_4164,In_123,In_199);
and U4165 (N_4165,In_687,In_511);
nor U4166 (N_4166,In_638,In_712);
nor U4167 (N_4167,In_225,In_189);
and U4168 (N_4168,In_411,In_629);
and U4169 (N_4169,In_430,In_422);
nor U4170 (N_4170,In_36,In_492);
nand U4171 (N_4171,In_452,In_496);
or U4172 (N_4172,In_39,In_966);
and U4173 (N_4173,In_997,In_394);
and U4174 (N_4174,In_960,In_398);
or U4175 (N_4175,In_151,In_166);
or U4176 (N_4176,In_939,In_643);
nand U4177 (N_4177,In_987,In_875);
nor U4178 (N_4178,In_929,In_51);
nand U4179 (N_4179,In_506,In_349);
nor U4180 (N_4180,In_337,In_27);
nor U4181 (N_4181,In_684,In_121);
and U4182 (N_4182,In_966,In_299);
xor U4183 (N_4183,In_270,In_525);
nor U4184 (N_4184,In_386,In_788);
nor U4185 (N_4185,In_233,In_670);
nor U4186 (N_4186,In_693,In_156);
nor U4187 (N_4187,In_568,In_856);
nor U4188 (N_4188,In_468,In_659);
xor U4189 (N_4189,In_297,In_473);
xor U4190 (N_4190,In_92,In_141);
nor U4191 (N_4191,In_433,In_577);
and U4192 (N_4192,In_308,In_8);
and U4193 (N_4193,In_921,In_884);
and U4194 (N_4194,In_656,In_897);
nand U4195 (N_4195,In_193,In_759);
or U4196 (N_4196,In_139,In_776);
or U4197 (N_4197,In_63,In_698);
and U4198 (N_4198,In_568,In_689);
or U4199 (N_4199,In_517,In_153);
nand U4200 (N_4200,In_214,In_0);
and U4201 (N_4201,In_66,In_578);
nor U4202 (N_4202,In_98,In_312);
nor U4203 (N_4203,In_886,In_489);
nor U4204 (N_4204,In_776,In_200);
and U4205 (N_4205,In_160,In_251);
and U4206 (N_4206,In_942,In_622);
or U4207 (N_4207,In_179,In_607);
nor U4208 (N_4208,In_198,In_654);
or U4209 (N_4209,In_145,In_758);
or U4210 (N_4210,In_267,In_906);
nand U4211 (N_4211,In_820,In_626);
nor U4212 (N_4212,In_971,In_993);
and U4213 (N_4213,In_511,In_164);
and U4214 (N_4214,In_925,In_788);
nor U4215 (N_4215,In_553,In_923);
nor U4216 (N_4216,In_304,In_645);
nor U4217 (N_4217,In_469,In_837);
and U4218 (N_4218,In_894,In_303);
xor U4219 (N_4219,In_902,In_362);
xor U4220 (N_4220,In_743,In_836);
or U4221 (N_4221,In_212,In_433);
nand U4222 (N_4222,In_357,In_515);
nor U4223 (N_4223,In_607,In_42);
nor U4224 (N_4224,In_765,In_352);
nand U4225 (N_4225,In_21,In_652);
nor U4226 (N_4226,In_345,In_9);
or U4227 (N_4227,In_867,In_87);
nand U4228 (N_4228,In_915,In_433);
nand U4229 (N_4229,In_653,In_270);
and U4230 (N_4230,In_58,In_399);
xnor U4231 (N_4231,In_316,In_177);
xor U4232 (N_4232,In_384,In_716);
and U4233 (N_4233,In_537,In_326);
or U4234 (N_4234,In_291,In_226);
nand U4235 (N_4235,In_240,In_967);
xor U4236 (N_4236,In_162,In_931);
and U4237 (N_4237,In_2,In_16);
nand U4238 (N_4238,In_669,In_815);
nand U4239 (N_4239,In_715,In_91);
or U4240 (N_4240,In_914,In_213);
nand U4241 (N_4241,In_881,In_604);
nand U4242 (N_4242,In_634,In_767);
and U4243 (N_4243,In_454,In_658);
nand U4244 (N_4244,In_296,In_470);
nor U4245 (N_4245,In_489,In_913);
nor U4246 (N_4246,In_412,In_299);
nor U4247 (N_4247,In_349,In_215);
and U4248 (N_4248,In_557,In_988);
nor U4249 (N_4249,In_268,In_471);
and U4250 (N_4250,In_706,In_276);
and U4251 (N_4251,In_111,In_916);
and U4252 (N_4252,In_687,In_578);
and U4253 (N_4253,In_594,In_758);
or U4254 (N_4254,In_467,In_695);
nand U4255 (N_4255,In_969,In_278);
nand U4256 (N_4256,In_724,In_576);
nand U4257 (N_4257,In_71,In_943);
or U4258 (N_4258,In_41,In_525);
and U4259 (N_4259,In_664,In_807);
nor U4260 (N_4260,In_113,In_410);
or U4261 (N_4261,In_500,In_4);
nor U4262 (N_4262,In_468,In_52);
or U4263 (N_4263,In_963,In_268);
nand U4264 (N_4264,In_581,In_352);
xnor U4265 (N_4265,In_153,In_708);
nor U4266 (N_4266,In_310,In_340);
or U4267 (N_4267,In_656,In_667);
nand U4268 (N_4268,In_147,In_828);
or U4269 (N_4269,In_377,In_962);
nand U4270 (N_4270,In_129,In_575);
nand U4271 (N_4271,In_445,In_178);
nand U4272 (N_4272,In_589,In_180);
or U4273 (N_4273,In_15,In_270);
and U4274 (N_4274,In_500,In_822);
xor U4275 (N_4275,In_631,In_292);
xnor U4276 (N_4276,In_181,In_824);
or U4277 (N_4277,In_371,In_246);
and U4278 (N_4278,In_909,In_308);
or U4279 (N_4279,In_122,In_234);
nand U4280 (N_4280,In_795,In_381);
or U4281 (N_4281,In_239,In_460);
or U4282 (N_4282,In_225,In_847);
and U4283 (N_4283,In_613,In_905);
nand U4284 (N_4284,In_486,In_680);
and U4285 (N_4285,In_980,In_630);
nand U4286 (N_4286,In_44,In_381);
and U4287 (N_4287,In_229,In_315);
or U4288 (N_4288,In_236,In_490);
nor U4289 (N_4289,In_354,In_850);
xor U4290 (N_4290,In_628,In_163);
or U4291 (N_4291,In_980,In_18);
xor U4292 (N_4292,In_107,In_587);
nor U4293 (N_4293,In_294,In_276);
and U4294 (N_4294,In_780,In_890);
nand U4295 (N_4295,In_204,In_302);
or U4296 (N_4296,In_786,In_95);
xnor U4297 (N_4297,In_634,In_287);
and U4298 (N_4298,In_681,In_922);
xnor U4299 (N_4299,In_110,In_278);
nor U4300 (N_4300,In_578,In_49);
nand U4301 (N_4301,In_184,In_360);
and U4302 (N_4302,In_216,In_743);
or U4303 (N_4303,In_919,In_575);
and U4304 (N_4304,In_327,In_3);
nand U4305 (N_4305,In_506,In_833);
or U4306 (N_4306,In_157,In_414);
nor U4307 (N_4307,In_999,In_315);
nor U4308 (N_4308,In_895,In_118);
nor U4309 (N_4309,In_141,In_346);
nor U4310 (N_4310,In_68,In_432);
or U4311 (N_4311,In_57,In_393);
nand U4312 (N_4312,In_826,In_166);
or U4313 (N_4313,In_321,In_698);
and U4314 (N_4314,In_701,In_895);
and U4315 (N_4315,In_986,In_430);
nor U4316 (N_4316,In_501,In_853);
or U4317 (N_4317,In_658,In_564);
and U4318 (N_4318,In_609,In_231);
nor U4319 (N_4319,In_894,In_685);
nand U4320 (N_4320,In_994,In_145);
nor U4321 (N_4321,In_553,In_745);
or U4322 (N_4322,In_637,In_287);
and U4323 (N_4323,In_394,In_117);
nor U4324 (N_4324,In_350,In_215);
or U4325 (N_4325,In_656,In_234);
or U4326 (N_4326,In_819,In_658);
nor U4327 (N_4327,In_234,In_430);
and U4328 (N_4328,In_110,In_558);
or U4329 (N_4329,In_38,In_374);
nand U4330 (N_4330,In_866,In_931);
nor U4331 (N_4331,In_747,In_197);
or U4332 (N_4332,In_603,In_199);
nand U4333 (N_4333,In_637,In_102);
nor U4334 (N_4334,In_925,In_765);
nor U4335 (N_4335,In_232,In_748);
xnor U4336 (N_4336,In_551,In_138);
and U4337 (N_4337,In_457,In_702);
and U4338 (N_4338,In_969,In_932);
nor U4339 (N_4339,In_703,In_56);
or U4340 (N_4340,In_740,In_698);
nor U4341 (N_4341,In_869,In_439);
or U4342 (N_4342,In_3,In_773);
nor U4343 (N_4343,In_482,In_67);
nor U4344 (N_4344,In_526,In_665);
nor U4345 (N_4345,In_991,In_457);
or U4346 (N_4346,In_145,In_225);
or U4347 (N_4347,In_333,In_575);
nand U4348 (N_4348,In_370,In_906);
nand U4349 (N_4349,In_752,In_19);
xor U4350 (N_4350,In_839,In_629);
or U4351 (N_4351,In_47,In_172);
nor U4352 (N_4352,In_306,In_327);
and U4353 (N_4353,In_586,In_570);
nand U4354 (N_4354,In_620,In_931);
and U4355 (N_4355,In_460,In_889);
nand U4356 (N_4356,In_495,In_728);
nand U4357 (N_4357,In_465,In_742);
or U4358 (N_4358,In_314,In_882);
xor U4359 (N_4359,In_860,In_358);
nor U4360 (N_4360,In_75,In_383);
xnor U4361 (N_4361,In_631,In_891);
or U4362 (N_4362,In_332,In_93);
nor U4363 (N_4363,In_63,In_746);
nand U4364 (N_4364,In_390,In_526);
and U4365 (N_4365,In_188,In_529);
nand U4366 (N_4366,In_253,In_188);
or U4367 (N_4367,In_873,In_21);
or U4368 (N_4368,In_509,In_497);
or U4369 (N_4369,In_706,In_505);
nand U4370 (N_4370,In_48,In_274);
xnor U4371 (N_4371,In_858,In_597);
or U4372 (N_4372,In_94,In_311);
or U4373 (N_4373,In_633,In_752);
or U4374 (N_4374,In_442,In_559);
nor U4375 (N_4375,In_632,In_727);
nor U4376 (N_4376,In_535,In_681);
nand U4377 (N_4377,In_834,In_67);
and U4378 (N_4378,In_575,In_473);
nor U4379 (N_4379,In_851,In_696);
nor U4380 (N_4380,In_536,In_85);
and U4381 (N_4381,In_186,In_440);
nand U4382 (N_4382,In_391,In_721);
nand U4383 (N_4383,In_257,In_771);
or U4384 (N_4384,In_261,In_3);
nand U4385 (N_4385,In_791,In_519);
or U4386 (N_4386,In_493,In_785);
nand U4387 (N_4387,In_512,In_471);
nor U4388 (N_4388,In_54,In_587);
nor U4389 (N_4389,In_792,In_677);
and U4390 (N_4390,In_649,In_129);
and U4391 (N_4391,In_735,In_971);
nand U4392 (N_4392,In_207,In_186);
nand U4393 (N_4393,In_158,In_38);
nor U4394 (N_4394,In_470,In_764);
nor U4395 (N_4395,In_728,In_664);
nor U4396 (N_4396,In_369,In_22);
or U4397 (N_4397,In_257,In_368);
or U4398 (N_4398,In_853,In_316);
or U4399 (N_4399,In_668,In_245);
and U4400 (N_4400,In_390,In_213);
or U4401 (N_4401,In_474,In_660);
nand U4402 (N_4402,In_328,In_966);
or U4403 (N_4403,In_395,In_219);
or U4404 (N_4404,In_751,In_365);
or U4405 (N_4405,In_231,In_52);
nand U4406 (N_4406,In_334,In_873);
nand U4407 (N_4407,In_862,In_174);
nor U4408 (N_4408,In_412,In_839);
or U4409 (N_4409,In_251,In_261);
or U4410 (N_4410,In_951,In_945);
and U4411 (N_4411,In_528,In_504);
nor U4412 (N_4412,In_897,In_654);
nand U4413 (N_4413,In_494,In_393);
and U4414 (N_4414,In_619,In_122);
xor U4415 (N_4415,In_583,In_468);
xnor U4416 (N_4416,In_417,In_597);
nand U4417 (N_4417,In_573,In_492);
and U4418 (N_4418,In_754,In_537);
nand U4419 (N_4419,In_921,In_63);
or U4420 (N_4420,In_580,In_674);
or U4421 (N_4421,In_228,In_550);
nand U4422 (N_4422,In_459,In_552);
nand U4423 (N_4423,In_65,In_512);
or U4424 (N_4424,In_731,In_392);
and U4425 (N_4425,In_5,In_918);
nand U4426 (N_4426,In_740,In_24);
and U4427 (N_4427,In_44,In_135);
nor U4428 (N_4428,In_316,In_628);
or U4429 (N_4429,In_161,In_751);
nand U4430 (N_4430,In_266,In_840);
nor U4431 (N_4431,In_362,In_4);
or U4432 (N_4432,In_424,In_667);
nand U4433 (N_4433,In_707,In_287);
or U4434 (N_4434,In_225,In_419);
nand U4435 (N_4435,In_981,In_152);
nor U4436 (N_4436,In_463,In_76);
or U4437 (N_4437,In_882,In_410);
or U4438 (N_4438,In_458,In_403);
nor U4439 (N_4439,In_411,In_873);
or U4440 (N_4440,In_80,In_434);
xnor U4441 (N_4441,In_878,In_331);
or U4442 (N_4442,In_70,In_783);
nand U4443 (N_4443,In_750,In_647);
and U4444 (N_4444,In_738,In_989);
nand U4445 (N_4445,In_5,In_488);
xnor U4446 (N_4446,In_610,In_786);
and U4447 (N_4447,In_985,In_365);
or U4448 (N_4448,In_545,In_29);
or U4449 (N_4449,In_76,In_834);
or U4450 (N_4450,In_726,In_68);
or U4451 (N_4451,In_197,In_970);
or U4452 (N_4452,In_25,In_5);
and U4453 (N_4453,In_211,In_245);
nand U4454 (N_4454,In_886,In_469);
and U4455 (N_4455,In_173,In_184);
nor U4456 (N_4456,In_946,In_720);
nand U4457 (N_4457,In_559,In_406);
and U4458 (N_4458,In_733,In_514);
or U4459 (N_4459,In_430,In_31);
nand U4460 (N_4460,In_402,In_535);
nand U4461 (N_4461,In_655,In_359);
and U4462 (N_4462,In_779,In_313);
nand U4463 (N_4463,In_928,In_234);
xor U4464 (N_4464,In_298,In_164);
or U4465 (N_4465,In_256,In_394);
or U4466 (N_4466,In_556,In_136);
or U4467 (N_4467,In_319,In_376);
or U4468 (N_4468,In_278,In_216);
or U4469 (N_4469,In_726,In_985);
or U4470 (N_4470,In_905,In_809);
nor U4471 (N_4471,In_941,In_258);
nand U4472 (N_4472,In_198,In_430);
or U4473 (N_4473,In_942,In_790);
nand U4474 (N_4474,In_985,In_463);
and U4475 (N_4475,In_609,In_281);
nor U4476 (N_4476,In_213,In_841);
nand U4477 (N_4477,In_626,In_62);
nor U4478 (N_4478,In_332,In_908);
and U4479 (N_4479,In_571,In_671);
or U4480 (N_4480,In_425,In_430);
or U4481 (N_4481,In_169,In_29);
and U4482 (N_4482,In_264,In_153);
or U4483 (N_4483,In_564,In_844);
and U4484 (N_4484,In_501,In_605);
or U4485 (N_4485,In_835,In_962);
nor U4486 (N_4486,In_295,In_550);
xnor U4487 (N_4487,In_839,In_21);
or U4488 (N_4488,In_346,In_675);
or U4489 (N_4489,In_560,In_792);
xnor U4490 (N_4490,In_81,In_551);
xnor U4491 (N_4491,In_93,In_947);
and U4492 (N_4492,In_115,In_636);
nor U4493 (N_4493,In_106,In_581);
nand U4494 (N_4494,In_392,In_378);
xor U4495 (N_4495,In_596,In_959);
nor U4496 (N_4496,In_10,In_262);
nand U4497 (N_4497,In_38,In_810);
nand U4498 (N_4498,In_368,In_342);
or U4499 (N_4499,In_86,In_353);
xnor U4500 (N_4500,In_505,In_834);
and U4501 (N_4501,In_116,In_765);
or U4502 (N_4502,In_206,In_334);
or U4503 (N_4503,In_10,In_173);
nand U4504 (N_4504,In_832,In_525);
nand U4505 (N_4505,In_4,In_535);
or U4506 (N_4506,In_400,In_305);
nand U4507 (N_4507,In_377,In_932);
or U4508 (N_4508,In_428,In_953);
or U4509 (N_4509,In_232,In_506);
and U4510 (N_4510,In_628,In_673);
xor U4511 (N_4511,In_343,In_165);
nor U4512 (N_4512,In_373,In_893);
nor U4513 (N_4513,In_566,In_168);
nand U4514 (N_4514,In_114,In_846);
nand U4515 (N_4515,In_201,In_649);
nor U4516 (N_4516,In_827,In_302);
and U4517 (N_4517,In_647,In_340);
nor U4518 (N_4518,In_986,In_340);
or U4519 (N_4519,In_22,In_682);
or U4520 (N_4520,In_278,In_484);
nand U4521 (N_4521,In_68,In_299);
xnor U4522 (N_4522,In_165,In_27);
or U4523 (N_4523,In_159,In_296);
or U4524 (N_4524,In_969,In_83);
nand U4525 (N_4525,In_498,In_979);
and U4526 (N_4526,In_952,In_366);
and U4527 (N_4527,In_729,In_316);
and U4528 (N_4528,In_377,In_867);
nand U4529 (N_4529,In_134,In_561);
nor U4530 (N_4530,In_147,In_275);
and U4531 (N_4531,In_981,In_439);
or U4532 (N_4532,In_834,In_14);
nand U4533 (N_4533,In_325,In_414);
nor U4534 (N_4534,In_674,In_388);
nand U4535 (N_4535,In_334,In_205);
and U4536 (N_4536,In_92,In_37);
xor U4537 (N_4537,In_358,In_338);
nor U4538 (N_4538,In_148,In_956);
and U4539 (N_4539,In_556,In_441);
xnor U4540 (N_4540,In_161,In_185);
nor U4541 (N_4541,In_728,In_226);
nand U4542 (N_4542,In_970,In_388);
or U4543 (N_4543,In_768,In_593);
xor U4544 (N_4544,In_232,In_215);
and U4545 (N_4545,In_284,In_637);
xnor U4546 (N_4546,In_629,In_666);
xor U4547 (N_4547,In_656,In_868);
and U4548 (N_4548,In_784,In_276);
or U4549 (N_4549,In_358,In_14);
nand U4550 (N_4550,In_440,In_751);
nand U4551 (N_4551,In_298,In_182);
or U4552 (N_4552,In_533,In_464);
and U4553 (N_4553,In_850,In_996);
and U4554 (N_4554,In_929,In_400);
or U4555 (N_4555,In_842,In_277);
and U4556 (N_4556,In_590,In_756);
or U4557 (N_4557,In_283,In_544);
and U4558 (N_4558,In_360,In_214);
and U4559 (N_4559,In_185,In_229);
and U4560 (N_4560,In_98,In_685);
or U4561 (N_4561,In_23,In_249);
nand U4562 (N_4562,In_380,In_313);
nand U4563 (N_4563,In_232,In_693);
or U4564 (N_4564,In_577,In_493);
and U4565 (N_4565,In_234,In_199);
nand U4566 (N_4566,In_898,In_468);
and U4567 (N_4567,In_912,In_378);
nor U4568 (N_4568,In_593,In_297);
nor U4569 (N_4569,In_505,In_423);
and U4570 (N_4570,In_260,In_230);
nand U4571 (N_4571,In_621,In_312);
nand U4572 (N_4572,In_395,In_893);
nor U4573 (N_4573,In_946,In_588);
or U4574 (N_4574,In_554,In_975);
or U4575 (N_4575,In_610,In_23);
nor U4576 (N_4576,In_195,In_87);
or U4577 (N_4577,In_53,In_665);
and U4578 (N_4578,In_621,In_601);
xor U4579 (N_4579,In_814,In_941);
nor U4580 (N_4580,In_659,In_126);
nand U4581 (N_4581,In_895,In_877);
nor U4582 (N_4582,In_512,In_660);
or U4583 (N_4583,In_647,In_119);
or U4584 (N_4584,In_618,In_152);
or U4585 (N_4585,In_972,In_773);
or U4586 (N_4586,In_93,In_751);
nand U4587 (N_4587,In_993,In_6);
and U4588 (N_4588,In_83,In_316);
or U4589 (N_4589,In_77,In_891);
xor U4590 (N_4590,In_330,In_684);
nor U4591 (N_4591,In_783,In_746);
or U4592 (N_4592,In_310,In_413);
nor U4593 (N_4593,In_847,In_878);
and U4594 (N_4594,In_924,In_306);
nand U4595 (N_4595,In_735,In_779);
xnor U4596 (N_4596,In_673,In_384);
and U4597 (N_4597,In_840,In_403);
nand U4598 (N_4598,In_466,In_899);
nor U4599 (N_4599,In_928,In_30);
or U4600 (N_4600,In_320,In_648);
or U4601 (N_4601,In_491,In_777);
and U4602 (N_4602,In_63,In_918);
nand U4603 (N_4603,In_496,In_622);
nand U4604 (N_4604,In_160,In_466);
nand U4605 (N_4605,In_139,In_706);
or U4606 (N_4606,In_41,In_989);
or U4607 (N_4607,In_401,In_961);
nor U4608 (N_4608,In_129,In_935);
nor U4609 (N_4609,In_683,In_303);
nor U4610 (N_4610,In_849,In_178);
nand U4611 (N_4611,In_274,In_794);
xor U4612 (N_4612,In_583,In_47);
and U4613 (N_4613,In_882,In_250);
nor U4614 (N_4614,In_419,In_194);
and U4615 (N_4615,In_29,In_618);
nor U4616 (N_4616,In_223,In_599);
nand U4617 (N_4617,In_531,In_188);
nor U4618 (N_4618,In_996,In_706);
and U4619 (N_4619,In_782,In_895);
or U4620 (N_4620,In_198,In_138);
nand U4621 (N_4621,In_174,In_114);
nor U4622 (N_4622,In_791,In_65);
or U4623 (N_4623,In_904,In_710);
nand U4624 (N_4624,In_627,In_731);
xnor U4625 (N_4625,In_785,In_114);
or U4626 (N_4626,In_661,In_302);
xor U4627 (N_4627,In_277,In_89);
and U4628 (N_4628,In_366,In_626);
xnor U4629 (N_4629,In_692,In_141);
or U4630 (N_4630,In_975,In_717);
nand U4631 (N_4631,In_795,In_458);
or U4632 (N_4632,In_207,In_509);
nand U4633 (N_4633,In_473,In_391);
xor U4634 (N_4634,In_261,In_404);
xor U4635 (N_4635,In_956,In_294);
xor U4636 (N_4636,In_531,In_979);
and U4637 (N_4637,In_372,In_200);
nand U4638 (N_4638,In_632,In_379);
nor U4639 (N_4639,In_531,In_954);
nand U4640 (N_4640,In_76,In_875);
and U4641 (N_4641,In_949,In_699);
and U4642 (N_4642,In_883,In_950);
nor U4643 (N_4643,In_388,In_182);
nand U4644 (N_4644,In_40,In_481);
or U4645 (N_4645,In_245,In_935);
nor U4646 (N_4646,In_224,In_757);
and U4647 (N_4647,In_830,In_902);
xor U4648 (N_4648,In_809,In_632);
xor U4649 (N_4649,In_952,In_49);
and U4650 (N_4650,In_589,In_983);
or U4651 (N_4651,In_673,In_590);
nor U4652 (N_4652,In_422,In_661);
nor U4653 (N_4653,In_443,In_407);
or U4654 (N_4654,In_118,In_858);
and U4655 (N_4655,In_953,In_919);
or U4656 (N_4656,In_271,In_890);
nor U4657 (N_4657,In_327,In_688);
or U4658 (N_4658,In_311,In_536);
nor U4659 (N_4659,In_240,In_540);
and U4660 (N_4660,In_453,In_655);
and U4661 (N_4661,In_342,In_106);
or U4662 (N_4662,In_910,In_38);
or U4663 (N_4663,In_110,In_116);
or U4664 (N_4664,In_568,In_871);
or U4665 (N_4665,In_433,In_261);
or U4666 (N_4666,In_714,In_607);
and U4667 (N_4667,In_606,In_144);
or U4668 (N_4668,In_7,In_785);
or U4669 (N_4669,In_611,In_826);
or U4670 (N_4670,In_795,In_670);
and U4671 (N_4671,In_46,In_442);
nor U4672 (N_4672,In_64,In_360);
xor U4673 (N_4673,In_506,In_404);
or U4674 (N_4674,In_572,In_97);
nor U4675 (N_4675,In_394,In_8);
nor U4676 (N_4676,In_581,In_291);
and U4677 (N_4677,In_183,In_636);
nand U4678 (N_4678,In_843,In_417);
nand U4679 (N_4679,In_865,In_482);
xor U4680 (N_4680,In_529,In_746);
nand U4681 (N_4681,In_419,In_483);
nand U4682 (N_4682,In_797,In_191);
and U4683 (N_4683,In_932,In_348);
or U4684 (N_4684,In_478,In_252);
and U4685 (N_4685,In_941,In_717);
xnor U4686 (N_4686,In_618,In_879);
xnor U4687 (N_4687,In_763,In_222);
and U4688 (N_4688,In_18,In_789);
and U4689 (N_4689,In_736,In_793);
or U4690 (N_4690,In_579,In_365);
nand U4691 (N_4691,In_650,In_912);
nor U4692 (N_4692,In_84,In_669);
nand U4693 (N_4693,In_176,In_170);
nand U4694 (N_4694,In_709,In_35);
or U4695 (N_4695,In_561,In_866);
and U4696 (N_4696,In_941,In_606);
nor U4697 (N_4697,In_914,In_786);
or U4698 (N_4698,In_325,In_940);
nor U4699 (N_4699,In_574,In_343);
and U4700 (N_4700,In_219,In_794);
nor U4701 (N_4701,In_85,In_272);
and U4702 (N_4702,In_420,In_22);
and U4703 (N_4703,In_931,In_818);
or U4704 (N_4704,In_774,In_275);
xnor U4705 (N_4705,In_384,In_614);
or U4706 (N_4706,In_426,In_751);
nand U4707 (N_4707,In_26,In_333);
nor U4708 (N_4708,In_807,In_21);
xnor U4709 (N_4709,In_913,In_431);
nor U4710 (N_4710,In_4,In_29);
and U4711 (N_4711,In_892,In_948);
nand U4712 (N_4712,In_995,In_676);
xnor U4713 (N_4713,In_227,In_936);
and U4714 (N_4714,In_338,In_47);
nand U4715 (N_4715,In_756,In_820);
and U4716 (N_4716,In_217,In_543);
nand U4717 (N_4717,In_832,In_547);
or U4718 (N_4718,In_773,In_758);
nor U4719 (N_4719,In_75,In_563);
xor U4720 (N_4720,In_837,In_751);
and U4721 (N_4721,In_912,In_494);
nor U4722 (N_4722,In_266,In_363);
or U4723 (N_4723,In_702,In_565);
nor U4724 (N_4724,In_692,In_709);
or U4725 (N_4725,In_205,In_273);
nor U4726 (N_4726,In_328,In_357);
nor U4727 (N_4727,In_233,In_535);
or U4728 (N_4728,In_894,In_127);
or U4729 (N_4729,In_395,In_54);
nor U4730 (N_4730,In_685,In_425);
nor U4731 (N_4731,In_488,In_765);
or U4732 (N_4732,In_845,In_804);
nand U4733 (N_4733,In_919,In_279);
or U4734 (N_4734,In_793,In_935);
or U4735 (N_4735,In_395,In_57);
nand U4736 (N_4736,In_510,In_755);
and U4737 (N_4737,In_334,In_370);
or U4738 (N_4738,In_4,In_613);
nor U4739 (N_4739,In_316,In_380);
and U4740 (N_4740,In_739,In_990);
or U4741 (N_4741,In_99,In_601);
nor U4742 (N_4742,In_477,In_522);
and U4743 (N_4743,In_742,In_343);
and U4744 (N_4744,In_199,In_568);
xnor U4745 (N_4745,In_952,In_971);
nor U4746 (N_4746,In_435,In_550);
xnor U4747 (N_4747,In_338,In_678);
nand U4748 (N_4748,In_289,In_844);
and U4749 (N_4749,In_446,In_251);
and U4750 (N_4750,In_687,In_253);
or U4751 (N_4751,In_453,In_599);
or U4752 (N_4752,In_686,In_377);
xor U4753 (N_4753,In_52,In_40);
nor U4754 (N_4754,In_286,In_431);
xnor U4755 (N_4755,In_140,In_475);
or U4756 (N_4756,In_821,In_308);
xor U4757 (N_4757,In_288,In_974);
nand U4758 (N_4758,In_319,In_16);
or U4759 (N_4759,In_945,In_108);
nor U4760 (N_4760,In_287,In_204);
nor U4761 (N_4761,In_144,In_663);
nor U4762 (N_4762,In_305,In_606);
and U4763 (N_4763,In_374,In_394);
xnor U4764 (N_4764,In_672,In_497);
or U4765 (N_4765,In_803,In_497);
nand U4766 (N_4766,In_352,In_279);
nand U4767 (N_4767,In_828,In_876);
and U4768 (N_4768,In_906,In_841);
nand U4769 (N_4769,In_953,In_301);
or U4770 (N_4770,In_946,In_6);
or U4771 (N_4771,In_910,In_888);
or U4772 (N_4772,In_894,In_190);
or U4773 (N_4773,In_223,In_457);
nor U4774 (N_4774,In_512,In_682);
or U4775 (N_4775,In_884,In_561);
or U4776 (N_4776,In_617,In_41);
xor U4777 (N_4777,In_585,In_926);
or U4778 (N_4778,In_269,In_663);
nor U4779 (N_4779,In_311,In_90);
or U4780 (N_4780,In_626,In_389);
nand U4781 (N_4781,In_822,In_988);
or U4782 (N_4782,In_966,In_432);
and U4783 (N_4783,In_375,In_274);
nor U4784 (N_4784,In_140,In_521);
xor U4785 (N_4785,In_209,In_182);
nand U4786 (N_4786,In_769,In_217);
nor U4787 (N_4787,In_812,In_664);
nor U4788 (N_4788,In_525,In_485);
nor U4789 (N_4789,In_953,In_760);
nor U4790 (N_4790,In_535,In_534);
nand U4791 (N_4791,In_801,In_679);
nor U4792 (N_4792,In_4,In_942);
nand U4793 (N_4793,In_177,In_536);
and U4794 (N_4794,In_184,In_448);
or U4795 (N_4795,In_254,In_788);
or U4796 (N_4796,In_315,In_825);
nor U4797 (N_4797,In_418,In_752);
and U4798 (N_4798,In_98,In_349);
or U4799 (N_4799,In_859,In_58);
or U4800 (N_4800,In_830,In_540);
nor U4801 (N_4801,In_990,In_985);
xor U4802 (N_4802,In_839,In_856);
xor U4803 (N_4803,In_603,In_566);
and U4804 (N_4804,In_36,In_874);
and U4805 (N_4805,In_981,In_692);
and U4806 (N_4806,In_645,In_34);
nor U4807 (N_4807,In_555,In_15);
nor U4808 (N_4808,In_291,In_111);
nor U4809 (N_4809,In_251,In_81);
xnor U4810 (N_4810,In_866,In_120);
xor U4811 (N_4811,In_703,In_938);
or U4812 (N_4812,In_26,In_421);
and U4813 (N_4813,In_239,In_866);
nor U4814 (N_4814,In_240,In_516);
nand U4815 (N_4815,In_838,In_344);
nand U4816 (N_4816,In_812,In_543);
nor U4817 (N_4817,In_278,In_105);
nor U4818 (N_4818,In_683,In_553);
nor U4819 (N_4819,In_47,In_30);
and U4820 (N_4820,In_878,In_966);
and U4821 (N_4821,In_71,In_742);
xnor U4822 (N_4822,In_396,In_121);
or U4823 (N_4823,In_943,In_124);
nor U4824 (N_4824,In_539,In_322);
nand U4825 (N_4825,In_592,In_494);
and U4826 (N_4826,In_43,In_438);
nand U4827 (N_4827,In_566,In_727);
nor U4828 (N_4828,In_314,In_512);
xnor U4829 (N_4829,In_107,In_829);
nor U4830 (N_4830,In_802,In_155);
or U4831 (N_4831,In_899,In_610);
nand U4832 (N_4832,In_700,In_912);
nor U4833 (N_4833,In_407,In_403);
nand U4834 (N_4834,In_84,In_336);
nor U4835 (N_4835,In_360,In_578);
nand U4836 (N_4836,In_473,In_676);
and U4837 (N_4837,In_622,In_6);
or U4838 (N_4838,In_470,In_990);
and U4839 (N_4839,In_138,In_679);
or U4840 (N_4840,In_680,In_564);
or U4841 (N_4841,In_964,In_427);
nand U4842 (N_4842,In_935,In_316);
nand U4843 (N_4843,In_233,In_999);
nand U4844 (N_4844,In_350,In_861);
nand U4845 (N_4845,In_296,In_110);
nand U4846 (N_4846,In_517,In_838);
or U4847 (N_4847,In_570,In_280);
or U4848 (N_4848,In_872,In_455);
or U4849 (N_4849,In_180,In_649);
nor U4850 (N_4850,In_851,In_479);
or U4851 (N_4851,In_468,In_157);
and U4852 (N_4852,In_365,In_660);
and U4853 (N_4853,In_464,In_32);
or U4854 (N_4854,In_8,In_798);
nor U4855 (N_4855,In_318,In_999);
xnor U4856 (N_4856,In_263,In_759);
nand U4857 (N_4857,In_67,In_241);
nor U4858 (N_4858,In_566,In_776);
nor U4859 (N_4859,In_380,In_196);
nor U4860 (N_4860,In_723,In_958);
xor U4861 (N_4861,In_436,In_524);
nand U4862 (N_4862,In_149,In_827);
nor U4863 (N_4863,In_682,In_229);
nand U4864 (N_4864,In_954,In_158);
and U4865 (N_4865,In_159,In_56);
and U4866 (N_4866,In_396,In_36);
nand U4867 (N_4867,In_6,In_32);
nor U4868 (N_4868,In_300,In_534);
nand U4869 (N_4869,In_253,In_240);
nand U4870 (N_4870,In_666,In_487);
and U4871 (N_4871,In_778,In_559);
xnor U4872 (N_4872,In_898,In_783);
nand U4873 (N_4873,In_227,In_959);
xnor U4874 (N_4874,In_174,In_372);
or U4875 (N_4875,In_688,In_564);
xnor U4876 (N_4876,In_780,In_672);
nand U4877 (N_4877,In_819,In_182);
nand U4878 (N_4878,In_469,In_582);
nor U4879 (N_4879,In_546,In_196);
or U4880 (N_4880,In_693,In_594);
xnor U4881 (N_4881,In_754,In_264);
nor U4882 (N_4882,In_422,In_111);
nor U4883 (N_4883,In_1,In_827);
nand U4884 (N_4884,In_217,In_302);
and U4885 (N_4885,In_274,In_294);
nand U4886 (N_4886,In_907,In_598);
nand U4887 (N_4887,In_79,In_749);
nand U4888 (N_4888,In_196,In_467);
nand U4889 (N_4889,In_741,In_428);
nor U4890 (N_4890,In_429,In_828);
or U4891 (N_4891,In_807,In_737);
and U4892 (N_4892,In_731,In_29);
nand U4893 (N_4893,In_171,In_310);
nor U4894 (N_4894,In_138,In_705);
nand U4895 (N_4895,In_323,In_751);
nor U4896 (N_4896,In_267,In_635);
nor U4897 (N_4897,In_296,In_628);
or U4898 (N_4898,In_602,In_953);
or U4899 (N_4899,In_629,In_298);
nand U4900 (N_4900,In_3,In_855);
and U4901 (N_4901,In_303,In_975);
or U4902 (N_4902,In_158,In_852);
xor U4903 (N_4903,In_563,In_850);
and U4904 (N_4904,In_574,In_295);
xor U4905 (N_4905,In_94,In_729);
xor U4906 (N_4906,In_295,In_499);
and U4907 (N_4907,In_8,In_356);
and U4908 (N_4908,In_924,In_826);
nand U4909 (N_4909,In_204,In_317);
xor U4910 (N_4910,In_133,In_194);
xnor U4911 (N_4911,In_148,In_40);
xor U4912 (N_4912,In_190,In_634);
xnor U4913 (N_4913,In_18,In_113);
and U4914 (N_4914,In_31,In_157);
or U4915 (N_4915,In_20,In_132);
nor U4916 (N_4916,In_662,In_475);
and U4917 (N_4917,In_617,In_775);
or U4918 (N_4918,In_800,In_985);
nand U4919 (N_4919,In_475,In_344);
and U4920 (N_4920,In_683,In_212);
nor U4921 (N_4921,In_758,In_332);
and U4922 (N_4922,In_644,In_554);
or U4923 (N_4923,In_907,In_996);
xor U4924 (N_4924,In_653,In_999);
nor U4925 (N_4925,In_541,In_405);
or U4926 (N_4926,In_13,In_490);
nor U4927 (N_4927,In_844,In_944);
nand U4928 (N_4928,In_815,In_29);
and U4929 (N_4929,In_326,In_566);
nand U4930 (N_4930,In_681,In_300);
nand U4931 (N_4931,In_366,In_239);
nand U4932 (N_4932,In_789,In_269);
and U4933 (N_4933,In_10,In_354);
xnor U4934 (N_4934,In_60,In_686);
or U4935 (N_4935,In_189,In_740);
nor U4936 (N_4936,In_274,In_185);
or U4937 (N_4937,In_191,In_49);
nand U4938 (N_4938,In_428,In_490);
nor U4939 (N_4939,In_443,In_337);
and U4940 (N_4940,In_536,In_126);
or U4941 (N_4941,In_715,In_347);
xnor U4942 (N_4942,In_357,In_513);
or U4943 (N_4943,In_262,In_249);
nand U4944 (N_4944,In_215,In_212);
nor U4945 (N_4945,In_683,In_367);
and U4946 (N_4946,In_518,In_7);
nand U4947 (N_4947,In_267,In_196);
or U4948 (N_4948,In_565,In_836);
nor U4949 (N_4949,In_597,In_324);
and U4950 (N_4950,In_963,In_574);
nand U4951 (N_4951,In_541,In_336);
xor U4952 (N_4952,In_493,In_855);
nor U4953 (N_4953,In_447,In_129);
or U4954 (N_4954,In_562,In_45);
xor U4955 (N_4955,In_516,In_103);
or U4956 (N_4956,In_715,In_109);
nor U4957 (N_4957,In_294,In_280);
nor U4958 (N_4958,In_801,In_63);
and U4959 (N_4959,In_953,In_917);
and U4960 (N_4960,In_148,In_57);
xnor U4961 (N_4961,In_554,In_939);
or U4962 (N_4962,In_651,In_40);
nor U4963 (N_4963,In_528,In_69);
and U4964 (N_4964,In_722,In_447);
nor U4965 (N_4965,In_658,In_465);
nand U4966 (N_4966,In_62,In_181);
or U4967 (N_4967,In_887,In_0);
nand U4968 (N_4968,In_475,In_623);
nor U4969 (N_4969,In_940,In_409);
and U4970 (N_4970,In_237,In_412);
or U4971 (N_4971,In_85,In_902);
and U4972 (N_4972,In_71,In_87);
nand U4973 (N_4973,In_904,In_553);
or U4974 (N_4974,In_579,In_513);
and U4975 (N_4975,In_780,In_683);
and U4976 (N_4976,In_717,In_934);
nor U4977 (N_4977,In_948,In_409);
nand U4978 (N_4978,In_728,In_346);
or U4979 (N_4979,In_146,In_10);
or U4980 (N_4980,In_598,In_379);
or U4981 (N_4981,In_23,In_807);
or U4982 (N_4982,In_663,In_418);
nor U4983 (N_4983,In_895,In_843);
or U4984 (N_4984,In_329,In_875);
nand U4985 (N_4985,In_182,In_80);
xor U4986 (N_4986,In_971,In_283);
or U4987 (N_4987,In_192,In_124);
xnor U4988 (N_4988,In_628,In_357);
nand U4989 (N_4989,In_937,In_62);
xor U4990 (N_4990,In_1,In_732);
nor U4991 (N_4991,In_926,In_114);
xor U4992 (N_4992,In_859,In_150);
nand U4993 (N_4993,In_938,In_709);
and U4994 (N_4994,In_801,In_494);
and U4995 (N_4995,In_39,In_577);
or U4996 (N_4996,In_659,In_29);
nor U4997 (N_4997,In_931,In_170);
nand U4998 (N_4998,In_46,In_329);
and U4999 (N_4999,In_335,In_869);
or U5000 (N_5000,N_1088,N_2849);
nor U5001 (N_5001,N_3423,N_449);
or U5002 (N_5002,N_4924,N_3578);
or U5003 (N_5003,N_4886,N_3594);
xnor U5004 (N_5004,N_1610,N_2370);
nand U5005 (N_5005,N_3428,N_2567);
nand U5006 (N_5006,N_1710,N_516);
nand U5007 (N_5007,N_1437,N_68);
nand U5008 (N_5008,N_4976,N_2205);
nor U5009 (N_5009,N_4680,N_3012);
and U5010 (N_5010,N_1826,N_4714);
and U5011 (N_5011,N_4136,N_1213);
and U5012 (N_5012,N_1691,N_353);
and U5013 (N_5013,N_4440,N_3288);
nor U5014 (N_5014,N_384,N_542);
nor U5015 (N_5015,N_1686,N_284);
and U5016 (N_5016,N_4177,N_4259);
nand U5017 (N_5017,N_2990,N_4222);
or U5018 (N_5018,N_332,N_2197);
nand U5019 (N_5019,N_1505,N_4786);
or U5020 (N_5020,N_3113,N_3373);
nor U5021 (N_5021,N_4605,N_4404);
or U5022 (N_5022,N_3268,N_4415);
nand U5023 (N_5023,N_2681,N_2314);
xor U5024 (N_5024,N_2328,N_1201);
nor U5025 (N_5025,N_1083,N_2794);
nor U5026 (N_5026,N_4422,N_3009);
nor U5027 (N_5027,N_2626,N_1108);
or U5028 (N_5028,N_4070,N_4048);
or U5029 (N_5029,N_4014,N_3456);
and U5030 (N_5030,N_3172,N_1488);
nand U5031 (N_5031,N_2699,N_374);
or U5032 (N_5032,N_3842,N_530);
nor U5033 (N_5033,N_4783,N_2540);
and U5034 (N_5034,N_4215,N_4956);
nand U5035 (N_5035,N_1314,N_2896);
or U5036 (N_5036,N_3753,N_1582);
and U5037 (N_5037,N_3967,N_495);
or U5038 (N_5038,N_2444,N_403);
nand U5039 (N_5039,N_2694,N_598);
nor U5040 (N_5040,N_510,N_716);
or U5041 (N_5041,N_921,N_3675);
nor U5042 (N_5042,N_3650,N_3345);
nand U5043 (N_5043,N_448,N_4472);
xor U5044 (N_5044,N_351,N_4116);
and U5045 (N_5045,N_55,N_764);
or U5046 (N_5046,N_1172,N_3623);
nor U5047 (N_5047,N_3700,N_3777);
nor U5048 (N_5048,N_2143,N_4474);
nand U5049 (N_5049,N_2703,N_459);
nor U5050 (N_5050,N_320,N_1198);
nand U5051 (N_5051,N_4616,N_976);
nand U5052 (N_5052,N_4436,N_2165);
xor U5053 (N_5053,N_807,N_2604);
or U5054 (N_5054,N_2901,N_1212);
nor U5055 (N_5055,N_4258,N_4851);
and U5056 (N_5056,N_2904,N_896);
or U5057 (N_5057,N_605,N_3786);
nor U5058 (N_5058,N_597,N_3391);
nand U5059 (N_5059,N_3244,N_4842);
nand U5060 (N_5060,N_945,N_1350);
xor U5061 (N_5061,N_835,N_1590);
nand U5062 (N_5062,N_537,N_22);
or U5063 (N_5063,N_4207,N_1336);
nand U5064 (N_5064,N_538,N_4279);
nand U5065 (N_5065,N_65,N_411);
and U5066 (N_5066,N_2474,N_3778);
and U5067 (N_5067,N_4109,N_540);
nor U5068 (N_5068,N_2520,N_1459);
nand U5069 (N_5069,N_1440,N_3323);
nand U5070 (N_5070,N_2397,N_2051);
xor U5071 (N_5071,N_738,N_3496);
or U5072 (N_5072,N_3211,N_1022);
nor U5073 (N_5073,N_382,N_4528);
nand U5074 (N_5074,N_2019,N_3875);
or U5075 (N_5075,N_4683,N_4500);
and U5076 (N_5076,N_2006,N_1103);
and U5077 (N_5077,N_4503,N_2677);
or U5078 (N_5078,N_4719,N_1567);
nor U5079 (N_5079,N_1176,N_2309);
nand U5080 (N_5080,N_1792,N_577);
nor U5081 (N_5081,N_2909,N_4064);
nor U5082 (N_5082,N_1099,N_1308);
nor U5083 (N_5083,N_1701,N_4774);
and U5084 (N_5084,N_2610,N_4505);
nor U5085 (N_5085,N_1704,N_3503);
nor U5086 (N_5086,N_4379,N_1355);
or U5087 (N_5087,N_155,N_1873);
nor U5088 (N_5088,N_1092,N_1476);
and U5089 (N_5089,N_418,N_1422);
nand U5090 (N_5090,N_35,N_518);
and U5091 (N_5091,N_1141,N_4891);
nor U5092 (N_5092,N_2706,N_2163);
and U5093 (N_5093,N_953,N_475);
nor U5094 (N_5094,N_2044,N_256);
or U5095 (N_5095,N_1556,N_792);
nand U5096 (N_5096,N_1418,N_2082);
nor U5097 (N_5097,N_3961,N_507);
or U5098 (N_5098,N_1205,N_4334);
and U5099 (N_5099,N_4321,N_130);
nand U5100 (N_5100,N_4547,N_955);
xnor U5101 (N_5101,N_4370,N_830);
nor U5102 (N_5102,N_2218,N_3067);
and U5103 (N_5103,N_1206,N_3595);
or U5104 (N_5104,N_2176,N_650);
xor U5105 (N_5105,N_975,N_293);
nand U5106 (N_5106,N_840,N_1927);
and U5107 (N_5107,N_2934,N_4834);
nand U5108 (N_5108,N_3591,N_298);
nor U5109 (N_5109,N_188,N_2511);
nor U5110 (N_5110,N_4923,N_1491);
nor U5111 (N_5111,N_4368,N_474);
xor U5112 (N_5112,N_4659,N_1664);
nand U5113 (N_5113,N_4942,N_2382);
nor U5114 (N_5114,N_1045,N_3965);
or U5115 (N_5115,N_684,N_961);
nor U5116 (N_5116,N_1294,N_972);
and U5117 (N_5117,N_4911,N_338);
and U5118 (N_5118,N_87,N_3597);
nand U5119 (N_5119,N_4726,N_1681);
nor U5120 (N_5120,N_4339,N_1279);
nor U5121 (N_5121,N_1102,N_2765);
and U5122 (N_5122,N_436,N_3713);
nor U5123 (N_5123,N_4543,N_2568);
nand U5124 (N_5124,N_360,N_2425);
xor U5125 (N_5125,N_460,N_2977);
and U5126 (N_5126,N_3133,N_671);
and U5127 (N_5127,N_1218,N_949);
or U5128 (N_5128,N_107,N_219);
and U5129 (N_5129,N_2277,N_4099);
nand U5130 (N_5130,N_4179,N_3197);
nor U5131 (N_5131,N_2516,N_1508);
and U5132 (N_5132,N_2641,N_2895);
nor U5133 (N_5133,N_3654,N_2938);
nand U5134 (N_5134,N_124,N_2409);
and U5135 (N_5135,N_3624,N_2774);
and U5136 (N_5136,N_3564,N_2858);
and U5137 (N_5137,N_3586,N_1276);
nand U5138 (N_5138,N_4518,N_3604);
nor U5139 (N_5139,N_349,N_3673);
nand U5140 (N_5140,N_4088,N_1760);
or U5141 (N_5141,N_3033,N_914);
nand U5142 (N_5142,N_4905,N_3336);
nand U5143 (N_5143,N_4311,N_4153);
nand U5144 (N_5144,N_4254,N_2480);
or U5145 (N_5145,N_435,N_29);
or U5146 (N_5146,N_1529,N_3402);
and U5147 (N_5147,N_3412,N_86);
nor U5148 (N_5148,N_1665,N_3659);
nand U5149 (N_5149,N_2380,N_3555);
nor U5150 (N_5150,N_454,N_2431);
nand U5151 (N_5151,N_311,N_2814);
nand U5152 (N_5152,N_1384,N_1601);
and U5153 (N_5153,N_3910,N_15);
nand U5154 (N_5154,N_3638,N_3621);
and U5155 (N_5155,N_3499,N_3683);
nand U5156 (N_5156,N_4283,N_4508);
and U5157 (N_5157,N_1475,N_1893);
nand U5158 (N_5158,N_243,N_2253);
and U5159 (N_5159,N_1140,N_3732);
nor U5160 (N_5160,N_4054,N_4164);
or U5161 (N_5161,N_1284,N_3854);
or U5162 (N_5162,N_3204,N_3494);
nand U5163 (N_5163,N_169,N_3188);
and U5164 (N_5164,N_4425,N_4243);
nand U5165 (N_5165,N_626,N_2771);
and U5166 (N_5166,N_3246,N_3461);
or U5167 (N_5167,N_1327,N_2209);
nand U5168 (N_5168,N_2462,N_3301);
or U5169 (N_5169,N_2929,N_1639);
or U5170 (N_5170,N_487,N_4560);
nor U5171 (N_5171,N_1097,N_1799);
and U5172 (N_5172,N_214,N_4042);
and U5173 (N_5173,N_1546,N_1771);
and U5174 (N_5174,N_4702,N_4183);
nand U5175 (N_5175,N_4374,N_2869);
nand U5176 (N_5176,N_1095,N_1575);
or U5177 (N_5177,N_1076,N_4304);
nand U5178 (N_5178,N_4507,N_3874);
nor U5179 (N_5179,N_37,N_3250);
nand U5180 (N_5180,N_2149,N_1400);
and U5181 (N_5181,N_343,N_3648);
or U5182 (N_5182,N_2288,N_4402);
nand U5183 (N_5183,N_4408,N_4716);
or U5184 (N_5184,N_765,N_581);
or U5185 (N_5185,N_3386,N_4821);
nand U5186 (N_5186,N_1419,N_1887);
nand U5187 (N_5187,N_1896,N_2062);
nor U5188 (N_5188,N_958,N_3319);
and U5189 (N_5189,N_3598,N_3614);
and U5190 (N_5190,N_2999,N_1617);
nor U5191 (N_5191,N_888,N_2112);
and U5192 (N_5192,N_3697,N_630);
nand U5193 (N_5193,N_3862,N_2490);
xnor U5194 (N_5194,N_4718,N_1146);
or U5195 (N_5195,N_140,N_2061);
xnor U5196 (N_5196,N_1075,N_1660);
and U5197 (N_5197,N_2427,N_2278);
and U5198 (N_5198,N_488,N_3796);
nor U5199 (N_5199,N_4953,N_4214);
and U5200 (N_5200,N_4754,N_1395);
nor U5201 (N_5201,N_3734,N_4388);
nand U5202 (N_5202,N_39,N_2730);
and U5203 (N_5203,N_162,N_873);
and U5204 (N_5204,N_3596,N_2429);
and U5205 (N_5205,N_1458,N_1871);
and U5206 (N_5206,N_1862,N_450);
xor U5207 (N_5207,N_4029,N_3532);
xor U5208 (N_5208,N_1137,N_1456);
or U5209 (N_5209,N_2147,N_1521);
nand U5210 (N_5210,N_612,N_920);
nand U5211 (N_5211,N_1714,N_4535);
nand U5212 (N_5212,N_4649,N_1929);
nor U5213 (N_5213,N_1132,N_3240);
or U5214 (N_5214,N_782,N_296);
and U5215 (N_5215,N_2925,N_3921);
and U5216 (N_5216,N_3147,N_845);
nand U5217 (N_5217,N_3587,N_0);
or U5218 (N_5218,N_4655,N_1415);
nand U5219 (N_5219,N_1585,N_3685);
nor U5220 (N_5220,N_3677,N_368);
nor U5221 (N_5221,N_1939,N_4701);
nand U5222 (N_5222,N_1588,N_1461);
xnor U5223 (N_5223,N_4584,N_4077);
nor U5224 (N_5224,N_3031,N_3138);
and U5225 (N_5225,N_3607,N_1436);
and U5226 (N_5226,N_2942,N_1775);
nor U5227 (N_5227,N_2401,N_3665);
and U5228 (N_5228,N_4089,N_752);
and U5229 (N_5229,N_3210,N_2827);
nand U5230 (N_5230,N_1304,N_3696);
nand U5231 (N_5231,N_3892,N_1693);
nor U5232 (N_5232,N_2748,N_4926);
nand U5233 (N_5233,N_1010,N_1913);
and U5234 (N_5234,N_512,N_1646);
xor U5235 (N_5235,N_4372,N_4004);
nor U5236 (N_5236,N_32,N_20);
xnor U5237 (N_5237,N_3284,N_4712);
nand U5238 (N_5238,N_4181,N_472);
or U5239 (N_5239,N_3296,N_1290);
xnor U5240 (N_5240,N_2248,N_1044);
or U5241 (N_5241,N_3377,N_2060);
xnor U5242 (N_5242,N_365,N_3452);
or U5243 (N_5243,N_4228,N_527);
or U5244 (N_5244,N_4567,N_962);
nand U5245 (N_5245,N_2717,N_3905);
nor U5246 (N_5246,N_2832,N_327);
xor U5247 (N_5247,N_3370,N_3759);
nand U5248 (N_5248,N_2598,N_1298);
or U5249 (N_5249,N_2788,N_4600);
nand U5250 (N_5250,N_3046,N_3127);
or U5251 (N_5251,N_1840,N_1204);
and U5252 (N_5252,N_4652,N_2530);
and U5253 (N_5253,N_359,N_4144);
and U5254 (N_5254,N_2004,N_319);
nand U5255 (N_5255,N_153,N_744);
nor U5256 (N_5256,N_3833,N_4050);
nand U5257 (N_5257,N_4271,N_543);
nor U5258 (N_5258,N_2737,N_3821);
nand U5259 (N_5259,N_3567,N_1560);
or U5260 (N_5260,N_3937,N_4628);
nor U5261 (N_5261,N_3890,N_2536);
and U5262 (N_5262,N_2663,N_1173);
nor U5263 (N_5263,N_4841,N_251);
nor U5264 (N_5264,N_2271,N_4142);
and U5265 (N_5265,N_1725,N_600);
and U5266 (N_5266,N_2624,N_261);
and U5267 (N_5267,N_3415,N_4951);
nand U5268 (N_5268,N_4693,N_1853);
nand U5269 (N_5269,N_3084,N_2643);
nand U5270 (N_5270,N_3514,N_4689);
or U5271 (N_5271,N_4172,N_508);
or U5272 (N_5272,N_3626,N_2813);
xor U5273 (N_5273,N_4594,N_1071);
or U5274 (N_5274,N_1987,N_2291);
nor U5275 (N_5275,N_805,N_3077);
nand U5276 (N_5276,N_2825,N_726);
or U5277 (N_5277,N_4987,N_615);
or U5278 (N_5278,N_3312,N_4313);
or U5279 (N_5279,N_4333,N_4103);
nand U5280 (N_5280,N_3531,N_4631);
and U5281 (N_5281,N_4804,N_1907);
and U5282 (N_5282,N_2662,N_795);
nand U5283 (N_5283,N_3277,N_1248);
and U5284 (N_5284,N_2974,N_2495);
nor U5285 (N_5285,N_811,N_1427);
nor U5286 (N_5286,N_2582,N_582);
or U5287 (N_5287,N_2809,N_2222);
and U5288 (N_5288,N_1729,N_2948);
xnor U5289 (N_5289,N_3105,N_4364);
nand U5290 (N_5290,N_1448,N_484);
or U5291 (N_5291,N_4908,N_3422);
nand U5292 (N_5292,N_101,N_4565);
nand U5293 (N_5293,N_3966,N_4041);
and U5294 (N_5294,N_899,N_1420);
xor U5295 (N_5295,N_115,N_2816);
nor U5296 (N_5296,N_2894,N_610);
and U5297 (N_5297,N_3995,N_3305);
nor U5298 (N_5298,N_3027,N_637);
or U5299 (N_5299,N_1550,N_2908);
or U5300 (N_5300,N_3234,N_2408);
or U5301 (N_5301,N_4520,N_3475);
nor U5302 (N_5302,N_3987,N_4833);
or U5303 (N_5303,N_2965,N_4371);
or U5304 (N_5304,N_1159,N_1531);
or U5305 (N_5305,N_3181,N_159);
and U5306 (N_5306,N_4295,N_864);
or U5307 (N_5307,N_2068,N_4767);
and U5308 (N_5308,N_1313,N_1905);
nand U5309 (N_5309,N_4017,N_3157);
or U5310 (N_5310,N_1779,N_1796);
and U5311 (N_5311,N_1062,N_2998);
nand U5312 (N_5312,N_3397,N_2808);
nor U5313 (N_5313,N_657,N_2295);
or U5314 (N_5314,N_1877,N_4133);
or U5315 (N_5315,N_2340,N_4185);
xnor U5316 (N_5316,N_3958,N_2870);
nor U5317 (N_5317,N_1202,N_3752);
and U5318 (N_5318,N_1101,N_3363);
or U5319 (N_5319,N_554,N_4820);
and U5320 (N_5320,N_4145,N_2014);
or U5321 (N_5321,N_861,N_266);
and U5322 (N_5322,N_4984,N_2466);
and U5323 (N_5323,N_2233,N_2400);
or U5324 (N_5324,N_2220,N_2763);
nor U5325 (N_5325,N_2216,N_1100);
nand U5326 (N_5326,N_1481,N_2415);
and U5327 (N_5327,N_2919,N_2056);
nand U5328 (N_5328,N_3886,N_642);
nor U5329 (N_5329,N_1995,N_4630);
xor U5330 (N_5330,N_3471,N_1018);
nand U5331 (N_5331,N_437,N_3693);
and U5332 (N_5332,N_3898,N_951);
or U5333 (N_5333,N_1744,N_427);
and U5334 (N_5334,N_3346,N_3448);
or U5335 (N_5335,N_971,N_3791);
nand U5336 (N_5336,N_171,N_1362);
and U5337 (N_5337,N_1372,N_205);
or U5338 (N_5338,N_370,N_2967);
nor U5339 (N_5339,N_245,N_1688);
and U5340 (N_5340,N_4843,N_1680);
nand U5341 (N_5341,N_4173,N_3913);
nand U5342 (N_5342,N_2432,N_1605);
xor U5343 (N_5343,N_3110,N_4865);
or U5344 (N_5344,N_3276,N_392);
or U5345 (N_5345,N_1397,N_851);
or U5346 (N_5346,N_1787,N_679);
or U5347 (N_5347,N_4491,N_838);
and U5348 (N_5348,N_3573,N_3477);
or U5349 (N_5349,N_2261,N_4779);
and U5350 (N_5350,N_2399,N_2489);
or U5351 (N_5351,N_1662,N_948);
nor U5352 (N_5352,N_2879,N_555);
nor U5353 (N_5353,N_4129,N_3869);
or U5354 (N_5354,N_2971,N_2544);
nor U5355 (N_5355,N_656,N_1453);
nor U5356 (N_5356,N_2303,N_99);
and U5357 (N_5357,N_4239,N_978);
and U5358 (N_5358,N_1906,N_3837);
nor U5359 (N_5359,N_2124,N_3652);
nor U5360 (N_5360,N_786,N_889);
and U5361 (N_5361,N_3960,N_341);
or U5362 (N_5362,N_578,N_2921);
nand U5363 (N_5363,N_3949,N_2607);
nand U5364 (N_5364,N_78,N_2933);
nand U5365 (N_5365,N_4000,N_2543);
and U5366 (N_5366,N_687,N_4894);
or U5367 (N_5367,N_1558,N_2649);
and U5368 (N_5368,N_4375,N_3727);
and U5369 (N_5369,N_2365,N_2029);
nor U5370 (N_5370,N_3616,N_4195);
nor U5371 (N_5371,N_4893,N_4967);
xor U5372 (N_5372,N_3316,N_4949);
xnor U5373 (N_5373,N_2549,N_4575);
nor U5374 (N_5374,N_526,N_1914);
xnor U5375 (N_5375,N_501,N_4853);
nand U5376 (N_5376,N_1300,N_399);
nor U5377 (N_5377,N_2606,N_2752);
nand U5378 (N_5378,N_3381,N_806);
nand U5379 (N_5379,N_4350,N_1207);
nor U5380 (N_5380,N_1940,N_878);
or U5381 (N_5381,N_1403,N_2134);
nand U5382 (N_5382,N_1330,N_2105);
nor U5383 (N_5383,N_439,N_3457);
nor U5384 (N_5384,N_3389,N_935);
xor U5385 (N_5385,N_3146,N_4939);
nor U5386 (N_5386,N_2012,N_706);
and U5387 (N_5387,N_3203,N_2089);
or U5388 (N_5388,N_4531,N_4648);
nor U5389 (N_5389,N_514,N_317);
and U5390 (N_5390,N_347,N_2636);
or U5391 (N_5391,N_2043,N_663);
nor U5392 (N_5392,N_1839,N_2762);
or U5393 (N_5393,N_2113,N_2839);
or U5394 (N_5394,N_16,N_1255);
nor U5395 (N_5395,N_4309,N_2426);
or U5396 (N_5396,N_762,N_4272);
xor U5397 (N_5397,N_768,N_886);
nand U5398 (N_5398,N_4387,N_952);
nand U5399 (N_5399,N_1769,N_4378);
nor U5400 (N_5400,N_3804,N_1346);
and U5401 (N_5401,N_865,N_3259);
nand U5402 (N_5402,N_932,N_3429);
and U5403 (N_5403,N_2665,N_1450);
nor U5404 (N_5404,N_2375,N_2414);
or U5405 (N_5405,N_2026,N_312);
and U5406 (N_5406,N_429,N_4685);
or U5407 (N_5407,N_1183,N_4502);
and U5408 (N_5408,N_2407,N_1916);
xnor U5409 (N_5409,N_4935,N_357);
xnor U5410 (N_5410,N_1162,N_992);
nand U5411 (N_5411,N_1563,N_2321);
nor U5412 (N_5412,N_2411,N_192);
or U5413 (N_5413,N_784,N_2419);
nand U5414 (N_5414,N_2772,N_239);
and U5415 (N_5415,N_2349,N_4204);
xnor U5416 (N_5416,N_4263,N_3201);
nor U5417 (N_5417,N_2308,N_2951);
and U5418 (N_5418,N_500,N_3800);
nand U5419 (N_5419,N_3577,N_371);
nand U5420 (N_5420,N_1741,N_2270);
nor U5421 (N_5421,N_1363,N_4592);
nor U5422 (N_5422,N_3534,N_4169);
nand U5423 (N_5423,N_4517,N_999);
nor U5424 (N_5424,N_4982,N_569);
nand U5425 (N_5425,N_217,N_940);
nand U5426 (N_5426,N_4098,N_1502);
and U5427 (N_5427,N_2650,N_3168);
nor U5428 (N_5428,N_4848,N_4051);
nand U5429 (N_5429,N_1245,N_3171);
xor U5430 (N_5430,N_4538,N_1874);
and U5431 (N_5431,N_1539,N_3006);
nand U5432 (N_5432,N_3334,N_236);
or U5433 (N_5433,N_1265,N_2387);
and U5434 (N_5434,N_2221,N_3841);
nor U5435 (N_5435,N_3055,N_4542);
and U5436 (N_5436,N_4020,N_2344);
xnor U5437 (N_5437,N_379,N_4997);
or U5438 (N_5438,N_3065,N_2651);
and U5439 (N_5439,N_4721,N_2484);
nand U5440 (N_5440,N_3088,N_3450);
nand U5441 (N_5441,N_3969,N_2383);
and U5442 (N_5442,N_4396,N_789);
nand U5443 (N_5443,N_4369,N_3142);
nor U5444 (N_5444,N_257,N_787);
xor U5445 (N_5445,N_660,N_3207);
and U5446 (N_5446,N_3897,N_2857);
nand U5447 (N_5447,N_3001,N_2889);
nand U5448 (N_5448,N_4147,N_3134);
nand U5449 (N_5449,N_4094,N_4138);
or U5450 (N_5450,N_1707,N_56);
or U5451 (N_5451,N_413,N_2041);
and U5452 (N_5452,N_3335,N_3498);
nor U5453 (N_5453,N_640,N_2562);
nor U5454 (N_5454,N_4019,N_2276);
nand U5455 (N_5455,N_592,N_3882);
xnor U5456 (N_5456,N_4516,N_903);
nand U5457 (N_5457,N_4838,N_4551);
and U5458 (N_5458,N_3900,N_2880);
nor U5459 (N_5459,N_4078,N_1910);
or U5460 (N_5460,N_2196,N_1636);
nor U5461 (N_5461,N_994,N_2623);
nand U5462 (N_5462,N_3689,N_2232);
or U5463 (N_5463,N_2773,N_4130);
nor U5464 (N_5464,N_2726,N_2701);
or U5465 (N_5465,N_2286,N_119);
xor U5466 (N_5466,N_2517,N_4969);
and U5467 (N_5467,N_4665,N_2842);
nor U5468 (N_5468,N_1150,N_3431);
or U5469 (N_5469,N_2445,N_3658);
nor U5470 (N_5470,N_1226,N_2733);
and U5471 (N_5471,N_2692,N_1003);
or U5472 (N_5472,N_3014,N_1193);
nor U5473 (N_5473,N_57,N_2787);
or U5474 (N_5474,N_203,N_925);
nor U5475 (N_5475,N_3580,N_2843);
xnor U5476 (N_5476,N_2352,N_2173);
or U5477 (N_5477,N_4522,N_653);
and U5478 (N_5478,N_3656,N_2900);
or U5479 (N_5479,N_799,N_639);
xor U5480 (N_5480,N_2053,N_2674);
nand U5481 (N_5481,N_4105,N_1780);
nand U5482 (N_5482,N_47,N_1865);
xor U5483 (N_5483,N_3979,N_4900);
or U5484 (N_5484,N_446,N_2386);
nor U5485 (N_5485,N_560,N_34);
nand U5486 (N_5486,N_4610,N_2910);
or U5487 (N_5487,N_4634,N_506);
or U5488 (N_5488,N_3694,N_3372);
nor U5489 (N_5489,N_4571,N_1609);
nor U5490 (N_5490,N_4977,N_4564);
or U5491 (N_5491,N_1053,N_1122);
and U5492 (N_5492,N_361,N_1698);
xnor U5493 (N_5493,N_1517,N_1189);
and U5494 (N_5494,N_1394,N_348);
xnor U5495 (N_5495,N_2793,N_3779);
and U5496 (N_5496,N_4839,N_2659);
and U5497 (N_5497,N_4810,N_550);
xor U5498 (N_5498,N_149,N_4373);
nand U5499 (N_5499,N_2855,N_3215);
and U5500 (N_5500,N_3068,N_2625);
and U5501 (N_5501,N_1953,N_2767);
xor U5502 (N_5502,N_2059,N_3283);
and U5503 (N_5503,N_3470,N_4161);
and U5504 (N_5504,N_4979,N_1264);
nand U5505 (N_5505,N_2478,N_559);
and U5506 (N_5506,N_3636,N_3628);
and U5507 (N_5507,N_897,N_2437);
and U5508 (N_5508,N_51,N_27);
and U5509 (N_5509,N_3893,N_822);
and U5510 (N_5510,N_2362,N_2577);
and U5511 (N_5511,N_3836,N_4134);
and U5512 (N_5512,N_1977,N_295);
or U5513 (N_5513,N_941,N_3540);
nand U5514 (N_5514,N_4148,N_1960);
nand U5515 (N_5515,N_1723,N_4018);
or U5516 (N_5516,N_1922,N_1990);
nand U5517 (N_5517,N_4947,N_2704);
nand U5518 (N_5518,N_2410,N_2956);
or U5519 (N_5519,N_520,N_1899);
and U5520 (N_5520,N_815,N_4081);
nor U5521 (N_5521,N_1217,N_1890);
nor U5522 (N_5522,N_3169,N_1435);
nand U5523 (N_5523,N_850,N_19);
and U5524 (N_5524,N_3563,N_3630);
xor U5525 (N_5525,N_1889,N_4242);
nand U5526 (N_5526,N_233,N_1036);
nor U5527 (N_5527,N_1370,N_3092);
xor U5528 (N_5528,N_3165,N_4732);
nor U5529 (N_5529,N_3343,N_4731);
nor U5530 (N_5530,N_3416,N_2137);
and U5531 (N_5531,N_2280,N_1802);
or U5532 (N_5532,N_4290,N_2509);
nor U5533 (N_5533,N_2175,N_2453);
nand U5534 (N_5534,N_3187,N_4430);
nand U5535 (N_5535,N_4460,N_184);
and U5536 (N_5536,N_536,N_3376);
xor U5537 (N_5537,N_2472,N_67);
nor U5538 (N_5538,N_3123,N_885);
and U5539 (N_5539,N_4326,N_1894);
nor U5540 (N_5540,N_1465,N_2713);
nor U5541 (N_5541,N_901,N_4510);
nor U5542 (N_5542,N_4633,N_1593);
xnor U5543 (N_5543,N_4559,N_1087);
or U5544 (N_5544,N_643,N_1188);
or U5545 (N_5545,N_737,N_386);
and U5546 (N_5546,N_441,N_4359);
and U5547 (N_5547,N_3091,N_1559);
and U5548 (N_5548,N_3190,N_699);
xnor U5549 (N_5549,N_2388,N_421);
nor U5550 (N_5550,N_1497,N_1528);
xor U5551 (N_5551,N_206,N_3390);
nor U5552 (N_5552,N_731,N_3755);
and U5553 (N_5553,N_4638,N_4598);
or U5554 (N_5554,N_2817,N_3660);
nor U5555 (N_5555,N_2807,N_834);
nor U5556 (N_5556,N_1014,N_3844);
nand U5557 (N_5557,N_3029,N_528);
and U5558 (N_5558,N_4798,N_1325);
xor U5559 (N_5559,N_3468,N_1446);
and U5560 (N_5560,N_4724,N_4027);
or U5561 (N_5561,N_3795,N_142);
nand U5562 (N_5562,N_267,N_2104);
and U5563 (N_5563,N_1342,N_4845);
nand U5564 (N_5564,N_4624,N_517);
or U5565 (N_5565,N_2348,N_3380);
nand U5566 (N_5566,N_2668,N_2497);
or U5567 (N_5567,N_1892,N_2768);
and U5568 (N_5568,N_867,N_3999);
xor U5569 (N_5569,N_4395,N_3909);
xnor U5570 (N_5570,N_3294,N_1032);
or U5571 (N_5571,N_808,N_2742);
and U5572 (N_5572,N_4858,N_4753);
nand U5573 (N_5573,N_4730,N_3249);
or U5574 (N_5574,N_3863,N_2202);
xnor U5575 (N_5575,N_1788,N_2036);
nand U5576 (N_5576,N_4080,N_3359);
nor U5577 (N_5577,N_2682,N_4938);
and U5578 (N_5578,N_3112,N_727);
nand U5579 (N_5579,N_674,N_76);
xor U5580 (N_5580,N_4962,N_1982);
nand U5581 (N_5581,N_1257,N_3691);
and U5582 (N_5582,N_4632,N_4645);
xor U5583 (N_5583,N_2574,N_2169);
xnor U5584 (N_5584,N_2501,N_1026);
or U5585 (N_5585,N_3255,N_4646);
nor U5586 (N_5586,N_2770,N_1282);
nor U5587 (N_5587,N_4619,N_4818);
nor U5588 (N_5588,N_1612,N_1514);
nand U5589 (N_5589,N_1349,N_2783);
and U5590 (N_5590,N_1085,N_1167);
or U5591 (N_5591,N_4096,N_12);
nor U5592 (N_5592,N_1523,N_933);
nor U5593 (N_5593,N_4699,N_2395);
nand U5594 (N_5594,N_3538,N_2091);
or U5595 (N_5595,N_1113,N_1711);
and U5596 (N_5596,N_3050,N_4189);
and U5597 (N_5597,N_38,N_496);
or U5598 (N_5598,N_4761,N_1970);
nor U5599 (N_5599,N_4793,N_1042);
nand U5600 (N_5600,N_1604,N_860);
and U5601 (N_5601,N_2116,N_1114);
and U5602 (N_5602,N_4265,N_4284);
or U5603 (N_5603,N_3045,N_4506);
nor U5604 (N_5604,N_1965,N_1552);
or U5605 (N_5605,N_2158,N_2024);
or U5606 (N_5606,N_1107,N_4409);
and U5607 (N_5607,N_2250,N_204);
xor U5608 (N_5608,N_2944,N_2049);
or U5609 (N_5609,N_3899,N_2323);
or U5610 (N_5610,N_1270,N_94);
xnor U5611 (N_5611,N_2596,N_2066);
or U5612 (N_5612,N_4015,N_61);
nor U5613 (N_5613,N_4097,N_4879);
and U5614 (N_5614,N_1829,N_3985);
nand U5615 (N_5615,N_2905,N_1216);
nor U5616 (N_5616,N_227,N_3823);
or U5617 (N_5617,N_4376,N_2247);
and U5618 (N_5618,N_1407,N_3198);
nand U5619 (N_5619,N_1624,N_469);
nand U5620 (N_5620,N_1947,N_2657);
or U5621 (N_5621,N_3264,N_729);
and U5622 (N_5622,N_2629,N_701);
and U5623 (N_5623,N_4238,N_72);
nor U5624 (N_5624,N_1904,N_633);
nand U5625 (N_5625,N_1589,N_682);
nand U5626 (N_5626,N_2826,N_1962);
nor U5627 (N_5627,N_3356,N_1699);
and U5628 (N_5628,N_1241,N_1396);
or U5629 (N_5629,N_3850,N_4250);
nand U5630 (N_5630,N_1119,N_857);
nand U5631 (N_5631,N_2957,N_3612);
nand U5632 (N_5632,N_4473,N_1510);
nand U5633 (N_5633,N_108,N_1574);
or U5634 (N_5634,N_1485,N_2950);
nor U5635 (N_5635,N_2099,N_4556);
or U5636 (N_5636,N_2390,N_1469);
or U5637 (N_5637,N_44,N_1256);
and U5638 (N_5638,N_2570,N_4209);
nor U5639 (N_5639,N_4684,N_2481);
nor U5640 (N_5640,N_524,N_3436);
nand U5641 (N_5641,N_2877,N_1561);
nor U5642 (N_5642,N_599,N_604);
or U5643 (N_5643,N_390,N_1057);
nor U5644 (N_5644,N_1078,N_4674);
and U5645 (N_5645,N_934,N_440);
nor U5646 (N_5646,N_3159,N_211);
nor U5647 (N_5647,N_801,N_4515);
xor U5648 (N_5648,N_75,N_2500);
nor U5649 (N_5649,N_1038,N_3367);
nand U5650 (N_5650,N_3097,N_2505);
or U5651 (N_5651,N_4044,N_292);
nor U5652 (N_5652,N_4533,N_2376);
nand U5653 (N_5653,N_2851,N_3024);
nor U5654 (N_5654,N_2789,N_3653);
and U5655 (N_5655,N_1633,N_1677);
and U5656 (N_5656,N_1816,N_152);
nand U5657 (N_5657,N_4887,N_2363);
nor U5658 (N_5658,N_1918,N_1676);
nor U5659 (N_5659,N_3655,N_1748);
nand U5660 (N_5660,N_3669,N_646);
nand U5661 (N_5661,N_259,N_2535);
and U5662 (N_5662,N_74,N_4807);
nand U5663 (N_5663,N_918,N_4480);
or U5664 (N_5664,N_739,N_4756);
and U5665 (N_5665,N_4868,N_215);
and U5666 (N_5666,N_3393,N_4345);
and U5667 (N_5667,N_2640,N_2553);
nand U5668 (N_5668,N_1428,N_2255);
or U5669 (N_5669,N_817,N_2360);
and U5670 (N_5670,N_52,N_594);
xor U5671 (N_5671,N_1039,N_3051);
or U5672 (N_5672,N_963,N_3);
nand U5673 (N_5673,N_2527,N_2368);
nor U5674 (N_5674,N_2424,N_2154);
or U5675 (N_5675,N_3179,N_3287);
nor U5676 (N_5676,N_2080,N_4846);
nor U5677 (N_5677,N_62,N_2680);
or U5678 (N_5678,N_1320,N_907);
nand U5679 (N_5679,N_2537,N_2614);
nor U5680 (N_5680,N_4047,N_1600);
and U5681 (N_5681,N_2738,N_777);
nor U5682 (N_5682,N_1161,N_158);
nand U5683 (N_5683,N_4291,N_3492);
or U5684 (N_5684,N_3839,N_3522);
xor U5685 (N_5685,N_2476,N_4590);
and U5686 (N_5686,N_1269,N_451);
or U5687 (N_5687,N_2023,N_2978);
and U5688 (N_5688,N_1489,N_165);
and U5689 (N_5689,N_1817,N_2985);
nor U5690 (N_5690,N_1885,N_186);
nand U5691 (N_5691,N_3042,N_1002);
nand U5692 (N_5692,N_1361,N_1006);
and U5693 (N_5693,N_139,N_1825);
nor U5694 (N_5694,N_1926,N_3990);
and U5695 (N_5695,N_1192,N_1105);
nand U5696 (N_5696,N_1357,N_1160);
nor U5697 (N_5697,N_4114,N_2404);
xor U5698 (N_5698,N_4104,N_4666);
nor U5699 (N_5699,N_4040,N_3383);
nand U5700 (N_5700,N_2013,N_4423);
and U5701 (N_5701,N_3644,N_709);
and U5702 (N_5702,N_1626,N_1157);
or U5703 (N_5703,N_3355,N_1319);
and U5704 (N_5704,N_1726,N_3449);
and U5705 (N_5705,N_877,N_3954);
or U5706 (N_5706,N_990,N_3501);
or U5707 (N_5707,N_2725,N_2402);
or U5708 (N_5708,N_2499,N_1640);
nand U5709 (N_5709,N_4039,N_1655);
or U5710 (N_5710,N_3743,N_4202);
nor U5711 (N_5711,N_2715,N_163);
nand U5712 (N_5712,N_80,N_4860);
nor U5713 (N_5713,N_3010,N_3723);
and U5714 (N_5714,N_2296,N_3827);
or U5715 (N_5715,N_1694,N_4660);
xnor U5716 (N_5716,N_1730,N_3666);
and U5717 (N_5717,N_3720,N_2403);
or U5718 (N_5718,N_2996,N_1818);
and U5719 (N_5719,N_2238,N_1875);
nand U5720 (N_5720,N_4813,N_634);
nor U5721 (N_5721,N_2760,N_3625);
or U5722 (N_5722,N_3482,N_1292);
or U5723 (N_5723,N_4030,N_1359);
xor U5724 (N_5724,N_4157,N_2204);
nand U5725 (N_5725,N_3868,N_2379);
nor U5726 (N_5726,N_1133,N_4262);
nand U5727 (N_5727,N_1430,N_3239);
nor U5728 (N_5728,N_3273,N_3489);
nor U5729 (N_5729,N_164,N_1713);
or U5730 (N_5730,N_534,N_229);
nand U5731 (N_5731,N_1936,N_2786);
or U5732 (N_5732,N_4031,N_4917);
and U5733 (N_5733,N_3940,N_3400);
nor U5734 (N_5734,N_3189,N_2334);
nor U5735 (N_5735,N_111,N_1747);
nand U5736 (N_5736,N_2145,N_302);
or U5737 (N_5737,N_4286,N_3619);
nor U5738 (N_5738,N_3831,N_3308);
nor U5739 (N_5739,N_4943,N_1536);
nand U5740 (N_5740,N_3038,N_4486);
nand U5741 (N_5741,N_4618,N_2769);
or U5742 (N_5742,N_3260,N_2868);
nor U5743 (N_5743,N_3816,N_3003);
nor U5744 (N_5744,N_1089,N_4410);
and U5745 (N_5745,N_3943,N_4599);
and U5746 (N_5746,N_2094,N_4419);
or U5747 (N_5747,N_750,N_1293);
and U5748 (N_5748,N_3344,N_675);
nand U5749 (N_5749,N_4260,N_4431);
nor U5750 (N_5750,N_3870,N_1841);
and U5751 (N_5751,N_1001,N_3620);
nand U5752 (N_5752,N_3221,N_434);
nand U5753 (N_5753,N_1291,N_3409);
nand U5754 (N_5754,N_3139,N_1244);
nor U5755 (N_5755,N_1804,N_770);
and U5756 (N_5756,N_909,N_2836);
and U5757 (N_5757,N_2777,N_2744);
nand U5758 (N_5758,N_485,N_2155);
nor U5759 (N_5759,N_3307,N_2798);
and U5760 (N_5760,N_532,N_1577);
nor U5761 (N_5761,N_3552,N_1271);
nor U5762 (N_5762,N_14,N_3873);
or U5763 (N_5763,N_1675,N_1414);
or U5764 (N_5764,N_1806,N_2459);
nand U5765 (N_5765,N_2063,N_4509);
or U5766 (N_5766,N_151,N_4916);
and U5767 (N_5767,N_4927,N_333);
and U5768 (N_5768,N_6,N_4413);
nand U5769 (N_5769,N_4058,N_974);
nand U5770 (N_5770,N_4954,N_4065);
nand U5771 (N_5771,N_3466,N_3519);
and U5772 (N_5772,N_2982,N_3136);
nand U5773 (N_5773,N_1219,N_841);
and U5774 (N_5774,N_2320,N_3382);
and U5775 (N_5775,N_4661,N_4417);
nor U5776 (N_5776,N_137,N_2829);
or U5777 (N_5777,N_232,N_2103);
nor U5778 (N_5778,N_1373,N_4775);
nand U5779 (N_5779,N_797,N_339);
xnor U5780 (N_5780,N_776,N_1242);
or U5781 (N_5781,N_3848,N_905);
nand U5782 (N_5782,N_3023,N_4708);
or U5783 (N_5783,N_291,N_3182);
nor U5784 (N_5784,N_2090,N_1870);
and U5785 (N_5785,N_502,N_4715);
and U5786 (N_5786,N_4667,N_2183);
and U5787 (N_5787,N_3131,N_748);
nand U5788 (N_5788,N_4074,N_1004);
nor U5789 (N_5789,N_4585,N_1471);
or U5790 (N_5790,N_715,N_3878);
nor U5791 (N_5791,N_2669,N_3408);
or U5792 (N_5792,N_2559,N_2194);
nand U5793 (N_5793,N_2750,N_344);
nand U5794 (N_5794,N_4449,N_3922);
nor U5795 (N_5795,N_1374,N_432);
and U5796 (N_5796,N_109,N_3037);
nor U5797 (N_5797,N_3889,N_1227);
and U5798 (N_5798,N_92,N_2761);
or U5799 (N_5799,N_3879,N_135);
nor U5800 (N_5800,N_1229,N_3270);
nand U5801 (N_5801,N_2185,N_2199);
and U5802 (N_5802,N_4323,N_4815);
nand U5803 (N_5803,N_1742,N_2312);
nor U5804 (N_5804,N_4566,N_308);
or U5805 (N_5805,N_4688,N_3923);
nand U5806 (N_5806,N_1049,N_1911);
nor U5807 (N_5807,N_1700,N_387);
or U5808 (N_5808,N_4925,N_1236);
or U5809 (N_5809,N_4698,N_3686);
nor U5810 (N_5810,N_672,N_26);
nor U5811 (N_5811,N_3769,N_2420);
or U5812 (N_5812,N_1421,N_4941);
or U5813 (N_5813,N_2893,N_480);
nor U5814 (N_5814,N_117,N_4992);
nor U5815 (N_5815,N_1743,N_196);
or U5816 (N_5816,N_59,N_891);
or U5817 (N_5817,N_4822,N_1565);
and U5818 (N_5818,N_1941,N_2672);
or U5819 (N_5819,N_2048,N_4615);
and U5820 (N_5820,N_1120,N_4817);
nand U5821 (N_5821,N_1484,N_4406);
and U5822 (N_5822,N_4971,N_3931);
nor U5823 (N_5823,N_3749,N_3592);
nor U5824 (N_5824,N_3867,N_2927);
nand U5825 (N_5825,N_2754,N_1312);
and U5826 (N_5826,N_1976,N_4391);
or U5827 (N_5827,N_2241,N_1368);
and U5828 (N_5828,N_118,N_445);
nor U5829 (N_5829,N_2588,N_4795);
or U5830 (N_5830,N_4218,N_1377);
nand U5831 (N_5831,N_571,N_3703);
and U5832 (N_5832,N_3664,N_1878);
or U5833 (N_5833,N_194,N_1203);
or U5834 (N_5834,N_401,N_2618);
and U5835 (N_5835,N_3549,N_2532);
xor U5836 (N_5836,N_405,N_3738);
and U5837 (N_5837,N_4211,N_617);
and U5838 (N_5838,N_1220,N_1123);
nand U5839 (N_5839,N_1619,N_3550);
and U5840 (N_5840,N_2987,N_3845);
nand U5841 (N_5841,N_1669,N_3760);
nand U5842 (N_5842,N_4240,N_3481);
and U5843 (N_5843,N_4768,N_4152);
nor U5844 (N_5844,N_2446,N_3434);
or U5845 (N_5845,N_309,N_1369);
nand U5846 (N_5846,N_1786,N_3774);
nor U5847 (N_5847,N_3736,N_4945);
xnor U5848 (N_5848,N_996,N_4675);
nor U5849 (N_5849,N_3695,N_3405);
and U5850 (N_5850,N_697,N_4878);
nand U5851 (N_5851,N_1064,N_3811);
or U5852 (N_5852,N_1959,N_2939);
and U5853 (N_5853,N_2700,N_852);
nor U5854 (N_5854,N_248,N_837);
and U5855 (N_5855,N_4792,N_1756);
nand U5856 (N_5856,N_3196,N_2174);
or U5857 (N_5857,N_3193,N_2764);
or U5858 (N_5858,N_4223,N_3311);
nand U5859 (N_5859,N_3290,N_4582);
or U5860 (N_5860,N_4901,N_1393);
and U5861 (N_5861,N_7,N_3232);
or U5862 (N_5862,N_2976,N_4483);
nand U5863 (N_5863,N_1499,N_4389);
or U5864 (N_5864,N_1568,N_3908);
xnor U5865 (N_5865,N_4060,N_4397);
or U5866 (N_5866,N_4914,N_3536);
or U5867 (N_5867,N_3447,N_4664);
xnor U5868 (N_5868,N_1772,N_220);
nand U5869 (N_5869,N_1823,N_2720);
and U5870 (N_5870,N_1807,N_2488);
and U5871 (N_5871,N_1261,N_3776);
xnor U5872 (N_5872,N_1687,N_1880);
and U5873 (N_5873,N_2766,N_1079);
and U5874 (N_5874,N_1854,N_2141);
nand U5875 (N_5875,N_1819,N_1275);
or U5876 (N_5876,N_2351,N_3585);
and U5877 (N_5877,N_2911,N_4307);
and U5878 (N_5878,N_3135,N_1280);
nor U5879 (N_5879,N_1067,N_2125);
xor U5880 (N_5880,N_2084,N_3074);
or U5881 (N_5881,N_1272,N_3740);
or U5882 (N_5882,N_4332,N_988);
or U5883 (N_5883,N_2696,N_3053);
nand U5884 (N_5884,N_3775,N_4100);
nor U5885 (N_5885,N_1500,N_4722);
nor U5886 (N_5886,N_161,N_410);
and U5887 (N_5887,N_105,N_3635);
and U5888 (N_5888,N_574,N_1833);
and U5889 (N_5889,N_289,N_1503);
or U5890 (N_5890,N_4450,N_669);
and U5891 (N_5891,N_4814,N_1155);
or U5892 (N_5892,N_4007,N_3989);
and U5893 (N_5893,N_521,N_4544);
and U5894 (N_5894,N_602,N_4340);
or U5895 (N_5895,N_1738,N_2922);
nor U5896 (N_5896,N_4355,N_1040);
and U5897 (N_5897,N_1883,N_4348);
nor U5898 (N_5898,N_419,N_2799);
nor U5899 (N_5899,N_2358,N_3392);
and U5900 (N_5900,N_4163,N_859);
xor U5901 (N_5901,N_168,N_2191);
nor U5902 (N_5902,N_2438,N_4146);
and U5903 (N_5903,N_3137,N_3440);
nor U5904 (N_5904,N_977,N_77);
or U5905 (N_5905,N_2398,N_601);
nand U5906 (N_5906,N_179,N_49);
xnor U5907 (N_5907,N_1656,N_4203);
and U5908 (N_5908,N_4005,N_4489);
and U5909 (N_5909,N_2384,N_1978);
nor U5910 (N_5910,N_511,N_4789);
xor U5911 (N_5911,N_4837,N_876);
and U5912 (N_5912,N_191,N_1326);
xor U5913 (N_5913,N_242,N_1354);
nand U5914 (N_5914,N_4787,N_1632);
nand U5915 (N_5915,N_4760,N_3173);
nor U5916 (N_5916,N_4964,N_3454);
and U5917 (N_5917,N_1028,N_3310);
or U5918 (N_5918,N_3951,N_2695);
and U5919 (N_5919,N_4257,N_790);
and U5920 (N_5920,N_2731,N_4448);
or U5921 (N_5921,N_4682,N_898);
or U5922 (N_5922,N_583,N_3304);
or U5923 (N_5923,N_693,N_2422);
and U5924 (N_5924,N_4973,N_1805);
and U5925 (N_5925,N_3075,N_1673);
xnor U5926 (N_5926,N_231,N_2357);
and U5927 (N_5927,N_4143,N_4539);
nand U5928 (N_5928,N_2718,N_2322);
nor U5929 (N_5929,N_3089,N_3751);
nor U5930 (N_5930,N_3912,N_2040);
or U5931 (N_5931,N_3572,N_1318);
or U5932 (N_5932,N_1984,N_1135);
or U5933 (N_5933,N_1943,N_4119);
nor U5934 (N_5934,N_3865,N_1025);
and U5935 (N_5935,N_3071,N_1591);
and U5936 (N_5936,N_3757,N_785);
nor U5937 (N_5937,N_4225,N_1752);
or U5938 (N_5938,N_4552,N_2545);
nor U5939 (N_5939,N_2980,N_1148);
and U5940 (N_5940,N_4275,N_1920);
nand U5941 (N_5941,N_1776,N_793);
xor U5942 (N_5942,N_1382,N_3692);
or U5943 (N_5943,N_1734,N_4289);
and U5944 (N_5944,N_2678,N_4493);
nand U5945 (N_5945,N_1988,N_41);
and U5946 (N_5946,N_2200,N_3668);
nor U5947 (N_5947,N_443,N_4626);
nand U5948 (N_5948,N_1544,N_4303);
and U5949 (N_5949,N_66,N_3357);
or U5950 (N_5950,N_1697,N_2902);
nor U5951 (N_5951,N_1925,N_3099);
nand U5952 (N_5952,N_2045,N_659);
nor U5953 (N_5953,N_4863,N_4466);
and U5954 (N_5954,N_4771,N_4650);
nor U5955 (N_5955,N_2430,N_4075);
xor U5956 (N_5956,N_4330,N_1917);
and U5957 (N_5957,N_4965,N_3047);
or U5958 (N_5958,N_4830,N_2917);
nand U5959 (N_5959,N_3642,N_960);
or U5960 (N_5960,N_1915,N_1731);
and U5961 (N_5961,N_3515,N_1955);
or U5962 (N_5962,N_3826,N_4091);
nand U5963 (N_5963,N_3970,N_328);
and U5964 (N_5964,N_145,N_2697);
nor U5965 (N_5965,N_922,N_2152);
nand U5966 (N_5966,N_1835,N_2937);
nor U5967 (N_5967,N_937,N_547);
or U5968 (N_5968,N_3420,N_4588);
nand U5969 (N_5969,N_3318,N_2001);
and U5970 (N_5970,N_4386,N_2110);
xnor U5971 (N_5971,N_3609,N_4705);
and U5972 (N_5972,N_4110,N_613);
nor U5973 (N_5973,N_3072,N_3584);
and U5974 (N_5974,N_4968,N_1979);
xor U5975 (N_5975,N_4249,N_4452);
nor U5976 (N_5976,N_1386,N_552);
nand U5977 (N_5977,N_1706,N_1149);
xor U5978 (N_5978,N_912,N_4499);
or U5979 (N_5979,N_755,N_3403);
nor U5980 (N_5980,N_3004,N_89);
nor U5981 (N_5981,N_3528,N_926);
nand U5982 (N_5982,N_1863,N_3143);
nor U5983 (N_5983,N_4414,N_4468);
nand U5984 (N_5984,N_4694,N_1163);
xor U5985 (N_5985,N_4246,N_2413);
nand U5986 (N_5986,N_628,N_1215);
nand U5987 (N_5987,N_2747,N_2316);
and U5988 (N_5988,N_766,N_2042);
nand U5989 (N_5989,N_1935,N_4407);
nand U5990 (N_5990,N_1846,N_1247);
nor U5991 (N_5991,N_1755,N_4519);
and U5992 (N_5992,N_2975,N_3388);
nand U5993 (N_5993,N_775,N_3787);
or U5994 (N_5994,N_4208,N_4435);
nand U5995 (N_5995,N_3439,N_4874);
and U5996 (N_5996,N_1961,N_3571);
xnor U5997 (N_5997,N_736,N_1413);
and U5998 (N_5998,N_1380,N_3930);
xnor U5999 (N_5999,N_228,N_1963);
or U6000 (N_6000,N_995,N_4032);
nor U6001 (N_6001,N_2335,N_498);
nor U6002 (N_6002,N_1487,N_1551);
and U6003 (N_6003,N_3226,N_246);
or U6004 (N_6004,N_4463,N_3219);
and U6005 (N_6005,N_3634,N_1716);
nor U6006 (N_6006,N_2755,N_4061);
nand U6007 (N_6007,N_4671,N_2600);
nand U6008 (N_6008,N_2955,N_3822);
and U6009 (N_6009,N_1331,N_4919);
or U6010 (N_6010,N_1838,N_887);
or U6011 (N_6011,N_2246,N_4046);
nand U6012 (N_6012,N_2666,N_1631);
nand U6013 (N_6013,N_1524,N_4611);
and U6014 (N_6014,N_2872,N_2960);
nor U6015 (N_6015,N_3435,N_337);
nor U6016 (N_6016,N_195,N_2947);
nor U6017 (N_6017,N_2721,N_177);
and U6018 (N_6018,N_3852,N_13);
nor U6019 (N_6019,N_3662,N_3761);
nand U6020 (N_6020,N_3698,N_4182);
nor U6021 (N_6021,N_4206,N_244);
and U6022 (N_6022,N_3484,N_4412);
and U6023 (N_6023,N_1992,N_2153);
nor U6024 (N_6024,N_4224,N_3511);
xor U6025 (N_6025,N_3216,N_2447);
nor U6026 (N_6026,N_1513,N_4749);
xor U6027 (N_6027,N_719,N_1378);
nor U6028 (N_6028,N_1366,N_2391);
or U6029 (N_6029,N_2589,N_1296);
or U6030 (N_6030,N_621,N_297);
nor U6031 (N_6031,N_1690,N_1996);
nor U6032 (N_6032,N_4139,N_4957);
xnor U6033 (N_6033,N_3741,N_4991);
nor U6034 (N_6034,N_226,N_2210);
or U6035 (N_6035,N_1048,N_4056);
nand U6036 (N_6036,N_4034,N_4151);
nand U6037 (N_6037,N_2118,N_4922);
nor U6038 (N_6038,N_2389,N_1110);
xor U6039 (N_6039,N_1441,N_4336);
nor U6040 (N_6040,N_4707,N_1358);
nand U6041 (N_6041,N_1872,N_2522);
or U6042 (N_6042,N_4270,N_4563);
nand U6043 (N_6043,N_4940,N_1375);
and U6044 (N_6044,N_2838,N_1196);
nand U6045 (N_6045,N_1310,N_584);
nand U6046 (N_6046,N_4458,N_1246);
or U6047 (N_6047,N_3589,N_2416);
and U6048 (N_6048,N_1117,N_1952);
nand U6049 (N_6049,N_1492,N_1228);
nand U6050 (N_6050,N_4233,N_924);
and U6051 (N_6051,N_2310,N_4536);
nor U6052 (N_6052,N_1719,N_180);
nor U6053 (N_6053,N_3748,N_3282);
or U6054 (N_6054,N_2354,N_844);
nand U6055 (N_6055,N_931,N_1460);
nand U6056 (N_6056,N_545,N_1351);
xnor U6057 (N_6057,N_3114,N_1545);
and U6058 (N_6058,N_3818,N_2576);
xnor U6059 (N_6059,N_3744,N_2712);
and U6060 (N_6060,N_4653,N_1168);
nor U6061 (N_6061,N_722,N_1065);
nor U6062 (N_6062,N_1781,N_688);
nor U6063 (N_6063,N_2751,N_3901);
or U6064 (N_6064,N_3407,N_4140);
nand U6065 (N_6065,N_1757,N_3238);
nand U6066 (N_6066,N_2030,N_1527);
nor U6067 (N_6067,N_3030,N_3166);
and U6068 (N_6068,N_2969,N_1391);
or U6069 (N_6069,N_3224,N_4366);
xnor U6070 (N_6070,N_4230,N_1184);
nand U6071 (N_6071,N_3254,N_1353);
nand U6072 (N_6072,N_842,N_3328);
xnor U6073 (N_6073,N_3019,N_717);
or U6074 (N_6074,N_10,N_3128);
or U6075 (N_6075,N_839,N_553);
nand U6076 (N_6076,N_3338,N_2791);
nand U6077 (N_6077,N_2243,N_2039);
and U6078 (N_6078,N_1784,N_1297);
nand U6079 (N_6079,N_3980,N_1142);
and U6080 (N_6080,N_1641,N_3504);
or U6081 (N_6081,N_3469,N_746);
nor U6082 (N_6082,N_1147,N_2906);
or U6083 (N_6083,N_2585,N_655);
and U6084 (N_6084,N_2299,N_3281);
nor U6085 (N_6085,N_4416,N_2069);
nor U6086 (N_6086,N_1134,N_3085);
or U6087 (N_6087,N_2298,N_3502);
and U6088 (N_6088,N_3766,N_2602);
nor U6089 (N_6089,N_1061,N_1199);
nand U6090 (N_6090,N_1611,N_3018);
nor U6091 (N_6091,N_4312,N_3360);
and U6092 (N_6092,N_1177,N_2235);
xnor U6093 (N_6093,N_2329,N_4796);
or U6094 (N_6094,N_335,N_3843);
or U6095 (N_6095,N_4062,N_3798);
nor U6096 (N_6096,N_420,N_2201);
nor U6097 (N_6097,N_4864,N_2339);
and U6098 (N_6098,N_2274,N_216);
xnor U6099 (N_6099,N_263,N_4862);
nand U6100 (N_6100,N_869,N_4931);
or U6101 (N_6101,N_3082,N_3887);
nand U6102 (N_6102,N_611,N_4426);
or U6103 (N_6103,N_4456,N_2418);
nand U6104 (N_6104,N_4780,N_596);
nor U6105 (N_6105,N_649,N_2635);
and U6106 (N_6106,N_4621,N_3525);
nor U6107 (N_6107,N_42,N_4226);
nor U6108 (N_6108,N_3057,N_2644);
nor U6109 (N_6109,N_3902,N_3952);
and U6110 (N_6110,N_1136,N_1063);
or U6111 (N_6111,N_1474,N_4073);
or U6112 (N_6112,N_733,N_477);
or U6113 (N_6113,N_3505,N_740);
and U6114 (N_6114,N_4640,N_225);
nor U6115 (N_6115,N_2722,N_590);
xor U6116 (N_6116,N_1884,N_2292);
nor U6117 (N_6117,N_1867,N_2055);
or U6118 (N_6118,N_2634,N_3474);
nand U6119 (N_6119,N_1530,N_2561);
nor U6120 (N_6120,N_4036,N_2867);
and U6121 (N_6121,N_1324,N_1638);
nor U6122 (N_6122,N_1041,N_1607);
or U6123 (N_6123,N_3605,N_2102);
and U6124 (N_6124,N_4357,N_1277);
nor U6125 (N_6125,N_3939,N_1468);
nor U6126 (N_6126,N_3932,N_1130);
nand U6127 (N_6127,N_3613,N_3286);
nand U6128 (N_6128,N_2008,N_4959);
or U6129 (N_6129,N_2690,N_3996);
nand U6130 (N_6130,N_4548,N_4437);
nor U6131 (N_6131,N_3674,N_2136);
nor U6132 (N_6132,N_3756,N_141);
xor U6133 (N_6133,N_4532,N_2442);
nor U6134 (N_6134,N_3858,N_2935);
and U6135 (N_6135,N_3963,N_36);
nand U6136 (N_6136,N_3263,N_3846);
and U6137 (N_6137,N_1654,N_306);
xor U6138 (N_6138,N_1498,N_2861);
nand U6139 (N_6139,N_4763,N_2361);
or U6140 (N_6140,N_4686,N_1770);
xor U6141 (N_6141,N_4999,N_548);
or U6142 (N_6142,N_1283,N_489);
nor U6143 (N_6143,N_3279,N_1912);
and U6144 (N_6144,N_3861,N_2519);
nand U6145 (N_6145,N_150,N_4481);
and U6146 (N_6146,N_3411,N_2095);
and U6147 (N_6147,N_832,N_928);
or U6148 (N_6148,N_3546,N_2854);
xnor U6149 (N_6149,N_725,N_783);
nor U6150 (N_6150,N_1836,N_3303);
or U6151 (N_6151,N_2645,N_2759);
xnor U6152 (N_6152,N_4487,N_2686);
nor U6153 (N_6153,N_1821,N_1127);
or U6154 (N_6154,N_3350,N_4338);
or U6155 (N_6155,N_1126,N_250);
and U6156 (N_6156,N_2676,N_4809);
and U6157 (N_6157,N_1449,N_2702);
xnor U6158 (N_6158,N_4026,N_2856);
xnor U6159 (N_6159,N_3918,N_4432);
and U6160 (N_6160,N_2258,N_3754);
or U6161 (N_6161,N_1223,N_4274);
nor U6162 (N_6162,N_3547,N_2583);
xnor U6163 (N_6163,N_3789,N_4052);
or U6164 (N_6164,N_1209,N_3353);
and U6165 (N_6165,N_1423,N_316);
nand U6166 (N_6166,N_4654,N_132);
nor U6167 (N_6167,N_3418,N_4823);
or U6168 (N_6168,N_771,N_4411);
or U6169 (N_6169,N_3976,N_4302);
nor U6170 (N_6170,N_2529,N_769);
or U6171 (N_6171,N_4876,N_1124);
or U6172 (N_6172,N_2632,N_2612);
or U6173 (N_6173,N_531,N_4108);
nand U6174 (N_6174,N_93,N_283);
or U6175 (N_6175,N_4141,N_2903);
nor U6176 (N_6176,N_2973,N_2984);
or U6177 (N_6177,N_2096,N_2620);
or U6178 (N_6178,N_2364,N_3767);
nor U6179 (N_6179,N_2884,N_3054);
nor U6180 (N_6180,N_1439,N_3864);
and U6181 (N_6181,N_2555,N_4673);
nand U6182 (N_6182,N_4057,N_1506);
and U6183 (N_6183,N_1239,N_3002);
or U6184 (N_6184,N_2687,N_1909);
or U6185 (N_6185,N_201,N_3115);
xor U6186 (N_6186,N_4639,N_1125);
and U6187 (N_6187,N_2888,N_2343);
nor U6188 (N_6188,N_73,N_631);
xor U6189 (N_6189,N_3840,N_3622);
nand U6190 (N_6190,N_707,N_4729);
nor U6191 (N_6191,N_692,N_4241);
xor U6192 (N_6192,N_4022,N_2371);
xnor U6193 (N_6193,N_3445,N_2198);
or U6194 (N_6194,N_2015,N_1647);
nor U6195 (N_6195,N_606,N_4614);
xnor U6196 (N_6196,N_476,N_2684);
and U6197 (N_6197,N_3322,N_1843);
nor U6198 (N_6198,N_3331,N_3925);
and U6199 (N_6199,N_710,N_2507);
or U6200 (N_6200,N_2780,N_636);
or U6201 (N_6201,N_3782,N_3541);
nand U6202 (N_6202,N_4679,N_2660);
or U6203 (N_6203,N_3903,N_1059);
nand U6204 (N_6204,N_2050,N_1009);
and U6205 (N_6205,N_1967,N_2150);
and U6206 (N_6206,N_2436,N_2057);
nor U6207 (N_6207,N_2458,N_567);
and U6208 (N_6208,N_1728,N_2127);
xor U6209 (N_6209,N_1068,N_1516);
xnor U6210 (N_6210,N_3994,N_4546);
nand U6211 (N_6211,N_3222,N_4113);
nand U6212 (N_6212,N_2502,N_1285);
nor U6213 (N_6213,N_4343,N_3746);
or U6214 (N_6214,N_791,N_1329);
or U6215 (N_6215,N_3508,N_352);
and U6216 (N_6216,N_4827,N_1851);
nor U6217 (N_6217,N_1571,N_1017);
nor U6218 (N_6218,N_685,N_1858);
and U6219 (N_6219,N_4285,N_299);
or U6220 (N_6220,N_3632,N_3368);
or U6221 (N_6221,N_651,N_281);
or U6222 (N_6222,N_1629,N_3299);
nor U6223 (N_6223,N_1086,N_3298);
and U6224 (N_6224,N_2037,N_4469);
nand U6225 (N_6225,N_1586,N_3520);
and U6226 (N_6226,N_4857,N_4580);
nand U6227 (N_6227,N_102,N_1179);
nand U6228 (N_6228,N_3705,N_2336);
nor U6229 (N_6229,N_3100,N_3735);
and U6230 (N_6230,N_2992,N_1399);
nor U6231 (N_6231,N_1708,N_4328);
and U6232 (N_6232,N_2518,N_3762);
or U6233 (N_6233,N_1968,N_3558);
nand U6234 (N_6234,N_2997,N_1861);
nand U6235 (N_6235,N_3860,N_1131);
nor U6236 (N_6236,N_3794,N_2554);
or U6237 (N_6237,N_3302,N_4676);
nand U6238 (N_6238,N_4928,N_1652);
nand U6239 (N_6239,N_2795,N_4554);
or U6240 (N_6240,N_619,N_4165);
nor U6241 (N_6241,N_1595,N_4902);
or U6242 (N_6242,N_4803,N_4111);
or U6243 (N_6243,N_4738,N_4603);
nor U6244 (N_6244,N_4210,N_3140);
nand U6245 (N_6245,N_4989,N_4958);
xnor U6246 (N_6246,N_1031,N_1994);
nand U6247 (N_6247,N_147,N_268);
and U6248 (N_6248,N_3293,N_2122);
nand U6249 (N_6249,N_3337,N_2208);
nor U6250 (N_6250,N_4960,N_1554);
and U6251 (N_6251,N_3069,N_264);
or U6252 (N_6252,N_3529,N_4083);
nand U6253 (N_6253,N_90,N_4816);
nand U6254 (N_6254,N_3855,N_4199);
xnor U6255 (N_6255,N_2304,N_1486);
nand U6256 (N_6256,N_3485,N_721);
nand U6257 (N_6257,N_2556,N_1658);
and U6258 (N_6258,N_4276,N_1263);
nor U6259 (N_6259,N_2450,N_1964);
or U6260 (N_6260,N_1634,N_1302);
or U6261 (N_6261,N_858,N_3441);
nand U6262 (N_6262,N_395,N_743);
or U6263 (N_6263,N_3225,N_1021);
nor U6264 (N_6264,N_570,N_1596);
nand U6265 (N_6265,N_1337,N_2162);
or U6266 (N_6266,N_2355,N_4003);
nand U6267 (N_6267,N_3227,N_415);
and U6268 (N_6268,N_1727,N_3565);
and U6269 (N_6269,N_4442,N_1392);
and U6270 (N_6270,N_2129,N_751);
xnor U6271 (N_6271,N_300,N_4212);
nand U6272 (N_6272,N_2796,N_2736);
nor U6273 (N_6273,N_2018,N_325);
or U6274 (N_6274,N_2192,N_3883);
xor U6275 (N_6275,N_1238,N_1709);
nor U6276 (N_6276,N_4550,N_70);
or U6277 (N_6277,N_2236,N_4072);
or U6278 (N_6278,N_3406,N_644);
nor U6279 (N_6279,N_4424,N_1975);
or U6280 (N_6280,N_1934,N_3444);
or U6281 (N_6281,N_4898,N_479);
or U6282 (N_6282,N_2301,N_3247);
or U6283 (N_6283,N_2106,N_2067);
xnor U6284 (N_6284,N_3035,N_2477);
nand U6285 (N_6285,N_2569,N_1763);
nand U6286 (N_6286,N_1519,N_478);
and U6287 (N_6287,N_3516,N_3646);
nand U6288 (N_6288,N_1511,N_366);
nor U6289 (N_6289,N_4244,N_916);
xor U6290 (N_6290,N_2108,N_4586);
and U6291 (N_6291,N_2560,N_3817);
xnor U6292 (N_6292,N_2268,N_3459);
xnor U6293 (N_6293,N_4351,N_3545);
and U6294 (N_6294,N_4418,N_3094);
nand U6295 (N_6295,N_3417,N_1623);
nor U6296 (N_6296,N_2932,N_3681);
xor U6297 (N_6297,N_3828,N_620);
nor U6298 (N_6298,N_4657,N_3458);
xor U6299 (N_6299,N_122,N_4994);
nand U6300 (N_6300,N_1620,N_3394);
nand U6301 (N_6301,N_187,N_704);
nor U6302 (N_6302,N_1143,N_2180);
nor U6303 (N_6303,N_1081,N_1791);
or U6304 (N_6304,N_3490,N_3278);
or U6305 (N_6305,N_720,N_1030);
and U6306 (N_6306,N_3601,N_2423);
and U6307 (N_6307,N_4453,N_2966);
nor U6308 (N_6308,N_661,N_4192);
or U6309 (N_6309,N_1645,N_2251);
nand U6310 (N_6310,N_4184,N_930);
xor U6311 (N_6311,N_493,N_564);
or U6312 (N_6312,N_2989,N_2723);
and U6313 (N_6313,N_3195,N_3633);
nand U6314 (N_6314,N_3347,N_3857);
xnor U6315 (N_6315,N_4069,N_4537);
xnor U6316 (N_6316,N_1557,N_1642);
nand U6317 (N_6317,N_4053,N_778);
nand U6318 (N_6318,N_1000,N_1027);
nand U6319 (N_6319,N_2898,N_3453);
or U6320 (N_6320,N_700,N_1573);
and U6321 (N_6321,N_286,N_377);
xnor U6322 (N_6322,N_686,N_464);
or U6323 (N_6323,N_2590,N_519);
and U6324 (N_6324,N_2848,N_848);
and U6325 (N_6325,N_2471,N_310);
xnor U6326 (N_6326,N_3629,N_4555);
nand U6327 (N_6327,N_3803,N_4512);
and U6328 (N_6328,N_3032,N_2609);
nor U6329 (N_6329,N_2075,N_3291);
xor U6330 (N_6330,N_2128,N_481);
xor U6331 (N_6331,N_2311,N_2009);
nor U6332 (N_6332,N_1761,N_104);
nor U6333 (N_6333,N_683,N_3313);
nor U6334 (N_6334,N_96,N_3568);
or U6335 (N_6335,N_2302,N_4910);
or U6336 (N_6336,N_88,N_3396);
and U6337 (N_6337,N_608,N_222);
or U6338 (N_6338,N_703,N_664);
nand U6339 (N_6339,N_3888,N_3824);
nand U6340 (N_6340,N_2281,N_2378);
and U6341 (N_6341,N_3981,N_1740);
nor U6342 (N_6342,N_2058,N_223);
and U6343 (N_6343,N_1187,N_558);
nor U6344 (N_6344,N_4390,N_544);
nor U6345 (N_6345,N_1008,N_2491);
or U6346 (N_6346,N_1303,N_629);
or U6347 (N_6347,N_3111,N_843);
and U6348 (N_6348,N_3710,N_2031);
or U6349 (N_6349,N_3500,N_175);
or U6350 (N_6350,N_781,N_1417);
and U6351 (N_6351,N_1402,N_2874);
nor U6352 (N_6352,N_2876,N_4071);
and U6353 (N_6353,N_1811,N_3473);
nand U6354 (N_6354,N_814,N_3684);
nor U6355 (N_6355,N_423,N_3667);
or U6356 (N_6356,N_4918,N_1856);
and U6357 (N_6357,N_4464,N_3233);
or U6358 (N_6358,N_18,N_1993);
nand U6359 (N_6359,N_2131,N_4095);
nor U6360 (N_6360,N_3708,N_467);
and U6361 (N_6361,N_4354,N_2866);
nor U6362 (N_6362,N_4188,N_2580);
nand U6363 (N_6363,N_4178,N_4651);
and U6364 (N_6364,N_3825,N_3911);
or U6365 (N_6365,N_3451,N_2033);
and U6366 (N_6366,N_4377,N_565);
and U6367 (N_6367,N_3745,N_2923);
or U6368 (N_6368,N_1093,N_3993);
nor U6369 (N_6369,N_3928,N_3885);
or U6370 (N_6370,N_3361,N_2785);
and U6371 (N_6371,N_2121,N_425);
or U6372 (N_6372,N_4852,N_128);
or U6373 (N_6373,N_4948,N_3699);
xor U6374 (N_6374,N_4273,N_849);
nand U6375 (N_6375,N_2709,N_2613);
nor U6376 (N_6376,N_1670,N_4812);
nand U6377 (N_6377,N_2443,N_3476);
and U6378 (N_6378,N_3414,N_4385);
or U6379 (N_6379,N_4191,N_1281);
nor U6380 (N_6380,N_1891,N_2551);
or U6381 (N_6381,N_2710,N_4829);
and U6382 (N_6382,N_3936,N_2078);
nand U6383 (N_6383,N_2603,N_2526);
nand U6384 (N_6384,N_2052,N_3289);
nor U6385 (N_6385,N_4765,N_2406);
or U6386 (N_6386,N_2504,N_2812);
or U6387 (N_6387,N_2993,N_1800);
and U6388 (N_6388,N_3711,N_4023);
nor U6389 (N_6389,N_1754,N_2249);
or U6390 (N_6390,N_3101,N_2739);
or U6391 (N_6391,N_1011,N_2756);
nor U6392 (N_6392,N_3806,N_563);
nand U6393 (N_6393,N_4772,N_2294);
nand U6394 (N_6394,N_1844,N_3108);
nand U6395 (N_6395,N_3243,N_362);
nand U6396 (N_6396,N_3788,N_3896);
nor U6397 (N_6397,N_4035,N_2005);
and U6398 (N_6398,N_3962,N_1859);
nor U6399 (N_6399,N_2330,N_3716);
and U6400 (N_6400,N_113,N_1200);
nor U6401 (N_6401,N_452,N_803);
and U6402 (N_6402,N_760,N_4445);
and U6403 (N_6403,N_2217,N_2638);
and U6404 (N_6404,N_3000,N_2936);
or U6405 (N_6405,N_4764,N_1902);
or U6406 (N_6406,N_3569,N_749);
nand U6407 (N_6407,N_1928,N_278);
or U6408 (N_6408,N_1949,N_2074);
nand U6409 (N_6409,N_3321,N_4595);
xnor U6410 (N_6410,N_3213,N_4079);
nor U6411 (N_6411,N_3701,N_458);
nand U6412 (N_6412,N_3121,N_4467);
or U6413 (N_6413,N_3771,N_1749);
or U6414 (N_6414,N_2245,N_3013);
or U6415 (N_6415,N_1750,N_728);
and U6416 (N_6416,N_3467,N_2622);
or U6417 (N_6417,N_668,N_2916);
nand U6418 (N_6418,N_3919,N_3938);
xor U6419 (N_6419,N_1774,N_2862);
or U6420 (N_6420,N_3348,N_2986);
nand U6421 (N_6421,N_1737,N_1705);
nand U6422 (N_6422,N_4504,N_2824);
and U6423 (N_6423,N_2837,N_3926);
nor U6424 (N_6424,N_2027,N_1322);
and U6425 (N_6425,N_632,N_2503);
nand U6426 (N_6426,N_4723,N_466);
or U6427 (N_6427,N_4963,N_4985);
and U6428 (N_6428,N_2465,N_4335);
nor U6429 (N_6429,N_1347,N_2891);
and U6430 (N_6430,N_1956,N_417);
nand U6431 (N_6431,N_3432,N_1933);
nand U6432 (N_6432,N_1684,N_4319);
and U6433 (N_6433,N_4255,N_2860);
and U6434 (N_6434,N_3365,N_252);
nor U6435 (N_6435,N_28,N_1315);
nor U6436 (N_6436,N_3834,N_46);
nand U6437 (N_6437,N_4872,N_522);
xor U6438 (N_6438,N_1250,N_1608);
or U6439 (N_6439,N_874,N_1431);
and U6440 (N_6440,N_3041,N_855);
nor U6441 (N_6441,N_1931,N_4356);
nor U6442 (N_6442,N_315,N_3582);
or U6443 (N_6443,N_4433,N_1208);
nand U6444 (N_6444,N_4855,N_4266);
or U6445 (N_6445,N_2719,N_1152);
or U6446 (N_6446,N_585,N_4490);
and U6447 (N_6447,N_4154,N_1074);
and U6448 (N_6448,N_4479,N_4320);
nor U6449 (N_6449,N_2035,N_1278);
nor U6450 (N_6450,N_2319,N_3618);
nand U6451 (N_6451,N_3523,N_1983);
nor U6452 (N_6452,N_2493,N_2954);
xnor U6453 (N_6453,N_396,N_1768);
nor U6454 (N_6454,N_4635,N_4066);
or U6455 (N_6455,N_3230,N_3807);
nand U6456 (N_6456,N_3983,N_391);
nand U6457 (N_6457,N_3208,N_2341);
nor U6458 (N_6458,N_2107,N_3947);
nor U6459 (N_6459,N_2581,N_3150);
and U6460 (N_6460,N_723,N_2593);
xnor U6461 (N_6461,N_1622,N_276);
nor U6462 (N_6462,N_4844,N_2290);
nor U6463 (N_6463,N_4678,N_238);
or U6464 (N_6464,N_3237,N_936);
and U6465 (N_6465,N_120,N_4068);
and U6466 (N_6466,N_3258,N_1852);
or U6467 (N_6467,N_4043,N_4380);
or U6468 (N_6468,N_3805,N_812);
and U6469 (N_6469,N_4785,N_2381);
xnor U6470 (N_6470,N_2392,N_523);
nand U6471 (N_6471,N_375,N_181);
and U6472 (N_6472,N_63,N_2784);
and U6473 (N_6473,N_2776,N_4308);
and U6474 (N_6474,N_3581,N_4623);
nand U6475 (N_6475,N_919,N_4086);
or U6476 (N_6476,N_4790,N_2714);
nand U6477 (N_6477,N_1253,N_3763);
nand U6478 (N_6478,N_154,N_3274);
or U6479 (N_6479,N_2374,N_4921);
or U6480 (N_6480,N_1405,N_2508);
nor U6481 (N_6481,N_3830,N_2887);
nor U6482 (N_6482,N_3231,N_3374);
nor U6483 (N_6483,N_3320,N_4750);
nand U6484 (N_6484,N_4617,N_4277);
nand U6485 (N_6485,N_3419,N_4836);
and U6486 (N_6486,N_3663,N_982);
nand U6487 (N_6487,N_1169,N_1651);
or U6488 (N_6488,N_4568,N_121);
nand U6489 (N_6489,N_2661,N_4367);
or U6490 (N_6490,N_4236,N_4735);
nand U6491 (N_6491,N_2628,N_4087);
xor U6492 (N_6492,N_4253,N_4441);
or U6493 (N_6493,N_3647,N_773);
or U6494 (N_6494,N_3829,N_1535);
and U6495 (N_6495,N_2405,N_3056);
nand U6496 (N_6496,N_2647,N_3465);
nor U6497 (N_6497,N_3044,N_3153);
nor U6498 (N_6498,N_1809,N_1689);
nand U6499 (N_6499,N_1569,N_2533);
and U6500 (N_6500,N_3463,N_1434);
and U6501 (N_6501,N_4322,N_2578);
xor U6502 (N_6502,N_872,N_1104);
xor U6503 (N_6503,N_4341,N_1855);
nor U6504 (N_6504,N_4826,N_1803);
nand U6505 (N_6505,N_2170,N_2315);
nand U6506 (N_6506,N_4166,N_3942);
nand U6507 (N_6507,N_2758,N_1733);
or U6508 (N_6508,N_2983,N_618);
or U6509 (N_6509,N_3413,N_473);
nand U6510 (N_6510,N_3241,N_4256);
and U6511 (N_6511,N_1692,N_2563);
nor U6512 (N_6512,N_761,N_1564);
or U6513 (N_6513,N_4033,N_269);
xnor U6514 (N_6514,N_2333,N_2749);
nor U6515 (N_6515,N_4471,N_322);
nand U6516 (N_6516,N_4126,N_758);
and U6517 (N_6517,N_1908,N_3574);
and U6518 (N_6518,N_3362,N_911);
or U6519 (N_6519,N_1778,N_562);
nor U6520 (N_6520,N_4315,N_2451);
nand U6521 (N_6521,N_3491,N_4747);
or U6522 (N_6522,N_3603,N_408);
and U6523 (N_6523,N_3090,N_406);
nand U6524 (N_6524,N_4261,N_393);
nor U6525 (N_6525,N_3530,N_2223);
nor U6526 (N_6526,N_3183,N_3507);
or U6527 (N_6527,N_2988,N_103);
and U6528 (N_6528,N_4082,N_2213);
nor U6529 (N_6529,N_862,N_4602);
nand U6530 (N_6530,N_1230,N_3610);
or U6531 (N_6531,N_2961,N_3917);
nor U6532 (N_6532,N_2306,N_779);
and U6533 (N_6533,N_4287,N_2514);
nor U6534 (N_6534,N_4197,N_4662);
nand U6535 (N_6535,N_4405,N_2534);
and U6536 (N_6536,N_3292,N_2428);
nor U6537 (N_6537,N_3941,N_3351);
or U6538 (N_6538,N_3191,N_1695);
nand U6539 (N_6539,N_3866,N_4180);
and U6540 (N_6540,N_884,N_4400);
and U6541 (N_6541,N_4981,N_503);
and U6542 (N_6542,N_3218,N_273);
nand U6543 (N_6543,N_3161,N_143);
nor U6544 (N_6544,N_1381,N_3124);
or U6545 (N_6545,N_209,N_2148);
and U6546 (N_6546,N_587,N_763);
or U6547 (N_6547,N_4447,N_2970);
xnor U6548 (N_6548,N_1479,N_904);
and U6549 (N_6549,N_200,N_4847);
nand U6550 (N_6550,N_4028,N_968);
or U6551 (N_6551,N_875,N_172);
nor U6552 (N_6552,N_4403,N_3799);
xor U6553 (N_6553,N_372,N_2467);
nor U6554 (N_6554,N_2548,N_1703);
or U6555 (N_6555,N_4808,N_970);
xor U6556 (N_6556,N_556,N_3206);
xnor U6557 (N_6557,N_3682,N_2531);
nor U6558 (N_6558,N_2835,N_4394);
nand U6559 (N_6559,N_819,N_1389);
or U6560 (N_6560,N_1023,N_3790);
or U6561 (N_6561,N_1345,N_2345);
nor U6562 (N_6562,N_1543,N_2346);
or U6563 (N_6563,N_3387,N_2133);
nor U6564 (N_6564,N_3497,N_2237);
nor U6565 (N_6565,N_4734,N_1980);
or U6566 (N_6566,N_2264,N_1842);
xor U6567 (N_6567,N_3729,N_4881);
and U6568 (N_6568,N_1060,N_1249);
or U6569 (N_6569,N_407,N_1679);
and U6570 (N_6570,N_3315,N_3426);
or U6571 (N_6571,N_4342,N_695);
or U6572 (N_6572,N_2088,N_4896);
nor U6573 (N_6573,N_4013,N_4477);
and U6574 (N_6574,N_442,N_1789);
nand U6575 (N_6575,N_4581,N_2617);
xor U6576 (N_6576,N_4561,N_1661);
and U6577 (N_6577,N_2729,N_3371);
or U6578 (N_6578,N_4150,N_2664);
or U6579 (N_6579,N_1231,N_2873);
xor U6580 (N_6580,N_4527,N_2151);
nor U6581 (N_6581,N_1837,N_4883);
nand U6582 (N_6582,N_2833,N_1151);
nor U6583 (N_6583,N_471,N_2038);
and U6584 (N_6584,N_4717,N_983);
or U6585 (N_6585,N_4668,N_3815);
nand U6586 (N_6586,N_2289,N_942);
or U6587 (N_6587,N_3810,N_2195);
nand U6588 (N_6588,N_714,N_3487);
nor U6589 (N_6589,N_3155,N_809);
or U6590 (N_6590,N_4782,N_2667);
or U6591 (N_6591,N_831,N_2190);
nor U6592 (N_6592,N_4001,N_1522);
and U6593 (N_6593,N_1773,N_3641);
and U6594 (N_6594,N_4627,N_2571);
and U6595 (N_6595,N_1758,N_4587);
nor U6596 (N_6596,N_4762,N_3649);
or U6597 (N_6597,N_1409,N_525);
nand U6598 (N_6598,N_240,N_4806);
nor U6599 (N_6599,N_2566,N_2313);
nor U6600 (N_6600,N_2234,N_50);
and U6601 (N_6601,N_759,N_2778);
nand U6602 (N_6602,N_698,N_635);
nor U6603 (N_6603,N_31,N_1333);
or U6604 (N_6604,N_4892,N_4451);
and U6605 (N_6605,N_800,N_4687);
nor U6606 (N_6606,N_1094,N_3562);
nor U6607 (N_6607,N_3608,N_2254);
xor U6608 (N_6608,N_3425,N_4012);
nand U6609 (N_6609,N_4247,N_3907);
xor U6610 (N_6610,N_2698,N_4545);
or U6611 (N_6611,N_3076,N_1834);
nand U6612 (N_6612,N_3160,N_2601);
and U6613 (N_6613,N_3058,N_1410);
and U6614 (N_6614,N_2523,N_1566);
or U6615 (N_6615,N_2656,N_2433);
nand U6616 (N_6616,N_4727,N_3758);
nor U6617 (N_6617,N_1144,N_1070);
and U6618 (N_6618,N_4292,N_997);
nand U6619 (N_6619,N_1234,N_3553);
nand U6620 (N_6620,N_1412,N_3856);
and U6621 (N_6621,N_3186,N_1109);
xnor U6622 (N_6622,N_2273,N_1653);
and U6623 (N_6623,N_2890,N_1547);
nor U6624 (N_6624,N_3957,N_3784);
and U6625 (N_6625,N_303,N_3548);
and U6626 (N_6626,N_3267,N_355);
and U6627 (N_6627,N_3510,N_2946);
xor U6628 (N_6628,N_1946,N_2840);
nor U6629 (N_6629,N_3542,N_193);
nor U6630 (N_6630,N_2449,N_3721);
nand U6631 (N_6631,N_735,N_3945);
nor U6632 (N_6632,N_1115,N_2394);
nor U6633 (N_6633,N_1383,N_4870);
or U6634 (N_6634,N_1668,N_4641);
xor U6635 (N_6635,N_3039,N_4866);
nor U6636 (N_6636,N_1235,N_2435);
or U6637 (N_6637,N_3098,N_3154);
nand U6638 (N_6638,N_4465,N_4427);
nand U6639 (N_6639,N_3271,N_1793);
xor U6640 (N_6640,N_3036,N_3948);
and U6641 (N_6641,N_2968,N_1463);
or U6642 (N_6642,N_1578,N_2745);
and U6643 (N_6643,N_826,N_3164);
nor U6644 (N_6644,N_4897,N_1341);
nor U6645 (N_6645,N_1630,N_3719);
or U6646 (N_6646,N_1470,N_3025);
nor U6647 (N_6647,N_2797,N_4974);
nand U6648 (N_6648,N_2482,N_3575);
and U6649 (N_6649,N_3726,N_3148);
nand U6650 (N_6650,N_1584,N_2792);
xnor U6651 (N_6651,N_1289,N_3851);
nor U6652 (N_6652,N_944,N_4755);
or U6653 (N_6653,N_1814,N_3369);
and U6654 (N_6654,N_689,N_2003);
nand U6655 (N_6655,N_2727,N_1845);
nor U6656 (N_6656,N_3627,N_457);
and U6657 (N_6657,N_369,N_272);
nor U6658 (N_6658,N_4221,N_3733);
and U6659 (N_6659,N_4229,N_4106);
nor U6660 (N_6660,N_350,N_24);
nand U6661 (N_6661,N_1457,N_3378);
or U6662 (N_6662,N_4955,N_1016);
nand U6663 (N_6663,N_389,N_4703);
xor U6664 (N_6664,N_1478,N_732);
nor U6665 (N_6665,N_1736,N_913);
and U6666 (N_6666,N_1360,N_4049);
nor U6667 (N_6667,N_3986,N_1233);
xnor U6668 (N_6668,N_2850,N_1534);
and U6669 (N_6669,N_1820,N_1674);
and U6670 (N_6670,N_3690,N_3078);
xor U6671 (N_6671,N_3780,N_1951);
or U6672 (N_6672,N_3462,N_4788);
or U6673 (N_6673,N_1348,N_4620);
or U6674 (N_6674,N_1267,N_2675);
nand U6675 (N_6675,N_3174,N_385);
or U6676 (N_6676,N_2513,N_4219);
nor U6677 (N_6677,N_97,N_373);
nor U6678 (N_6678,N_207,N_1035);
nor U6679 (N_6679,N_4849,N_870);
and U6680 (N_6680,N_3016,N_3984);
or U6681 (N_6681,N_2724,N_609);
nand U6682 (N_6682,N_199,N_4399);
or U6683 (N_6683,N_1850,N_4231);
nor U6684 (N_6684,N_380,N_894);
nand U6685 (N_6685,N_3772,N_2552);
xor U6686 (N_6686,N_4529,N_2852);
or U6687 (N_6687,N_2109,N_3750);
nand U6688 (N_6688,N_221,N_4102);
nor U6689 (N_6689,N_2886,N_984);
xnor U6690 (N_6690,N_2806,N_4462);
nand U6691 (N_6691,N_1881,N_4205);
and U6692 (N_6692,N_3978,N_1046);
nor U6693 (N_6693,N_3015,N_1762);
and U6694 (N_6694,N_1540,N_662);
nand U6695 (N_6695,N_2907,N_1429);
or U6696 (N_6696,N_1637,N_4118);
nor U6697 (N_6697,N_3040,N_4736);
nor U6698 (N_6698,N_1685,N_422);
nand U6699 (N_6699,N_4541,N_652);
nor U6700 (N_6700,N_3935,N_2804);
nor U6701 (N_6701,N_2331,N_4895);
nand U6702 (N_6702,N_4930,N_202);
and U6703 (N_6703,N_4010,N_665);
and U6704 (N_6704,N_3175,N_2356);
or U6705 (N_6705,N_3083,N_197);
and U6706 (N_6706,N_4744,N_1307);
nand U6707 (N_6707,N_3637,N_4107);
xnor U6708 (N_6708,N_3342,N_2619);
nand U6709 (N_6709,N_1210,N_1323);
xor U6710 (N_6710,N_4950,N_767);
and U6711 (N_6711,N_4802,N_780);
nand U6712 (N_6712,N_5,N_2541);
nor U6713 (N_6713,N_2679,N_1182);
and U6714 (N_6714,N_1832,N_1013);
and U6715 (N_6715,N_2456,N_3670);
xor U6716 (N_6716,N_1764,N_4583);
and U6717 (N_6717,N_1398,N_513);
xor U6718 (N_6718,N_3877,N_4597);
nor U6719 (N_6719,N_3518,N_586);
and U6720 (N_6720,N_1886,N_4572);
or U6721 (N_6721,N_3007,N_21);
xor U6722 (N_6722,N_2396,N_4840);
nor U6723 (N_6723,N_3061,N_4248);
or U6724 (N_6724,N_3714,N_2605);
and U6725 (N_6725,N_2224,N_593);
nand U6726 (N_6726,N_1232,N_2144);
nand U6727 (N_6727,N_3149,N_3972);
xnor U6728 (N_6728,N_463,N_535);
or U6729 (N_6729,N_1581,N_1287);
nor U6730 (N_6730,N_638,N_1583);
and U6731 (N_6731,N_1473,N_4622);
nor U6732 (N_6732,N_3162,N_680);
nand U6733 (N_6733,N_1957,N_4875);
nand U6734 (N_6734,N_2475,N_2092);
nor U6735 (N_6735,N_2156,N_4282);
or U6736 (N_6736,N_4280,N_1999);
nor U6737 (N_6737,N_923,N_1882);
nor U6738 (N_6738,N_4360,N_1919);
or U6739 (N_6739,N_1164,N_2653);
or U6740 (N_6740,N_2924,N_3950);
nor U6741 (N_6741,N_2800,N_4758);
nor U6742 (N_6742,N_4382,N_378);
nand U6743 (N_6743,N_4123,N_2463);
nor U6744 (N_6744,N_2805,N_3599);
or U6745 (N_6745,N_2608,N_4972);
or U6746 (N_6746,N_2046,N_1525);
and U6747 (N_6747,N_367,N_1317);
and U6748 (N_6748,N_705,N_4899);
nor U6749 (N_6749,N_1783,N_3096);
and U6750 (N_6750,N_4361,N_4381);
nor U6751 (N_6751,N_741,N_2486);
nor U6752 (N_6752,N_3512,N_456);
or U6753 (N_6753,N_270,N_381);
nand U6754 (N_6754,N_4672,N_492);
or U6755 (N_6755,N_3570,N_3728);
nor U6756 (N_6756,N_313,N_1518);
and U6757 (N_6757,N_591,N_1156);
nand U6758 (N_6758,N_1254,N_4558);
nor U6759 (N_6759,N_499,N_1580);
or U6760 (N_6760,N_4961,N_4484);
nor U6761 (N_6761,N_54,N_340);
and U6762 (N_6762,N_2591,N_2558);
xnor U6763 (N_6763,N_2741,N_694);
nand U6764 (N_6764,N_1240,N_847);
nor U6765 (N_6765,N_3339,N_323);
xor U6766 (N_6766,N_4363,N_2461);
or U6767 (N_6767,N_3229,N_2963);
xnor U6768 (N_6768,N_4281,N_1998);
or U6769 (N_6769,N_1966,N_277);
nand U6770 (N_6770,N_426,N_4305);
or U6771 (N_6771,N_4392,N_957);
nand U6772 (N_6772,N_1408,N_2469);
or U6773 (N_6773,N_991,N_1625);
or U6774 (N_6774,N_1371,N_213);
nor U6775 (N_6775,N_2912,N_81);
nand U6776 (N_6776,N_2161,N_2528);
nor U6777 (N_6777,N_4008,N_1462);
nor U6778 (N_6778,N_4799,N_3527);
and U6779 (N_6779,N_987,N_3438);
nand U6780 (N_6780,N_2307,N_1937);
and U6781 (N_6781,N_2524,N_4420);
nand U6782 (N_6782,N_329,N_1387);
and U6783 (N_6783,N_691,N_1007);
nand U6784 (N_6784,N_4310,N_4885);
and U6785 (N_6785,N_4485,N_3561);
or U6786 (N_6786,N_2655,N_756);
xnor U6787 (N_6787,N_3341,N_1751);
or U6788 (N_6788,N_1592,N_3332);
nand U6789 (N_6789,N_3920,N_2631);
or U6790 (N_6790,N_4995,N_1224);
or U6791 (N_6791,N_1153,N_2086);
xnor U6792 (N_6792,N_589,N_2979);
and U6793 (N_6793,N_3464,N_4850);
nand U6794 (N_6794,N_4252,N_4167);
or U6795 (N_6795,N_724,N_572);
nand U6796 (N_6796,N_2550,N_3676);
and U6797 (N_6797,N_3151,N_127);
and U6798 (N_6798,N_4801,N_23);
nor U6799 (N_6799,N_1493,N_4016);
nand U6800 (N_6800,N_3176,N_1526);
and U6801 (N_6801,N_2047,N_1944);
or U6802 (N_6802,N_4871,N_3688);
nor U6803 (N_6803,N_125,N_2325);
xor U6804 (N_6804,N_1411,N_4811);
nor U6805 (N_6805,N_2757,N_3678);
xor U6806 (N_6806,N_2599,N_3178);
nand U6807 (N_6807,N_677,N_3959);
and U6808 (N_6808,N_2206,N_4636);
or U6809 (N_6809,N_1997,N_3483);
or U6810 (N_6810,N_2512,N_1033);
or U6811 (N_6811,N_2830,N_1069);
xor U6812 (N_6812,N_2164,N_2);
and U6813 (N_6813,N_2991,N_1548);
nor U6814 (N_6814,N_3731,N_1306);
nand U6815 (N_6815,N_1260,N_2801);
and U6816 (N_6816,N_3835,N_3615);
xor U6817 (N_6817,N_2845,N_4797);
or U6818 (N_6818,N_4742,N_1401);
or U6819 (N_6819,N_796,N_1542);
nor U6820 (N_6820,N_2881,N_3117);
nor U6821 (N_6821,N_4092,N_4476);
and U6822 (N_6822,N_4781,N_1745);
or U6823 (N_6823,N_4704,N_2670);
nor U6824 (N_6824,N_825,N_4828);
xnor U6825 (N_6825,N_3205,N_157);
nor U6826 (N_6826,N_1798,N_4006);
nand U6827 (N_6827,N_2448,N_1678);
and U6828 (N_6828,N_950,N_2181);
nor U6829 (N_6829,N_465,N_1672);
or U6830 (N_6830,N_2875,N_2865);
nand U6831 (N_6831,N_627,N_3602);
or U6832 (N_6832,N_4824,N_483);
nor U6833 (N_6833,N_1452,N_131);
and U6834 (N_6834,N_2262,N_711);
xor U6835 (N_6835,N_3132,N_3026);
nor U6836 (N_6836,N_4904,N_3060);
nand U6837 (N_6837,N_3793,N_4269);
or U6838 (N_6838,N_4201,N_2790);
nor U6839 (N_6839,N_4794,N_3158);
nand U6840 (N_6840,N_1252,N_3295);
or U6841 (N_6841,N_4643,N_1969);
nand U6842 (N_6842,N_4946,N_3145);
nand U6843 (N_6843,N_1739,N_2615);
nor U6844 (N_6844,N_4658,N_3129);
or U6845 (N_6845,N_4213,N_3513);
xnor U6846 (N_6846,N_69,N_1985);
nor U6847 (N_6847,N_4234,N_2353);
or U6848 (N_6848,N_4737,N_1618);
xnor U6849 (N_6849,N_1847,N_1864);
xnor U6850 (N_6850,N_383,N_4906);
or U6851 (N_6851,N_212,N_324);
or U6852 (N_6852,N_3679,N_431);
xor U6853 (N_6853,N_2525,N_4059);
or U6854 (N_6854,N_2781,N_1444);
xnor U6855 (N_6855,N_4297,N_2138);
nand U6856 (N_6856,N_1627,N_3401);
nand U6857 (N_6857,N_4187,N_1785);
nand U6858 (N_6858,N_2952,N_579);
or U6859 (N_6859,N_3262,N_3395);
and U6860 (N_6860,N_3554,N_2347);
nand U6861 (N_6861,N_1237,N_3488);
nor U6862 (N_6862,N_3087,N_3809);
and U6863 (N_6863,N_2627,N_4149);
or U6864 (N_6864,N_3737,N_3521);
nand U6865 (N_6865,N_2287,N_4190);
nand U6866 (N_6866,N_305,N_2119);
and U6867 (N_6867,N_114,N_846);
or U6868 (N_6868,N_2266,N_1849);
xnor U6869 (N_6869,N_1175,N_810);
and U6870 (N_6870,N_254,N_4496);
nand U6871 (N_6871,N_2367,N_4037);
and U6872 (N_6872,N_4346,N_1214);
or U6873 (N_6873,N_539,N_943);
xnor U6874 (N_6874,N_1735,N_2820);
and U6875 (N_6875,N_4728,N_2652);
nand U6876 (N_6876,N_1376,N_533);
nand U6877 (N_6877,N_470,N_3924);
nand U6878 (N_6878,N_4825,N_2646);
nor U6879 (N_6879,N_4021,N_2455);
or U6880 (N_6880,N_2732,N_3560);
and U6881 (N_6881,N_2914,N_2159);
nor U6882 (N_6882,N_1732,N_927);
xnor U6883 (N_6883,N_2972,N_2100);
nand U6884 (N_6884,N_4882,N_2487);
nor U6885 (N_6885,N_1553,N_2579);
or U6886 (N_6886,N_3643,N_4903);
nor U6887 (N_6887,N_1295,N_893);
xnor U6888 (N_6888,N_4697,N_2648);
nand U6889 (N_6889,N_973,N_1496);
nor U6890 (N_6890,N_2642,N_3352);
or U6891 (N_6891,N_3192,N_915);
and U6892 (N_6892,N_2538,N_1603);
or U6893 (N_6893,N_4478,N_424);
and U6894 (N_6894,N_985,N_551);
and U6895 (N_6895,N_1466,N_2267);
nor U6896 (N_6896,N_576,N_3326);
nor U6897 (N_6897,N_2300,N_2918);
or U6898 (N_6898,N_3170,N_2417);
and U6899 (N_6899,N_4492,N_3812);
xnor U6900 (N_6900,N_2187,N_1989);
or U6901 (N_6901,N_4800,N_8);
xor U6902 (N_6902,N_3049,N_3687);
or U6903 (N_6903,N_314,N_1056);
nor U6904 (N_6904,N_2457,N_3493);
and U6905 (N_6905,N_4245,N_2539);
and U6906 (N_6906,N_1043,N_1);
nand U6907 (N_6907,N_4444,N_1051);
nor U6908 (N_6908,N_3217,N_4944);
xor U6909 (N_6909,N_2028,N_287);
or U6910 (N_6910,N_1406,N_2111);
nor U6911 (N_6911,N_2073,N_444);
nor U6912 (N_6912,N_4076,N_1671);
nor U6913 (N_6913,N_566,N_3640);
or U6914 (N_6914,N_1447,N_2847);
or U6915 (N_6915,N_890,N_3043);
nor U6916 (N_6916,N_3557,N_2081);
nand U6917 (N_6917,N_1037,N_4344);
or U6918 (N_6918,N_824,N_1767);
xnor U6919 (N_6919,N_2229,N_2244);
nand U6920 (N_6920,N_1616,N_237);
and U6921 (N_6921,N_863,N_3974);
and U6922 (N_6922,N_1090,N_100);
nor U6923 (N_6923,N_4482,N_3838);
nand U6924 (N_6924,N_3103,N_486);
or U6925 (N_6925,N_3202,N_4316);
nand U6926 (N_6926,N_3048,N_1599);
and U6927 (N_6927,N_2815,N_146);
or U6928 (N_6928,N_4725,N_4511);
nor U6929 (N_6929,N_1024,N_614);
or U6930 (N_6930,N_3712,N_241);
and U6931 (N_6931,N_3764,N_2123);
nand U6932 (N_6932,N_1648,N_1311);
nor U6933 (N_6933,N_156,N_1753);
or U6934 (N_6934,N_1482,N_1831);
and U6935 (N_6935,N_490,N_3251);
or U6936 (N_6936,N_1869,N_404);
nor U6937 (N_6937,N_2157,N_2565);
nor U6938 (N_6938,N_1129,N_3242);
or U6939 (N_6939,N_4993,N_412);
xor U6940 (N_6940,N_568,N_4494);
and U6941 (N_6941,N_2705,N_2633);
nor U6942 (N_6942,N_1876,N_880);
or U6943 (N_6943,N_1812,N_1116);
and U6944 (N_6944,N_3265,N_3008);
and U6945 (N_6945,N_43,N_198);
nand U6946 (N_6946,N_1520,N_4124);
or U6947 (N_6947,N_1174,N_255);
nor U6948 (N_6948,N_1424,N_1299);
nand U6949 (N_6949,N_2115,N_2240);
nand U6950 (N_6950,N_1549,N_1790);
nor U6951 (N_6951,N_3266,N_1587);
and U6952 (N_6952,N_4952,N_624);
nand U6953 (N_6953,N_3768,N_1047);
or U6954 (N_6954,N_2393,N_4232);
nand U6955 (N_6955,N_1356,N_4352);
and U6956 (N_6956,N_900,N_1194);
nand U6957 (N_6957,N_4220,N_2160);
nor U6958 (N_6958,N_25,N_409);
and U6959 (N_6959,N_573,N_4353);
xor U6960 (N_6960,N_30,N_2188);
nor U6961 (N_6961,N_3680,N_4743);
and U6962 (N_6962,N_183,N_4365);
xnor U6963 (N_6963,N_208,N_1942);
and U6964 (N_6964,N_4324,N_2454);
nand U6965 (N_6965,N_79,N_3248);
and U6966 (N_6966,N_4831,N_260);
and U6967 (N_6967,N_3122,N_275);
nand U6968 (N_6968,N_4637,N_4983);
and U6969 (N_6969,N_1718,N_2225);
and U6970 (N_6970,N_2831,N_742);
nand U6971 (N_6971,N_2032,N_4401);
nand U6972 (N_6972,N_956,N_4121);
nor U6973 (N_6973,N_641,N_2803);
nor U6974 (N_6974,N_4,N_294);
nor U6975 (N_6975,N_1765,N_882);
and U6976 (N_6976,N_148,N_2338);
nand U6977 (N_6977,N_966,N_2385);
nor U6978 (N_6978,N_2332,N_1766);
nand U6979 (N_6979,N_1185,N_4525);
xor U6980 (N_6980,N_3306,N_3881);
nand U6981 (N_6981,N_3437,N_1195);
and U6982 (N_6982,N_234,N_2452);
and U6983 (N_6983,N_4294,N_4122);
nand U6984 (N_6984,N_98,N_2412);
and U6985 (N_6985,N_4877,N_4739);
xor U6986 (N_6986,N_1903,N_2257);
or U6987 (N_6987,N_2671,N_1058);
nand U6988 (N_6988,N_4601,N_2468);
nand U6989 (N_6989,N_3253,N_326);
or U6990 (N_6990,N_4596,N_4880);
nand U6991 (N_6991,N_3364,N_3066);
nor U6992 (N_6992,N_2318,N_85);
and U6993 (N_6993,N_4740,N_2892);
and U6994 (N_6994,N_2272,N_3739);
nand U6995 (N_6995,N_2434,N_58);
nand U6996 (N_6996,N_3819,N_4690);
nand U6997 (N_6997,N_2178,N_4237);
or U6998 (N_6998,N_833,N_3539);
nor U6999 (N_6999,N_3946,N_4752);
nor U7000 (N_7000,N_2931,N_402);
nand U7001 (N_7001,N_358,N_4131);
nand U7002 (N_7002,N_2140,N_280);
or U7003 (N_7003,N_4306,N_3104);
nand U7004 (N_7004,N_4038,N_1570);
and U7005 (N_7005,N_3933,N_2584);
and U7006 (N_7006,N_2166,N_575);
nor U7007 (N_7007,N_4349,N_2953);
xnor U7008 (N_7008,N_2269,N_1898);
nand U7009 (N_7009,N_1606,N_4347);
or U7010 (N_7010,N_4194,N_2637);
nor U7011 (N_7011,N_84,N_4159);
nor U7012 (N_7012,N_4856,N_3256);
and U7013 (N_7013,N_2685,N_2284);
and U7014 (N_7014,N_4986,N_4300);
nor U7015 (N_7015,N_2994,N_745);
and U7016 (N_7016,N_2981,N_1722);
and U7017 (N_7017,N_2142,N_2172);
nor U7018 (N_7018,N_2959,N_2920);
or U7019 (N_7019,N_2734,N_3551);
or U7020 (N_7020,N_2743,N_4093);
xnor U7021 (N_7021,N_33,N_3017);
nor U7022 (N_7022,N_3535,N_133);
or U7023 (N_7023,N_2819,N_1888);
nor U7024 (N_7024,N_4884,N_4115);
nand U7025 (N_7025,N_1334,N_4578);
or U7026 (N_7026,N_588,N_3583);
nor U7027 (N_7027,N_262,N_3080);
and U7028 (N_7028,N_2728,N_3524);
or U7029 (N_7029,N_1879,N_3781);
or U7030 (N_7030,N_182,N_1635);
and U7031 (N_7031,N_1901,N_4155);
nor U7032 (N_7032,N_2373,N_4861);
nand U7033 (N_7033,N_1801,N_2775);
or U7034 (N_7034,N_2473,N_854);
nor U7035 (N_7035,N_4301,N_2864);
and U7036 (N_7036,N_681,N_4613);
xnor U7037 (N_7037,N_398,N_346);
nor U7038 (N_7038,N_3443,N_2740);
nand U7039 (N_7039,N_929,N_3955);
nor U7040 (N_7040,N_2716,N_696);
and U7041 (N_7041,N_1286,N_430);
nor U7042 (N_7042,N_1860,N_4171);
or U7043 (N_7043,N_3730,N_3717);
nand U7044 (N_7044,N_2130,N_271);
or U7045 (N_7045,N_2025,N_3773);
and U7046 (N_7046,N_129,N_173);
nand U7047 (N_7047,N_3971,N_967);
and U7048 (N_7048,N_3576,N_2265);
xnor U7049 (N_7049,N_871,N_4835);
or U7050 (N_7050,N_1338,N_1158);
or U7051 (N_7051,N_3194,N_331);
nand U7052 (N_7052,N_1827,N_3801);
or U7053 (N_7053,N_4549,N_1562);
or U7054 (N_7054,N_4428,N_4318);
or U7055 (N_7055,N_4063,N_3704);
nand U7056 (N_7056,N_713,N_1170);
or U7057 (N_7057,N_1828,N_2016);
and U7058 (N_7058,N_509,N_1251);
nand U7059 (N_7059,N_2186,N_144);
and U7060 (N_7060,N_747,N_3724);
nand U7061 (N_7061,N_433,N_4934);
or U7062 (N_7062,N_1098,N_4757);
and U7063 (N_7063,N_4156,N_279);
and U7064 (N_7064,N_3813,N_462);
or U7065 (N_7065,N_4296,N_2587);
nor U7066 (N_7066,N_2691,N_45);
xnor U7067 (N_7067,N_1084,N_4216);
xor U7068 (N_7068,N_828,N_1991);
nor U7069 (N_7069,N_4607,N_2275);
and U7070 (N_7070,N_356,N_3715);
or U7071 (N_7071,N_3125,N_4776);
xor U7072 (N_7072,N_1715,N_2823);
nand U7073 (N_7073,N_3354,N_1112);
nor U7074 (N_7074,N_2871,N_4475);
nor U7075 (N_7075,N_4888,N_1455);
and U7076 (N_7076,N_2515,N_529);
or U7077 (N_7077,N_397,N_4526);
and U7078 (N_7078,N_3070,N_4970);
or U7079 (N_7079,N_2485,N_4577);
xor U7080 (N_7080,N_2227,N_4160);
and U7081 (N_7081,N_3223,N_3375);
nand U7082 (N_7082,N_2621,N_1824);
nand U7083 (N_7083,N_166,N_1615);
and U7084 (N_7084,N_2592,N_1128);
xor U7085 (N_7085,N_895,N_1190);
nand U7086 (N_7086,N_2546,N_1222);
nor U7087 (N_7087,N_4691,N_1015);
and U7088 (N_7088,N_1451,N_1178);
nor U7089 (N_7089,N_3209,N_4625);
and U7090 (N_7090,N_879,N_1332);
and U7091 (N_7091,N_3116,N_2252);
or U7092 (N_7092,N_3410,N_2167);
nor U7093 (N_7093,N_1954,N_1657);
nor U7094 (N_7094,N_2327,N_2279);
and U7095 (N_7095,N_1077,N_3929);
or U7096 (N_7096,N_3533,N_190);
and U7097 (N_7097,N_2782,N_676);
nand U7098 (N_7098,N_3544,N_189);
or U7099 (N_7099,N_1480,N_2828);
nor U7100 (N_7100,N_95,N_1197);
nor U7101 (N_7101,N_3880,N_3747);
and U7102 (N_7102,N_1379,N_4135);
xnor U7103 (N_7103,N_902,N_3657);
nand U7104 (N_7104,N_2542,N_3849);
or U7105 (N_7105,N_802,N_2479);
nor U7106 (N_7106,N_416,N_1186);
xor U7107 (N_7107,N_4045,N_247);
nor U7108 (N_7108,N_388,N_1029);
or U7109 (N_7109,N_3095,N_1900);
nand U7110 (N_7110,N_1613,N_2708);
nor U7111 (N_7111,N_2853,N_4025);
nand U7112 (N_7112,N_3606,N_2834);
nor U7113 (N_7113,N_83,N_2846);
nand U7114 (N_7114,N_71,N_3914);
or U7115 (N_7115,N_2885,N_3661);
nor U7116 (N_7116,N_4162,N_304);
nor U7117 (N_7117,N_3245,N_708);
and U7118 (N_7118,N_3314,N_2064);
nand U7119 (N_7119,N_2928,N_2293);
or U7120 (N_7120,N_321,N_2189);
and U7121 (N_7121,N_4751,N_3964);
and U7122 (N_7122,N_3702,N_3891);
nor U7123 (N_7123,N_1180,N_4978);
or U7124 (N_7124,N_2683,N_1897);
or U7125 (N_7125,N_4912,N_2305);
and U7126 (N_7126,N_4117,N_112);
nor U7127 (N_7127,N_1696,N_3792);
xor U7128 (N_7128,N_4217,N_938);
nor U7129 (N_7129,N_4913,N_265);
or U7130 (N_7130,N_1106,N_2494);
xnor U7131 (N_7131,N_1274,N_4175);
xnor U7132 (N_7132,N_134,N_718);
nor U7133 (N_7133,N_3433,N_4327);
nor U7134 (N_7134,N_4642,N_1344);
nand U7135 (N_7135,N_3968,N_3853);
and U7136 (N_7136,N_2658,N_4530);
nand U7137 (N_7137,N_3953,N_3236);
xor U7138 (N_7138,N_1930,N_1659);
and U7139 (N_7139,N_3651,N_494);
and U7140 (N_7140,N_376,N_4438);
nand U7141 (N_7141,N_4186,N_1830);
and U7142 (N_7142,N_4501,N_4867);
nor U7143 (N_7143,N_330,N_3141);
nor U7144 (N_7144,N_603,N_4198);
xor U7145 (N_7145,N_60,N_1259);
and U7146 (N_7146,N_4454,N_4534);
nand U7147 (N_7147,N_3021,N_2616);
or U7148 (N_7148,N_288,N_616);
or U7149 (N_7149,N_1921,N_3379);
and U7150 (N_7150,N_4593,N_1154);
or U7151 (N_7151,N_670,N_3086);
xor U7152 (N_7152,N_2882,N_1052);
and U7153 (N_7153,N_4176,N_4746);
nand U7154 (N_7154,N_1512,N_1868);
nor U7155 (N_7155,N_3820,N_623);
or U7156 (N_7156,N_174,N_3645);
or U7157 (N_7157,N_1621,N_4090);
or U7158 (N_7158,N_3975,N_3814);
and U7159 (N_7159,N_3200,N_2230);
nand U7160 (N_7160,N_1746,N_4278);
nand U7161 (N_7161,N_883,N_4692);
and U7162 (N_7162,N_4024,N_3916);
nor U7163 (N_7163,N_3588,N_2093);
nor U7164 (N_7164,N_4393,N_3785);
nand U7165 (N_7165,N_40,N_1650);
xor U7166 (N_7166,N_453,N_1139);
nor U7167 (N_7167,N_2863,N_2260);
or U7168 (N_7168,N_3062,N_253);
nand U7169 (N_7169,N_1301,N_3430);
xor U7170 (N_7170,N_2707,N_4909);
nor U7171 (N_7171,N_1572,N_3479);
nand U7172 (N_7172,N_3275,N_1328);
and U7173 (N_7173,N_2735,N_1683);
nand U7174 (N_7174,N_1082,N_3093);
or U7175 (N_7175,N_4268,N_2256);
and U7176 (N_7176,N_666,N_4819);
nand U7177 (N_7177,N_2087,N_4267);
and U7178 (N_7178,N_818,N_4429);
and U7179 (N_7179,N_3252,N_400);
and U7180 (N_7180,N_116,N_2818);
nor U7181 (N_7181,N_4227,N_647);
and U7182 (N_7182,N_4562,N_1533);
nand U7183 (N_7183,N_622,N_4009);
nand U7184 (N_7184,N_4773,N_2926);
nor U7185 (N_7185,N_1795,N_3718);
nand U7186 (N_7186,N_2211,N_892);
and U7187 (N_7187,N_645,N_4990);
and U7188 (N_7188,N_4988,N_856);
nor U7189 (N_7189,N_1948,N_3904);
and U7190 (N_7190,N_2421,N_1073);
or U7191 (N_7191,N_2193,N_1364);
and U7192 (N_7192,N_1268,N_4777);
nand U7193 (N_7193,N_2117,N_4859);
nor U7194 (N_7194,N_3808,N_138);
and U7195 (N_7195,N_1507,N_4569);
and U7196 (N_7196,N_2483,N_4656);
and U7197 (N_7197,N_1243,N_2000);
nand U7198 (N_7198,N_1432,N_2177);
and U7199 (N_7199,N_2746,N_4937);
and U7200 (N_7200,N_3709,N_4907);
nor U7201 (N_7201,N_249,N_2859);
and U7202 (N_7202,N_4251,N_2753);
and U7203 (N_7203,N_2259,N_798);
and U7204 (N_7204,N_959,N_505);
nor U7205 (N_7205,N_1597,N_3765);
or U7206 (N_7206,N_829,N_3537);
nor U7207 (N_7207,N_1425,N_2510);
and U7208 (N_7208,N_3309,N_821);
nor U7209 (N_7209,N_3220,N_2132);
and U7210 (N_7210,N_1981,N_1111);
xor U7211 (N_7211,N_3199,N_2171);
nand U7212 (N_7212,N_2711,N_1628);
and U7213 (N_7213,N_2083,N_64);
nand U7214 (N_7214,N_1594,N_2572);
nand U7215 (N_7215,N_4002,N_2586);
nand U7216 (N_7216,N_4677,N_3895);
and U7217 (N_7217,N_170,N_4778);
or U7218 (N_7218,N_4720,N_2878);
nor U7219 (N_7219,N_1388,N_3725);
nor U7220 (N_7220,N_2179,N_2440);
nand U7221 (N_7221,N_1171,N_3102);
or U7222 (N_7222,N_2139,N_1932);
and U7223 (N_7223,N_3109,N_1262);
and U7224 (N_7224,N_491,N_3404);
xor U7225 (N_7225,N_3063,N_2342);
or U7226 (N_7226,N_3366,N_730);
nor U7227 (N_7227,N_2811,N_2226);
xor U7228 (N_7228,N_3472,N_4713);
and U7229 (N_7229,N_342,N_1339);
or U7230 (N_7230,N_2688,N_167);
and U7231 (N_7231,N_1822,N_4398);
nor U7232 (N_7232,N_2941,N_4112);
nor U7233 (N_7233,N_48,N_3163);
nand U7234 (N_7234,N_2168,N_258);
or U7235 (N_7235,N_1054,N_307);
nor U7236 (N_7236,N_4629,N_3421);
nand U7237 (N_7237,N_4514,N_794);
or U7238 (N_7238,N_4929,N_3358);
or U7239 (N_7239,N_455,N_210);
xnor U7240 (N_7240,N_4383,N_2943);
nand U7241 (N_7241,N_673,N_3956);
nand U7242 (N_7242,N_2231,N_910);
and U7243 (N_7243,N_2126,N_4745);
or U7244 (N_7244,N_3297,N_3871);
or U7245 (N_7245,N_3832,N_2945);
nor U7246 (N_7246,N_2597,N_2350);
nand U7247 (N_7247,N_2958,N_1404);
nor U7248 (N_7248,N_4770,N_3285);
nand U7249 (N_7249,N_2326,N_1181);
nor U7250 (N_7250,N_3876,N_2212);
nand U7251 (N_7251,N_4137,N_4443);
and U7252 (N_7252,N_836,N_1759);
nand U7253 (N_7253,N_4647,N_110);
nor U7254 (N_7254,N_753,N_1923);
nor U7255 (N_7255,N_4710,N_2557);
xnor U7256 (N_7256,N_1810,N_3706);
nor U7257 (N_7257,N_774,N_3872);
and U7258 (N_7258,N_4920,N_2366);
and U7259 (N_7259,N_3797,N_3340);
or U7260 (N_7260,N_1433,N_3398);
and U7261 (N_7261,N_2844,N_3455);
xor U7262 (N_7262,N_1720,N_3184);
nand U7263 (N_7263,N_2899,N_1483);
or U7264 (N_7264,N_1958,N_2297);
and U7265 (N_7265,N_1895,N_1848);
nor U7266 (N_7266,N_4832,N_1221);
nand U7267 (N_7267,N_4293,N_2070);
or U7268 (N_7268,N_906,N_3543);
or U7269 (N_7269,N_3427,N_3327);
and U7270 (N_7270,N_4362,N_868);
or U7271 (N_7271,N_468,N_178);
nor U7272 (N_7272,N_3152,N_1416);
and U7273 (N_7273,N_2547,N_230);
and U7274 (N_7274,N_1973,N_702);
nand U7275 (N_7275,N_3859,N_1986);
nor U7276 (N_7276,N_4996,N_2324);
nor U7277 (N_7277,N_2098,N_1537);
and U7278 (N_7278,N_3460,N_3992);
nand U7279 (N_7279,N_3997,N_3118);
or U7280 (N_7280,N_4805,N_4434);
and U7281 (N_7281,N_3052,N_1426);
nand U7282 (N_7282,N_4521,N_3495);
and U7283 (N_7283,N_2897,N_1367);
or U7284 (N_7284,N_3185,N_1019);
xor U7285 (N_7285,N_4325,N_4579);
nor U7286 (N_7286,N_4540,N_2215);
or U7287 (N_7287,N_11,N_4011);
and U7288 (N_7288,N_607,N_3617);
or U7289 (N_7289,N_2810,N_2022);
nand U7290 (N_7290,N_1445,N_4733);
and U7291 (N_7291,N_1777,N_4998);
or U7292 (N_7292,N_2521,N_3556);
nand U7293 (N_7293,N_881,N_965);
and U7294 (N_7294,N_3034,N_285);
or U7295 (N_7295,N_1494,N_2841);
xnor U7296 (N_7296,N_2964,N_1495);
nand U7297 (N_7297,N_667,N_2595);
nor U7298 (N_7298,N_1509,N_3944);
xnor U7299 (N_7299,N_4741,N_1598);
nor U7300 (N_7300,N_2359,N_4589);
or U7301 (N_7301,N_2995,N_993);
and U7302 (N_7302,N_1490,N_274);
nand U7303 (N_7303,N_3144,N_866);
or U7304 (N_7304,N_980,N_3611);
xnor U7305 (N_7305,N_1343,N_964);
and U7306 (N_7306,N_1012,N_3988);
and U7307 (N_7307,N_2184,N_3167);
nand U7308 (N_7308,N_981,N_4120);
or U7309 (N_7309,N_282,N_2470);
xor U7310 (N_7310,N_1390,N_3005);
and U7311 (N_7311,N_1066,N_2054);
nand U7312 (N_7312,N_4573,N_354);
or U7313 (N_7313,N_3228,N_648);
nand U7314 (N_7314,N_4127,N_4854);
or U7315 (N_7315,N_235,N_123);
nor U7316 (N_7316,N_2654,N_4513);
and U7317 (N_7317,N_3884,N_1273);
and U7318 (N_7318,N_2077,N_3022);
and U7319 (N_7319,N_2377,N_4314);
and U7320 (N_7320,N_989,N_2822);
nor U7321 (N_7321,N_947,N_1165);
nor U7322 (N_7322,N_3214,N_345);
and U7323 (N_7323,N_757,N_4459);
xor U7324 (N_7324,N_106,N_4644);
or U7325 (N_7325,N_2076,N_1258);
and U7326 (N_7326,N_939,N_3349);
nand U7327 (N_7327,N_2821,N_1866);
nor U7328 (N_7328,N_804,N_2263);
nor U7329 (N_7329,N_438,N_4709);
xnor U7330 (N_7330,N_3257,N_3915);
nor U7331 (N_7331,N_1717,N_4869);
or U7332 (N_7332,N_218,N_1504);
nand U7333 (N_7333,N_82,N_4329);
nor U7334 (N_7334,N_17,N_1538);
nor U7335 (N_7335,N_3509,N_2317);
nand U7336 (N_7336,N_504,N_3934);
nand U7337 (N_7337,N_2097,N_1316);
nand U7338 (N_7338,N_3478,N_1813);
nand U7339 (N_7339,N_3707,N_2242);
nand U7340 (N_7340,N_4766,N_3280);
nand U7341 (N_7341,N_3081,N_4235);
or U7342 (N_7342,N_4457,N_3329);
nand U7343 (N_7343,N_3590,N_497);
nor U7344 (N_7344,N_4498,N_515);
or U7345 (N_7345,N_1794,N_1663);
or U7346 (N_7346,N_1288,N_2630);
nor U7347 (N_7347,N_4553,N_712);
nand U7348 (N_7348,N_2214,N_3130);
nor U7349 (N_7349,N_2182,N_549);
and U7350 (N_7350,N_1145,N_3261);
or U7351 (N_7351,N_734,N_2285);
and U7352 (N_7352,N_4524,N_1191);
xnor U7353 (N_7353,N_290,N_1974);
or U7354 (N_7354,N_4101,N_9);
or U7355 (N_7355,N_1797,N_4497);
and U7356 (N_7356,N_2146,N_2492);
nand U7357 (N_7357,N_4606,N_1602);
nor U7358 (N_7358,N_4193,N_1080);
nand U7359 (N_7359,N_2460,N_4681);
nand U7360 (N_7360,N_4696,N_1782);
nand U7361 (N_7361,N_2017,N_1464);
nand U7362 (N_7362,N_4125,N_4384);
nand U7363 (N_7363,N_4706,N_1305);
or U7364 (N_7364,N_3177,N_3982);
nor U7365 (N_7365,N_3672,N_3977);
and U7366 (N_7366,N_1266,N_1649);
nor U7367 (N_7367,N_546,N_2079);
and U7368 (N_7368,N_979,N_1321);
xnor U7369 (N_7369,N_3317,N_3272);
nand U7370 (N_7370,N_2010,N_813);
xnor U7371 (N_7371,N_4791,N_3399);
nor U7372 (N_7372,N_1950,N_2071);
nand U7373 (N_7373,N_1365,N_4170);
and U7374 (N_7374,N_2207,N_827);
and U7375 (N_7375,N_3998,N_1096);
nand U7376 (N_7376,N_2611,N_2575);
nand U7377 (N_7377,N_3506,N_3446);
or U7378 (N_7378,N_2496,N_1352);
and U7379 (N_7379,N_1050,N_1118);
nand U7380 (N_7380,N_3802,N_541);
or U7381 (N_7381,N_2135,N_414);
xnor U7382 (N_7382,N_4557,N_1138);
or U7383 (N_7383,N_2372,N_2034);
nor U7384 (N_7384,N_3906,N_969);
nand U7385 (N_7385,N_1515,N_3639);
and U7386 (N_7386,N_3442,N_461);
nand U7387 (N_7387,N_4132,N_3333);
nand U7388 (N_7388,N_301,N_3486);
and U7389 (N_7389,N_3894,N_318);
nand U7390 (N_7390,N_3269,N_2673);
and U7391 (N_7391,N_3385,N_1532);
nor U7392 (N_7392,N_2639,N_2962);
nor U7393 (N_7393,N_4298,N_4591);
nand U7394 (N_7394,N_2802,N_1072);
and U7395 (N_7395,N_986,N_176);
xor U7396 (N_7396,N_4200,N_3579);
nand U7397 (N_7397,N_2573,N_4748);
and U7398 (N_7398,N_1091,N_1501);
or U7399 (N_7399,N_2498,N_823);
or U7400 (N_7400,N_1442,N_2239);
nor U7401 (N_7401,N_1971,N_4439);
or U7402 (N_7402,N_3212,N_2065);
or U7403 (N_7403,N_2282,N_561);
and U7404 (N_7404,N_482,N_2439);
or U7405 (N_7405,N_788,N_4609);
nor U7406 (N_7406,N_816,N_3330);
and U7407 (N_7407,N_3126,N_3079);
nand U7408 (N_7408,N_447,N_1815);
and U7409 (N_7409,N_754,N_3180);
nand U7410 (N_7410,N_4670,N_4523);
nor U7411 (N_7411,N_3020,N_3783);
and U7412 (N_7412,N_3120,N_2021);
nand U7413 (N_7413,N_3480,N_4711);
nor U7414 (N_7414,N_908,N_2228);
and U7415 (N_7415,N_4331,N_4612);
nand U7416 (N_7416,N_1335,N_3156);
nor U7417 (N_7417,N_4358,N_4085);
and U7418 (N_7418,N_4570,N_1938);
and U7419 (N_7419,N_4488,N_4784);
nand U7420 (N_7420,N_2101,N_4975);
and U7421 (N_7421,N_136,N_1225);
nand U7422 (N_7422,N_946,N_4455);
xor U7423 (N_7423,N_4608,N_1712);
and U7424 (N_7424,N_2219,N_2120);
nand U7425 (N_7425,N_625,N_3631);
and U7426 (N_7426,N_954,N_1702);
xor U7427 (N_7427,N_1472,N_4055);
and U7428 (N_7428,N_998,N_1211);
or U7429 (N_7429,N_1555,N_1721);
nand U7430 (N_7430,N_3847,N_4669);
nor U7431 (N_7431,N_1644,N_2203);
or U7432 (N_7432,N_2930,N_2283);
xor U7433 (N_7433,N_2594,N_595);
nand U7434 (N_7434,N_3119,N_4936);
and U7435 (N_7435,N_336,N_4174);
xnor U7436 (N_7436,N_4873,N_3059);
nand U7437 (N_7437,N_1340,N_3927);
or U7438 (N_7438,N_4966,N_4446);
nand U7439 (N_7439,N_3011,N_4695);
and U7440 (N_7440,N_3235,N_4663);
and U7441 (N_7441,N_3973,N_1034);
nand U7442 (N_7442,N_160,N_4461);
xnor U7443 (N_7443,N_4495,N_1666);
nand U7444 (N_7444,N_4932,N_4421);
nor U7445 (N_7445,N_3671,N_2940);
or U7446 (N_7446,N_917,N_1857);
nand U7447 (N_7447,N_185,N_2949);
nor U7448 (N_7448,N_2564,N_2007);
nor U7449 (N_7449,N_2913,N_4158);
and U7450 (N_7450,N_2085,N_334);
and U7451 (N_7451,N_1541,N_4915);
nor U7452 (N_7452,N_126,N_3028);
nor U7453 (N_7453,N_4084,N_658);
nand U7454 (N_7454,N_678,N_2072);
xor U7455 (N_7455,N_1166,N_3526);
nor U7456 (N_7456,N_2337,N_820);
xor U7457 (N_7457,N_364,N_3722);
or U7458 (N_7458,N_53,N_1477);
or U7459 (N_7459,N_4889,N_2441);
or U7460 (N_7460,N_4576,N_1309);
nand U7461 (N_7461,N_3324,N_2883);
nand U7462 (N_7462,N_4759,N_853);
nand U7463 (N_7463,N_2779,N_394);
nor U7464 (N_7464,N_3107,N_3064);
nor U7465 (N_7465,N_4067,N_3600);
or U7466 (N_7466,N_654,N_2464);
or U7467 (N_7467,N_580,N_428);
nand U7468 (N_7468,N_4700,N_2011);
or U7469 (N_7469,N_1972,N_4317);
and U7470 (N_7470,N_4264,N_1005);
nor U7471 (N_7471,N_1724,N_1945);
nand U7472 (N_7472,N_1579,N_4769);
nand U7473 (N_7473,N_1385,N_2114);
nand U7474 (N_7474,N_4604,N_3559);
and U7475 (N_7475,N_1467,N_3770);
nor U7476 (N_7476,N_4574,N_2506);
or U7477 (N_7477,N_4288,N_2693);
xor U7478 (N_7478,N_3424,N_4933);
and U7479 (N_7479,N_4196,N_4470);
nand U7480 (N_7480,N_2020,N_4337);
or U7481 (N_7481,N_91,N_1020);
nand U7482 (N_7482,N_2369,N_3566);
xnor U7483 (N_7483,N_1438,N_3517);
or U7484 (N_7484,N_772,N_1576);
nor U7485 (N_7485,N_3742,N_3593);
or U7486 (N_7486,N_4980,N_1055);
nor U7487 (N_7487,N_690,N_1667);
nand U7488 (N_7488,N_3325,N_557);
xnor U7489 (N_7489,N_1454,N_224);
nor U7490 (N_7490,N_3300,N_4890);
or U7491 (N_7491,N_3106,N_1643);
nor U7492 (N_7492,N_1614,N_3073);
and U7493 (N_7493,N_1924,N_1121);
nand U7494 (N_7494,N_2002,N_1443);
nand U7495 (N_7495,N_363,N_4168);
or U7496 (N_7496,N_1682,N_3991);
nor U7497 (N_7497,N_3384,N_2915);
nand U7498 (N_7498,N_2689,N_4299);
nor U7499 (N_7499,N_4128,N_1808);
nand U7500 (N_7500,N_1855,N_217);
and U7501 (N_7501,N_1778,N_3869);
nand U7502 (N_7502,N_3800,N_2144);
or U7503 (N_7503,N_2878,N_265);
or U7504 (N_7504,N_1563,N_3958);
and U7505 (N_7505,N_1517,N_3102);
or U7506 (N_7506,N_3037,N_3210);
nor U7507 (N_7507,N_4108,N_951);
and U7508 (N_7508,N_1473,N_2460);
nand U7509 (N_7509,N_2387,N_1645);
or U7510 (N_7510,N_2915,N_4181);
nor U7511 (N_7511,N_2509,N_1115);
and U7512 (N_7512,N_883,N_4547);
or U7513 (N_7513,N_4413,N_1143);
nand U7514 (N_7514,N_1878,N_3431);
nor U7515 (N_7515,N_4346,N_4499);
and U7516 (N_7516,N_3386,N_122);
and U7517 (N_7517,N_1394,N_2395);
or U7518 (N_7518,N_2949,N_1384);
and U7519 (N_7519,N_746,N_175);
and U7520 (N_7520,N_1028,N_2471);
nor U7521 (N_7521,N_1145,N_3990);
or U7522 (N_7522,N_2037,N_2607);
xnor U7523 (N_7523,N_3862,N_1962);
nor U7524 (N_7524,N_1193,N_305);
xor U7525 (N_7525,N_1109,N_2272);
and U7526 (N_7526,N_3860,N_4443);
and U7527 (N_7527,N_4318,N_4706);
nand U7528 (N_7528,N_2783,N_4595);
and U7529 (N_7529,N_1033,N_2817);
nand U7530 (N_7530,N_1688,N_4626);
or U7531 (N_7531,N_4698,N_1583);
and U7532 (N_7532,N_4100,N_694);
nor U7533 (N_7533,N_1536,N_1634);
nor U7534 (N_7534,N_2524,N_484);
nand U7535 (N_7535,N_1256,N_753);
nor U7536 (N_7536,N_1813,N_3558);
and U7537 (N_7537,N_4789,N_3531);
nor U7538 (N_7538,N_2857,N_2998);
nand U7539 (N_7539,N_1366,N_4307);
nor U7540 (N_7540,N_871,N_2330);
nand U7541 (N_7541,N_610,N_2771);
nor U7542 (N_7542,N_905,N_2552);
and U7543 (N_7543,N_4977,N_4950);
or U7544 (N_7544,N_2704,N_4810);
or U7545 (N_7545,N_583,N_4515);
xor U7546 (N_7546,N_435,N_4249);
xor U7547 (N_7547,N_464,N_3074);
and U7548 (N_7548,N_1714,N_924);
nor U7549 (N_7549,N_115,N_194);
or U7550 (N_7550,N_661,N_378);
or U7551 (N_7551,N_2932,N_2432);
or U7552 (N_7552,N_712,N_609);
and U7553 (N_7553,N_2372,N_554);
or U7554 (N_7554,N_92,N_1300);
nand U7555 (N_7555,N_2811,N_4710);
and U7556 (N_7556,N_3866,N_960);
and U7557 (N_7557,N_2013,N_1257);
nor U7558 (N_7558,N_3273,N_1671);
and U7559 (N_7559,N_2230,N_2213);
nand U7560 (N_7560,N_3135,N_3577);
and U7561 (N_7561,N_306,N_2969);
nor U7562 (N_7562,N_2948,N_1362);
nor U7563 (N_7563,N_325,N_2609);
or U7564 (N_7564,N_1844,N_3031);
or U7565 (N_7565,N_1101,N_2329);
nand U7566 (N_7566,N_1704,N_893);
nand U7567 (N_7567,N_4628,N_1751);
or U7568 (N_7568,N_1361,N_3039);
or U7569 (N_7569,N_3754,N_940);
nor U7570 (N_7570,N_4664,N_1423);
nand U7571 (N_7571,N_1203,N_3113);
nor U7572 (N_7572,N_4037,N_3584);
nor U7573 (N_7573,N_4750,N_606);
nor U7574 (N_7574,N_4926,N_4781);
or U7575 (N_7575,N_4198,N_4970);
nor U7576 (N_7576,N_1293,N_465);
or U7577 (N_7577,N_2728,N_4995);
and U7578 (N_7578,N_2945,N_4388);
nand U7579 (N_7579,N_1818,N_2964);
nand U7580 (N_7580,N_3705,N_4056);
nor U7581 (N_7581,N_4594,N_3542);
or U7582 (N_7582,N_3969,N_954);
nor U7583 (N_7583,N_762,N_3652);
nand U7584 (N_7584,N_4128,N_4720);
xnor U7585 (N_7585,N_2832,N_1391);
or U7586 (N_7586,N_3774,N_119);
xor U7587 (N_7587,N_1828,N_4907);
nand U7588 (N_7588,N_438,N_2043);
nor U7589 (N_7589,N_1248,N_1020);
xnor U7590 (N_7590,N_2946,N_829);
nor U7591 (N_7591,N_1688,N_1740);
or U7592 (N_7592,N_3111,N_423);
xor U7593 (N_7593,N_3057,N_2804);
or U7594 (N_7594,N_2909,N_3192);
nor U7595 (N_7595,N_1646,N_4823);
nand U7596 (N_7596,N_632,N_520);
and U7597 (N_7597,N_3532,N_16);
and U7598 (N_7598,N_2506,N_1491);
nor U7599 (N_7599,N_2423,N_3015);
or U7600 (N_7600,N_3756,N_3794);
xnor U7601 (N_7601,N_642,N_3301);
and U7602 (N_7602,N_2801,N_4280);
xor U7603 (N_7603,N_3190,N_3527);
and U7604 (N_7604,N_642,N_371);
nand U7605 (N_7605,N_110,N_151);
and U7606 (N_7606,N_2583,N_3466);
nor U7607 (N_7607,N_784,N_29);
or U7608 (N_7608,N_3113,N_1015);
and U7609 (N_7609,N_1050,N_3038);
nand U7610 (N_7610,N_3365,N_4613);
nor U7611 (N_7611,N_4822,N_3517);
and U7612 (N_7612,N_3730,N_4330);
nand U7613 (N_7613,N_3359,N_1360);
and U7614 (N_7614,N_896,N_970);
and U7615 (N_7615,N_2689,N_637);
nand U7616 (N_7616,N_402,N_449);
and U7617 (N_7617,N_1376,N_2716);
nor U7618 (N_7618,N_2067,N_3674);
nand U7619 (N_7619,N_4569,N_3446);
and U7620 (N_7620,N_1865,N_4442);
and U7621 (N_7621,N_3446,N_4921);
nor U7622 (N_7622,N_724,N_615);
nand U7623 (N_7623,N_211,N_4204);
or U7624 (N_7624,N_153,N_3448);
xnor U7625 (N_7625,N_4505,N_2477);
or U7626 (N_7626,N_1378,N_3932);
xnor U7627 (N_7627,N_1408,N_2989);
xor U7628 (N_7628,N_866,N_3258);
and U7629 (N_7629,N_160,N_1567);
xor U7630 (N_7630,N_1874,N_1579);
and U7631 (N_7631,N_665,N_3262);
nand U7632 (N_7632,N_1728,N_2309);
and U7633 (N_7633,N_860,N_2717);
nor U7634 (N_7634,N_4764,N_3886);
or U7635 (N_7635,N_502,N_2050);
nand U7636 (N_7636,N_2468,N_4497);
nand U7637 (N_7637,N_4423,N_2730);
or U7638 (N_7638,N_4127,N_63);
or U7639 (N_7639,N_2086,N_880);
or U7640 (N_7640,N_3118,N_3759);
nor U7641 (N_7641,N_326,N_1687);
nand U7642 (N_7642,N_1965,N_4420);
or U7643 (N_7643,N_2821,N_1022);
or U7644 (N_7644,N_243,N_3131);
or U7645 (N_7645,N_66,N_71);
nand U7646 (N_7646,N_4689,N_1809);
nand U7647 (N_7647,N_3225,N_4898);
xor U7648 (N_7648,N_4253,N_3682);
xor U7649 (N_7649,N_1742,N_1797);
xnor U7650 (N_7650,N_4952,N_3189);
nand U7651 (N_7651,N_3042,N_2073);
nor U7652 (N_7652,N_2001,N_3915);
or U7653 (N_7653,N_4994,N_4690);
xor U7654 (N_7654,N_1592,N_3750);
or U7655 (N_7655,N_4312,N_4012);
and U7656 (N_7656,N_3665,N_4265);
xnor U7657 (N_7657,N_3258,N_3250);
or U7658 (N_7658,N_411,N_792);
and U7659 (N_7659,N_804,N_2999);
and U7660 (N_7660,N_3826,N_2473);
nor U7661 (N_7661,N_1677,N_4593);
or U7662 (N_7662,N_1409,N_952);
nand U7663 (N_7663,N_2679,N_3252);
xor U7664 (N_7664,N_4253,N_3111);
nand U7665 (N_7665,N_4881,N_712);
nand U7666 (N_7666,N_3241,N_4392);
or U7667 (N_7667,N_828,N_3168);
nand U7668 (N_7668,N_1148,N_626);
nand U7669 (N_7669,N_381,N_3957);
nor U7670 (N_7670,N_3400,N_4633);
and U7671 (N_7671,N_2757,N_4168);
and U7672 (N_7672,N_4445,N_1805);
or U7673 (N_7673,N_3857,N_2158);
nand U7674 (N_7674,N_1250,N_1876);
nor U7675 (N_7675,N_4783,N_3025);
or U7676 (N_7676,N_1194,N_3841);
and U7677 (N_7677,N_1068,N_570);
or U7678 (N_7678,N_493,N_2482);
and U7679 (N_7679,N_2090,N_2105);
nor U7680 (N_7680,N_1027,N_2647);
or U7681 (N_7681,N_222,N_1476);
nor U7682 (N_7682,N_4280,N_1603);
and U7683 (N_7683,N_2596,N_514);
and U7684 (N_7684,N_1820,N_1602);
or U7685 (N_7685,N_2605,N_3606);
and U7686 (N_7686,N_3859,N_2375);
nand U7687 (N_7687,N_2540,N_246);
nor U7688 (N_7688,N_340,N_4367);
and U7689 (N_7689,N_4941,N_3471);
xor U7690 (N_7690,N_4026,N_1154);
xor U7691 (N_7691,N_2965,N_2783);
and U7692 (N_7692,N_281,N_4506);
or U7693 (N_7693,N_752,N_4358);
or U7694 (N_7694,N_81,N_4868);
nand U7695 (N_7695,N_3284,N_825);
nor U7696 (N_7696,N_4379,N_4955);
nor U7697 (N_7697,N_1594,N_2392);
and U7698 (N_7698,N_4384,N_3747);
nand U7699 (N_7699,N_560,N_3660);
xor U7700 (N_7700,N_801,N_670);
nand U7701 (N_7701,N_106,N_1223);
nand U7702 (N_7702,N_781,N_1243);
nand U7703 (N_7703,N_204,N_976);
nor U7704 (N_7704,N_1874,N_3388);
or U7705 (N_7705,N_4041,N_737);
and U7706 (N_7706,N_370,N_1949);
nand U7707 (N_7707,N_1497,N_1186);
nand U7708 (N_7708,N_727,N_2376);
nand U7709 (N_7709,N_1787,N_1642);
nor U7710 (N_7710,N_529,N_1490);
nand U7711 (N_7711,N_4227,N_1216);
xnor U7712 (N_7712,N_4498,N_808);
or U7713 (N_7713,N_4512,N_2113);
and U7714 (N_7714,N_3299,N_1642);
and U7715 (N_7715,N_2196,N_726);
nor U7716 (N_7716,N_1154,N_1420);
or U7717 (N_7717,N_835,N_2037);
or U7718 (N_7718,N_2857,N_2574);
xnor U7719 (N_7719,N_3810,N_1911);
nand U7720 (N_7720,N_3041,N_258);
and U7721 (N_7721,N_1894,N_4436);
and U7722 (N_7722,N_903,N_1920);
or U7723 (N_7723,N_809,N_2315);
nor U7724 (N_7724,N_3813,N_3673);
xnor U7725 (N_7725,N_373,N_4197);
nand U7726 (N_7726,N_3587,N_409);
nor U7727 (N_7727,N_226,N_3820);
nor U7728 (N_7728,N_1278,N_842);
nor U7729 (N_7729,N_1875,N_1766);
nor U7730 (N_7730,N_1638,N_4762);
and U7731 (N_7731,N_664,N_639);
nand U7732 (N_7732,N_517,N_1486);
and U7733 (N_7733,N_2220,N_450);
and U7734 (N_7734,N_1982,N_1220);
or U7735 (N_7735,N_2350,N_2889);
or U7736 (N_7736,N_1575,N_2911);
nor U7737 (N_7737,N_3325,N_2887);
nand U7738 (N_7738,N_2073,N_511);
nand U7739 (N_7739,N_256,N_1172);
nor U7740 (N_7740,N_4104,N_1631);
nand U7741 (N_7741,N_3691,N_1790);
nor U7742 (N_7742,N_2772,N_4543);
nor U7743 (N_7743,N_4213,N_31);
or U7744 (N_7744,N_4334,N_2671);
and U7745 (N_7745,N_4121,N_3816);
nand U7746 (N_7746,N_4135,N_4284);
nand U7747 (N_7747,N_1149,N_1441);
nor U7748 (N_7748,N_1671,N_2176);
or U7749 (N_7749,N_1354,N_2585);
and U7750 (N_7750,N_279,N_346);
and U7751 (N_7751,N_2470,N_3223);
or U7752 (N_7752,N_2528,N_1254);
nor U7753 (N_7753,N_1561,N_4269);
or U7754 (N_7754,N_2688,N_3109);
or U7755 (N_7755,N_611,N_892);
nor U7756 (N_7756,N_1105,N_2504);
and U7757 (N_7757,N_3819,N_1151);
nor U7758 (N_7758,N_2305,N_1411);
nor U7759 (N_7759,N_3651,N_1844);
and U7760 (N_7760,N_151,N_1771);
nor U7761 (N_7761,N_656,N_3839);
and U7762 (N_7762,N_1845,N_3579);
and U7763 (N_7763,N_3529,N_4946);
nor U7764 (N_7764,N_4811,N_160);
or U7765 (N_7765,N_1945,N_234);
nand U7766 (N_7766,N_4974,N_4610);
and U7767 (N_7767,N_1643,N_205);
nor U7768 (N_7768,N_1424,N_4478);
xor U7769 (N_7769,N_798,N_3881);
nor U7770 (N_7770,N_2929,N_355);
or U7771 (N_7771,N_1891,N_1183);
nor U7772 (N_7772,N_2549,N_1266);
xnor U7773 (N_7773,N_454,N_2929);
nor U7774 (N_7774,N_4130,N_1544);
nor U7775 (N_7775,N_2871,N_3835);
nor U7776 (N_7776,N_1868,N_1929);
xor U7777 (N_7777,N_3052,N_4165);
nand U7778 (N_7778,N_1992,N_949);
xor U7779 (N_7779,N_3352,N_4894);
or U7780 (N_7780,N_4468,N_2816);
or U7781 (N_7781,N_3347,N_841);
and U7782 (N_7782,N_949,N_1718);
nor U7783 (N_7783,N_1762,N_4169);
or U7784 (N_7784,N_851,N_555);
nor U7785 (N_7785,N_3021,N_180);
nand U7786 (N_7786,N_2073,N_4299);
nand U7787 (N_7787,N_143,N_549);
xor U7788 (N_7788,N_3708,N_4267);
and U7789 (N_7789,N_1257,N_3971);
and U7790 (N_7790,N_4797,N_3086);
and U7791 (N_7791,N_3159,N_4634);
xor U7792 (N_7792,N_2132,N_3924);
or U7793 (N_7793,N_3515,N_2032);
nand U7794 (N_7794,N_3419,N_1307);
or U7795 (N_7795,N_4837,N_2354);
nand U7796 (N_7796,N_844,N_3236);
nor U7797 (N_7797,N_3209,N_2162);
nand U7798 (N_7798,N_593,N_1485);
nor U7799 (N_7799,N_2191,N_89);
nand U7800 (N_7800,N_1305,N_816);
nand U7801 (N_7801,N_2289,N_739);
or U7802 (N_7802,N_3226,N_2593);
and U7803 (N_7803,N_688,N_1193);
and U7804 (N_7804,N_1317,N_3547);
or U7805 (N_7805,N_4733,N_4049);
and U7806 (N_7806,N_4977,N_229);
or U7807 (N_7807,N_754,N_1724);
xor U7808 (N_7808,N_2699,N_3629);
or U7809 (N_7809,N_1891,N_3933);
and U7810 (N_7810,N_363,N_3089);
nand U7811 (N_7811,N_4217,N_2838);
or U7812 (N_7812,N_2869,N_3633);
or U7813 (N_7813,N_889,N_2850);
and U7814 (N_7814,N_2193,N_1962);
xor U7815 (N_7815,N_188,N_944);
nor U7816 (N_7816,N_2853,N_2327);
nor U7817 (N_7817,N_1977,N_2975);
nor U7818 (N_7818,N_1866,N_2375);
nor U7819 (N_7819,N_1908,N_3940);
or U7820 (N_7820,N_3997,N_4695);
nor U7821 (N_7821,N_1189,N_2958);
or U7822 (N_7822,N_2336,N_4883);
nand U7823 (N_7823,N_4640,N_2960);
or U7824 (N_7824,N_4229,N_4757);
and U7825 (N_7825,N_4852,N_2989);
nor U7826 (N_7826,N_337,N_2286);
xnor U7827 (N_7827,N_1841,N_925);
or U7828 (N_7828,N_84,N_4396);
and U7829 (N_7829,N_1064,N_3295);
and U7830 (N_7830,N_2226,N_2143);
nand U7831 (N_7831,N_2372,N_2993);
nor U7832 (N_7832,N_38,N_2128);
and U7833 (N_7833,N_689,N_3613);
nand U7834 (N_7834,N_2603,N_4185);
or U7835 (N_7835,N_4922,N_2030);
nand U7836 (N_7836,N_2492,N_4833);
and U7837 (N_7837,N_1615,N_720);
nor U7838 (N_7838,N_3043,N_3285);
nand U7839 (N_7839,N_150,N_1745);
nor U7840 (N_7840,N_2812,N_2950);
nor U7841 (N_7841,N_1991,N_1876);
nor U7842 (N_7842,N_4715,N_2894);
nor U7843 (N_7843,N_4663,N_2641);
nor U7844 (N_7844,N_1247,N_4996);
nand U7845 (N_7845,N_2007,N_2175);
nand U7846 (N_7846,N_3499,N_1244);
or U7847 (N_7847,N_4207,N_963);
nor U7848 (N_7848,N_3071,N_2084);
or U7849 (N_7849,N_2369,N_192);
xnor U7850 (N_7850,N_1760,N_1358);
nor U7851 (N_7851,N_3318,N_1207);
and U7852 (N_7852,N_1184,N_1119);
and U7853 (N_7853,N_1566,N_2531);
and U7854 (N_7854,N_737,N_1849);
and U7855 (N_7855,N_3957,N_1524);
and U7856 (N_7856,N_521,N_869);
or U7857 (N_7857,N_2809,N_3547);
nor U7858 (N_7858,N_990,N_315);
nor U7859 (N_7859,N_4252,N_4481);
nor U7860 (N_7860,N_1684,N_3370);
nor U7861 (N_7861,N_347,N_4440);
and U7862 (N_7862,N_1485,N_1867);
nor U7863 (N_7863,N_3431,N_2917);
nor U7864 (N_7864,N_186,N_1967);
nor U7865 (N_7865,N_4766,N_2966);
and U7866 (N_7866,N_327,N_1459);
xnor U7867 (N_7867,N_4234,N_2911);
nand U7868 (N_7868,N_4722,N_4844);
nand U7869 (N_7869,N_427,N_2845);
nand U7870 (N_7870,N_4387,N_3077);
xor U7871 (N_7871,N_124,N_2336);
or U7872 (N_7872,N_4618,N_1566);
and U7873 (N_7873,N_2694,N_400);
or U7874 (N_7874,N_3053,N_971);
nand U7875 (N_7875,N_1719,N_1434);
and U7876 (N_7876,N_1355,N_2030);
and U7877 (N_7877,N_754,N_931);
and U7878 (N_7878,N_4691,N_4957);
nor U7879 (N_7879,N_2864,N_569);
or U7880 (N_7880,N_4268,N_1259);
nor U7881 (N_7881,N_4468,N_4350);
or U7882 (N_7882,N_6,N_4096);
xor U7883 (N_7883,N_2068,N_818);
nor U7884 (N_7884,N_3680,N_3787);
and U7885 (N_7885,N_2167,N_2679);
and U7886 (N_7886,N_3818,N_1518);
nor U7887 (N_7887,N_381,N_4599);
xor U7888 (N_7888,N_2470,N_1943);
nand U7889 (N_7889,N_4668,N_857);
or U7890 (N_7890,N_1354,N_2066);
nand U7891 (N_7891,N_2544,N_1485);
nand U7892 (N_7892,N_2118,N_2527);
or U7893 (N_7893,N_4558,N_1740);
or U7894 (N_7894,N_179,N_2578);
nand U7895 (N_7895,N_276,N_4366);
and U7896 (N_7896,N_1203,N_4086);
xnor U7897 (N_7897,N_456,N_1929);
and U7898 (N_7898,N_2666,N_2114);
nor U7899 (N_7899,N_2068,N_2776);
or U7900 (N_7900,N_1330,N_62);
or U7901 (N_7901,N_2109,N_1580);
or U7902 (N_7902,N_121,N_4814);
and U7903 (N_7903,N_1212,N_522);
nand U7904 (N_7904,N_3888,N_4329);
and U7905 (N_7905,N_50,N_4519);
nor U7906 (N_7906,N_4213,N_4992);
nand U7907 (N_7907,N_1314,N_3195);
or U7908 (N_7908,N_2646,N_2520);
and U7909 (N_7909,N_3748,N_2202);
nor U7910 (N_7910,N_1729,N_459);
xor U7911 (N_7911,N_1289,N_4054);
nor U7912 (N_7912,N_1049,N_4204);
or U7913 (N_7913,N_4248,N_2269);
xnor U7914 (N_7914,N_4993,N_1279);
or U7915 (N_7915,N_760,N_5);
nand U7916 (N_7916,N_1144,N_2413);
nor U7917 (N_7917,N_98,N_2196);
and U7918 (N_7918,N_4366,N_1404);
or U7919 (N_7919,N_4555,N_3346);
and U7920 (N_7920,N_276,N_1921);
nand U7921 (N_7921,N_4692,N_1715);
nand U7922 (N_7922,N_3254,N_1432);
xor U7923 (N_7923,N_323,N_1760);
nand U7924 (N_7924,N_67,N_732);
and U7925 (N_7925,N_2751,N_3529);
and U7926 (N_7926,N_4224,N_2038);
nand U7927 (N_7927,N_1284,N_4520);
nand U7928 (N_7928,N_4499,N_4430);
nand U7929 (N_7929,N_1819,N_837);
nor U7930 (N_7930,N_119,N_4187);
or U7931 (N_7931,N_1290,N_2783);
and U7932 (N_7932,N_2368,N_1687);
nor U7933 (N_7933,N_1348,N_1701);
nand U7934 (N_7934,N_954,N_703);
and U7935 (N_7935,N_4366,N_344);
nor U7936 (N_7936,N_607,N_1898);
and U7937 (N_7937,N_527,N_1372);
nor U7938 (N_7938,N_4995,N_4362);
nand U7939 (N_7939,N_1125,N_2621);
nand U7940 (N_7940,N_4661,N_3483);
nor U7941 (N_7941,N_2881,N_1888);
or U7942 (N_7942,N_3626,N_744);
nand U7943 (N_7943,N_441,N_1233);
nand U7944 (N_7944,N_2490,N_1288);
and U7945 (N_7945,N_4463,N_536);
nand U7946 (N_7946,N_2634,N_793);
and U7947 (N_7947,N_3486,N_2480);
and U7948 (N_7948,N_813,N_4244);
nor U7949 (N_7949,N_4275,N_2143);
and U7950 (N_7950,N_3148,N_5);
nor U7951 (N_7951,N_606,N_1572);
or U7952 (N_7952,N_376,N_3223);
and U7953 (N_7953,N_4559,N_3447);
xnor U7954 (N_7954,N_2654,N_4887);
nor U7955 (N_7955,N_3962,N_2067);
xor U7956 (N_7956,N_783,N_2941);
or U7957 (N_7957,N_4034,N_4548);
or U7958 (N_7958,N_4453,N_3820);
nor U7959 (N_7959,N_201,N_937);
or U7960 (N_7960,N_4767,N_2885);
and U7961 (N_7961,N_4351,N_964);
and U7962 (N_7962,N_1628,N_3610);
and U7963 (N_7963,N_2233,N_2820);
and U7964 (N_7964,N_3690,N_3949);
xnor U7965 (N_7965,N_2374,N_1703);
nand U7966 (N_7966,N_83,N_4875);
and U7967 (N_7967,N_2267,N_3761);
and U7968 (N_7968,N_671,N_1853);
nand U7969 (N_7969,N_4826,N_2156);
or U7970 (N_7970,N_2326,N_4902);
nor U7971 (N_7971,N_3829,N_572);
or U7972 (N_7972,N_633,N_575);
and U7973 (N_7973,N_2929,N_2422);
or U7974 (N_7974,N_2807,N_8);
and U7975 (N_7975,N_2935,N_4146);
nor U7976 (N_7976,N_3475,N_1209);
or U7977 (N_7977,N_2501,N_3777);
and U7978 (N_7978,N_240,N_2496);
nand U7979 (N_7979,N_4493,N_1659);
and U7980 (N_7980,N_1574,N_2941);
or U7981 (N_7981,N_4393,N_4389);
or U7982 (N_7982,N_3685,N_4996);
and U7983 (N_7983,N_2347,N_1022);
nand U7984 (N_7984,N_2265,N_3318);
or U7985 (N_7985,N_4340,N_2847);
nand U7986 (N_7986,N_423,N_124);
nor U7987 (N_7987,N_3088,N_3086);
nor U7988 (N_7988,N_4099,N_1277);
xnor U7989 (N_7989,N_3085,N_1806);
and U7990 (N_7990,N_390,N_1037);
or U7991 (N_7991,N_2830,N_3739);
xor U7992 (N_7992,N_2347,N_1220);
nand U7993 (N_7993,N_3118,N_3792);
or U7994 (N_7994,N_3690,N_3713);
xor U7995 (N_7995,N_3324,N_32);
nand U7996 (N_7996,N_3201,N_1861);
xnor U7997 (N_7997,N_2554,N_2551);
nor U7998 (N_7998,N_889,N_1370);
and U7999 (N_7999,N_346,N_4572);
nand U8000 (N_8000,N_3115,N_513);
nor U8001 (N_8001,N_4072,N_334);
nor U8002 (N_8002,N_3272,N_2542);
nand U8003 (N_8003,N_3118,N_3);
nor U8004 (N_8004,N_962,N_1460);
or U8005 (N_8005,N_1332,N_568);
nor U8006 (N_8006,N_3284,N_2283);
or U8007 (N_8007,N_660,N_3163);
and U8008 (N_8008,N_387,N_3563);
and U8009 (N_8009,N_211,N_257);
nor U8010 (N_8010,N_3922,N_3791);
xnor U8011 (N_8011,N_4935,N_3755);
nor U8012 (N_8012,N_4767,N_4803);
and U8013 (N_8013,N_2704,N_526);
and U8014 (N_8014,N_3320,N_593);
nor U8015 (N_8015,N_9,N_1589);
and U8016 (N_8016,N_1221,N_1402);
or U8017 (N_8017,N_1847,N_496);
nand U8018 (N_8018,N_1101,N_3117);
nand U8019 (N_8019,N_2201,N_3996);
and U8020 (N_8020,N_2471,N_314);
nand U8021 (N_8021,N_2785,N_4223);
nor U8022 (N_8022,N_2676,N_2642);
or U8023 (N_8023,N_4340,N_4515);
xnor U8024 (N_8024,N_3711,N_2346);
and U8025 (N_8025,N_2853,N_2270);
or U8026 (N_8026,N_3425,N_3061);
nor U8027 (N_8027,N_255,N_858);
xnor U8028 (N_8028,N_4247,N_2318);
nor U8029 (N_8029,N_3790,N_4156);
nand U8030 (N_8030,N_1580,N_2249);
nor U8031 (N_8031,N_934,N_3879);
nor U8032 (N_8032,N_3555,N_4981);
nand U8033 (N_8033,N_1639,N_1239);
nand U8034 (N_8034,N_968,N_2006);
nor U8035 (N_8035,N_654,N_4179);
xor U8036 (N_8036,N_3490,N_1340);
and U8037 (N_8037,N_2773,N_4121);
and U8038 (N_8038,N_1392,N_2740);
xnor U8039 (N_8039,N_2502,N_1769);
nand U8040 (N_8040,N_2441,N_4508);
nand U8041 (N_8041,N_2367,N_1174);
nand U8042 (N_8042,N_127,N_4785);
nor U8043 (N_8043,N_2626,N_3781);
nor U8044 (N_8044,N_2847,N_3333);
or U8045 (N_8045,N_217,N_113);
nand U8046 (N_8046,N_298,N_429);
nand U8047 (N_8047,N_4819,N_241);
and U8048 (N_8048,N_4428,N_4597);
nor U8049 (N_8049,N_798,N_2587);
and U8050 (N_8050,N_2703,N_3403);
or U8051 (N_8051,N_4787,N_2662);
and U8052 (N_8052,N_1350,N_3928);
and U8053 (N_8053,N_171,N_4963);
nand U8054 (N_8054,N_624,N_2464);
xor U8055 (N_8055,N_48,N_2513);
nand U8056 (N_8056,N_1688,N_3537);
or U8057 (N_8057,N_756,N_2257);
nor U8058 (N_8058,N_1400,N_2331);
or U8059 (N_8059,N_475,N_3011);
nand U8060 (N_8060,N_3125,N_1898);
nor U8061 (N_8061,N_2918,N_2824);
xor U8062 (N_8062,N_585,N_4354);
nor U8063 (N_8063,N_945,N_2117);
or U8064 (N_8064,N_3577,N_903);
or U8065 (N_8065,N_2035,N_4645);
nor U8066 (N_8066,N_2330,N_1563);
nand U8067 (N_8067,N_725,N_1927);
and U8068 (N_8068,N_1966,N_880);
or U8069 (N_8069,N_4215,N_3935);
nor U8070 (N_8070,N_1836,N_2623);
nor U8071 (N_8071,N_4106,N_4623);
and U8072 (N_8072,N_3868,N_2654);
xnor U8073 (N_8073,N_2142,N_2851);
or U8074 (N_8074,N_1644,N_4832);
nand U8075 (N_8075,N_775,N_695);
and U8076 (N_8076,N_720,N_4659);
and U8077 (N_8077,N_44,N_903);
nor U8078 (N_8078,N_3015,N_1954);
xor U8079 (N_8079,N_298,N_4809);
nor U8080 (N_8080,N_666,N_4667);
nor U8081 (N_8081,N_2385,N_1823);
xor U8082 (N_8082,N_4433,N_1148);
or U8083 (N_8083,N_1970,N_4533);
and U8084 (N_8084,N_3889,N_4415);
nand U8085 (N_8085,N_927,N_2291);
nor U8086 (N_8086,N_2576,N_56);
nor U8087 (N_8087,N_4088,N_1581);
nand U8088 (N_8088,N_3522,N_2101);
and U8089 (N_8089,N_3882,N_4109);
nor U8090 (N_8090,N_3472,N_3587);
or U8091 (N_8091,N_2092,N_4511);
xnor U8092 (N_8092,N_2877,N_3846);
or U8093 (N_8093,N_1472,N_294);
and U8094 (N_8094,N_302,N_3183);
and U8095 (N_8095,N_3208,N_3585);
or U8096 (N_8096,N_2328,N_1588);
nor U8097 (N_8097,N_1150,N_25);
xnor U8098 (N_8098,N_2449,N_182);
and U8099 (N_8099,N_2379,N_2449);
or U8100 (N_8100,N_3296,N_4407);
nor U8101 (N_8101,N_1826,N_2230);
or U8102 (N_8102,N_2964,N_1251);
or U8103 (N_8103,N_3040,N_2766);
nand U8104 (N_8104,N_3151,N_1558);
and U8105 (N_8105,N_1308,N_151);
nand U8106 (N_8106,N_4340,N_2425);
or U8107 (N_8107,N_2824,N_3961);
nor U8108 (N_8108,N_4489,N_923);
xnor U8109 (N_8109,N_1461,N_2811);
nand U8110 (N_8110,N_2747,N_2491);
and U8111 (N_8111,N_538,N_1383);
xor U8112 (N_8112,N_3620,N_1493);
or U8113 (N_8113,N_1816,N_4745);
nand U8114 (N_8114,N_3146,N_737);
nand U8115 (N_8115,N_1494,N_1896);
and U8116 (N_8116,N_597,N_3649);
nor U8117 (N_8117,N_1868,N_3918);
and U8118 (N_8118,N_4639,N_516);
nor U8119 (N_8119,N_1791,N_3212);
nand U8120 (N_8120,N_2031,N_4742);
nor U8121 (N_8121,N_3035,N_4324);
or U8122 (N_8122,N_3905,N_4783);
and U8123 (N_8123,N_3047,N_1193);
and U8124 (N_8124,N_1021,N_730);
and U8125 (N_8125,N_4926,N_184);
or U8126 (N_8126,N_4557,N_219);
nand U8127 (N_8127,N_4944,N_3637);
nor U8128 (N_8128,N_4644,N_2372);
nand U8129 (N_8129,N_193,N_2744);
nand U8130 (N_8130,N_1412,N_4692);
and U8131 (N_8131,N_4012,N_3819);
and U8132 (N_8132,N_4416,N_4690);
nand U8133 (N_8133,N_1934,N_969);
or U8134 (N_8134,N_4264,N_4230);
nor U8135 (N_8135,N_4619,N_4583);
or U8136 (N_8136,N_1509,N_4640);
xor U8137 (N_8137,N_993,N_4932);
nor U8138 (N_8138,N_2221,N_1563);
nor U8139 (N_8139,N_1564,N_4465);
nor U8140 (N_8140,N_2758,N_401);
and U8141 (N_8141,N_2299,N_4981);
nor U8142 (N_8142,N_563,N_3819);
nand U8143 (N_8143,N_2755,N_4451);
nand U8144 (N_8144,N_773,N_3325);
nand U8145 (N_8145,N_3897,N_2154);
nand U8146 (N_8146,N_2080,N_4756);
nand U8147 (N_8147,N_346,N_1820);
and U8148 (N_8148,N_3011,N_4519);
or U8149 (N_8149,N_536,N_1347);
nand U8150 (N_8150,N_3582,N_3141);
nor U8151 (N_8151,N_3193,N_4032);
nor U8152 (N_8152,N_3596,N_611);
nor U8153 (N_8153,N_1300,N_1555);
and U8154 (N_8154,N_3977,N_3275);
nand U8155 (N_8155,N_1428,N_1383);
or U8156 (N_8156,N_3431,N_4262);
nor U8157 (N_8157,N_2873,N_4900);
or U8158 (N_8158,N_3563,N_3604);
nor U8159 (N_8159,N_718,N_2696);
or U8160 (N_8160,N_2411,N_608);
nor U8161 (N_8161,N_174,N_409);
or U8162 (N_8162,N_3591,N_4494);
and U8163 (N_8163,N_2943,N_4841);
and U8164 (N_8164,N_4376,N_3241);
nand U8165 (N_8165,N_2206,N_2112);
nor U8166 (N_8166,N_4620,N_3514);
or U8167 (N_8167,N_371,N_996);
xnor U8168 (N_8168,N_291,N_471);
nand U8169 (N_8169,N_1964,N_2233);
or U8170 (N_8170,N_3619,N_784);
nor U8171 (N_8171,N_504,N_2856);
nor U8172 (N_8172,N_3555,N_3659);
nor U8173 (N_8173,N_503,N_2834);
or U8174 (N_8174,N_2861,N_2212);
nand U8175 (N_8175,N_1496,N_3615);
nor U8176 (N_8176,N_860,N_3305);
or U8177 (N_8177,N_1538,N_3658);
xor U8178 (N_8178,N_2643,N_4836);
and U8179 (N_8179,N_984,N_2519);
nor U8180 (N_8180,N_2623,N_1507);
or U8181 (N_8181,N_3393,N_617);
nor U8182 (N_8182,N_3504,N_1710);
nor U8183 (N_8183,N_2195,N_3397);
nor U8184 (N_8184,N_2674,N_4607);
xnor U8185 (N_8185,N_1812,N_1029);
or U8186 (N_8186,N_2193,N_1232);
and U8187 (N_8187,N_2626,N_4150);
nor U8188 (N_8188,N_1967,N_1936);
or U8189 (N_8189,N_4074,N_1531);
nand U8190 (N_8190,N_755,N_2503);
and U8191 (N_8191,N_292,N_1233);
or U8192 (N_8192,N_2419,N_4930);
xnor U8193 (N_8193,N_4032,N_2426);
or U8194 (N_8194,N_192,N_3676);
xor U8195 (N_8195,N_2446,N_2064);
xor U8196 (N_8196,N_4726,N_181);
nor U8197 (N_8197,N_93,N_4142);
nand U8198 (N_8198,N_178,N_4664);
and U8199 (N_8199,N_3410,N_4908);
or U8200 (N_8200,N_4329,N_2891);
or U8201 (N_8201,N_2462,N_1797);
nor U8202 (N_8202,N_3493,N_110);
xor U8203 (N_8203,N_2985,N_290);
nand U8204 (N_8204,N_4490,N_3287);
or U8205 (N_8205,N_3021,N_3512);
nor U8206 (N_8206,N_415,N_2143);
xor U8207 (N_8207,N_727,N_3404);
or U8208 (N_8208,N_944,N_539);
xnor U8209 (N_8209,N_2113,N_409);
nand U8210 (N_8210,N_1301,N_1158);
nand U8211 (N_8211,N_3521,N_867);
nor U8212 (N_8212,N_1306,N_1153);
nor U8213 (N_8213,N_1176,N_468);
or U8214 (N_8214,N_3236,N_4719);
nor U8215 (N_8215,N_4890,N_2106);
nor U8216 (N_8216,N_2855,N_535);
or U8217 (N_8217,N_580,N_308);
nor U8218 (N_8218,N_1279,N_4626);
or U8219 (N_8219,N_3550,N_1373);
nor U8220 (N_8220,N_1100,N_1045);
or U8221 (N_8221,N_2711,N_4459);
or U8222 (N_8222,N_4103,N_4805);
nand U8223 (N_8223,N_4160,N_2113);
nor U8224 (N_8224,N_628,N_589);
or U8225 (N_8225,N_4968,N_4426);
nand U8226 (N_8226,N_2652,N_4940);
nor U8227 (N_8227,N_2963,N_1894);
and U8228 (N_8228,N_2667,N_3258);
nor U8229 (N_8229,N_2925,N_3489);
nor U8230 (N_8230,N_3053,N_2608);
and U8231 (N_8231,N_4129,N_2754);
and U8232 (N_8232,N_2292,N_4287);
and U8233 (N_8233,N_2604,N_275);
or U8234 (N_8234,N_1362,N_1049);
nor U8235 (N_8235,N_3095,N_3428);
or U8236 (N_8236,N_3593,N_2752);
nor U8237 (N_8237,N_3526,N_1670);
nand U8238 (N_8238,N_191,N_4753);
or U8239 (N_8239,N_4543,N_864);
and U8240 (N_8240,N_811,N_2213);
nand U8241 (N_8241,N_1418,N_3495);
or U8242 (N_8242,N_2491,N_4403);
and U8243 (N_8243,N_2693,N_4400);
and U8244 (N_8244,N_3918,N_32);
nor U8245 (N_8245,N_3347,N_2676);
or U8246 (N_8246,N_4403,N_3891);
and U8247 (N_8247,N_495,N_1391);
nor U8248 (N_8248,N_4356,N_358);
nand U8249 (N_8249,N_876,N_4616);
or U8250 (N_8250,N_4446,N_2112);
and U8251 (N_8251,N_749,N_4312);
or U8252 (N_8252,N_3140,N_2734);
and U8253 (N_8253,N_4469,N_3607);
and U8254 (N_8254,N_1131,N_357);
xnor U8255 (N_8255,N_580,N_1831);
or U8256 (N_8256,N_2404,N_3803);
and U8257 (N_8257,N_1225,N_3115);
and U8258 (N_8258,N_2341,N_1011);
or U8259 (N_8259,N_3530,N_113);
and U8260 (N_8260,N_3051,N_3898);
nor U8261 (N_8261,N_4823,N_3076);
nor U8262 (N_8262,N_2932,N_1318);
xnor U8263 (N_8263,N_811,N_629);
xnor U8264 (N_8264,N_362,N_3648);
and U8265 (N_8265,N_1113,N_300);
nand U8266 (N_8266,N_1099,N_1622);
xnor U8267 (N_8267,N_275,N_1805);
or U8268 (N_8268,N_2700,N_4405);
or U8269 (N_8269,N_1410,N_1885);
nor U8270 (N_8270,N_3508,N_2657);
xor U8271 (N_8271,N_1699,N_3220);
nor U8272 (N_8272,N_557,N_2686);
and U8273 (N_8273,N_200,N_984);
nand U8274 (N_8274,N_4247,N_983);
xnor U8275 (N_8275,N_2860,N_94);
or U8276 (N_8276,N_2085,N_2533);
nor U8277 (N_8277,N_1205,N_2068);
nor U8278 (N_8278,N_3619,N_1190);
or U8279 (N_8279,N_2918,N_2568);
nand U8280 (N_8280,N_4410,N_2396);
or U8281 (N_8281,N_4659,N_4775);
or U8282 (N_8282,N_3941,N_2952);
and U8283 (N_8283,N_329,N_772);
or U8284 (N_8284,N_2356,N_4708);
xnor U8285 (N_8285,N_280,N_3620);
or U8286 (N_8286,N_52,N_4498);
or U8287 (N_8287,N_376,N_2070);
or U8288 (N_8288,N_4014,N_1421);
or U8289 (N_8289,N_1323,N_2417);
xor U8290 (N_8290,N_2026,N_4655);
or U8291 (N_8291,N_4813,N_2284);
and U8292 (N_8292,N_3862,N_2175);
and U8293 (N_8293,N_1598,N_1501);
or U8294 (N_8294,N_1530,N_4509);
or U8295 (N_8295,N_2208,N_23);
or U8296 (N_8296,N_2760,N_3459);
or U8297 (N_8297,N_1198,N_2645);
nand U8298 (N_8298,N_3476,N_1815);
nor U8299 (N_8299,N_286,N_1598);
nand U8300 (N_8300,N_2254,N_351);
nor U8301 (N_8301,N_909,N_1760);
or U8302 (N_8302,N_3505,N_4096);
and U8303 (N_8303,N_1938,N_4480);
and U8304 (N_8304,N_2720,N_3658);
nand U8305 (N_8305,N_2166,N_3755);
nand U8306 (N_8306,N_367,N_1030);
and U8307 (N_8307,N_3957,N_3561);
nor U8308 (N_8308,N_2042,N_1937);
or U8309 (N_8309,N_2029,N_565);
nor U8310 (N_8310,N_4806,N_61);
or U8311 (N_8311,N_947,N_4115);
and U8312 (N_8312,N_3928,N_3356);
nand U8313 (N_8313,N_345,N_332);
nand U8314 (N_8314,N_600,N_2625);
nor U8315 (N_8315,N_865,N_3290);
xnor U8316 (N_8316,N_4576,N_4802);
nand U8317 (N_8317,N_4231,N_3637);
nor U8318 (N_8318,N_4880,N_2419);
nor U8319 (N_8319,N_1662,N_4982);
nand U8320 (N_8320,N_4122,N_2086);
nand U8321 (N_8321,N_4468,N_4346);
or U8322 (N_8322,N_4046,N_1994);
nand U8323 (N_8323,N_4671,N_4959);
nor U8324 (N_8324,N_3282,N_1950);
xnor U8325 (N_8325,N_3691,N_4384);
and U8326 (N_8326,N_1620,N_2191);
xor U8327 (N_8327,N_1721,N_963);
nor U8328 (N_8328,N_4015,N_1826);
nor U8329 (N_8329,N_4421,N_1912);
or U8330 (N_8330,N_4888,N_20);
nor U8331 (N_8331,N_2226,N_1197);
and U8332 (N_8332,N_2909,N_1849);
and U8333 (N_8333,N_4327,N_2576);
nor U8334 (N_8334,N_3862,N_3011);
nor U8335 (N_8335,N_664,N_4274);
nand U8336 (N_8336,N_4730,N_2884);
or U8337 (N_8337,N_4425,N_3353);
xnor U8338 (N_8338,N_2709,N_4598);
nor U8339 (N_8339,N_1950,N_455);
xnor U8340 (N_8340,N_613,N_2966);
or U8341 (N_8341,N_3484,N_1590);
xnor U8342 (N_8342,N_4027,N_3414);
nand U8343 (N_8343,N_44,N_2594);
nand U8344 (N_8344,N_3943,N_1117);
and U8345 (N_8345,N_4746,N_98);
nand U8346 (N_8346,N_4255,N_4666);
and U8347 (N_8347,N_4494,N_3296);
nand U8348 (N_8348,N_1128,N_4765);
nand U8349 (N_8349,N_622,N_2909);
nor U8350 (N_8350,N_3623,N_3296);
nor U8351 (N_8351,N_1845,N_897);
nor U8352 (N_8352,N_4218,N_2088);
and U8353 (N_8353,N_2130,N_3512);
nor U8354 (N_8354,N_1500,N_4347);
or U8355 (N_8355,N_1543,N_2873);
nand U8356 (N_8356,N_313,N_64);
nand U8357 (N_8357,N_4104,N_269);
or U8358 (N_8358,N_2831,N_3941);
or U8359 (N_8359,N_3889,N_3269);
nand U8360 (N_8360,N_3172,N_4474);
xor U8361 (N_8361,N_2845,N_1920);
nor U8362 (N_8362,N_4606,N_1363);
nand U8363 (N_8363,N_3930,N_3821);
or U8364 (N_8364,N_1854,N_780);
and U8365 (N_8365,N_362,N_2569);
and U8366 (N_8366,N_4296,N_2671);
nand U8367 (N_8367,N_4758,N_2915);
or U8368 (N_8368,N_1832,N_4016);
nor U8369 (N_8369,N_4466,N_3002);
nand U8370 (N_8370,N_2743,N_822);
nor U8371 (N_8371,N_4988,N_4580);
and U8372 (N_8372,N_3723,N_971);
or U8373 (N_8373,N_2725,N_1224);
and U8374 (N_8374,N_2105,N_1489);
xor U8375 (N_8375,N_2069,N_3485);
nor U8376 (N_8376,N_3604,N_4669);
and U8377 (N_8377,N_955,N_503);
and U8378 (N_8378,N_1428,N_2278);
nand U8379 (N_8379,N_4392,N_1762);
and U8380 (N_8380,N_1712,N_3804);
and U8381 (N_8381,N_466,N_346);
and U8382 (N_8382,N_646,N_2973);
or U8383 (N_8383,N_900,N_402);
xor U8384 (N_8384,N_3791,N_1470);
nand U8385 (N_8385,N_1591,N_1518);
or U8386 (N_8386,N_4696,N_746);
nand U8387 (N_8387,N_2868,N_1232);
or U8388 (N_8388,N_4279,N_2463);
or U8389 (N_8389,N_23,N_3466);
nand U8390 (N_8390,N_3555,N_1377);
or U8391 (N_8391,N_3233,N_3481);
and U8392 (N_8392,N_1308,N_815);
nor U8393 (N_8393,N_4376,N_3877);
or U8394 (N_8394,N_1741,N_3829);
and U8395 (N_8395,N_869,N_824);
and U8396 (N_8396,N_1686,N_3962);
or U8397 (N_8397,N_1419,N_1396);
and U8398 (N_8398,N_1459,N_2674);
nor U8399 (N_8399,N_2682,N_86);
nand U8400 (N_8400,N_2489,N_4810);
nand U8401 (N_8401,N_4656,N_3653);
or U8402 (N_8402,N_4274,N_1334);
xnor U8403 (N_8403,N_2770,N_2268);
or U8404 (N_8404,N_1752,N_4509);
nand U8405 (N_8405,N_3360,N_628);
or U8406 (N_8406,N_1449,N_2811);
xor U8407 (N_8407,N_1502,N_167);
nor U8408 (N_8408,N_2583,N_4552);
nand U8409 (N_8409,N_501,N_3454);
nor U8410 (N_8410,N_1549,N_1443);
and U8411 (N_8411,N_2932,N_1149);
nor U8412 (N_8412,N_3594,N_4261);
and U8413 (N_8413,N_2101,N_917);
nor U8414 (N_8414,N_3117,N_835);
nor U8415 (N_8415,N_2669,N_3956);
or U8416 (N_8416,N_2692,N_361);
xnor U8417 (N_8417,N_3383,N_778);
and U8418 (N_8418,N_4404,N_283);
or U8419 (N_8419,N_3361,N_3092);
and U8420 (N_8420,N_3993,N_3595);
nor U8421 (N_8421,N_1182,N_292);
and U8422 (N_8422,N_4385,N_4734);
xor U8423 (N_8423,N_3894,N_4838);
and U8424 (N_8424,N_3399,N_4814);
nand U8425 (N_8425,N_2753,N_1636);
nor U8426 (N_8426,N_4464,N_3473);
and U8427 (N_8427,N_3883,N_3833);
nand U8428 (N_8428,N_1223,N_2550);
nor U8429 (N_8429,N_3789,N_446);
and U8430 (N_8430,N_1121,N_1479);
xor U8431 (N_8431,N_502,N_3285);
xor U8432 (N_8432,N_4745,N_1422);
nand U8433 (N_8433,N_2307,N_1406);
or U8434 (N_8434,N_3488,N_2649);
nor U8435 (N_8435,N_553,N_1154);
and U8436 (N_8436,N_2150,N_4647);
and U8437 (N_8437,N_2046,N_1554);
or U8438 (N_8438,N_4295,N_1262);
nand U8439 (N_8439,N_2522,N_1369);
nor U8440 (N_8440,N_4975,N_3459);
or U8441 (N_8441,N_1763,N_3274);
and U8442 (N_8442,N_4342,N_3162);
nor U8443 (N_8443,N_1904,N_649);
nand U8444 (N_8444,N_4775,N_3420);
or U8445 (N_8445,N_4943,N_3187);
nor U8446 (N_8446,N_1415,N_956);
nand U8447 (N_8447,N_4243,N_258);
nand U8448 (N_8448,N_4757,N_3531);
nor U8449 (N_8449,N_963,N_679);
nor U8450 (N_8450,N_3552,N_2686);
or U8451 (N_8451,N_4229,N_4521);
or U8452 (N_8452,N_4547,N_2485);
nor U8453 (N_8453,N_971,N_2136);
or U8454 (N_8454,N_3756,N_4473);
or U8455 (N_8455,N_3742,N_2851);
nand U8456 (N_8456,N_4901,N_595);
nor U8457 (N_8457,N_3867,N_3188);
and U8458 (N_8458,N_2658,N_199);
nor U8459 (N_8459,N_4308,N_3797);
and U8460 (N_8460,N_4428,N_324);
nand U8461 (N_8461,N_721,N_4007);
nor U8462 (N_8462,N_4049,N_4699);
nor U8463 (N_8463,N_4966,N_1081);
nor U8464 (N_8464,N_2321,N_1638);
nor U8465 (N_8465,N_1510,N_469);
or U8466 (N_8466,N_3820,N_1926);
xor U8467 (N_8467,N_2328,N_874);
and U8468 (N_8468,N_15,N_3399);
nor U8469 (N_8469,N_3807,N_1228);
or U8470 (N_8470,N_2561,N_4284);
nor U8471 (N_8471,N_1169,N_4027);
or U8472 (N_8472,N_3159,N_3864);
nor U8473 (N_8473,N_240,N_1055);
or U8474 (N_8474,N_4931,N_15);
nand U8475 (N_8475,N_3292,N_2000);
xnor U8476 (N_8476,N_2961,N_2173);
nand U8477 (N_8477,N_2182,N_1394);
and U8478 (N_8478,N_1668,N_1849);
nand U8479 (N_8479,N_3849,N_816);
and U8480 (N_8480,N_2108,N_4980);
or U8481 (N_8481,N_1666,N_1264);
nand U8482 (N_8482,N_2382,N_2687);
or U8483 (N_8483,N_1378,N_2916);
nand U8484 (N_8484,N_1081,N_1896);
xor U8485 (N_8485,N_1039,N_840);
or U8486 (N_8486,N_4960,N_4588);
and U8487 (N_8487,N_4612,N_3848);
or U8488 (N_8488,N_1610,N_4114);
or U8489 (N_8489,N_1840,N_4241);
or U8490 (N_8490,N_478,N_3037);
and U8491 (N_8491,N_183,N_2619);
or U8492 (N_8492,N_1267,N_3397);
nand U8493 (N_8493,N_3375,N_169);
nor U8494 (N_8494,N_1788,N_2185);
and U8495 (N_8495,N_4354,N_1046);
nand U8496 (N_8496,N_4854,N_1625);
or U8497 (N_8497,N_4895,N_1344);
and U8498 (N_8498,N_2702,N_0);
xnor U8499 (N_8499,N_3974,N_4662);
and U8500 (N_8500,N_4446,N_3929);
and U8501 (N_8501,N_2875,N_3136);
xor U8502 (N_8502,N_1814,N_1489);
nand U8503 (N_8503,N_2391,N_4351);
xor U8504 (N_8504,N_2609,N_1246);
nor U8505 (N_8505,N_395,N_1731);
nand U8506 (N_8506,N_3903,N_4511);
and U8507 (N_8507,N_2213,N_3903);
and U8508 (N_8508,N_4489,N_2580);
or U8509 (N_8509,N_1694,N_3139);
nand U8510 (N_8510,N_1045,N_4782);
or U8511 (N_8511,N_2042,N_1474);
and U8512 (N_8512,N_3846,N_372);
or U8513 (N_8513,N_4937,N_1753);
or U8514 (N_8514,N_3334,N_173);
or U8515 (N_8515,N_1323,N_894);
nand U8516 (N_8516,N_4769,N_2564);
or U8517 (N_8517,N_3965,N_1954);
or U8518 (N_8518,N_4673,N_3012);
and U8519 (N_8519,N_1160,N_4156);
and U8520 (N_8520,N_3874,N_4964);
nand U8521 (N_8521,N_2852,N_2586);
xor U8522 (N_8522,N_3431,N_1915);
xnor U8523 (N_8523,N_452,N_3894);
nor U8524 (N_8524,N_4807,N_3284);
nor U8525 (N_8525,N_3577,N_4088);
and U8526 (N_8526,N_4475,N_1440);
or U8527 (N_8527,N_4725,N_4241);
nor U8528 (N_8528,N_4048,N_1512);
and U8529 (N_8529,N_3436,N_1565);
or U8530 (N_8530,N_2014,N_827);
nor U8531 (N_8531,N_2440,N_3666);
nor U8532 (N_8532,N_3597,N_2769);
nand U8533 (N_8533,N_3551,N_4587);
nor U8534 (N_8534,N_2381,N_685);
xor U8535 (N_8535,N_884,N_441);
nand U8536 (N_8536,N_4989,N_1254);
nor U8537 (N_8537,N_4172,N_2603);
or U8538 (N_8538,N_2683,N_206);
nor U8539 (N_8539,N_3411,N_1231);
or U8540 (N_8540,N_642,N_2496);
xor U8541 (N_8541,N_2525,N_1509);
nor U8542 (N_8542,N_4273,N_2415);
or U8543 (N_8543,N_2874,N_3088);
nor U8544 (N_8544,N_3505,N_3245);
nand U8545 (N_8545,N_528,N_2066);
nand U8546 (N_8546,N_1775,N_836);
nand U8547 (N_8547,N_3878,N_2796);
nor U8548 (N_8548,N_1248,N_3593);
nor U8549 (N_8549,N_4230,N_821);
and U8550 (N_8550,N_3388,N_1999);
or U8551 (N_8551,N_440,N_176);
nand U8552 (N_8552,N_2720,N_1369);
or U8553 (N_8553,N_234,N_4908);
and U8554 (N_8554,N_932,N_3614);
or U8555 (N_8555,N_4421,N_3939);
xor U8556 (N_8556,N_1683,N_2196);
nor U8557 (N_8557,N_1852,N_4391);
nand U8558 (N_8558,N_647,N_2684);
or U8559 (N_8559,N_314,N_1565);
and U8560 (N_8560,N_3347,N_4709);
or U8561 (N_8561,N_409,N_1095);
nand U8562 (N_8562,N_1771,N_779);
nor U8563 (N_8563,N_3981,N_3966);
and U8564 (N_8564,N_1576,N_4392);
xor U8565 (N_8565,N_370,N_3244);
and U8566 (N_8566,N_3110,N_2381);
nand U8567 (N_8567,N_596,N_4560);
nand U8568 (N_8568,N_4167,N_2759);
and U8569 (N_8569,N_4874,N_4752);
nor U8570 (N_8570,N_1581,N_1533);
or U8571 (N_8571,N_952,N_1576);
or U8572 (N_8572,N_1136,N_772);
nand U8573 (N_8573,N_2763,N_1116);
and U8574 (N_8574,N_2273,N_969);
and U8575 (N_8575,N_2973,N_2197);
xnor U8576 (N_8576,N_4076,N_1151);
nor U8577 (N_8577,N_3519,N_4286);
or U8578 (N_8578,N_3693,N_1251);
nor U8579 (N_8579,N_4491,N_1326);
nand U8580 (N_8580,N_1436,N_353);
or U8581 (N_8581,N_4257,N_406);
xnor U8582 (N_8582,N_2129,N_2974);
or U8583 (N_8583,N_588,N_378);
or U8584 (N_8584,N_4248,N_3118);
or U8585 (N_8585,N_1923,N_578);
and U8586 (N_8586,N_2825,N_3377);
or U8587 (N_8587,N_790,N_4757);
nand U8588 (N_8588,N_3105,N_2779);
xor U8589 (N_8589,N_255,N_3894);
nand U8590 (N_8590,N_777,N_486);
xor U8591 (N_8591,N_4163,N_1866);
nor U8592 (N_8592,N_82,N_1747);
nand U8593 (N_8593,N_1253,N_1351);
nor U8594 (N_8594,N_138,N_2848);
nor U8595 (N_8595,N_2706,N_4861);
and U8596 (N_8596,N_1290,N_3727);
nor U8597 (N_8597,N_281,N_3546);
nor U8598 (N_8598,N_464,N_215);
and U8599 (N_8599,N_335,N_3511);
xnor U8600 (N_8600,N_1752,N_3778);
or U8601 (N_8601,N_3027,N_4455);
and U8602 (N_8602,N_3384,N_921);
nor U8603 (N_8603,N_101,N_2946);
and U8604 (N_8604,N_2908,N_3141);
xnor U8605 (N_8605,N_4757,N_2610);
and U8606 (N_8606,N_3639,N_2734);
and U8607 (N_8607,N_1445,N_1950);
and U8608 (N_8608,N_824,N_1159);
nor U8609 (N_8609,N_828,N_1187);
or U8610 (N_8610,N_3930,N_4585);
xnor U8611 (N_8611,N_523,N_1470);
or U8612 (N_8612,N_3092,N_3201);
or U8613 (N_8613,N_4798,N_4391);
nand U8614 (N_8614,N_658,N_4637);
or U8615 (N_8615,N_3895,N_2296);
nor U8616 (N_8616,N_159,N_1401);
nand U8617 (N_8617,N_4733,N_2547);
nand U8618 (N_8618,N_1394,N_349);
nor U8619 (N_8619,N_3390,N_4044);
or U8620 (N_8620,N_2891,N_4997);
nand U8621 (N_8621,N_2750,N_1546);
xor U8622 (N_8622,N_1204,N_3205);
nor U8623 (N_8623,N_2995,N_652);
or U8624 (N_8624,N_2785,N_1854);
xor U8625 (N_8625,N_1319,N_4017);
nand U8626 (N_8626,N_3115,N_3840);
or U8627 (N_8627,N_415,N_3028);
and U8628 (N_8628,N_812,N_4744);
nor U8629 (N_8629,N_2370,N_1366);
and U8630 (N_8630,N_1457,N_1051);
nor U8631 (N_8631,N_4673,N_697);
nand U8632 (N_8632,N_770,N_345);
nor U8633 (N_8633,N_3284,N_4524);
nor U8634 (N_8634,N_3146,N_2720);
and U8635 (N_8635,N_906,N_125);
nor U8636 (N_8636,N_4379,N_4270);
and U8637 (N_8637,N_3866,N_265);
xor U8638 (N_8638,N_3467,N_2731);
and U8639 (N_8639,N_3086,N_1732);
or U8640 (N_8640,N_166,N_4374);
xnor U8641 (N_8641,N_3730,N_599);
nand U8642 (N_8642,N_2189,N_3776);
and U8643 (N_8643,N_3943,N_1547);
and U8644 (N_8644,N_2058,N_219);
nand U8645 (N_8645,N_1445,N_4129);
or U8646 (N_8646,N_2882,N_323);
or U8647 (N_8647,N_1663,N_2802);
and U8648 (N_8648,N_3728,N_2345);
xnor U8649 (N_8649,N_698,N_681);
nand U8650 (N_8650,N_1103,N_2455);
nor U8651 (N_8651,N_497,N_91);
nor U8652 (N_8652,N_2812,N_204);
nor U8653 (N_8653,N_1894,N_4931);
and U8654 (N_8654,N_4225,N_3793);
nor U8655 (N_8655,N_3957,N_3035);
or U8656 (N_8656,N_4588,N_2326);
or U8657 (N_8657,N_252,N_3936);
or U8658 (N_8658,N_1736,N_1976);
nand U8659 (N_8659,N_105,N_3034);
nand U8660 (N_8660,N_3275,N_2438);
nand U8661 (N_8661,N_1568,N_2492);
nor U8662 (N_8662,N_2452,N_162);
nor U8663 (N_8663,N_4224,N_803);
or U8664 (N_8664,N_1893,N_1941);
xnor U8665 (N_8665,N_1378,N_2220);
nand U8666 (N_8666,N_1052,N_3985);
or U8667 (N_8667,N_3195,N_1362);
and U8668 (N_8668,N_1949,N_4376);
nor U8669 (N_8669,N_313,N_2251);
nand U8670 (N_8670,N_2656,N_883);
or U8671 (N_8671,N_3445,N_227);
or U8672 (N_8672,N_3902,N_3852);
nand U8673 (N_8673,N_126,N_2767);
and U8674 (N_8674,N_2381,N_2344);
and U8675 (N_8675,N_3368,N_3152);
nor U8676 (N_8676,N_4583,N_1212);
nor U8677 (N_8677,N_9,N_4333);
or U8678 (N_8678,N_66,N_3479);
nor U8679 (N_8679,N_832,N_787);
nor U8680 (N_8680,N_3470,N_3225);
nand U8681 (N_8681,N_4965,N_4146);
and U8682 (N_8682,N_2169,N_2675);
or U8683 (N_8683,N_3373,N_2149);
or U8684 (N_8684,N_4249,N_466);
nor U8685 (N_8685,N_895,N_365);
and U8686 (N_8686,N_19,N_2706);
nand U8687 (N_8687,N_2443,N_498);
and U8688 (N_8688,N_4450,N_3466);
or U8689 (N_8689,N_1370,N_1196);
or U8690 (N_8690,N_4639,N_1594);
nor U8691 (N_8691,N_2258,N_3309);
and U8692 (N_8692,N_3814,N_4096);
nor U8693 (N_8693,N_404,N_4485);
or U8694 (N_8694,N_3900,N_543);
nor U8695 (N_8695,N_3903,N_1772);
nand U8696 (N_8696,N_4808,N_1572);
nand U8697 (N_8697,N_3168,N_2174);
or U8698 (N_8698,N_1953,N_4909);
and U8699 (N_8699,N_3613,N_3125);
nand U8700 (N_8700,N_621,N_764);
nor U8701 (N_8701,N_2394,N_2628);
and U8702 (N_8702,N_2397,N_4133);
nor U8703 (N_8703,N_3814,N_4873);
nor U8704 (N_8704,N_3292,N_183);
and U8705 (N_8705,N_1849,N_3897);
or U8706 (N_8706,N_4877,N_3513);
and U8707 (N_8707,N_3610,N_1416);
or U8708 (N_8708,N_3305,N_3811);
nor U8709 (N_8709,N_424,N_476);
nor U8710 (N_8710,N_1033,N_4003);
nor U8711 (N_8711,N_2960,N_832);
or U8712 (N_8712,N_3117,N_3895);
nor U8713 (N_8713,N_2444,N_1408);
or U8714 (N_8714,N_2201,N_2798);
or U8715 (N_8715,N_2734,N_3608);
xnor U8716 (N_8716,N_2295,N_1541);
and U8717 (N_8717,N_3036,N_575);
nor U8718 (N_8718,N_2231,N_148);
nand U8719 (N_8719,N_106,N_3006);
or U8720 (N_8720,N_2469,N_3456);
xnor U8721 (N_8721,N_4433,N_3882);
or U8722 (N_8722,N_734,N_3098);
nand U8723 (N_8723,N_4513,N_238);
nand U8724 (N_8724,N_3212,N_640);
or U8725 (N_8725,N_25,N_2797);
xor U8726 (N_8726,N_225,N_1989);
nand U8727 (N_8727,N_2335,N_3428);
nor U8728 (N_8728,N_2875,N_3161);
nand U8729 (N_8729,N_4025,N_4857);
and U8730 (N_8730,N_2587,N_3889);
nand U8731 (N_8731,N_758,N_4101);
nand U8732 (N_8732,N_4750,N_4466);
nor U8733 (N_8733,N_484,N_2525);
or U8734 (N_8734,N_4312,N_776);
or U8735 (N_8735,N_1909,N_4254);
and U8736 (N_8736,N_369,N_3874);
and U8737 (N_8737,N_2037,N_4037);
xnor U8738 (N_8738,N_4661,N_1202);
and U8739 (N_8739,N_2723,N_1471);
and U8740 (N_8740,N_1567,N_3189);
or U8741 (N_8741,N_665,N_758);
or U8742 (N_8742,N_4068,N_345);
nand U8743 (N_8743,N_3934,N_4659);
nand U8744 (N_8744,N_33,N_2352);
nand U8745 (N_8745,N_438,N_3375);
nand U8746 (N_8746,N_979,N_264);
and U8747 (N_8747,N_1581,N_424);
nand U8748 (N_8748,N_3397,N_4581);
and U8749 (N_8749,N_814,N_4004);
nand U8750 (N_8750,N_4954,N_913);
or U8751 (N_8751,N_4197,N_4472);
or U8752 (N_8752,N_2314,N_695);
nand U8753 (N_8753,N_2967,N_1143);
nand U8754 (N_8754,N_1468,N_3793);
nand U8755 (N_8755,N_259,N_1033);
and U8756 (N_8756,N_4308,N_2998);
or U8757 (N_8757,N_1001,N_2055);
nor U8758 (N_8758,N_482,N_3302);
nor U8759 (N_8759,N_1259,N_2944);
nand U8760 (N_8760,N_4061,N_1600);
or U8761 (N_8761,N_557,N_3290);
and U8762 (N_8762,N_2970,N_76);
or U8763 (N_8763,N_1574,N_2981);
nor U8764 (N_8764,N_3378,N_2072);
nand U8765 (N_8765,N_3130,N_4288);
nor U8766 (N_8766,N_3365,N_4419);
nor U8767 (N_8767,N_1723,N_3266);
and U8768 (N_8768,N_4656,N_3849);
or U8769 (N_8769,N_1583,N_887);
nand U8770 (N_8770,N_2977,N_2156);
xnor U8771 (N_8771,N_1358,N_27);
or U8772 (N_8772,N_3510,N_4888);
nor U8773 (N_8773,N_1745,N_3113);
nor U8774 (N_8774,N_4873,N_879);
nand U8775 (N_8775,N_3322,N_1278);
or U8776 (N_8776,N_4748,N_4168);
nor U8777 (N_8777,N_441,N_2813);
nor U8778 (N_8778,N_153,N_1088);
or U8779 (N_8779,N_2302,N_192);
or U8780 (N_8780,N_1227,N_2490);
nand U8781 (N_8781,N_3313,N_3196);
and U8782 (N_8782,N_3526,N_1739);
xor U8783 (N_8783,N_415,N_4746);
or U8784 (N_8784,N_924,N_548);
and U8785 (N_8785,N_3142,N_2695);
or U8786 (N_8786,N_732,N_10);
nor U8787 (N_8787,N_3522,N_2043);
nand U8788 (N_8788,N_2365,N_1463);
and U8789 (N_8789,N_839,N_4312);
or U8790 (N_8790,N_684,N_1969);
or U8791 (N_8791,N_2557,N_1236);
xor U8792 (N_8792,N_2461,N_1671);
nand U8793 (N_8793,N_85,N_2700);
xnor U8794 (N_8794,N_4834,N_4242);
nor U8795 (N_8795,N_1011,N_4917);
or U8796 (N_8796,N_87,N_899);
nor U8797 (N_8797,N_3490,N_4396);
nor U8798 (N_8798,N_896,N_928);
xnor U8799 (N_8799,N_200,N_326);
nand U8800 (N_8800,N_4040,N_3021);
nand U8801 (N_8801,N_667,N_4024);
or U8802 (N_8802,N_1746,N_1213);
or U8803 (N_8803,N_1746,N_3000);
or U8804 (N_8804,N_1180,N_2255);
nand U8805 (N_8805,N_970,N_3055);
nand U8806 (N_8806,N_2190,N_3217);
nor U8807 (N_8807,N_3955,N_3287);
nand U8808 (N_8808,N_4465,N_802);
nand U8809 (N_8809,N_1602,N_4351);
nor U8810 (N_8810,N_1727,N_2224);
nor U8811 (N_8811,N_4021,N_2701);
nor U8812 (N_8812,N_2427,N_4888);
nor U8813 (N_8813,N_4238,N_3352);
and U8814 (N_8814,N_3231,N_653);
xor U8815 (N_8815,N_4503,N_4213);
nand U8816 (N_8816,N_989,N_746);
or U8817 (N_8817,N_807,N_2906);
nand U8818 (N_8818,N_504,N_2677);
or U8819 (N_8819,N_1184,N_1581);
or U8820 (N_8820,N_4488,N_2175);
nor U8821 (N_8821,N_1764,N_4151);
nand U8822 (N_8822,N_4435,N_3698);
nand U8823 (N_8823,N_4130,N_3853);
nand U8824 (N_8824,N_1759,N_4807);
and U8825 (N_8825,N_4639,N_721);
nand U8826 (N_8826,N_4823,N_2333);
nand U8827 (N_8827,N_4464,N_3484);
or U8828 (N_8828,N_1416,N_2771);
and U8829 (N_8829,N_260,N_4297);
nor U8830 (N_8830,N_4844,N_656);
xnor U8831 (N_8831,N_1705,N_2318);
or U8832 (N_8832,N_4313,N_631);
nand U8833 (N_8833,N_270,N_1705);
xor U8834 (N_8834,N_3508,N_3217);
and U8835 (N_8835,N_4987,N_2147);
nand U8836 (N_8836,N_1725,N_2167);
nor U8837 (N_8837,N_3462,N_3634);
nand U8838 (N_8838,N_12,N_2095);
or U8839 (N_8839,N_1067,N_4471);
and U8840 (N_8840,N_180,N_4405);
nand U8841 (N_8841,N_1154,N_3939);
or U8842 (N_8842,N_4111,N_365);
nand U8843 (N_8843,N_3084,N_2907);
xnor U8844 (N_8844,N_2275,N_1386);
and U8845 (N_8845,N_4741,N_2830);
xor U8846 (N_8846,N_1706,N_121);
nand U8847 (N_8847,N_64,N_3359);
and U8848 (N_8848,N_2849,N_2884);
nor U8849 (N_8849,N_4705,N_738);
or U8850 (N_8850,N_2759,N_3273);
and U8851 (N_8851,N_1019,N_4223);
and U8852 (N_8852,N_156,N_2394);
or U8853 (N_8853,N_3195,N_51);
nand U8854 (N_8854,N_1984,N_1068);
and U8855 (N_8855,N_3556,N_663);
xnor U8856 (N_8856,N_3586,N_2354);
nand U8857 (N_8857,N_547,N_4316);
nand U8858 (N_8858,N_552,N_3009);
nand U8859 (N_8859,N_304,N_3035);
and U8860 (N_8860,N_2586,N_840);
nand U8861 (N_8861,N_1787,N_3061);
nor U8862 (N_8862,N_203,N_3464);
and U8863 (N_8863,N_1966,N_2572);
or U8864 (N_8864,N_3451,N_829);
nor U8865 (N_8865,N_3508,N_3125);
and U8866 (N_8866,N_4165,N_3087);
and U8867 (N_8867,N_2498,N_2702);
nand U8868 (N_8868,N_2834,N_274);
and U8869 (N_8869,N_970,N_3468);
or U8870 (N_8870,N_2850,N_127);
nand U8871 (N_8871,N_3898,N_3160);
nand U8872 (N_8872,N_3443,N_2479);
and U8873 (N_8873,N_4175,N_727);
xor U8874 (N_8874,N_679,N_4017);
nand U8875 (N_8875,N_1524,N_56);
nand U8876 (N_8876,N_155,N_2877);
nand U8877 (N_8877,N_1815,N_474);
or U8878 (N_8878,N_248,N_4744);
xor U8879 (N_8879,N_2607,N_1187);
nand U8880 (N_8880,N_3595,N_4509);
nor U8881 (N_8881,N_1592,N_3926);
and U8882 (N_8882,N_842,N_2290);
and U8883 (N_8883,N_469,N_2065);
or U8884 (N_8884,N_2799,N_1642);
xnor U8885 (N_8885,N_2176,N_4483);
and U8886 (N_8886,N_4042,N_1382);
and U8887 (N_8887,N_883,N_1647);
nor U8888 (N_8888,N_3244,N_448);
nand U8889 (N_8889,N_1349,N_1681);
and U8890 (N_8890,N_3546,N_4039);
and U8891 (N_8891,N_1849,N_486);
nand U8892 (N_8892,N_2609,N_3553);
nand U8893 (N_8893,N_4470,N_2840);
nor U8894 (N_8894,N_3962,N_2390);
or U8895 (N_8895,N_4902,N_2498);
nor U8896 (N_8896,N_1983,N_3020);
nor U8897 (N_8897,N_1883,N_2222);
or U8898 (N_8898,N_1124,N_2293);
nor U8899 (N_8899,N_744,N_1663);
nor U8900 (N_8900,N_4426,N_4050);
nand U8901 (N_8901,N_1249,N_1121);
and U8902 (N_8902,N_1155,N_3769);
or U8903 (N_8903,N_2755,N_2327);
nor U8904 (N_8904,N_1678,N_4515);
nand U8905 (N_8905,N_244,N_2326);
or U8906 (N_8906,N_1341,N_2941);
nor U8907 (N_8907,N_3536,N_2407);
and U8908 (N_8908,N_780,N_2457);
nand U8909 (N_8909,N_4404,N_1779);
nor U8910 (N_8910,N_3190,N_3345);
nand U8911 (N_8911,N_1420,N_780);
and U8912 (N_8912,N_4708,N_2270);
and U8913 (N_8913,N_376,N_3375);
nand U8914 (N_8914,N_3078,N_3883);
and U8915 (N_8915,N_763,N_3998);
and U8916 (N_8916,N_157,N_1100);
nor U8917 (N_8917,N_2545,N_1243);
and U8918 (N_8918,N_1920,N_1236);
or U8919 (N_8919,N_721,N_4453);
nand U8920 (N_8920,N_4717,N_1430);
xor U8921 (N_8921,N_232,N_215);
and U8922 (N_8922,N_4849,N_348);
and U8923 (N_8923,N_2899,N_2554);
and U8924 (N_8924,N_1838,N_3070);
nand U8925 (N_8925,N_1936,N_3636);
and U8926 (N_8926,N_1076,N_2409);
and U8927 (N_8927,N_3287,N_3724);
nand U8928 (N_8928,N_2198,N_802);
or U8929 (N_8929,N_4428,N_3196);
nor U8930 (N_8930,N_1073,N_4568);
nand U8931 (N_8931,N_3853,N_3782);
nor U8932 (N_8932,N_2835,N_1783);
nand U8933 (N_8933,N_3881,N_3671);
nor U8934 (N_8934,N_2232,N_1530);
or U8935 (N_8935,N_2299,N_1923);
nand U8936 (N_8936,N_483,N_387);
xor U8937 (N_8937,N_2308,N_3031);
and U8938 (N_8938,N_2539,N_1993);
nor U8939 (N_8939,N_2858,N_3678);
nor U8940 (N_8940,N_167,N_4102);
and U8941 (N_8941,N_2248,N_4802);
nor U8942 (N_8942,N_2334,N_2749);
or U8943 (N_8943,N_3477,N_1573);
or U8944 (N_8944,N_3384,N_2028);
nand U8945 (N_8945,N_3750,N_1422);
nand U8946 (N_8946,N_391,N_899);
nor U8947 (N_8947,N_2400,N_303);
or U8948 (N_8948,N_4612,N_154);
and U8949 (N_8949,N_1326,N_2661);
nor U8950 (N_8950,N_836,N_1210);
or U8951 (N_8951,N_2042,N_2290);
or U8952 (N_8952,N_2459,N_2369);
or U8953 (N_8953,N_4350,N_1302);
nand U8954 (N_8954,N_3016,N_4156);
or U8955 (N_8955,N_3980,N_4006);
or U8956 (N_8956,N_3493,N_2388);
and U8957 (N_8957,N_1330,N_4267);
nor U8958 (N_8958,N_1663,N_317);
nand U8959 (N_8959,N_325,N_106);
xnor U8960 (N_8960,N_1737,N_2623);
and U8961 (N_8961,N_4496,N_3561);
nand U8962 (N_8962,N_4465,N_3867);
nand U8963 (N_8963,N_4574,N_806);
nand U8964 (N_8964,N_3127,N_4999);
or U8965 (N_8965,N_4031,N_2519);
and U8966 (N_8966,N_28,N_1258);
nor U8967 (N_8967,N_4233,N_475);
or U8968 (N_8968,N_2211,N_4890);
nand U8969 (N_8969,N_2897,N_1591);
nor U8970 (N_8970,N_4166,N_4260);
nor U8971 (N_8971,N_4847,N_3358);
or U8972 (N_8972,N_2062,N_3373);
or U8973 (N_8973,N_1248,N_499);
or U8974 (N_8974,N_1329,N_498);
or U8975 (N_8975,N_352,N_1299);
and U8976 (N_8976,N_2185,N_3575);
and U8977 (N_8977,N_4994,N_815);
or U8978 (N_8978,N_4116,N_227);
and U8979 (N_8979,N_4276,N_2404);
nor U8980 (N_8980,N_2247,N_4944);
and U8981 (N_8981,N_4406,N_730);
nand U8982 (N_8982,N_4959,N_2959);
nand U8983 (N_8983,N_80,N_888);
or U8984 (N_8984,N_1367,N_3633);
or U8985 (N_8985,N_2906,N_1076);
or U8986 (N_8986,N_2360,N_2828);
or U8987 (N_8987,N_2861,N_4668);
or U8988 (N_8988,N_4928,N_4579);
nand U8989 (N_8989,N_1408,N_4377);
nor U8990 (N_8990,N_2199,N_3446);
or U8991 (N_8991,N_2850,N_1000);
or U8992 (N_8992,N_1376,N_1968);
xor U8993 (N_8993,N_453,N_3810);
and U8994 (N_8994,N_2276,N_2094);
and U8995 (N_8995,N_4540,N_3657);
or U8996 (N_8996,N_2265,N_1112);
nor U8997 (N_8997,N_1383,N_1246);
and U8998 (N_8998,N_4086,N_2067);
or U8999 (N_8999,N_2093,N_3743);
or U9000 (N_9000,N_4731,N_1025);
xnor U9001 (N_9001,N_1808,N_247);
or U9002 (N_9002,N_1903,N_3063);
or U9003 (N_9003,N_917,N_1385);
xnor U9004 (N_9004,N_4451,N_3493);
or U9005 (N_9005,N_1751,N_1884);
nor U9006 (N_9006,N_2403,N_317);
xor U9007 (N_9007,N_3817,N_4604);
and U9008 (N_9008,N_3911,N_2662);
and U9009 (N_9009,N_4870,N_1522);
and U9010 (N_9010,N_970,N_2016);
nor U9011 (N_9011,N_3275,N_163);
or U9012 (N_9012,N_809,N_4655);
xor U9013 (N_9013,N_1683,N_2894);
nand U9014 (N_9014,N_3410,N_4129);
nor U9015 (N_9015,N_2859,N_3673);
xnor U9016 (N_9016,N_2960,N_1528);
or U9017 (N_9017,N_2238,N_1687);
nor U9018 (N_9018,N_4663,N_4340);
or U9019 (N_9019,N_3333,N_1606);
or U9020 (N_9020,N_1415,N_2814);
nor U9021 (N_9021,N_506,N_213);
or U9022 (N_9022,N_4984,N_13);
nor U9023 (N_9023,N_2113,N_3369);
nor U9024 (N_9024,N_510,N_1780);
nand U9025 (N_9025,N_4725,N_2120);
nand U9026 (N_9026,N_494,N_4385);
or U9027 (N_9027,N_3391,N_76);
nor U9028 (N_9028,N_2144,N_2722);
nand U9029 (N_9029,N_3496,N_3421);
xor U9030 (N_9030,N_3147,N_4181);
xor U9031 (N_9031,N_2569,N_3927);
or U9032 (N_9032,N_4377,N_1350);
or U9033 (N_9033,N_3277,N_1845);
and U9034 (N_9034,N_4734,N_1146);
and U9035 (N_9035,N_4617,N_2680);
and U9036 (N_9036,N_3621,N_1445);
xnor U9037 (N_9037,N_1451,N_4450);
and U9038 (N_9038,N_525,N_2909);
xor U9039 (N_9039,N_2747,N_2597);
and U9040 (N_9040,N_4831,N_2492);
or U9041 (N_9041,N_2596,N_971);
or U9042 (N_9042,N_3750,N_3177);
or U9043 (N_9043,N_4350,N_2255);
and U9044 (N_9044,N_3079,N_154);
and U9045 (N_9045,N_27,N_2381);
nand U9046 (N_9046,N_3622,N_2644);
or U9047 (N_9047,N_3379,N_220);
or U9048 (N_9048,N_809,N_819);
or U9049 (N_9049,N_3332,N_3608);
nand U9050 (N_9050,N_129,N_2726);
nor U9051 (N_9051,N_2542,N_1384);
nand U9052 (N_9052,N_4703,N_3385);
nor U9053 (N_9053,N_1901,N_3247);
and U9054 (N_9054,N_3988,N_167);
nand U9055 (N_9055,N_1449,N_4613);
or U9056 (N_9056,N_1367,N_3927);
nor U9057 (N_9057,N_1915,N_4446);
or U9058 (N_9058,N_4196,N_3535);
nand U9059 (N_9059,N_970,N_1903);
and U9060 (N_9060,N_1675,N_3954);
nand U9061 (N_9061,N_1806,N_1491);
or U9062 (N_9062,N_1131,N_4527);
nor U9063 (N_9063,N_563,N_4831);
and U9064 (N_9064,N_1778,N_3127);
or U9065 (N_9065,N_377,N_3605);
and U9066 (N_9066,N_3517,N_293);
xor U9067 (N_9067,N_3954,N_4155);
nor U9068 (N_9068,N_578,N_3070);
nand U9069 (N_9069,N_5,N_2951);
nor U9070 (N_9070,N_2802,N_739);
nor U9071 (N_9071,N_1824,N_1186);
or U9072 (N_9072,N_4913,N_1004);
or U9073 (N_9073,N_2600,N_1480);
nor U9074 (N_9074,N_4948,N_717);
and U9075 (N_9075,N_397,N_3354);
nand U9076 (N_9076,N_3866,N_3583);
nor U9077 (N_9077,N_629,N_273);
nand U9078 (N_9078,N_1017,N_4064);
nand U9079 (N_9079,N_4017,N_981);
and U9080 (N_9080,N_2244,N_2983);
and U9081 (N_9081,N_3282,N_3009);
or U9082 (N_9082,N_3574,N_212);
nor U9083 (N_9083,N_2965,N_3980);
or U9084 (N_9084,N_4727,N_3558);
nor U9085 (N_9085,N_573,N_3481);
xnor U9086 (N_9086,N_2747,N_821);
nor U9087 (N_9087,N_117,N_398);
and U9088 (N_9088,N_493,N_2823);
nor U9089 (N_9089,N_4220,N_2710);
or U9090 (N_9090,N_2689,N_294);
or U9091 (N_9091,N_3725,N_1116);
nor U9092 (N_9092,N_3809,N_4152);
nor U9093 (N_9093,N_1740,N_58);
or U9094 (N_9094,N_3100,N_1183);
nor U9095 (N_9095,N_2078,N_2444);
nor U9096 (N_9096,N_13,N_3617);
nand U9097 (N_9097,N_4669,N_1047);
nor U9098 (N_9098,N_2843,N_1636);
nand U9099 (N_9099,N_3859,N_1640);
and U9100 (N_9100,N_2624,N_3011);
nor U9101 (N_9101,N_613,N_4531);
and U9102 (N_9102,N_21,N_2062);
or U9103 (N_9103,N_322,N_3476);
nand U9104 (N_9104,N_3449,N_2231);
xnor U9105 (N_9105,N_4953,N_4441);
and U9106 (N_9106,N_4592,N_1520);
or U9107 (N_9107,N_1089,N_251);
and U9108 (N_9108,N_654,N_2299);
and U9109 (N_9109,N_3710,N_4282);
nand U9110 (N_9110,N_109,N_2572);
and U9111 (N_9111,N_3356,N_424);
and U9112 (N_9112,N_2518,N_4815);
nor U9113 (N_9113,N_1391,N_1263);
and U9114 (N_9114,N_4425,N_2975);
nor U9115 (N_9115,N_2625,N_3111);
nor U9116 (N_9116,N_2285,N_3837);
nand U9117 (N_9117,N_2061,N_227);
or U9118 (N_9118,N_2310,N_3447);
nor U9119 (N_9119,N_2346,N_1792);
nand U9120 (N_9120,N_724,N_2267);
or U9121 (N_9121,N_1097,N_283);
nand U9122 (N_9122,N_2389,N_4911);
nor U9123 (N_9123,N_3620,N_4488);
and U9124 (N_9124,N_1594,N_1073);
nand U9125 (N_9125,N_255,N_3805);
and U9126 (N_9126,N_2294,N_4712);
nand U9127 (N_9127,N_2034,N_3238);
and U9128 (N_9128,N_1588,N_3859);
nor U9129 (N_9129,N_90,N_2016);
nand U9130 (N_9130,N_4824,N_85);
and U9131 (N_9131,N_1225,N_809);
and U9132 (N_9132,N_680,N_1247);
nand U9133 (N_9133,N_2462,N_4076);
nor U9134 (N_9134,N_3147,N_3641);
nor U9135 (N_9135,N_1588,N_2355);
and U9136 (N_9136,N_1169,N_3973);
and U9137 (N_9137,N_1006,N_3781);
nor U9138 (N_9138,N_3705,N_3688);
xor U9139 (N_9139,N_3201,N_923);
and U9140 (N_9140,N_3880,N_3463);
nor U9141 (N_9141,N_3904,N_665);
and U9142 (N_9142,N_52,N_2352);
or U9143 (N_9143,N_2137,N_4943);
nor U9144 (N_9144,N_785,N_1271);
nor U9145 (N_9145,N_4092,N_3887);
nand U9146 (N_9146,N_2171,N_3731);
and U9147 (N_9147,N_2029,N_3992);
and U9148 (N_9148,N_3210,N_2933);
nor U9149 (N_9149,N_4946,N_2147);
or U9150 (N_9150,N_4071,N_348);
xnor U9151 (N_9151,N_78,N_448);
nor U9152 (N_9152,N_3438,N_732);
and U9153 (N_9153,N_3172,N_4941);
nand U9154 (N_9154,N_4664,N_1959);
and U9155 (N_9155,N_3052,N_3635);
nor U9156 (N_9156,N_1127,N_3413);
or U9157 (N_9157,N_2182,N_3252);
nand U9158 (N_9158,N_2477,N_3587);
or U9159 (N_9159,N_3564,N_2753);
and U9160 (N_9160,N_4780,N_755);
or U9161 (N_9161,N_2566,N_1937);
nand U9162 (N_9162,N_4086,N_1735);
or U9163 (N_9163,N_2875,N_1191);
nand U9164 (N_9164,N_4617,N_2105);
and U9165 (N_9165,N_238,N_1484);
and U9166 (N_9166,N_4218,N_1658);
or U9167 (N_9167,N_3682,N_4391);
or U9168 (N_9168,N_3876,N_4485);
and U9169 (N_9169,N_3949,N_4795);
nand U9170 (N_9170,N_424,N_2803);
or U9171 (N_9171,N_2458,N_2821);
or U9172 (N_9172,N_2368,N_363);
nand U9173 (N_9173,N_1339,N_832);
and U9174 (N_9174,N_3010,N_2859);
nor U9175 (N_9175,N_2992,N_4748);
and U9176 (N_9176,N_2941,N_1261);
nor U9177 (N_9177,N_3360,N_4206);
nor U9178 (N_9178,N_4232,N_91);
nand U9179 (N_9179,N_3800,N_2824);
or U9180 (N_9180,N_1521,N_1944);
and U9181 (N_9181,N_4493,N_3502);
and U9182 (N_9182,N_1668,N_3865);
or U9183 (N_9183,N_740,N_2265);
nor U9184 (N_9184,N_709,N_4791);
nor U9185 (N_9185,N_2058,N_3158);
or U9186 (N_9186,N_4635,N_3527);
nor U9187 (N_9187,N_698,N_2113);
and U9188 (N_9188,N_293,N_1514);
nor U9189 (N_9189,N_1547,N_860);
and U9190 (N_9190,N_805,N_3709);
nor U9191 (N_9191,N_4779,N_3794);
nand U9192 (N_9192,N_484,N_3910);
and U9193 (N_9193,N_329,N_4487);
or U9194 (N_9194,N_1457,N_3745);
and U9195 (N_9195,N_4799,N_4271);
or U9196 (N_9196,N_4469,N_1415);
or U9197 (N_9197,N_3573,N_1648);
xor U9198 (N_9198,N_4706,N_1511);
and U9199 (N_9199,N_2232,N_1518);
and U9200 (N_9200,N_1921,N_1940);
nand U9201 (N_9201,N_2900,N_4138);
and U9202 (N_9202,N_1820,N_1663);
xor U9203 (N_9203,N_2524,N_2773);
or U9204 (N_9204,N_4303,N_1792);
nor U9205 (N_9205,N_3073,N_2362);
and U9206 (N_9206,N_870,N_2577);
nor U9207 (N_9207,N_4361,N_1081);
or U9208 (N_9208,N_2208,N_816);
nor U9209 (N_9209,N_922,N_1251);
and U9210 (N_9210,N_596,N_2198);
and U9211 (N_9211,N_4307,N_2470);
and U9212 (N_9212,N_1990,N_3857);
or U9213 (N_9213,N_168,N_1933);
or U9214 (N_9214,N_4910,N_1617);
nor U9215 (N_9215,N_1938,N_3110);
nand U9216 (N_9216,N_1695,N_3501);
nor U9217 (N_9217,N_35,N_1620);
nor U9218 (N_9218,N_3513,N_1827);
or U9219 (N_9219,N_2523,N_1981);
nand U9220 (N_9220,N_1649,N_2934);
and U9221 (N_9221,N_1440,N_2318);
and U9222 (N_9222,N_2716,N_1237);
and U9223 (N_9223,N_4257,N_4783);
or U9224 (N_9224,N_2475,N_3560);
or U9225 (N_9225,N_4330,N_290);
nand U9226 (N_9226,N_4735,N_1769);
nand U9227 (N_9227,N_2028,N_111);
and U9228 (N_9228,N_1647,N_230);
or U9229 (N_9229,N_173,N_718);
or U9230 (N_9230,N_1621,N_4836);
nor U9231 (N_9231,N_3282,N_3643);
and U9232 (N_9232,N_3295,N_2009);
and U9233 (N_9233,N_72,N_962);
nand U9234 (N_9234,N_4965,N_4473);
or U9235 (N_9235,N_1526,N_3777);
or U9236 (N_9236,N_2719,N_4270);
nor U9237 (N_9237,N_4727,N_1920);
nor U9238 (N_9238,N_2864,N_256);
and U9239 (N_9239,N_4206,N_2745);
nand U9240 (N_9240,N_1184,N_1013);
nand U9241 (N_9241,N_658,N_3898);
nand U9242 (N_9242,N_1902,N_4744);
and U9243 (N_9243,N_4062,N_271);
and U9244 (N_9244,N_3154,N_2464);
and U9245 (N_9245,N_623,N_1567);
and U9246 (N_9246,N_3808,N_4925);
nand U9247 (N_9247,N_853,N_1190);
or U9248 (N_9248,N_3777,N_4183);
nor U9249 (N_9249,N_1240,N_1225);
nand U9250 (N_9250,N_1906,N_1970);
nand U9251 (N_9251,N_2213,N_470);
or U9252 (N_9252,N_1107,N_2881);
nor U9253 (N_9253,N_2802,N_2732);
nor U9254 (N_9254,N_2337,N_3883);
xor U9255 (N_9255,N_2057,N_4602);
and U9256 (N_9256,N_2870,N_70);
or U9257 (N_9257,N_3375,N_2268);
or U9258 (N_9258,N_1427,N_584);
or U9259 (N_9259,N_107,N_3625);
and U9260 (N_9260,N_4255,N_4993);
and U9261 (N_9261,N_844,N_3899);
or U9262 (N_9262,N_707,N_3951);
or U9263 (N_9263,N_2119,N_589);
and U9264 (N_9264,N_2285,N_3204);
nor U9265 (N_9265,N_3030,N_3024);
and U9266 (N_9266,N_856,N_4882);
nor U9267 (N_9267,N_163,N_4541);
or U9268 (N_9268,N_330,N_4612);
and U9269 (N_9269,N_484,N_123);
and U9270 (N_9270,N_2612,N_3986);
nand U9271 (N_9271,N_3080,N_2596);
and U9272 (N_9272,N_4189,N_3662);
nor U9273 (N_9273,N_3418,N_1124);
or U9274 (N_9274,N_3521,N_2025);
and U9275 (N_9275,N_763,N_3843);
or U9276 (N_9276,N_4964,N_1014);
nor U9277 (N_9277,N_4025,N_3837);
nor U9278 (N_9278,N_4496,N_3499);
nor U9279 (N_9279,N_751,N_1301);
nand U9280 (N_9280,N_57,N_4162);
and U9281 (N_9281,N_387,N_4539);
and U9282 (N_9282,N_1711,N_1540);
and U9283 (N_9283,N_3060,N_1336);
and U9284 (N_9284,N_1239,N_159);
nand U9285 (N_9285,N_230,N_1361);
nor U9286 (N_9286,N_212,N_1357);
xnor U9287 (N_9287,N_3791,N_1023);
xnor U9288 (N_9288,N_1794,N_1511);
nor U9289 (N_9289,N_1748,N_2462);
xor U9290 (N_9290,N_4169,N_3393);
and U9291 (N_9291,N_2135,N_4477);
nor U9292 (N_9292,N_1773,N_934);
nand U9293 (N_9293,N_2160,N_2133);
nand U9294 (N_9294,N_3037,N_3286);
or U9295 (N_9295,N_1898,N_2731);
nand U9296 (N_9296,N_4674,N_4885);
and U9297 (N_9297,N_3370,N_1510);
nand U9298 (N_9298,N_2862,N_2669);
nand U9299 (N_9299,N_767,N_1334);
xnor U9300 (N_9300,N_2840,N_1246);
nand U9301 (N_9301,N_1090,N_291);
and U9302 (N_9302,N_2128,N_3082);
or U9303 (N_9303,N_1205,N_3570);
nor U9304 (N_9304,N_3154,N_4878);
and U9305 (N_9305,N_3225,N_4098);
xor U9306 (N_9306,N_3754,N_649);
nand U9307 (N_9307,N_69,N_894);
and U9308 (N_9308,N_2654,N_1448);
and U9309 (N_9309,N_2453,N_4608);
and U9310 (N_9310,N_4998,N_2099);
nand U9311 (N_9311,N_424,N_2423);
nand U9312 (N_9312,N_1114,N_443);
xnor U9313 (N_9313,N_2620,N_1026);
nand U9314 (N_9314,N_944,N_1771);
xnor U9315 (N_9315,N_1250,N_1236);
nand U9316 (N_9316,N_1763,N_4425);
and U9317 (N_9317,N_3202,N_3320);
nor U9318 (N_9318,N_1986,N_30);
or U9319 (N_9319,N_3451,N_2716);
and U9320 (N_9320,N_3461,N_51);
or U9321 (N_9321,N_2797,N_3413);
nand U9322 (N_9322,N_3830,N_3618);
nand U9323 (N_9323,N_2904,N_299);
or U9324 (N_9324,N_4126,N_4765);
nand U9325 (N_9325,N_625,N_694);
or U9326 (N_9326,N_1432,N_318);
nand U9327 (N_9327,N_4398,N_1615);
or U9328 (N_9328,N_2683,N_3299);
nand U9329 (N_9329,N_1691,N_4054);
nor U9330 (N_9330,N_2024,N_1218);
and U9331 (N_9331,N_4241,N_2145);
nor U9332 (N_9332,N_3858,N_3672);
nand U9333 (N_9333,N_3406,N_2673);
or U9334 (N_9334,N_4071,N_4557);
and U9335 (N_9335,N_435,N_304);
nand U9336 (N_9336,N_478,N_3865);
nand U9337 (N_9337,N_594,N_4262);
or U9338 (N_9338,N_2483,N_1846);
and U9339 (N_9339,N_3678,N_4552);
or U9340 (N_9340,N_25,N_797);
nand U9341 (N_9341,N_2654,N_4514);
or U9342 (N_9342,N_638,N_923);
and U9343 (N_9343,N_258,N_465);
or U9344 (N_9344,N_2029,N_2769);
or U9345 (N_9345,N_1138,N_4314);
nand U9346 (N_9346,N_3066,N_2665);
or U9347 (N_9347,N_632,N_1948);
or U9348 (N_9348,N_4532,N_3519);
nor U9349 (N_9349,N_2740,N_1255);
or U9350 (N_9350,N_2012,N_4676);
nor U9351 (N_9351,N_864,N_4492);
nor U9352 (N_9352,N_98,N_477);
nand U9353 (N_9353,N_1366,N_3248);
or U9354 (N_9354,N_4708,N_4227);
nand U9355 (N_9355,N_1849,N_2259);
nand U9356 (N_9356,N_2874,N_761);
and U9357 (N_9357,N_1146,N_3725);
nor U9358 (N_9358,N_1077,N_1119);
nor U9359 (N_9359,N_1601,N_2283);
nand U9360 (N_9360,N_366,N_2188);
nor U9361 (N_9361,N_2749,N_2622);
and U9362 (N_9362,N_2878,N_2512);
and U9363 (N_9363,N_1797,N_4798);
or U9364 (N_9364,N_935,N_4714);
and U9365 (N_9365,N_559,N_2917);
nand U9366 (N_9366,N_2472,N_2667);
nand U9367 (N_9367,N_4569,N_4253);
and U9368 (N_9368,N_1037,N_2131);
and U9369 (N_9369,N_3841,N_1976);
or U9370 (N_9370,N_4943,N_1827);
nor U9371 (N_9371,N_1167,N_3339);
and U9372 (N_9372,N_2828,N_3983);
and U9373 (N_9373,N_1260,N_4314);
nor U9374 (N_9374,N_1140,N_2760);
and U9375 (N_9375,N_2824,N_4435);
nor U9376 (N_9376,N_985,N_2871);
or U9377 (N_9377,N_2972,N_1263);
nand U9378 (N_9378,N_1445,N_1934);
or U9379 (N_9379,N_3181,N_216);
nor U9380 (N_9380,N_3567,N_3710);
nor U9381 (N_9381,N_2698,N_1890);
and U9382 (N_9382,N_3007,N_1937);
xnor U9383 (N_9383,N_2545,N_3930);
nand U9384 (N_9384,N_1378,N_3124);
and U9385 (N_9385,N_3277,N_646);
and U9386 (N_9386,N_2281,N_1526);
xor U9387 (N_9387,N_54,N_2760);
and U9388 (N_9388,N_1287,N_3654);
and U9389 (N_9389,N_632,N_332);
and U9390 (N_9390,N_495,N_4160);
or U9391 (N_9391,N_2765,N_2554);
nand U9392 (N_9392,N_1368,N_1835);
and U9393 (N_9393,N_2668,N_2268);
or U9394 (N_9394,N_2107,N_2715);
or U9395 (N_9395,N_2606,N_3246);
nor U9396 (N_9396,N_403,N_2160);
or U9397 (N_9397,N_932,N_2566);
nor U9398 (N_9398,N_4979,N_2432);
nor U9399 (N_9399,N_3185,N_2688);
or U9400 (N_9400,N_1676,N_3915);
and U9401 (N_9401,N_1640,N_1051);
or U9402 (N_9402,N_1022,N_4291);
and U9403 (N_9403,N_53,N_2223);
and U9404 (N_9404,N_4714,N_1752);
nand U9405 (N_9405,N_1320,N_3005);
and U9406 (N_9406,N_4709,N_1558);
xnor U9407 (N_9407,N_12,N_2781);
nor U9408 (N_9408,N_4588,N_2892);
nand U9409 (N_9409,N_4081,N_3788);
xnor U9410 (N_9410,N_536,N_2269);
nor U9411 (N_9411,N_2893,N_774);
nand U9412 (N_9412,N_3116,N_3196);
nand U9413 (N_9413,N_4054,N_2853);
or U9414 (N_9414,N_3950,N_2747);
nand U9415 (N_9415,N_820,N_1116);
nor U9416 (N_9416,N_1622,N_1815);
or U9417 (N_9417,N_3413,N_4937);
nand U9418 (N_9418,N_2618,N_3997);
and U9419 (N_9419,N_4658,N_1435);
nand U9420 (N_9420,N_2976,N_4770);
xor U9421 (N_9421,N_3095,N_3875);
nor U9422 (N_9422,N_4428,N_115);
nand U9423 (N_9423,N_1746,N_4418);
nand U9424 (N_9424,N_3638,N_3596);
nand U9425 (N_9425,N_4099,N_520);
nor U9426 (N_9426,N_3291,N_677);
and U9427 (N_9427,N_4355,N_4256);
nand U9428 (N_9428,N_1603,N_2580);
and U9429 (N_9429,N_983,N_339);
and U9430 (N_9430,N_2054,N_4318);
or U9431 (N_9431,N_3413,N_3347);
and U9432 (N_9432,N_477,N_2358);
nor U9433 (N_9433,N_1372,N_2413);
and U9434 (N_9434,N_2969,N_3060);
and U9435 (N_9435,N_63,N_4966);
nand U9436 (N_9436,N_1473,N_3721);
and U9437 (N_9437,N_2637,N_1696);
or U9438 (N_9438,N_2687,N_4493);
nor U9439 (N_9439,N_4994,N_413);
and U9440 (N_9440,N_161,N_2638);
or U9441 (N_9441,N_4369,N_1179);
or U9442 (N_9442,N_1484,N_2499);
nor U9443 (N_9443,N_3923,N_166);
and U9444 (N_9444,N_2672,N_2957);
and U9445 (N_9445,N_3082,N_4963);
nor U9446 (N_9446,N_1181,N_3965);
nor U9447 (N_9447,N_1431,N_1335);
nor U9448 (N_9448,N_539,N_4782);
and U9449 (N_9449,N_3489,N_1733);
xor U9450 (N_9450,N_3253,N_3245);
xnor U9451 (N_9451,N_1839,N_2623);
nand U9452 (N_9452,N_4979,N_3055);
xnor U9453 (N_9453,N_3234,N_3078);
or U9454 (N_9454,N_3301,N_2664);
or U9455 (N_9455,N_3527,N_2128);
nand U9456 (N_9456,N_3148,N_1239);
nand U9457 (N_9457,N_4124,N_11);
nor U9458 (N_9458,N_3394,N_3828);
and U9459 (N_9459,N_4892,N_4622);
or U9460 (N_9460,N_4000,N_4551);
and U9461 (N_9461,N_1293,N_866);
and U9462 (N_9462,N_2481,N_2347);
nor U9463 (N_9463,N_3739,N_3797);
nor U9464 (N_9464,N_443,N_2480);
nand U9465 (N_9465,N_4810,N_3817);
nor U9466 (N_9466,N_3810,N_672);
nand U9467 (N_9467,N_4188,N_3405);
nand U9468 (N_9468,N_1818,N_3777);
or U9469 (N_9469,N_428,N_1347);
nor U9470 (N_9470,N_4638,N_4016);
nor U9471 (N_9471,N_3560,N_4488);
nor U9472 (N_9472,N_2810,N_991);
or U9473 (N_9473,N_1438,N_122);
xnor U9474 (N_9474,N_4818,N_3696);
or U9475 (N_9475,N_4120,N_3846);
and U9476 (N_9476,N_441,N_988);
nor U9477 (N_9477,N_2652,N_400);
and U9478 (N_9478,N_2778,N_2639);
xor U9479 (N_9479,N_2676,N_2416);
nand U9480 (N_9480,N_2444,N_4191);
nor U9481 (N_9481,N_497,N_3289);
nor U9482 (N_9482,N_2730,N_42);
and U9483 (N_9483,N_3689,N_1749);
or U9484 (N_9484,N_3272,N_646);
or U9485 (N_9485,N_3323,N_1236);
and U9486 (N_9486,N_3762,N_1040);
nor U9487 (N_9487,N_807,N_1760);
and U9488 (N_9488,N_715,N_4507);
nand U9489 (N_9489,N_4381,N_2730);
nand U9490 (N_9490,N_1536,N_1554);
and U9491 (N_9491,N_861,N_3039);
nand U9492 (N_9492,N_4451,N_4142);
or U9493 (N_9493,N_2129,N_4175);
and U9494 (N_9494,N_141,N_147);
xor U9495 (N_9495,N_2579,N_1923);
and U9496 (N_9496,N_212,N_924);
or U9497 (N_9497,N_3689,N_1914);
nor U9498 (N_9498,N_53,N_20);
and U9499 (N_9499,N_1130,N_395);
and U9500 (N_9500,N_1160,N_4707);
xnor U9501 (N_9501,N_3510,N_4440);
and U9502 (N_9502,N_1568,N_983);
and U9503 (N_9503,N_141,N_3742);
and U9504 (N_9504,N_1016,N_3729);
or U9505 (N_9505,N_4828,N_4106);
and U9506 (N_9506,N_4888,N_4014);
nor U9507 (N_9507,N_1081,N_716);
and U9508 (N_9508,N_1736,N_3264);
nand U9509 (N_9509,N_1041,N_4435);
xnor U9510 (N_9510,N_673,N_1637);
nor U9511 (N_9511,N_3654,N_1465);
or U9512 (N_9512,N_1492,N_2778);
nand U9513 (N_9513,N_830,N_2431);
nor U9514 (N_9514,N_4136,N_4443);
or U9515 (N_9515,N_4909,N_1981);
nor U9516 (N_9516,N_3969,N_2680);
or U9517 (N_9517,N_1324,N_2732);
nand U9518 (N_9518,N_3489,N_2531);
nor U9519 (N_9519,N_3665,N_3506);
nand U9520 (N_9520,N_1777,N_2952);
and U9521 (N_9521,N_2612,N_585);
nor U9522 (N_9522,N_560,N_4808);
nor U9523 (N_9523,N_30,N_2168);
xnor U9524 (N_9524,N_3361,N_3668);
nand U9525 (N_9525,N_3386,N_3044);
or U9526 (N_9526,N_1862,N_2831);
or U9527 (N_9527,N_1982,N_1578);
xor U9528 (N_9528,N_3801,N_2031);
or U9529 (N_9529,N_1263,N_2929);
nor U9530 (N_9530,N_122,N_278);
or U9531 (N_9531,N_4456,N_2818);
nand U9532 (N_9532,N_2250,N_4144);
nand U9533 (N_9533,N_4912,N_4306);
and U9534 (N_9534,N_2952,N_83);
nand U9535 (N_9535,N_1514,N_1805);
nand U9536 (N_9536,N_3091,N_782);
and U9537 (N_9537,N_811,N_3659);
nand U9538 (N_9538,N_2039,N_493);
xor U9539 (N_9539,N_4675,N_753);
or U9540 (N_9540,N_4510,N_110);
or U9541 (N_9541,N_2498,N_1145);
or U9542 (N_9542,N_3169,N_4611);
nor U9543 (N_9543,N_2028,N_1526);
and U9544 (N_9544,N_1332,N_2456);
and U9545 (N_9545,N_2483,N_1799);
nor U9546 (N_9546,N_4452,N_4726);
or U9547 (N_9547,N_4899,N_1097);
and U9548 (N_9548,N_961,N_3611);
and U9549 (N_9549,N_3577,N_4175);
or U9550 (N_9550,N_3738,N_2699);
nand U9551 (N_9551,N_1252,N_4456);
nand U9552 (N_9552,N_1878,N_1482);
and U9553 (N_9553,N_2494,N_3390);
and U9554 (N_9554,N_4330,N_1290);
and U9555 (N_9555,N_4618,N_4500);
xnor U9556 (N_9556,N_633,N_2178);
or U9557 (N_9557,N_3433,N_2113);
nand U9558 (N_9558,N_1259,N_3578);
and U9559 (N_9559,N_2154,N_452);
or U9560 (N_9560,N_1359,N_3708);
nor U9561 (N_9561,N_4656,N_2031);
xnor U9562 (N_9562,N_509,N_658);
and U9563 (N_9563,N_3490,N_4557);
and U9564 (N_9564,N_4601,N_3008);
or U9565 (N_9565,N_476,N_2958);
or U9566 (N_9566,N_2622,N_428);
or U9567 (N_9567,N_2736,N_3030);
and U9568 (N_9568,N_2398,N_2682);
and U9569 (N_9569,N_4772,N_1342);
or U9570 (N_9570,N_1985,N_4587);
nor U9571 (N_9571,N_4335,N_4552);
xnor U9572 (N_9572,N_1642,N_2837);
nor U9573 (N_9573,N_147,N_1252);
nor U9574 (N_9574,N_358,N_2699);
xnor U9575 (N_9575,N_1024,N_2365);
and U9576 (N_9576,N_1469,N_3087);
xor U9577 (N_9577,N_1195,N_1527);
nor U9578 (N_9578,N_3728,N_1253);
nand U9579 (N_9579,N_3920,N_2319);
nor U9580 (N_9580,N_3004,N_2076);
and U9581 (N_9581,N_3159,N_20);
nor U9582 (N_9582,N_3028,N_2440);
nand U9583 (N_9583,N_990,N_3682);
nor U9584 (N_9584,N_810,N_3490);
and U9585 (N_9585,N_4010,N_2770);
xnor U9586 (N_9586,N_3227,N_3338);
nor U9587 (N_9587,N_3809,N_1648);
nor U9588 (N_9588,N_3966,N_4561);
xnor U9589 (N_9589,N_3407,N_647);
or U9590 (N_9590,N_255,N_355);
nand U9591 (N_9591,N_4386,N_3211);
and U9592 (N_9592,N_2465,N_1511);
nor U9593 (N_9593,N_196,N_2863);
or U9594 (N_9594,N_3688,N_4444);
xnor U9595 (N_9595,N_4572,N_323);
or U9596 (N_9596,N_820,N_2127);
xor U9597 (N_9597,N_1841,N_101);
and U9598 (N_9598,N_2231,N_2262);
nor U9599 (N_9599,N_4606,N_4766);
and U9600 (N_9600,N_1951,N_3133);
and U9601 (N_9601,N_543,N_483);
xor U9602 (N_9602,N_2476,N_3408);
nor U9603 (N_9603,N_1799,N_1431);
nand U9604 (N_9604,N_2160,N_851);
nand U9605 (N_9605,N_2348,N_3838);
or U9606 (N_9606,N_4259,N_3175);
or U9607 (N_9607,N_568,N_274);
nand U9608 (N_9608,N_2299,N_740);
or U9609 (N_9609,N_975,N_1387);
or U9610 (N_9610,N_4209,N_1183);
nand U9611 (N_9611,N_3889,N_3593);
xor U9612 (N_9612,N_3046,N_2810);
nand U9613 (N_9613,N_4616,N_1059);
nand U9614 (N_9614,N_1658,N_576);
nor U9615 (N_9615,N_3230,N_2160);
and U9616 (N_9616,N_4933,N_1943);
and U9617 (N_9617,N_4036,N_626);
and U9618 (N_9618,N_772,N_2996);
and U9619 (N_9619,N_4251,N_3219);
nand U9620 (N_9620,N_2168,N_2659);
nor U9621 (N_9621,N_3316,N_1045);
and U9622 (N_9622,N_116,N_1669);
or U9623 (N_9623,N_4604,N_3378);
nand U9624 (N_9624,N_1982,N_2800);
nand U9625 (N_9625,N_3897,N_2037);
and U9626 (N_9626,N_3636,N_3384);
or U9627 (N_9627,N_1479,N_1026);
and U9628 (N_9628,N_1015,N_2440);
xor U9629 (N_9629,N_619,N_1059);
nand U9630 (N_9630,N_3625,N_1625);
xnor U9631 (N_9631,N_1613,N_2439);
nand U9632 (N_9632,N_316,N_2180);
and U9633 (N_9633,N_699,N_3233);
and U9634 (N_9634,N_3318,N_643);
nand U9635 (N_9635,N_4638,N_1193);
or U9636 (N_9636,N_2554,N_3131);
and U9637 (N_9637,N_209,N_472);
nand U9638 (N_9638,N_4887,N_1478);
or U9639 (N_9639,N_4913,N_17);
nand U9640 (N_9640,N_1670,N_4410);
and U9641 (N_9641,N_4745,N_1979);
nand U9642 (N_9642,N_981,N_608);
nand U9643 (N_9643,N_881,N_4796);
xnor U9644 (N_9644,N_2104,N_3220);
or U9645 (N_9645,N_577,N_3217);
or U9646 (N_9646,N_4461,N_1550);
and U9647 (N_9647,N_903,N_388);
or U9648 (N_9648,N_1737,N_4755);
nor U9649 (N_9649,N_3887,N_2944);
and U9650 (N_9650,N_6,N_572);
and U9651 (N_9651,N_3037,N_4324);
or U9652 (N_9652,N_442,N_2306);
nor U9653 (N_9653,N_2029,N_4827);
nand U9654 (N_9654,N_2722,N_1517);
nand U9655 (N_9655,N_2429,N_2757);
and U9656 (N_9656,N_1132,N_136);
nand U9657 (N_9657,N_4998,N_380);
nand U9658 (N_9658,N_542,N_395);
nor U9659 (N_9659,N_1262,N_4282);
xor U9660 (N_9660,N_2503,N_3274);
nor U9661 (N_9661,N_203,N_7);
or U9662 (N_9662,N_900,N_3481);
nand U9663 (N_9663,N_1372,N_731);
nand U9664 (N_9664,N_4598,N_3738);
xnor U9665 (N_9665,N_524,N_4069);
and U9666 (N_9666,N_4275,N_3346);
nand U9667 (N_9667,N_324,N_4906);
nor U9668 (N_9668,N_4784,N_4922);
nor U9669 (N_9669,N_4966,N_1169);
xnor U9670 (N_9670,N_3386,N_3207);
xnor U9671 (N_9671,N_4440,N_3561);
or U9672 (N_9672,N_2490,N_811);
xor U9673 (N_9673,N_1013,N_3970);
and U9674 (N_9674,N_3511,N_3655);
xnor U9675 (N_9675,N_3361,N_4733);
nor U9676 (N_9676,N_3833,N_2390);
nor U9677 (N_9677,N_3432,N_3350);
xnor U9678 (N_9678,N_4769,N_962);
and U9679 (N_9679,N_2092,N_2143);
and U9680 (N_9680,N_3510,N_2892);
nor U9681 (N_9681,N_1067,N_3132);
or U9682 (N_9682,N_180,N_718);
nor U9683 (N_9683,N_3189,N_4812);
nor U9684 (N_9684,N_2105,N_4046);
nor U9685 (N_9685,N_876,N_4857);
nand U9686 (N_9686,N_1407,N_344);
or U9687 (N_9687,N_4708,N_2925);
nor U9688 (N_9688,N_3130,N_3279);
nand U9689 (N_9689,N_1986,N_782);
or U9690 (N_9690,N_1317,N_3372);
and U9691 (N_9691,N_3543,N_3894);
nand U9692 (N_9692,N_503,N_1402);
nor U9693 (N_9693,N_2200,N_2527);
nand U9694 (N_9694,N_4311,N_3981);
and U9695 (N_9695,N_789,N_1265);
nand U9696 (N_9696,N_328,N_1296);
or U9697 (N_9697,N_2766,N_2901);
xnor U9698 (N_9698,N_634,N_855);
or U9699 (N_9699,N_137,N_4430);
nor U9700 (N_9700,N_1848,N_1642);
and U9701 (N_9701,N_2145,N_1401);
and U9702 (N_9702,N_3601,N_1412);
and U9703 (N_9703,N_943,N_1869);
nand U9704 (N_9704,N_3400,N_3701);
or U9705 (N_9705,N_2858,N_4434);
or U9706 (N_9706,N_903,N_4169);
nor U9707 (N_9707,N_1294,N_726);
and U9708 (N_9708,N_3214,N_3565);
and U9709 (N_9709,N_4904,N_1777);
nand U9710 (N_9710,N_3896,N_4102);
or U9711 (N_9711,N_733,N_4413);
and U9712 (N_9712,N_857,N_1402);
or U9713 (N_9713,N_3420,N_3918);
nor U9714 (N_9714,N_1697,N_3385);
or U9715 (N_9715,N_3200,N_1033);
xnor U9716 (N_9716,N_2544,N_2345);
nand U9717 (N_9717,N_4386,N_4997);
nor U9718 (N_9718,N_1452,N_2475);
nand U9719 (N_9719,N_526,N_990);
xor U9720 (N_9720,N_4296,N_3412);
nand U9721 (N_9721,N_291,N_3699);
xor U9722 (N_9722,N_4685,N_77);
nor U9723 (N_9723,N_213,N_3055);
or U9724 (N_9724,N_3365,N_1409);
or U9725 (N_9725,N_3548,N_1200);
or U9726 (N_9726,N_744,N_690);
nand U9727 (N_9727,N_1347,N_3481);
nor U9728 (N_9728,N_425,N_712);
xor U9729 (N_9729,N_584,N_1508);
nor U9730 (N_9730,N_4417,N_1382);
or U9731 (N_9731,N_752,N_3626);
nand U9732 (N_9732,N_330,N_2218);
and U9733 (N_9733,N_2623,N_2079);
and U9734 (N_9734,N_2459,N_2323);
nor U9735 (N_9735,N_74,N_2670);
or U9736 (N_9736,N_1292,N_739);
nand U9737 (N_9737,N_260,N_4151);
xnor U9738 (N_9738,N_781,N_3407);
xnor U9739 (N_9739,N_4681,N_611);
and U9740 (N_9740,N_4326,N_1746);
or U9741 (N_9741,N_843,N_4829);
and U9742 (N_9742,N_964,N_4363);
and U9743 (N_9743,N_4192,N_3918);
nor U9744 (N_9744,N_2044,N_4484);
and U9745 (N_9745,N_4223,N_4125);
or U9746 (N_9746,N_659,N_1560);
or U9747 (N_9747,N_3188,N_4435);
or U9748 (N_9748,N_1134,N_543);
nand U9749 (N_9749,N_2181,N_2729);
nor U9750 (N_9750,N_3589,N_620);
or U9751 (N_9751,N_2484,N_3121);
or U9752 (N_9752,N_2452,N_1614);
xor U9753 (N_9753,N_1003,N_2556);
or U9754 (N_9754,N_2437,N_3773);
nor U9755 (N_9755,N_2330,N_1219);
or U9756 (N_9756,N_3706,N_1516);
or U9757 (N_9757,N_2350,N_813);
nand U9758 (N_9758,N_4048,N_104);
or U9759 (N_9759,N_963,N_1587);
or U9760 (N_9760,N_1966,N_3139);
xor U9761 (N_9761,N_2160,N_2596);
or U9762 (N_9762,N_112,N_4255);
nor U9763 (N_9763,N_2159,N_2308);
xor U9764 (N_9764,N_1905,N_633);
and U9765 (N_9765,N_2133,N_3520);
or U9766 (N_9766,N_4814,N_1162);
nand U9767 (N_9767,N_2019,N_1766);
nand U9768 (N_9768,N_1158,N_1630);
or U9769 (N_9769,N_1596,N_1528);
or U9770 (N_9770,N_2813,N_3486);
nor U9771 (N_9771,N_3046,N_43);
or U9772 (N_9772,N_3171,N_1656);
or U9773 (N_9773,N_2093,N_4397);
nor U9774 (N_9774,N_4985,N_2341);
nor U9775 (N_9775,N_912,N_4155);
nor U9776 (N_9776,N_1193,N_395);
xor U9777 (N_9777,N_1538,N_381);
or U9778 (N_9778,N_4062,N_1860);
or U9779 (N_9779,N_4684,N_2068);
nand U9780 (N_9780,N_2078,N_2274);
and U9781 (N_9781,N_1535,N_2726);
and U9782 (N_9782,N_4026,N_2007);
xor U9783 (N_9783,N_4915,N_4576);
nand U9784 (N_9784,N_1178,N_2264);
or U9785 (N_9785,N_1868,N_4563);
nor U9786 (N_9786,N_1525,N_703);
xor U9787 (N_9787,N_316,N_1358);
nor U9788 (N_9788,N_2435,N_4970);
nand U9789 (N_9789,N_4137,N_1105);
nand U9790 (N_9790,N_4452,N_3327);
xnor U9791 (N_9791,N_4899,N_1242);
nor U9792 (N_9792,N_4930,N_1388);
nand U9793 (N_9793,N_3462,N_3352);
or U9794 (N_9794,N_913,N_4069);
nand U9795 (N_9795,N_4300,N_1349);
nor U9796 (N_9796,N_894,N_1560);
or U9797 (N_9797,N_210,N_4021);
nor U9798 (N_9798,N_176,N_3108);
and U9799 (N_9799,N_2682,N_1296);
and U9800 (N_9800,N_3052,N_2525);
or U9801 (N_9801,N_3661,N_1147);
nand U9802 (N_9802,N_782,N_676);
xor U9803 (N_9803,N_3504,N_4737);
nor U9804 (N_9804,N_2236,N_3960);
and U9805 (N_9805,N_963,N_906);
nand U9806 (N_9806,N_1222,N_315);
or U9807 (N_9807,N_4996,N_2606);
or U9808 (N_9808,N_1458,N_3643);
nor U9809 (N_9809,N_4344,N_1973);
nor U9810 (N_9810,N_1700,N_791);
or U9811 (N_9811,N_1671,N_2155);
nor U9812 (N_9812,N_4900,N_164);
nor U9813 (N_9813,N_1294,N_1078);
nand U9814 (N_9814,N_2380,N_4370);
and U9815 (N_9815,N_2686,N_3075);
or U9816 (N_9816,N_1755,N_3304);
nor U9817 (N_9817,N_4997,N_2449);
nand U9818 (N_9818,N_749,N_3442);
and U9819 (N_9819,N_4642,N_4602);
nand U9820 (N_9820,N_2558,N_4356);
nand U9821 (N_9821,N_1369,N_1871);
nand U9822 (N_9822,N_1250,N_1116);
or U9823 (N_9823,N_3732,N_1769);
or U9824 (N_9824,N_302,N_565);
nor U9825 (N_9825,N_307,N_1093);
nor U9826 (N_9826,N_1412,N_2394);
nand U9827 (N_9827,N_4473,N_2886);
and U9828 (N_9828,N_4916,N_3260);
nor U9829 (N_9829,N_1924,N_4280);
or U9830 (N_9830,N_1872,N_1415);
nor U9831 (N_9831,N_2577,N_2554);
or U9832 (N_9832,N_1743,N_3137);
or U9833 (N_9833,N_406,N_1144);
and U9834 (N_9834,N_191,N_3344);
nand U9835 (N_9835,N_822,N_4864);
or U9836 (N_9836,N_3874,N_1905);
nand U9837 (N_9837,N_674,N_3829);
nor U9838 (N_9838,N_3248,N_1757);
nand U9839 (N_9839,N_524,N_1512);
and U9840 (N_9840,N_1583,N_1623);
nand U9841 (N_9841,N_3352,N_4492);
or U9842 (N_9842,N_2111,N_1722);
nor U9843 (N_9843,N_1014,N_3913);
xnor U9844 (N_9844,N_1244,N_1428);
nor U9845 (N_9845,N_1883,N_656);
and U9846 (N_9846,N_2456,N_2914);
nor U9847 (N_9847,N_1399,N_4186);
nand U9848 (N_9848,N_1651,N_966);
nor U9849 (N_9849,N_4442,N_1388);
and U9850 (N_9850,N_2322,N_1469);
nor U9851 (N_9851,N_466,N_4809);
xnor U9852 (N_9852,N_3617,N_1202);
or U9853 (N_9853,N_3734,N_4126);
nor U9854 (N_9854,N_2519,N_4331);
or U9855 (N_9855,N_2780,N_3264);
and U9856 (N_9856,N_979,N_1991);
or U9857 (N_9857,N_1677,N_2176);
and U9858 (N_9858,N_1444,N_1320);
or U9859 (N_9859,N_4257,N_331);
xnor U9860 (N_9860,N_652,N_1527);
or U9861 (N_9861,N_1984,N_4905);
nor U9862 (N_9862,N_4864,N_480);
nor U9863 (N_9863,N_461,N_4764);
nand U9864 (N_9864,N_1379,N_2548);
or U9865 (N_9865,N_4479,N_2125);
nand U9866 (N_9866,N_4122,N_2598);
nand U9867 (N_9867,N_4090,N_1443);
or U9868 (N_9868,N_2608,N_4003);
nor U9869 (N_9869,N_2868,N_1531);
nor U9870 (N_9870,N_4288,N_4730);
or U9871 (N_9871,N_3108,N_2065);
nand U9872 (N_9872,N_1418,N_2392);
nand U9873 (N_9873,N_2144,N_54);
or U9874 (N_9874,N_50,N_939);
xnor U9875 (N_9875,N_37,N_1838);
and U9876 (N_9876,N_420,N_1074);
nor U9877 (N_9877,N_587,N_4502);
nand U9878 (N_9878,N_3382,N_1824);
nor U9879 (N_9879,N_562,N_1660);
and U9880 (N_9880,N_4920,N_121);
or U9881 (N_9881,N_170,N_1645);
nor U9882 (N_9882,N_2645,N_4612);
and U9883 (N_9883,N_1404,N_2966);
nor U9884 (N_9884,N_3252,N_1343);
nor U9885 (N_9885,N_4898,N_181);
or U9886 (N_9886,N_2229,N_3791);
nand U9887 (N_9887,N_2695,N_4786);
or U9888 (N_9888,N_4385,N_2648);
or U9889 (N_9889,N_3130,N_227);
or U9890 (N_9890,N_1756,N_1718);
and U9891 (N_9891,N_3360,N_654);
xnor U9892 (N_9892,N_1606,N_2056);
nand U9893 (N_9893,N_4826,N_1563);
and U9894 (N_9894,N_4614,N_1439);
nor U9895 (N_9895,N_4742,N_824);
nand U9896 (N_9896,N_3914,N_842);
xor U9897 (N_9897,N_2672,N_1180);
nor U9898 (N_9898,N_4278,N_4503);
nor U9899 (N_9899,N_3212,N_3571);
or U9900 (N_9900,N_4876,N_4157);
nor U9901 (N_9901,N_3049,N_2622);
nand U9902 (N_9902,N_3828,N_162);
or U9903 (N_9903,N_4219,N_571);
or U9904 (N_9904,N_3697,N_4062);
nand U9905 (N_9905,N_696,N_2944);
nand U9906 (N_9906,N_2920,N_586);
xor U9907 (N_9907,N_503,N_2561);
and U9908 (N_9908,N_3661,N_3031);
nor U9909 (N_9909,N_4166,N_2940);
nand U9910 (N_9910,N_160,N_1350);
and U9911 (N_9911,N_1717,N_3831);
and U9912 (N_9912,N_848,N_3760);
xor U9913 (N_9913,N_4113,N_1382);
or U9914 (N_9914,N_2479,N_3295);
xor U9915 (N_9915,N_4217,N_4939);
and U9916 (N_9916,N_3508,N_1746);
or U9917 (N_9917,N_2915,N_3166);
nor U9918 (N_9918,N_1105,N_4441);
nor U9919 (N_9919,N_850,N_4753);
or U9920 (N_9920,N_2720,N_3277);
xnor U9921 (N_9921,N_2758,N_4231);
or U9922 (N_9922,N_2028,N_1352);
xnor U9923 (N_9923,N_223,N_4864);
or U9924 (N_9924,N_3170,N_4596);
nand U9925 (N_9925,N_2070,N_2626);
or U9926 (N_9926,N_477,N_2444);
or U9927 (N_9927,N_3090,N_3577);
nand U9928 (N_9928,N_2951,N_1334);
or U9929 (N_9929,N_3914,N_4017);
nand U9930 (N_9930,N_657,N_1909);
nor U9931 (N_9931,N_785,N_679);
or U9932 (N_9932,N_4532,N_3642);
nor U9933 (N_9933,N_34,N_4712);
and U9934 (N_9934,N_4543,N_3482);
or U9935 (N_9935,N_198,N_159);
nor U9936 (N_9936,N_1458,N_1429);
xnor U9937 (N_9937,N_1763,N_879);
nand U9938 (N_9938,N_1613,N_3414);
or U9939 (N_9939,N_1084,N_3031);
nand U9940 (N_9940,N_838,N_1195);
nor U9941 (N_9941,N_2325,N_424);
and U9942 (N_9942,N_2993,N_1933);
nand U9943 (N_9943,N_4909,N_4826);
and U9944 (N_9944,N_814,N_1725);
and U9945 (N_9945,N_1829,N_949);
or U9946 (N_9946,N_1196,N_1125);
or U9947 (N_9947,N_3016,N_4544);
nor U9948 (N_9948,N_3806,N_2167);
or U9949 (N_9949,N_1432,N_142);
nand U9950 (N_9950,N_4374,N_3522);
nor U9951 (N_9951,N_1608,N_3930);
nor U9952 (N_9952,N_4786,N_1128);
and U9953 (N_9953,N_437,N_1463);
or U9954 (N_9954,N_3950,N_3241);
or U9955 (N_9955,N_3689,N_647);
nor U9956 (N_9956,N_682,N_1188);
or U9957 (N_9957,N_2220,N_4091);
or U9958 (N_9958,N_218,N_4887);
nand U9959 (N_9959,N_344,N_4363);
xnor U9960 (N_9960,N_362,N_2302);
and U9961 (N_9961,N_4998,N_1064);
nor U9962 (N_9962,N_4743,N_1458);
or U9963 (N_9963,N_3611,N_3007);
nand U9964 (N_9964,N_3852,N_3865);
nor U9965 (N_9965,N_3331,N_4829);
nand U9966 (N_9966,N_3193,N_513);
or U9967 (N_9967,N_2459,N_2507);
nand U9968 (N_9968,N_1779,N_4285);
nand U9969 (N_9969,N_2033,N_2856);
nor U9970 (N_9970,N_806,N_1963);
nand U9971 (N_9971,N_2567,N_3230);
nand U9972 (N_9972,N_3794,N_1622);
and U9973 (N_9973,N_4108,N_406);
and U9974 (N_9974,N_4854,N_1867);
and U9975 (N_9975,N_1410,N_3667);
nand U9976 (N_9976,N_1760,N_2740);
nand U9977 (N_9977,N_262,N_629);
nand U9978 (N_9978,N_1614,N_3490);
nand U9979 (N_9979,N_3190,N_2216);
xnor U9980 (N_9980,N_1992,N_2227);
nor U9981 (N_9981,N_3312,N_4990);
nand U9982 (N_9982,N_3408,N_504);
and U9983 (N_9983,N_655,N_951);
nand U9984 (N_9984,N_677,N_3814);
or U9985 (N_9985,N_2819,N_4408);
xnor U9986 (N_9986,N_4204,N_280);
and U9987 (N_9987,N_72,N_1797);
or U9988 (N_9988,N_74,N_799);
or U9989 (N_9989,N_2190,N_3812);
nor U9990 (N_9990,N_2965,N_1932);
or U9991 (N_9991,N_2826,N_862);
nor U9992 (N_9992,N_4607,N_4989);
nand U9993 (N_9993,N_862,N_1);
xor U9994 (N_9994,N_2264,N_3374);
nor U9995 (N_9995,N_1207,N_4865);
and U9996 (N_9996,N_2392,N_2656);
and U9997 (N_9997,N_1819,N_3090);
and U9998 (N_9998,N_737,N_2202);
nand U9999 (N_9999,N_1708,N_3751);
and UO_0 (O_0,N_8064,N_5279);
nor UO_1 (O_1,N_7738,N_7555);
xor UO_2 (O_2,N_6779,N_7352);
or UO_3 (O_3,N_6544,N_7953);
nor UO_4 (O_4,N_7875,N_5328);
nor UO_5 (O_5,N_7501,N_5566);
or UO_6 (O_6,N_8758,N_8749);
and UO_7 (O_7,N_8461,N_9187);
xnor UO_8 (O_8,N_9748,N_8504);
nand UO_9 (O_9,N_7526,N_6034);
nand UO_10 (O_10,N_6459,N_7083);
nand UO_11 (O_11,N_9809,N_6369);
or UO_12 (O_12,N_6193,N_7243);
nor UO_13 (O_13,N_8212,N_5579);
nor UO_14 (O_14,N_5795,N_5019);
or UO_15 (O_15,N_6377,N_9061);
nand UO_16 (O_16,N_5268,N_6026);
nor UO_17 (O_17,N_7760,N_9698);
nor UO_18 (O_18,N_5006,N_5562);
nor UO_19 (O_19,N_6027,N_5174);
nand UO_20 (O_20,N_7613,N_9463);
or UO_21 (O_21,N_5168,N_5335);
nor UO_22 (O_22,N_9108,N_8495);
nand UO_23 (O_23,N_8382,N_9749);
nand UO_24 (O_24,N_9130,N_5413);
or UO_25 (O_25,N_8457,N_6775);
or UO_26 (O_26,N_7683,N_8462);
nor UO_27 (O_27,N_7670,N_6317);
and UO_28 (O_28,N_6581,N_9740);
xor UO_29 (O_29,N_8409,N_7795);
nand UO_30 (O_30,N_8349,N_9140);
or UO_31 (O_31,N_8678,N_8522);
nor UO_32 (O_32,N_6441,N_9111);
or UO_33 (O_33,N_5702,N_5836);
nor UO_34 (O_34,N_9145,N_7354);
nor UO_35 (O_35,N_6298,N_6816);
or UO_36 (O_36,N_5839,N_8975);
and UO_37 (O_37,N_8022,N_6992);
nor UO_38 (O_38,N_8342,N_5851);
xnor UO_39 (O_39,N_9332,N_5911);
or UO_40 (O_40,N_7332,N_6944);
xor UO_41 (O_41,N_5528,N_7467);
or UO_42 (O_42,N_7866,N_6186);
nand UO_43 (O_43,N_9116,N_9169);
and UO_44 (O_44,N_8660,N_9669);
and UO_45 (O_45,N_9562,N_8588);
and UO_46 (O_46,N_8093,N_6991);
nor UO_47 (O_47,N_6077,N_5510);
nand UO_48 (O_48,N_9765,N_6085);
nand UO_49 (O_49,N_7029,N_7198);
nand UO_50 (O_50,N_8658,N_5339);
or UO_51 (O_51,N_9153,N_7168);
and UO_52 (O_52,N_5825,N_9189);
or UO_53 (O_53,N_5657,N_5861);
or UO_54 (O_54,N_9812,N_6577);
nand UO_55 (O_55,N_5197,N_9119);
xnor UO_56 (O_56,N_6154,N_7230);
nand UO_57 (O_57,N_9227,N_7099);
nand UO_58 (O_58,N_7408,N_5398);
or UO_59 (O_59,N_7711,N_7596);
nor UO_60 (O_60,N_9975,N_5214);
nand UO_61 (O_61,N_8401,N_6115);
nor UO_62 (O_62,N_9553,N_6379);
nand UO_63 (O_63,N_6660,N_7782);
nand UO_64 (O_64,N_9157,N_8331);
and UO_65 (O_65,N_6840,N_7398);
nor UO_66 (O_66,N_7406,N_7510);
or UO_67 (O_67,N_8154,N_7308);
nand UO_68 (O_68,N_5062,N_6198);
nor UO_69 (O_69,N_7434,N_6288);
and UO_70 (O_70,N_9896,N_5625);
or UO_71 (O_71,N_7878,N_9602);
and UO_72 (O_72,N_9185,N_8899);
nor UO_73 (O_73,N_6489,N_9272);
xnor UO_74 (O_74,N_5988,N_9107);
and UO_75 (O_75,N_6396,N_5204);
and UO_76 (O_76,N_9416,N_5491);
nand UO_77 (O_77,N_7787,N_5112);
or UO_78 (O_78,N_6265,N_5014);
and UO_79 (O_79,N_8556,N_6630);
and UO_80 (O_80,N_8627,N_8406);
or UO_81 (O_81,N_9077,N_9310);
or UO_82 (O_82,N_5842,N_8989);
nand UO_83 (O_83,N_7342,N_6218);
xnor UO_84 (O_84,N_5266,N_9033);
nand UO_85 (O_85,N_5121,N_7070);
and UO_86 (O_86,N_7946,N_5611);
nor UO_87 (O_87,N_9243,N_9003);
nor UO_88 (O_88,N_8779,N_9105);
and UO_89 (O_89,N_6296,N_8566);
xor UO_90 (O_90,N_5955,N_8884);
or UO_91 (O_91,N_7799,N_7572);
nand UO_92 (O_92,N_9404,N_8450);
nor UO_93 (O_93,N_5650,N_9832);
nor UO_94 (O_94,N_8568,N_8106);
nor UO_95 (O_95,N_9911,N_8309);
xnor UO_96 (O_96,N_6168,N_7331);
nor UO_97 (O_97,N_5455,N_8062);
nand UO_98 (O_98,N_6167,N_8105);
nand UO_99 (O_99,N_7836,N_7412);
nand UO_100 (O_100,N_6197,N_9659);
or UO_101 (O_101,N_6746,N_8468);
and UO_102 (O_102,N_7216,N_5743);
and UO_103 (O_103,N_9358,N_9924);
nor UO_104 (O_104,N_9475,N_8574);
nor UO_105 (O_105,N_5598,N_7197);
or UO_106 (O_106,N_9805,N_6422);
nor UO_107 (O_107,N_7717,N_9307);
nand UO_108 (O_108,N_6654,N_5231);
and UO_109 (O_109,N_7374,N_5042);
nor UO_110 (O_110,N_7266,N_7397);
and UO_111 (O_111,N_7653,N_9472);
nor UO_112 (O_112,N_8535,N_6004);
nor UO_113 (O_113,N_9953,N_5762);
xor UO_114 (O_114,N_7169,N_8870);
nand UO_115 (O_115,N_8742,N_5622);
nand UO_116 (O_116,N_9417,N_5325);
nand UO_117 (O_117,N_9010,N_6281);
and UO_118 (O_118,N_9387,N_5549);
nor UO_119 (O_119,N_6751,N_8737);
nand UO_120 (O_120,N_7806,N_7837);
nor UO_121 (O_121,N_7618,N_7036);
or UO_122 (O_122,N_7281,N_5661);
and UO_123 (O_123,N_7330,N_5544);
nor UO_124 (O_124,N_6339,N_5684);
nor UO_125 (O_125,N_6905,N_7270);
nor UO_126 (O_126,N_9082,N_5559);
or UO_127 (O_127,N_6821,N_9137);
xnor UO_128 (O_128,N_8005,N_7925);
nand UO_129 (O_129,N_5847,N_8030);
or UO_130 (O_130,N_5332,N_8199);
nand UO_131 (O_131,N_6545,N_7845);
or UO_132 (O_132,N_7887,N_9364);
nand UO_133 (O_133,N_5369,N_7239);
or UO_134 (O_134,N_8051,N_8042);
or UO_135 (O_135,N_6625,N_5664);
nand UO_136 (O_136,N_6081,N_7833);
nand UO_137 (O_137,N_9067,N_5930);
nor UO_138 (O_138,N_6615,N_9551);
or UO_139 (O_139,N_6829,N_8951);
or UO_140 (O_140,N_6929,N_9688);
and UO_141 (O_141,N_9980,N_5406);
and UO_142 (O_142,N_8286,N_5731);
nand UO_143 (O_143,N_9897,N_8897);
and UO_144 (O_144,N_8725,N_8127);
nand UO_145 (O_145,N_8455,N_9324);
and UO_146 (O_146,N_5086,N_9859);
nand UO_147 (O_147,N_5443,N_8232);
or UO_148 (O_148,N_6348,N_7646);
and UO_149 (O_149,N_8976,N_9423);
nand UO_150 (O_150,N_6790,N_6029);
or UO_151 (O_151,N_9302,N_5125);
and UO_152 (O_152,N_8819,N_5685);
nand UO_153 (O_153,N_9737,N_6608);
or UO_154 (O_154,N_6338,N_7346);
and UO_155 (O_155,N_9655,N_8335);
or UO_156 (O_156,N_6144,N_9907);
nor UO_157 (O_157,N_8711,N_7075);
nand UO_158 (O_158,N_5460,N_7989);
and UO_159 (O_159,N_6648,N_8084);
nand UO_160 (O_160,N_5931,N_9853);
nand UO_161 (O_161,N_8787,N_9965);
and UO_162 (O_162,N_6210,N_8430);
xor UO_163 (O_163,N_8463,N_5001);
or UO_164 (O_164,N_9758,N_9322);
nand UO_165 (O_165,N_7685,N_9340);
xnor UO_166 (O_166,N_8016,N_8380);
nand UO_167 (O_167,N_9004,N_7771);
nand UO_168 (O_168,N_6859,N_9595);
or UO_169 (O_169,N_5716,N_9470);
nor UO_170 (O_170,N_7707,N_8708);
nor UO_171 (O_171,N_8514,N_5752);
or UO_172 (O_172,N_6776,N_6242);
nor UO_173 (O_173,N_5555,N_6427);
and UO_174 (O_174,N_7570,N_5069);
nand UO_175 (O_175,N_6067,N_7933);
nor UO_176 (O_176,N_9906,N_9860);
or UO_177 (O_177,N_9142,N_6327);
xnor UO_178 (O_178,N_5954,N_9089);
nand UO_179 (O_179,N_6241,N_9667);
nand UO_180 (O_180,N_9776,N_6060);
nor UO_181 (O_181,N_6901,N_6870);
and UO_182 (O_182,N_9266,N_7494);
and UO_183 (O_183,N_5789,N_6656);
and UO_184 (O_184,N_5844,N_6563);
or UO_185 (O_185,N_8023,N_7460);
or UO_186 (O_186,N_9132,N_6058);
xor UO_187 (O_187,N_7114,N_6096);
and UO_188 (O_188,N_6925,N_7648);
and UO_189 (O_189,N_8702,N_8176);
nand UO_190 (O_190,N_6330,N_5302);
nand UO_191 (O_191,N_9982,N_6958);
nor UO_192 (O_192,N_5777,N_9007);
nor UO_193 (O_193,N_8783,N_7777);
nand UO_194 (O_194,N_6036,N_9276);
and UO_195 (O_195,N_8510,N_5553);
nor UO_196 (O_196,N_9828,N_6732);
or UO_197 (O_197,N_7165,N_8235);
and UO_198 (O_198,N_8276,N_9791);
nor UO_199 (O_199,N_7102,N_6409);
xnor UO_200 (O_200,N_5740,N_7359);
and UO_201 (O_201,N_9599,N_8958);
and UO_202 (O_202,N_5998,N_7662);
nand UO_203 (O_203,N_9676,N_6684);
and UO_204 (O_204,N_6028,N_5708);
or UO_205 (O_205,N_7812,N_8361);
or UO_206 (O_206,N_5849,N_7233);
and UO_207 (O_207,N_6150,N_9511);
or UO_208 (O_208,N_9124,N_8719);
nand UO_209 (O_209,N_9605,N_8037);
or UO_210 (O_210,N_6325,N_6996);
nand UO_211 (O_211,N_5415,N_5819);
or UO_212 (O_212,N_8004,N_6287);
and UO_213 (O_213,N_8720,N_5324);
and UO_214 (O_214,N_6472,N_6397);
nor UO_215 (O_215,N_7241,N_8765);
nand UO_216 (O_216,N_9448,N_9284);
nand UO_217 (O_217,N_5571,N_8133);
and UO_218 (O_218,N_7969,N_7750);
or UO_219 (O_219,N_7607,N_6579);
nand UO_220 (O_220,N_7615,N_8539);
nand UO_221 (O_221,N_6784,N_6827);
and UO_222 (O_222,N_8862,N_6432);
nor UO_223 (O_223,N_8563,N_6393);
or UO_224 (O_224,N_5918,N_5305);
or UO_225 (O_225,N_7027,N_7104);
xor UO_226 (O_226,N_9228,N_7227);
nor UO_227 (O_227,N_7868,N_5570);
and UO_228 (O_228,N_6069,N_7269);
nor UO_229 (O_229,N_7641,N_7926);
or UO_230 (O_230,N_8634,N_8540);
or UO_231 (O_231,N_8942,N_7992);
nor UO_232 (O_232,N_9192,N_7826);
or UO_233 (O_233,N_7502,N_6597);
or UO_234 (O_234,N_5452,N_6105);
nand UO_235 (O_235,N_6014,N_9995);
or UO_236 (O_236,N_8186,N_9051);
or UO_237 (O_237,N_5953,N_6117);
and UO_238 (O_238,N_8933,N_5993);
or UO_239 (O_239,N_9833,N_7417);
or UO_240 (O_240,N_6131,N_9764);
nor UO_241 (O_241,N_5935,N_8432);
or UO_242 (O_242,N_5144,N_5393);
nand UO_243 (O_243,N_9457,N_9296);
and UO_244 (O_244,N_5904,N_5936);
nand UO_245 (O_245,N_5768,N_5145);
nor UO_246 (O_246,N_5186,N_7049);
and UO_247 (O_247,N_8486,N_6051);
nor UO_248 (O_248,N_7538,N_9478);
nand UO_249 (O_249,N_5151,N_9537);
nand UO_250 (O_250,N_9646,N_9584);
nand UO_251 (O_251,N_6340,N_9580);
or UO_252 (O_252,N_9047,N_5627);
nor UO_253 (O_253,N_9733,N_8081);
and UO_254 (O_254,N_5782,N_9330);
nor UO_255 (O_255,N_9956,N_7333);
nor UO_256 (O_256,N_9435,N_7465);
or UO_257 (O_257,N_5900,N_6243);
nor UO_258 (O_258,N_7443,N_8520);
nand UO_259 (O_259,N_9120,N_8441);
nor UO_260 (O_260,N_7729,N_7073);
nand UO_261 (O_261,N_6054,N_7949);
nand UO_262 (O_262,N_7864,N_9175);
xnor UO_263 (O_263,N_6798,N_8739);
and UO_264 (O_264,N_5426,N_6479);
nor UO_265 (O_265,N_7181,N_8466);
or UO_266 (O_266,N_6213,N_8519);
nor UO_267 (O_267,N_7171,N_6043);
nand UO_268 (O_268,N_7437,N_7031);
xor UO_269 (O_269,N_8372,N_5869);
nor UO_270 (O_270,N_5690,N_6753);
or UO_271 (O_271,N_9413,N_6251);
and UO_272 (O_272,N_5390,N_8148);
and UO_273 (O_273,N_7234,N_5588);
nor UO_274 (O_274,N_5568,N_8251);
and UO_275 (O_275,N_7715,N_9856);
nor UO_276 (O_276,N_8122,N_9984);
nor UO_277 (O_277,N_6858,N_7663);
nor UO_278 (O_278,N_5671,N_9571);
nor UO_279 (O_279,N_5009,N_8333);
nor UO_280 (O_280,N_8423,N_5881);
or UO_281 (O_281,N_7880,N_9960);
nor UO_282 (O_282,N_8200,N_6245);
nand UO_283 (O_283,N_8650,N_8659);
or UO_284 (O_284,N_7739,N_7353);
and UO_285 (O_285,N_5886,N_9623);
nor UO_286 (O_286,N_6224,N_8070);
and UO_287 (O_287,N_7874,N_6989);
or UO_288 (O_288,N_6598,N_6617);
and UO_289 (O_289,N_6765,N_8880);
and UO_290 (O_290,N_8866,N_9957);
nand UO_291 (O_291,N_7003,N_6853);
or UO_292 (O_292,N_6607,N_7038);
or UO_293 (O_293,N_6374,N_8831);
or UO_294 (O_294,N_7654,N_7283);
xor UO_295 (O_295,N_9362,N_6578);
nor UO_296 (O_296,N_7774,N_9734);
nor UO_297 (O_297,N_8275,N_6739);
and UO_298 (O_298,N_7082,N_5974);
or UO_299 (O_299,N_6721,N_9123);
and UO_300 (O_300,N_5928,N_9869);
nor UO_301 (O_301,N_5534,N_9703);
and UO_302 (O_302,N_6297,N_9931);
nor UO_303 (O_303,N_5055,N_6543);
xnor UO_304 (O_304,N_9723,N_5806);
and UO_305 (O_305,N_7162,N_9938);
or UO_306 (O_306,N_8549,N_6201);
nand UO_307 (O_307,N_7513,N_5068);
and UO_308 (O_308,N_5164,N_8433);
and UO_309 (O_309,N_7495,N_9480);
and UO_310 (O_310,N_6585,N_7123);
nand UO_311 (O_311,N_5076,N_7871);
and UO_312 (O_312,N_5888,N_7847);
and UO_313 (O_313,N_7840,N_5447);
nor UO_314 (O_314,N_5940,N_6553);
nor UO_315 (O_315,N_9557,N_9760);
or UO_316 (O_316,N_5876,N_9280);
nor UO_317 (O_317,N_6667,N_9221);
or UO_318 (O_318,N_7537,N_6611);
nand UO_319 (O_319,N_6041,N_9333);
and UO_320 (O_320,N_6644,N_8611);
and UO_321 (O_321,N_6047,N_8923);
and UO_322 (O_322,N_6104,N_9411);
or UO_323 (O_323,N_7455,N_9675);
and UO_324 (O_324,N_9178,N_6985);
xnor UO_325 (O_325,N_8895,N_5310);
nor UO_326 (O_326,N_9244,N_8826);
and UO_327 (O_327,N_8931,N_5999);
or UO_328 (O_328,N_9492,N_7034);
or UO_329 (O_329,N_9513,N_8507);
nand UO_330 (O_330,N_9230,N_8655);
nor UO_331 (O_331,N_8652,N_6110);
nor UO_332 (O_332,N_9545,N_5858);
and UO_333 (O_333,N_6233,N_7207);
and UO_334 (O_334,N_5431,N_6621);
nand UO_335 (O_335,N_5937,N_8784);
nand UO_336 (O_336,N_6939,N_5547);
or UO_337 (O_337,N_5113,N_8515);
nor UO_338 (O_338,N_7789,N_7578);
nor UO_339 (O_339,N_5053,N_5527);
nand UO_340 (O_340,N_7192,N_6876);
nand UO_341 (O_341,N_9055,N_9813);
nand UO_342 (O_342,N_5691,N_7704);
or UO_343 (O_343,N_7334,N_7053);
nand UO_344 (O_344,N_7372,N_8334);
and UO_345 (O_345,N_8934,N_5639);
and UO_346 (O_346,N_8035,N_5137);
and UO_347 (O_347,N_9843,N_6045);
or UO_348 (O_348,N_9894,N_5599);
nor UO_349 (O_349,N_7280,N_8282);
nor UO_350 (O_350,N_5833,N_6783);
nand UO_351 (O_351,N_9918,N_6189);
nor UO_352 (O_352,N_9912,N_7008);
nor UO_353 (O_353,N_5264,N_9876);
nor UO_354 (O_354,N_5737,N_6674);
or UO_355 (O_355,N_7295,N_8196);
or UO_356 (O_356,N_6370,N_8304);
xnor UO_357 (O_357,N_9084,N_5383);
and UO_358 (O_358,N_8647,N_5356);
nor UO_359 (O_359,N_8644,N_7788);
nor UO_360 (O_360,N_7050,N_5025);
or UO_361 (O_361,N_6515,N_8633);
or UO_362 (O_362,N_9796,N_9775);
nor UO_363 (O_363,N_7575,N_8339);
and UO_364 (O_364,N_9292,N_9136);
or UO_365 (O_365,N_5285,N_9969);
xor UO_366 (O_366,N_6909,N_6863);
and UO_367 (O_367,N_6881,N_6208);
or UO_368 (O_368,N_7426,N_8236);
or UO_369 (O_369,N_9146,N_8575);
xnor UO_370 (O_370,N_9769,N_8590);
or UO_371 (O_371,N_8190,N_9155);
or UO_372 (O_372,N_8981,N_5963);
or UO_373 (O_373,N_5171,N_9589);
or UO_374 (O_374,N_5983,N_7156);
and UO_375 (O_375,N_7160,N_7065);
or UO_376 (O_376,N_7818,N_6070);
nand UO_377 (O_377,N_9134,N_9708);
nand UO_378 (O_378,N_9388,N_7107);
or UO_379 (O_379,N_6470,N_8370);
xnor UO_380 (O_380,N_7453,N_6789);
xor UO_381 (O_381,N_5400,N_7931);
or UO_382 (O_382,N_5992,N_8124);
nand UO_383 (O_383,N_9664,N_6316);
or UO_384 (O_384,N_9793,N_8775);
nor UO_385 (O_385,N_5978,N_9757);
nand UO_386 (O_386,N_7628,N_8695);
and UO_387 (O_387,N_8400,N_5256);
nor UO_388 (O_388,N_8859,N_6907);
or UO_389 (O_389,N_5536,N_9886);
and UO_390 (O_390,N_6938,N_7834);
and UO_391 (O_391,N_8919,N_6583);
nand UO_392 (O_392,N_9210,N_9471);
nand UO_393 (O_393,N_9059,N_6093);
or UO_394 (O_394,N_7547,N_5593);
and UO_395 (O_395,N_5065,N_7690);
or UO_396 (O_396,N_6999,N_6584);
nand UO_397 (O_397,N_9823,N_9390);
nand UO_398 (O_398,N_9196,N_9645);
xor UO_399 (O_399,N_8690,N_7480);
nor UO_400 (O_400,N_8926,N_6864);
nand UO_401 (O_401,N_6392,N_9485);
and UO_402 (O_402,N_9792,N_7487);
nor UO_403 (O_403,N_5933,N_5263);
or UO_404 (O_404,N_8523,N_9046);
nor UO_405 (O_405,N_5700,N_8714);
or UO_406 (O_406,N_9075,N_6586);
nand UO_407 (O_407,N_5091,N_9798);
or UO_408 (O_408,N_5697,N_6671);
or UO_409 (O_409,N_6285,N_8344);
and UO_410 (O_410,N_8213,N_5997);
xor UO_411 (O_411,N_7569,N_7457);
nor UO_412 (O_412,N_6449,N_7399);
or UO_413 (O_413,N_9406,N_5453);
xnor UO_414 (O_414,N_9392,N_8354);
nand UO_415 (O_415,N_8375,N_6118);
nand UO_416 (O_416,N_8233,N_6155);
or UO_417 (O_417,N_5665,N_8343);
and UO_418 (O_418,N_6098,N_9163);
and UO_419 (O_419,N_5399,N_7966);
and UO_420 (O_420,N_7898,N_7155);
nand UO_421 (O_421,N_6044,N_6526);
nand UO_422 (O_422,N_9453,N_7365);
nor UO_423 (O_423,N_7862,N_8823);
nor UO_424 (O_424,N_5360,N_6371);
or UO_425 (O_425,N_6426,N_9369);
and UO_426 (O_426,N_7877,N_9403);
or UO_427 (O_427,N_6972,N_9999);
nand UO_428 (O_428,N_8833,N_6643);
nor UO_429 (O_429,N_6177,N_7375);
xnor UO_430 (O_430,N_7580,N_7043);
and UO_431 (O_431,N_6078,N_9662);
and UO_432 (O_432,N_7164,N_9516);
nand UO_433 (O_433,N_5118,N_5628);
nand UO_434 (O_434,N_6493,N_5222);
or UO_435 (O_435,N_7635,N_8078);
or UO_436 (O_436,N_6813,N_5321);
nor UO_437 (O_437,N_6935,N_7606);
xnor UO_438 (O_438,N_9978,N_9032);
nor UO_439 (O_439,N_6178,N_8688);
and UO_440 (O_440,N_5459,N_5182);
and UO_441 (O_441,N_5388,N_9313);
and UO_442 (O_442,N_5159,N_8912);
or UO_443 (O_443,N_6452,N_9396);
and UO_444 (O_444,N_9690,N_8241);
nand UO_445 (O_445,N_6384,N_7028);
nand UO_446 (O_446,N_8219,N_5709);
xor UO_447 (O_447,N_6540,N_7976);
or UO_448 (O_448,N_6689,N_8597);
nand UO_449 (O_449,N_6582,N_9519);
xnor UO_450 (O_450,N_5387,N_8205);
nand UO_451 (O_451,N_9541,N_8825);
and UO_452 (O_452,N_6204,N_7219);
or UO_453 (O_453,N_5191,N_9290);
or UO_454 (O_454,N_8843,N_6712);
xor UO_455 (O_455,N_9722,N_6156);
nand UO_456 (O_456,N_8705,N_8589);
nor UO_457 (O_457,N_8263,N_9534);
nand UO_458 (O_458,N_6742,N_6668);
nor UO_459 (O_459,N_5891,N_9744);
and UO_460 (O_460,N_7135,N_5155);
and UO_461 (O_461,N_6716,N_5524);
and UO_462 (O_462,N_5132,N_9766);
nand UO_463 (O_463,N_8284,N_8807);
nand UO_464 (O_464,N_5587,N_9222);
or UO_465 (O_465,N_6273,N_5011);
nor UO_466 (O_466,N_6166,N_8987);
or UO_467 (O_467,N_6533,N_9042);
nor UO_468 (O_468,N_8502,N_9920);
xor UO_469 (O_469,N_9129,N_5093);
or UO_470 (O_470,N_6904,N_8669);
and UO_471 (O_471,N_6566,N_9908);
nand UO_472 (O_472,N_8099,N_9745);
nor UO_473 (O_473,N_7500,N_9342);
nor UO_474 (O_474,N_7475,N_9438);
or UO_475 (O_475,N_7968,N_8904);
nand UO_476 (O_476,N_8228,N_7865);
xor UO_477 (O_477,N_7894,N_5812);
nor UO_478 (O_478,N_9432,N_7336);
nand UO_479 (O_479,N_9346,N_6395);
or UO_480 (O_480,N_8104,N_5021);
nor UO_481 (O_481,N_6814,N_7870);
nor UO_482 (O_482,N_8140,N_9048);
nor UO_483 (O_483,N_6521,N_7228);
nand UO_484 (O_484,N_7705,N_7424);
nand UO_485 (O_485,N_5142,N_5530);
nand UO_486 (O_486,N_7791,N_8065);
nor UO_487 (O_487,N_9905,N_9425);
nor UO_488 (O_488,N_6824,N_5234);
or UO_489 (O_489,N_5496,N_8731);
or UO_490 (O_490,N_9782,N_9184);
and UO_491 (O_491,N_8876,N_6314);
xor UO_492 (O_492,N_8855,N_5834);
or UO_493 (O_493,N_8670,N_7328);
nand UO_494 (O_494,N_9014,N_5689);
nand UO_495 (O_495,N_5377,N_5470);
or UO_496 (O_496,N_8234,N_6079);
xor UO_497 (O_497,N_8570,N_7483);
nor UO_498 (O_498,N_8917,N_6300);
nor UO_499 (O_499,N_9408,N_8143);
nand UO_500 (O_500,N_6183,N_8996);
nor UO_501 (O_501,N_7252,N_5206);
nor UO_502 (O_502,N_5783,N_9997);
xnor UO_503 (O_503,N_5167,N_7535);
or UO_504 (O_504,N_7622,N_6013);
xor UO_505 (O_505,N_5706,N_5403);
xnor UO_506 (O_506,N_9610,N_7505);
or UO_507 (O_507,N_9182,N_6012);
and UO_508 (O_508,N_7360,N_6887);
nor UO_509 (O_509,N_7303,N_7153);
and UO_510 (O_510,N_9455,N_6261);
nand UO_511 (O_511,N_5735,N_5898);
nand UO_512 (O_512,N_8404,N_6031);
and UO_513 (O_513,N_9087,N_7282);
xnor UO_514 (O_514,N_5970,N_8155);
nor UO_515 (O_515,N_8617,N_8785);
nand UO_516 (O_516,N_9616,N_7433);
and UO_517 (O_517,N_7901,N_7665);
nor UO_518 (O_518,N_8312,N_9533);
or UO_519 (O_519,N_8326,N_8320);
nor UO_520 (O_520,N_8193,N_7756);
nand UO_521 (O_521,N_7285,N_6548);
nand UO_522 (O_522,N_9607,N_5910);
nor UO_523 (O_523,N_9458,N_6017);
xor UO_524 (O_524,N_9400,N_8314);
or UO_525 (O_525,N_5624,N_8204);
or UO_526 (O_526,N_6590,N_8603);
and UO_527 (O_527,N_5721,N_9606);
and UO_528 (O_528,N_6246,N_6456);
and UO_529 (O_529,N_7316,N_7598);
nand UO_530 (O_530,N_8900,N_6124);
or UO_531 (O_531,N_5666,N_5601);
and UO_532 (O_532,N_6429,N_5785);
and UO_533 (O_533,N_6690,N_5581);
and UO_534 (O_534,N_5194,N_8487);
nor UO_535 (O_535,N_8672,N_6698);
nor UO_536 (O_536,N_6128,N_7311);
nand UO_537 (O_537,N_6455,N_7805);
nor UO_538 (O_538,N_9762,N_7389);
and UO_539 (O_539,N_8422,N_6196);
and UO_540 (O_540,N_5394,N_9476);
nor UO_541 (O_541,N_8733,N_6699);
and UO_542 (O_542,N_7203,N_6556);
nand UO_543 (O_543,N_5728,N_7511);
or UO_544 (O_544,N_9728,N_9429);
or UO_545 (O_545,N_7416,N_9420);
and UO_546 (O_546,N_6046,N_6519);
or UO_547 (O_547,N_5516,N_5809);
or UO_548 (O_548,N_6922,N_6157);
nor UO_549 (O_549,N_6943,N_6795);
nand UO_550 (O_550,N_8560,N_7603);
nor UO_551 (O_551,N_9025,N_8518);
nand UO_552 (O_552,N_5660,N_9657);
nand UO_553 (O_553,N_9540,N_9229);
and UO_554 (O_554,N_8755,N_6373);
and UO_555 (O_555,N_7721,N_8129);
and UO_556 (O_556,N_9531,N_9495);
nand UO_557 (O_557,N_8082,N_6679);
and UO_558 (O_558,N_8152,N_6305);
xnor UO_559 (O_559,N_7206,N_9579);
or UO_560 (O_560,N_6320,N_5565);
xor UO_561 (O_561,N_7888,N_9523);
and UO_562 (O_562,N_7235,N_7960);
xnor UO_563 (O_563,N_7136,N_6534);
nand UO_564 (O_564,N_8451,N_5218);
and UO_565 (O_565,N_6346,N_5163);
and UO_566 (O_566,N_9011,N_8411);
nand UO_567 (O_567,N_7462,N_5675);
nand UO_568 (O_568,N_6931,N_9992);
nor UO_569 (O_569,N_8153,N_8316);
nand UO_570 (O_570,N_5987,N_5725);
xnor UO_571 (O_571,N_7425,N_9477);
nand UO_572 (O_572,N_6412,N_8681);
nor UO_573 (O_573,N_9903,N_8489);
nand UO_574 (O_574,N_5617,N_5345);
nor UO_575 (O_575,N_9875,N_5027);
nor UO_576 (O_576,N_9591,N_5572);
nand UO_577 (O_577,N_5347,N_9600);
and UO_578 (O_578,N_5673,N_9979);
xor UO_579 (O_579,N_8761,N_7436);
and UO_580 (O_580,N_7922,N_5450);
nor UO_581 (O_581,N_6978,N_9955);
and UO_582 (O_582,N_9743,N_7097);
nor UO_583 (O_583,N_7928,N_9684);
nor UO_584 (O_584,N_8446,N_5800);
nor UO_585 (O_585,N_5154,N_8764);
or UO_586 (O_586,N_5012,N_9974);
or UO_587 (O_587,N_5723,N_8759);
xnor UO_588 (O_588,N_7215,N_7669);
or UO_589 (O_589,N_6133,N_5781);
and UO_590 (O_590,N_9451,N_5212);
xnor UO_591 (O_591,N_6289,N_6596);
or UO_592 (O_592,N_9661,N_8762);
and UO_593 (O_593,N_9829,N_5084);
or UO_594 (O_594,N_9288,N_5313);
nand UO_595 (O_595,N_5958,N_8621);
and UO_596 (O_596,N_5733,N_9687);
nor UO_597 (O_597,N_5648,N_6830);
and UO_598 (O_598,N_8861,N_7813);
xnor UO_599 (O_599,N_7773,N_9939);
nor UO_600 (O_600,N_6365,N_9535);
and UO_601 (O_601,N_5209,N_6506);
nand UO_602 (O_602,N_9452,N_5149);
and UO_603 (O_603,N_6469,N_5126);
or UO_604 (O_604,N_5859,N_7488);
and UO_605 (O_605,N_5951,N_6971);
or UO_606 (O_606,N_6362,N_9091);
and UO_607 (O_607,N_5715,N_6796);
or UO_608 (O_608,N_5780,N_7786);
nor UO_609 (O_609,N_9524,N_9826);
and UO_610 (O_610,N_5701,N_9312);
xor UO_611 (O_611,N_7879,N_6328);
xnor UO_612 (O_612,N_6127,N_9842);
or UO_613 (O_613,N_8206,N_8239);
nor UO_614 (O_614,N_9267,N_7379);
xnor UO_615 (O_615,N_8494,N_7523);
xnor UO_616 (O_616,N_6755,N_7428);
nor UO_617 (O_617,N_6394,N_5329);
and UO_618 (O_618,N_6520,N_9658);
or UO_619 (O_619,N_6200,N_5778);
nor UO_620 (O_620,N_6477,N_9808);
nand UO_621 (O_621,N_6355,N_7349);
and UO_622 (O_622,N_6532,N_8249);
and UO_623 (O_623,N_8045,N_7548);
nor UO_624 (O_624,N_8738,N_9318);
nand UO_625 (O_625,N_5606,N_7832);
and UO_626 (O_626,N_7421,N_8091);
xor UO_627 (O_627,N_9943,N_9525);
nor UO_628 (O_628,N_5794,N_9294);
nand UO_629 (O_629,N_5397,N_6979);
or UO_630 (O_630,N_6257,N_9604);
nor UO_631 (O_631,N_7040,N_7867);
and UO_632 (O_632,N_6194,N_8116);
nand UO_633 (O_633,N_6324,N_8173);
xor UO_634 (O_634,N_6729,N_8192);
and UO_635 (O_635,N_8521,N_8110);
or UO_636 (O_636,N_7461,N_5283);
xnor UO_637 (O_637,N_9854,N_8417);
nand UO_638 (O_638,N_7212,N_7745);
and UO_639 (O_639,N_7558,N_7815);
xor UO_640 (O_640,N_5023,N_5801);
nand UO_641 (O_641,N_7620,N_6462);
nor UO_642 (O_642,N_5105,N_6003);
nor UO_643 (O_643,N_7148,N_9321);
nand UO_644 (O_644,N_7369,N_5575);
and UO_645 (O_645,N_6653,N_9668);
and UO_646 (O_646,N_7753,N_8366);
xor UO_647 (O_647,N_9015,N_8307);
and UO_648 (O_648,N_8420,N_8226);
or UO_649 (O_649,N_8419,N_9674);
nand UO_650 (O_650,N_6190,N_7147);
nand UO_651 (O_651,N_5022,N_7941);
or UO_652 (O_652,N_9301,N_6501);
nand UO_653 (O_653,N_7629,N_9643);
nand UO_654 (O_654,N_6757,N_8967);
or UO_655 (O_655,N_7770,N_5585);
nor UO_656 (O_656,N_8703,N_6220);
or UO_657 (O_657,N_8001,N_5043);
or UO_658 (O_658,N_6042,N_9804);
nor UO_659 (O_659,N_5591,N_6360);
and UO_660 (O_660,N_6588,N_8524);
xor UO_661 (O_661,N_5533,N_9215);
nor UO_662 (O_662,N_7058,N_9884);
or UO_663 (O_663,N_5966,N_8724);
nand UO_664 (O_664,N_6147,N_9277);
or UO_665 (O_665,N_9634,N_5323);
and UO_666 (O_666,N_8614,N_5338);
nand UO_667 (O_667,N_7950,N_6293);
nand UO_668 (O_668,N_7260,N_9577);
or UO_669 (O_669,N_6319,N_7130);
and UO_670 (O_670,N_7706,N_5309);
or UO_671 (O_671,N_6927,N_9270);
nor UO_672 (O_672,N_6567,N_6682);
and UO_673 (O_673,N_7191,N_5583);
xnor UO_674 (O_674,N_8428,N_5767);
and UO_675 (O_675,N_8049,N_9509);
xor UO_676 (O_676,N_8555,N_9325);
nand UO_677 (O_677,N_7087,N_6209);
nand UO_678 (O_678,N_6308,N_9747);
and UO_679 (O_679,N_9981,N_8797);
nand UO_680 (O_680,N_8794,N_8592);
nor UO_681 (O_681,N_6626,N_7021);
nand UO_682 (O_682,N_5196,N_9977);
or UO_683 (O_683,N_6344,N_8608);
or UO_684 (O_684,N_6263,N_7621);
and UO_685 (O_685,N_9214,N_7935);
nor UO_686 (O_686,N_9665,N_8340);
nand UO_687 (O_687,N_9154,N_7441);
and UO_688 (O_688,N_7205,N_8272);
and UO_689 (O_689,N_6800,N_7490);
xnor UO_690 (O_690,N_8243,N_7000);
nor UO_691 (O_691,N_6768,N_9268);
nor UO_692 (O_692,N_8854,N_7497);
nor UO_693 (O_693,N_6276,N_8265);
nand UO_694 (O_694,N_8580,N_5414);
or UO_695 (O_695,N_7988,N_5586);
xnor UO_696 (O_696,N_5255,N_6471);
or UO_697 (O_697,N_5960,N_7009);
nand UO_698 (O_698,N_8437,N_7910);
and UO_699 (O_699,N_7154,N_6860);
nor UO_700 (O_700,N_9637,N_6068);
or UO_701 (O_701,N_5448,N_6451);
nand UO_702 (O_702,N_7098,N_5771);
and UO_703 (O_703,N_6253,N_7719);
and UO_704 (O_704,N_5607,N_7368);
or UO_705 (O_705,N_9078,N_8216);
nand UO_706 (O_706,N_9239,N_7936);
xor UO_707 (O_707,N_9113,N_8632);
nor UO_708 (O_708,N_9468,N_8939);
and UO_709 (O_709,N_9681,N_7672);
or UO_710 (O_710,N_9857,N_8217);
nor UO_711 (O_711,N_8087,N_5745);
nand UO_712 (O_712,N_6683,N_6696);
nor UO_713 (O_713,N_8682,N_7447);
nor UO_714 (O_714,N_9323,N_7108);
nor UO_715 (O_715,N_9150,N_7121);
or UO_716 (O_716,N_7395,N_8172);
and UO_717 (O_717,N_6000,N_6899);
nor UO_718 (O_718,N_6160,N_5658);
nor UO_719 (O_719,N_6882,N_7987);
nor UO_720 (O_720,N_8541,N_5694);
nand UO_721 (O_721,N_7747,N_7673);
or UO_722 (O_722,N_9935,N_9001);
nor UO_723 (O_723,N_9019,N_6635);
nor UO_724 (O_724,N_7999,N_9874);
or UO_725 (O_725,N_6740,N_8503);
nand UO_726 (O_726,N_8665,N_6366);
and UO_727 (O_727,N_6833,N_8492);
nor UO_728 (O_728,N_9149,N_7007);
nor UO_729 (O_729,N_8548,N_8068);
or UO_730 (O_730,N_8285,N_9993);
and UO_731 (O_731,N_9785,N_6812);
and UO_732 (O_732,N_5463,N_9633);
nand UO_733 (O_733,N_6052,N_5950);
or UO_734 (O_734,N_8530,N_5823);
nor UO_735 (O_735,N_6890,N_5890);
or UO_736 (O_736,N_5726,N_9326);
and UO_737 (O_737,N_9121,N_9058);
nor UO_738 (O_738,N_8849,N_8469);
nand UO_739 (O_739,N_8318,N_9216);
xor UO_740 (O_740,N_5776,N_7117);
or UO_741 (O_741,N_6071,N_9917);
or UO_742 (O_742,N_6806,N_6398);
nand UO_743 (O_743,N_7856,N_7701);
nand UO_744 (O_744,N_7326,N_9506);
or UO_745 (O_745,N_7384,N_5501);
xnor UO_746 (O_746,N_6769,N_8768);
nor UO_747 (O_747,N_6122,N_9660);
nor UO_748 (O_748,N_6587,N_9647);
nor UO_749 (O_749,N_6512,N_9536);
nand UO_750 (O_750,N_5129,N_5763);
or UO_751 (O_751,N_5975,N_6793);
nand UO_752 (O_752,N_7722,N_8863);
or UO_753 (O_753,N_7792,N_9338);
and UO_754 (O_754,N_9922,N_7810);
or UO_755 (O_755,N_5130,N_7780);
nand UO_756 (O_756,N_8896,N_5766);
nand UO_757 (O_757,N_6088,N_9348);
and UO_758 (O_758,N_5317,N_8648);
nand UO_759 (O_759,N_7236,N_8500);
nor UO_760 (O_760,N_8144,N_7751);
and UO_761 (O_761,N_5727,N_7515);
nand UO_762 (O_762,N_5169,N_9497);
nand UO_763 (O_763,N_7390,N_9653);
nand UO_764 (O_764,N_7273,N_5122);
and UO_765 (O_765,N_8874,N_7419);
and UO_766 (O_766,N_7324,N_5220);
nand UO_767 (O_767,N_7307,N_5210);
or UO_768 (O_768,N_8587,N_8135);
and UO_769 (O_769,N_6715,N_5078);
nor UO_770 (O_770,N_6763,N_9278);
nand UO_771 (O_771,N_7403,N_8214);
nor UO_772 (O_772,N_7649,N_9836);
or UO_773 (O_773,N_7014,N_9799);
or UO_774 (O_774,N_5106,N_7261);
nor UO_775 (O_775,N_6097,N_7591);
nor UO_776 (O_776,N_7896,N_5832);
nand UO_777 (O_777,N_7470,N_8857);
or UO_778 (O_778,N_5311,N_8999);
or UO_779 (O_779,N_8125,N_9095);
xnor UO_780 (O_780,N_5535,N_6815);
nand UO_781 (O_781,N_9753,N_5686);
nor UO_782 (O_782,N_9552,N_7918);
nand UO_783 (O_783,N_9772,N_5538);
or UO_784 (O_784,N_9152,N_9919);
and UO_785 (O_785,N_7740,N_5295);
and UO_786 (O_786,N_9286,N_7594);
nor UO_787 (O_787,N_6282,N_6454);
nand UO_788 (O_788,N_9592,N_8606);
nor UO_789 (O_789,N_5747,N_9283);
nor UO_790 (O_790,N_6400,N_5427);
xnor UO_791 (O_791,N_9756,N_5848);
and UO_792 (O_792,N_6730,N_7716);
nand UO_793 (O_793,N_8387,N_9036);
or UO_794 (O_794,N_9071,N_9720);
and UO_795 (O_795,N_8145,N_5649);
or UO_796 (O_796,N_7843,N_6733);
nor UO_797 (O_797,N_5730,N_6254);
nor UO_798 (O_798,N_6143,N_8405);
or UO_799 (O_799,N_9648,N_7011);
nor UO_800 (O_800,N_5814,N_6403);
nand UO_801 (O_801,N_6059,N_6856);
nand UO_802 (O_802,N_6351,N_5957);
or UO_803 (O_803,N_9689,N_8248);
xor UO_804 (O_804,N_9309,N_9355);
nand UO_805 (O_805,N_7240,N_6311);
nor UO_806 (O_806,N_8815,N_7188);
nand UO_807 (O_807,N_6560,N_8726);
and UO_808 (O_808,N_6141,N_7149);
and UO_809 (O_809,N_6862,N_6505);
nand UO_810 (O_810,N_6606,N_7185);
xnor UO_811 (O_811,N_6787,N_7585);
xor UO_812 (O_812,N_9073,N_7784);
nor UO_813 (O_813,N_7068,N_6274);
nor UO_814 (O_814,N_7956,N_6321);
nand UO_815 (O_815,N_5034,N_7650);
or UO_816 (O_816,N_8024,N_8992);
and UO_817 (O_817,N_9012,N_7329);
and UO_818 (O_818,N_7568,N_9702);
or UO_819 (O_819,N_6458,N_9778);
and UO_820 (O_820,N_7695,N_5267);
nor UO_821 (O_821,N_6024,N_7838);
nand UO_822 (O_822,N_7446,N_8572);
xnor UO_823 (O_823,N_7137,N_5097);
and UO_824 (O_824,N_6116,N_6884);
nand UO_825 (O_825,N_5016,N_8848);
and UO_826 (O_826,N_8772,N_9693);
nor UO_827 (O_827,N_5850,N_9361);
nor UO_828 (O_828,N_8610,N_8834);
nor UO_829 (O_829,N_9391,N_6847);
nand UO_830 (O_830,N_7211,N_7195);
nand UO_831 (O_831,N_6411,N_8924);
xnor UO_832 (O_832,N_7981,N_7339);
xnor UO_833 (O_833,N_8668,N_9821);
or UO_834 (O_834,N_9251,N_7427);
and UO_835 (O_835,N_7358,N_9009);
xnor UO_836 (O_836,N_5198,N_6857);
or UO_837 (O_837,N_5124,N_8625);
and UO_838 (O_838,N_8769,N_7942);
xor UO_839 (O_839,N_5557,N_7226);
or UO_840 (O_840,N_7516,N_5343);
xor UO_841 (O_841,N_5687,N_7546);
and UO_842 (O_842,N_5410,N_9436);
and UO_843 (O_843,N_6217,N_7301);
and UO_844 (O_844,N_8657,N_7908);
nor UO_845 (O_845,N_9538,N_7376);
nand UO_846 (O_846,N_7017,N_9316);
or UO_847 (O_847,N_9002,N_6923);
xnor UO_848 (O_848,N_8802,N_8579);
and UO_849 (O_849,N_9751,N_6140);
nor UO_850 (O_850,N_5240,N_9017);
nor UO_851 (O_851,N_6777,N_9341);
or UO_852 (O_852,N_5364,N_8175);
and UO_853 (O_853,N_6386,N_8493);
xor UO_854 (O_854,N_9434,N_7553);
and UO_855 (O_855,N_8979,N_5089);
nor UO_856 (O_856,N_7903,N_7413);
and UO_857 (O_857,N_5504,N_7963);
xor UO_858 (O_858,N_6664,N_5749);
or UO_859 (O_859,N_9128,N_8806);
nor UO_860 (O_860,N_8346,N_9127);
nand UO_861 (O_861,N_5300,N_6271);
or UO_862 (O_862,N_9131,N_7974);
and UO_863 (O_863,N_8111,N_9881);
xnor UO_864 (O_864,N_7208,N_5797);
nand UO_865 (O_865,N_8687,N_6735);
and UO_866 (O_866,N_9848,N_9949);
nor UO_867 (O_867,N_8168,N_8264);
nand UO_868 (O_868,N_8128,N_9871);
nand UO_869 (O_869,N_8383,N_8932);
nor UO_870 (O_870,N_5556,N_7238);
nand UO_871 (O_871,N_7180,N_7420);
nor UO_872 (O_872,N_6175,N_9414);
nor UO_873 (O_873,N_5015,N_6278);
or UO_874 (O_874,N_7357,N_8698);
and UO_875 (O_875,N_9112,N_8258);
or UO_876 (O_876,N_5226,N_7166);
xnor UO_877 (O_877,N_8266,N_9697);
and UO_878 (O_878,N_5031,N_6181);
nand UO_879 (O_879,N_7566,N_5349);
nor UO_880 (O_880,N_7737,N_5802);
nor UO_881 (O_881,N_6357,N_5948);
or UO_882 (O_882,N_7825,N_6436);
and UO_883 (O_883,N_6011,N_5358);
or UO_884 (O_884,N_9770,N_5002);
xor UO_885 (O_885,N_5351,N_9818);
nand UO_886 (O_886,N_9247,N_7214);
and UO_887 (O_887,N_9972,N_8139);
and UO_888 (O_888,N_6444,N_6828);
xnor UO_889 (O_889,N_7914,N_9308);
and UO_890 (O_890,N_7489,N_7039);
or UO_891 (O_891,N_6255,N_9068);
or UO_892 (O_892,N_7076,N_8074);
xnor UO_893 (O_893,N_9433,N_7982);
nand UO_894 (O_894,N_7533,N_6188);
nand UO_895 (O_895,N_6385,N_8439);
xnor UO_896 (O_896,N_6524,N_6794);
nor UO_897 (O_897,N_5525,N_9529);
nor UO_898 (O_898,N_5616,N_5761);
and UO_899 (O_899,N_7666,N_5188);
nor UO_900 (O_900,N_8680,N_9985);
nand UO_901 (O_901,N_6952,N_9245);
and UO_902 (O_902,N_6531,N_7545);
nor UO_903 (O_903,N_6484,N_9563);
nor UO_904 (O_904,N_5934,N_9183);
or UO_905 (O_905,N_7442,N_6852);
and UO_906 (O_906,N_5271,N_7939);
nor UO_907 (O_907,N_8837,N_8210);
nand UO_908 (O_908,N_6759,N_7602);
nand UO_909 (O_909,N_9542,N_9079);
nand UO_910 (O_910,N_5495,N_6954);
nor UO_911 (O_911,N_9925,N_8811);
nor UO_912 (O_912,N_9279,N_9559);
and UO_913 (O_913,N_5094,N_7404);
or UO_914 (O_914,N_6490,N_6946);
nor UO_915 (O_915,N_7544,N_5367);
or UO_916 (O_916,N_9349,N_7559);
nor UO_917 (O_917,N_5245,N_9262);
xnor UO_918 (O_918,N_6692,N_5297);
nor UO_919 (O_919,N_6353,N_9608);
nand UO_920 (O_920,N_9915,N_8821);
nand UO_921 (O_921,N_5554,N_9705);
and UO_922 (O_922,N_6329,N_7869);
nor UO_923 (O_923,N_7218,N_5498);
nor UO_924 (O_924,N_7762,N_5444);
nand UO_925 (O_925,N_7536,N_6614);
or UO_926 (O_926,N_6185,N_9212);
nand UO_927 (O_927,N_8260,N_9663);
and UO_928 (O_928,N_8227,N_5114);
nand UO_929 (O_929,N_7640,N_6764);
xor UO_930 (O_930,N_6083,N_7004);
xor UO_931 (O_931,N_7508,N_5945);
nor UO_932 (O_932,N_8721,N_5037);
nand UO_933 (O_933,N_7196,N_8980);
nor UO_934 (O_934,N_7062,N_9170);
or UO_935 (O_935,N_6616,N_5773);
and UO_936 (O_936,N_8255,N_5569);
xnor UO_937 (O_937,N_5262,N_7052);
nor UO_938 (O_938,N_8161,N_5755);
and UO_939 (O_939,N_6841,N_6334);
nand UO_940 (O_940,N_9726,N_7085);
nand UO_941 (O_941,N_5230,N_6559);
or UO_942 (O_942,N_7611,N_5272);
or UO_943 (O_943,N_6180,N_7676);
nand UO_944 (O_944,N_7503,N_7176);
nor UO_945 (O_945,N_8269,N_5308);
or UO_946 (O_946,N_5941,N_7016);
nand UO_947 (O_947,N_7900,N_7682);
nor UO_948 (O_948,N_5079,N_7699);
and UO_949 (O_949,N_5051,N_9282);
nor UO_950 (O_950,N_5216,N_5748);
nand UO_951 (O_951,N_5636,N_6854);
or UO_952 (O_952,N_7290,N_8027);
xnor UO_953 (O_953,N_8986,N_6082);
nor UO_954 (O_954,N_8076,N_9625);
or UO_955 (O_955,N_9114,N_7199);
nand UO_956 (O_956,N_7857,N_7157);
nand UO_957 (O_957,N_8317,N_8119);
nor UO_958 (O_958,N_5877,N_9335);
nand UO_959 (O_959,N_5788,N_7775);
nor UO_960 (O_960,N_6416,N_6375);
and UO_961 (O_961,N_8547,N_7418);
nand UO_962 (O_962,N_6867,N_9909);
nand UO_963 (O_963,N_5301,N_6440);
or UO_964 (O_964,N_8982,N_6629);
nor UO_965 (O_965,N_6982,N_9198);
and UO_966 (O_966,N_7749,N_5791);
xor UO_967 (O_967,N_8550,N_9000);
and UO_968 (O_968,N_9795,N_6639);
and UO_969 (O_969,N_7758,N_6235);
nand UO_970 (O_970,N_7249,N_7860);
or UO_971 (O_971,N_8345,N_9904);
or UO_972 (O_972,N_7911,N_7094);
and UO_973 (O_973,N_5678,N_8292);
nand UO_974 (O_974,N_5104,N_8910);
xnor UO_975 (O_975,N_7820,N_7370);
or UO_976 (O_976,N_5242,N_9811);
and UO_977 (O_977,N_5341,N_8962);
nand UO_978 (O_978,N_5623,N_6997);
and UO_979 (O_979,N_8308,N_8407);
xor UO_980 (O_980,N_8166,N_9165);
nor UO_981 (O_981,N_8885,N_8571);
nand UO_982 (O_982,N_9902,N_6926);
nor UO_983 (O_983,N_7472,N_7069);
or UO_984 (O_984,N_9285,N_9373);
or UO_985 (O_985,N_9096,N_5720);
nand UO_986 (O_986,N_8352,N_7338);
and UO_987 (O_987,N_6781,N_7595);
or UO_988 (O_988,N_9696,N_7973);
nand UO_989 (O_989,N_6270,N_5732);
xor UO_990 (O_990,N_7492,N_9991);
nor UO_991 (O_991,N_9138,N_6499);
or UO_992 (O_992,N_6968,N_9503);
or UO_993 (O_993,N_7872,N_8674);
and UO_994 (O_994,N_9746,N_8997);
nor UO_995 (O_995,N_8701,N_6623);
nor UO_996 (O_996,N_5915,N_5286);
nor UO_997 (O_997,N_5925,N_9855);
and UO_998 (O_998,N_7623,N_7312);
nand UO_999 (O_999,N_9815,N_9830);
xor UO_1000 (O_1000,N_5885,N_5880);
and UO_1001 (O_1001,N_8183,N_6075);
and UO_1002 (O_1002,N_7800,N_6260);
or UO_1003 (O_1003,N_5085,N_5229);
xor UO_1004 (O_1004,N_9889,N_5499);
nand UO_1005 (O_1005,N_9986,N_7221);
nand UO_1006 (O_1006,N_7522,N_6618);
nor UO_1007 (O_1007,N_7054,N_5962);
nor UO_1008 (O_1008,N_7383,N_5445);
or UO_1009 (O_1009,N_9337,N_8666);
or UO_1010 (O_1010,N_6463,N_6447);
or UO_1011 (O_1011,N_5253,N_7245);
nand UO_1012 (O_1012,N_5247,N_5054);
nor UO_1013 (O_1013,N_5259,N_7972);
and UO_1014 (O_1014,N_9530,N_6258);
nor UO_1015 (O_1015,N_6100,N_6822);
or UO_1016 (O_1016,N_6676,N_5652);
xor UO_1017 (O_1017,N_6231,N_6424);
or UO_1018 (O_1018,N_8732,N_8586);
and UO_1019 (O_1019,N_8620,N_6161);
or UO_1020 (O_1020,N_6685,N_9736);
nor UO_1021 (O_1021,N_9063,N_6076);
or UO_1022 (O_1022,N_7517,N_6695);
xnor UO_1023 (O_1023,N_5380,N_7013);
nand UO_1024 (O_1024,N_7044,N_5291);
nor UO_1025 (O_1025,N_7886,N_8799);
or UO_1026 (O_1026,N_9217,N_6291);
nand UO_1027 (O_1027,N_6358,N_6771);
or UO_1028 (O_1028,N_8416,N_6810);
or UO_1029 (O_1029,N_9594,N_7345);
nor UO_1030 (O_1030,N_8020,N_6704);
or UO_1031 (O_1031,N_5883,N_7113);
and UO_1032 (O_1032,N_9711,N_6900);
nor UO_1033 (O_1033,N_8691,N_6211);
nand UO_1034 (O_1034,N_6920,N_9374);
nand UO_1035 (O_1035,N_9327,N_6169);
and UO_1036 (O_1036,N_9065,N_6908);
nand UO_1037 (O_1037,N_8748,N_9499);
and UO_1038 (O_1038,N_6673,N_5449);
nand UO_1039 (O_1039,N_9343,N_5352);
or UO_1040 (O_1040,N_6924,N_6843);
nor UO_1041 (O_1041,N_9093,N_8436);
and UO_1042 (O_1042,N_9927,N_7401);
nor UO_1043 (O_1043,N_8875,N_6749);
or UO_1044 (O_1044,N_6961,N_6609);
xor UO_1045 (O_1045,N_7674,N_6216);
or UO_1046 (O_1046,N_9256,N_8390);
nand UO_1047 (O_1047,N_5115,N_7979);
nor UO_1048 (O_1048,N_8873,N_8645);
and UO_1049 (O_1049,N_6146,N_6430);
nor UO_1050 (O_1050,N_5486,N_5298);
and UO_1051 (O_1051,N_7187,N_5667);
and UO_1052 (O_1052,N_7179,N_7634);
xor UO_1053 (O_1053,N_6980,N_5156);
nand UO_1054 (O_1054,N_8288,N_8306);
nor UO_1055 (O_1055,N_5252,N_7127);
nor UO_1056 (O_1056,N_5477,N_8134);
nor UO_1057 (O_1057,N_7581,N_8147);
xnor UO_1058 (O_1058,N_7975,N_8126);
nand UO_1059 (O_1059,N_5764,N_9727);
and UO_1060 (O_1060,N_7209,N_6483);
nor UO_1061 (O_1061,N_7952,N_6191);
nand UO_1062 (O_1062,N_6638,N_5605);
nand UO_1063 (O_1063,N_5662,N_6561);
xnor UO_1064 (O_1064,N_5314,N_5804);
or UO_1065 (O_1065,N_8677,N_6604);
nor UO_1066 (O_1066,N_6934,N_5087);
and UO_1067 (O_1067,N_9050,N_6574);
and UO_1068 (O_1068,N_8047,N_5938);
or UO_1069 (O_1069,N_5385,N_8189);
nand UO_1070 (O_1070,N_7550,N_7909);
or UO_1071 (O_1071,N_6514,N_8694);
and UO_1072 (O_1072,N_8477,N_9319);
xor UO_1073 (O_1073,N_5852,N_6006);
or UO_1074 (O_1074,N_9356,N_8809);
and UO_1075 (O_1075,N_8957,N_6089);
or UO_1076 (O_1076,N_7752,N_5907);
nand UO_1077 (O_1077,N_9948,N_5863);
nand UO_1078 (O_1078,N_7037,N_8676);
nand UO_1079 (O_1079,N_6306,N_7529);
or UO_1080 (O_1080,N_5175,N_8371);
nand UO_1081 (O_1081,N_9236,N_6244);
xor UO_1082 (O_1082,N_8452,N_5381);
and UO_1083 (O_1083,N_9518,N_9202);
or UO_1084 (O_1084,N_7732,N_5462);
xnor UO_1085 (O_1085,N_7576,N_6410);
nand UO_1086 (O_1086,N_6277,N_6072);
or UO_1087 (O_1087,N_9193,N_7725);
nor UO_1088 (O_1088,N_9431,N_8778);
nor UO_1089 (O_1089,N_6415,N_5110);
or UO_1090 (O_1090,N_5348,N_6283);
and UO_1091 (O_1091,N_6710,N_9716);
or UO_1092 (O_1092,N_7484,N_5567);
and UO_1093 (O_1093,N_8801,N_5818);
or UO_1094 (O_1094,N_6990,N_9739);
nand UO_1095 (O_1095,N_7476,N_6066);
nor UO_1096 (O_1096,N_8646,N_7146);
or UO_1097 (O_1097,N_7095,N_6825);
and UO_1098 (O_1098,N_5273,N_6678);
and UO_1099 (O_1099,N_6652,N_8341);
and UO_1100 (O_1100,N_9651,N_8743);
or UO_1101 (O_1101,N_5835,N_9947);
or UO_1102 (O_1102,N_7579,N_9735);
nand UO_1103 (O_1103,N_9496,N_7361);
nand UO_1104 (O_1104,N_6465,N_5595);
nand UO_1105 (O_1105,N_6111,N_8043);
or UO_1106 (O_1106,N_5303,N_5968);
and UO_1107 (O_1107,N_7920,N_9567);
and UO_1108 (O_1108,N_5292,N_8230);
or UO_1109 (O_1109,N_5074,N_7364);
xor UO_1110 (O_1110,N_6949,N_6569);
and UO_1111 (O_1111,N_6487,N_8516);
and UO_1112 (O_1112,N_5874,N_8864);
nor UO_1113 (O_1113,N_7022,N_8971);
and UO_1114 (O_1114,N_5096,N_9174);
or UO_1115 (O_1115,N_5922,N_7262);
and UO_1116 (O_1116,N_5704,N_8685);
and UO_1117 (O_1117,N_5905,N_8356);
nor UO_1118 (O_1118,N_7012,N_8925);
nor UO_1119 (O_1119,N_7090,N_6142);
nor UO_1120 (O_1120,N_9218,N_7122);
and UO_1121 (O_1121,N_8643,N_9427);
or UO_1122 (O_1122,N_8017,N_6138);
or UO_1123 (O_1123,N_7890,N_5312);
or UO_1124 (O_1124,N_8927,N_9725);
and UO_1125 (O_1125,N_5493,N_5075);
nand UO_1126 (O_1126,N_5919,N_7366);
nor UO_1127 (O_1127,N_7573,N_6713);
nor UO_1128 (O_1128,N_8220,N_9621);
or UO_1129 (O_1129,N_5867,N_6176);
xor UO_1130 (O_1130,N_7321,N_6570);
or UO_1131 (O_1131,N_9415,N_6669);
and UO_1132 (O_1132,N_7305,N_9181);
or UO_1133 (O_1133,N_8581,N_6681);
and UO_1134 (O_1134,N_7276,N_7904);
or UO_1135 (O_1135,N_5035,N_6661);
nand UO_1136 (O_1136,N_5635,N_9887);
nor UO_1137 (O_1137,N_7734,N_6610);
and UO_1138 (O_1138,N_9126,N_8488);
nor UO_1139 (O_1139,N_7439,N_8921);
nand UO_1140 (O_1140,N_9635,N_7746);
and UO_1141 (O_1141,N_5932,N_5211);
xor UO_1142 (O_1142,N_9510,N_7264);
and UO_1143 (O_1143,N_8641,N_7597);
and UO_1144 (O_1144,N_5734,N_8256);
or UO_1145 (O_1145,N_5870,N_6457);
nand UO_1146 (O_1146,N_5573,N_9188);
nand UO_1147 (O_1147,N_5676,N_7163);
or UO_1148 (O_1148,N_9449,N_9083);
or UO_1149 (O_1149,N_5318,N_9786);
or UO_1150 (O_1150,N_6378,N_6434);
nor UO_1151 (O_1151,N_8561,N_8546);
nor UO_1152 (O_1152,N_9964,N_5602);
nor UO_1153 (O_1153,N_5071,N_5003);
and UO_1154 (O_1154,N_7983,N_7861);
nand UO_1155 (O_1155,N_8368,N_7409);
and UO_1156 (O_1156,N_6516,N_7802);
nand UO_1157 (O_1157,N_9789,N_7093);
xnor UO_1158 (O_1158,N_8279,N_5710);
nor UO_1159 (O_1159,N_9564,N_9258);
nor UO_1160 (O_1160,N_7984,N_8337);
xor UO_1161 (O_1161,N_5432,N_7708);
nor UO_1162 (O_1162,N_8014,N_6986);
and UO_1163 (O_1163,N_7957,N_5875);
nor UO_1164 (O_1164,N_5215,N_6109);
or UO_1165 (O_1165,N_8978,N_6275);
nor UO_1166 (O_1166,N_9630,N_9546);
nor UO_1167 (O_1167,N_8839,N_8824);
nor UO_1168 (O_1168,N_9304,N_6094);
nand UO_1169 (O_1169,N_6998,N_5576);
nand UO_1170 (O_1170,N_9710,N_6542);
or UO_1171 (O_1171,N_9085,N_6565);
nand UO_1172 (O_1172,N_9644,N_7741);
nor UO_1173 (O_1173,N_6551,N_6136);
or UO_1174 (O_1174,N_8353,N_9489);
xnor UO_1175 (O_1175,N_7691,N_6921);
nor UO_1176 (O_1176,N_7552,N_7624);
and UO_1177 (O_1177,N_5376,N_6399);
nand UO_1178 (O_1178,N_9946,N_9257);
nor UO_1179 (O_1179,N_8692,N_6388);
and UO_1180 (O_1180,N_8973,N_9691);
nor UO_1181 (O_1181,N_5261,N_5640);
or UO_1182 (O_1182,N_8716,N_6528);
or UO_1183 (O_1183,N_6743,N_8810);
or UO_1184 (O_1184,N_5980,N_6101);
nand UO_1185 (O_1185,N_6199,N_7118);
or UO_1186 (O_1186,N_5160,N_5969);
xor UO_1187 (O_1187,N_5840,N_7327);
nand UO_1188 (O_1188,N_6889,N_6788);
and UO_1189 (O_1189,N_5473,N_7527);
and UO_1190 (O_1190,N_5633,N_5026);
and UO_1191 (O_1191,N_7084,N_7754);
nand UO_1192 (O_1192,N_7659,N_8771);
or UO_1193 (O_1193,N_5590,N_9424);
or UO_1194 (O_1194,N_6807,N_9070);
nor UO_1195 (O_1195,N_7932,N_6705);
xor UO_1196 (O_1196,N_8058,N_6309);
nand UO_1197 (O_1197,N_6546,N_7643);
or UO_1198 (O_1198,N_8920,N_7551);
or UO_1199 (O_1199,N_6091,N_6809);
nor UO_1200 (O_1200,N_5254,N_9952);
nor UO_1201 (O_1201,N_7694,N_7251);
and UO_1202 (O_1202,N_6401,N_7884);
nor UO_1203 (O_1203,N_7814,N_9741);
or UO_1204 (O_1204,N_5421,N_5117);
nand UO_1205 (O_1205,N_6125,N_9035);
nand UO_1206 (O_1206,N_5090,N_5098);
nand UO_1207 (O_1207,N_6523,N_5551);
and UO_1208 (O_1208,N_8756,N_7562);
xor UO_1209 (O_1209,N_7943,N_7077);
nand UO_1210 (O_1210,N_9888,N_5227);
nor UO_1211 (O_1211,N_8595,N_6861);
and UO_1212 (O_1212,N_6202,N_7571);
nor UO_1213 (O_1213,N_8551,N_6554);
nor UO_1214 (O_1214,N_8729,N_8639);
nor UO_1215 (O_1215,N_9622,N_6315);
or UO_1216 (O_1216,N_5580,N_6482);
nor UO_1217 (O_1217,N_9106,N_7183);
and UO_1218 (O_1218,N_7965,N_7554);
or UO_1219 (O_1219,N_6227,N_7491);
or UO_1220 (O_1220,N_7927,N_5507);
and UO_1221 (O_1221,N_7448,N_8905);
nand UO_1222 (O_1222,N_8327,N_9858);
and UO_1223 (O_1223,N_9483,N_6187);
or UO_1224 (O_1224,N_9493,N_8850);
nor UO_1225 (O_1225,N_8475,N_8745);
and UO_1226 (O_1226,N_6509,N_9086);
and UO_1227 (O_1227,N_5333,N_9714);
or UO_1228 (O_1228,N_7100,N_7675);
nor UO_1229 (O_1229,N_8019,N_7032);
nor UO_1230 (O_1230,N_7885,N_9940);
and UO_1231 (O_1231,N_5550,N_5792);
and UO_1232 (O_1232,N_5899,N_5985);
nand UO_1233 (O_1233,N_9197,N_8247);
xor UO_1234 (O_1234,N_9773,N_8533);
nand UO_1235 (O_1235,N_5529,N_6964);
and UO_1236 (O_1236,N_8803,N_9841);
nand UO_1237 (O_1237,N_9944,N_8208);
nand UO_1238 (O_1238,N_9713,N_9717);
nand UO_1239 (O_1239,N_7923,N_9892);
and UO_1240 (O_1240,N_9314,N_8160);
and UO_1241 (O_1241,N_6323,N_6279);
nor UO_1242 (O_1242,N_9914,N_6064);
or UO_1243 (O_1243,N_5682,N_8907);
xnor UO_1244 (O_1244,N_8103,N_8426);
nor UO_1245 (O_1245,N_9199,N_5007);
or UO_1246 (O_1246,N_5236,N_9334);
and UO_1247 (O_1247,N_8012,N_6803);
nor UO_1248 (O_1248,N_7463,N_6214);
or UO_1249 (O_1249,N_6304,N_7371);
and UO_1250 (O_1250,N_5195,N_7142);
nor UO_1251 (O_1251,N_9275,N_6651);
and UO_1252 (O_1252,N_9803,N_7259);
nor UO_1253 (O_1253,N_9581,N_7431);
nor UO_1254 (O_1254,N_7769,N_6752);
and UO_1255 (O_1255,N_5542,N_8619);
or UO_1256 (O_1256,N_5059,N_7667);
or UO_1257 (O_1257,N_8102,N_9817);
and UO_1258 (O_1258,N_7020,N_5060);
or UO_1259 (O_1259,N_5705,N_5013);
nand UO_1260 (O_1260,N_7514,N_7078);
nor UO_1261 (O_1261,N_6368,N_6503);
nand UO_1262 (O_1262,N_6727,N_6851);
or UO_1263 (O_1263,N_7759,N_9574);
and UO_1264 (O_1264,N_6855,N_5138);
and UO_1265 (O_1265,N_9913,N_8079);
and UO_1266 (O_1266,N_5472,N_9037);
nand UO_1267 (O_1267,N_9885,N_5483);
or UO_1268 (O_1268,N_6703,N_7468);
and UO_1269 (O_1269,N_8543,N_6496);
nand UO_1270 (O_1270,N_7680,N_8710);
nor UO_1271 (O_1271,N_7103,N_9191);
and UO_1272 (O_1272,N_7524,N_8618);
nand UO_1273 (O_1273,N_8321,N_6050);
nand UO_1274 (O_1274,N_7201,N_6172);
or UO_1275 (O_1275,N_8950,N_8829);
nand UO_1276 (O_1276,N_9117,N_5199);
or UO_1277 (O_1277,N_5337,N_9768);
or UO_1278 (O_1278,N_8622,N_5779);
nand UO_1279 (O_1279,N_5707,N_8915);
nand UO_1280 (O_1280,N_5131,N_8542);
nand UO_1281 (O_1281,N_9893,N_6249);
and UO_1282 (O_1282,N_7386,N_5233);
nand UO_1283 (O_1283,N_7018,N_9759);
xnor UO_1284 (O_1284,N_5063,N_9806);
or UO_1285 (O_1285,N_8448,N_8640);
nand UO_1286 (O_1286,N_9179,N_5816);
nor UO_1287 (O_1287,N_8626,N_8444);
or UO_1288 (O_1288,N_9099,N_8913);
nor UO_1289 (O_1289,N_8531,N_7846);
or UO_1290 (O_1290,N_8871,N_7605);
and UO_1291 (O_1291,N_8777,N_9601);
and UO_1292 (O_1292,N_5088,N_8582);
nand UO_1293 (O_1293,N_5760,N_5637);
xor UO_1294 (O_1294,N_8860,N_5471);
and UO_1295 (O_1295,N_6838,N_7348);
or UO_1296 (O_1296,N_6772,N_8046);
and UO_1297 (O_1297,N_8898,N_9397);
or UO_1298 (O_1298,N_6670,N_7469);
nor UO_1299 (O_1299,N_9219,N_7445);
nand UO_1300 (O_1300,N_6402,N_7478);
and UO_1301 (O_1301,N_5396,N_8242);
nor UO_1302 (O_1302,N_5995,N_9246);
or UO_1303 (O_1303,N_9053,N_5860);
and UO_1304 (O_1304,N_8086,N_5509);
nand UO_1305 (O_1305,N_9186,N_8922);
or UO_1306 (O_1306,N_5289,N_5672);
nand UO_1307 (O_1307,N_7839,N_7913);
nor UO_1308 (O_1308,N_6015,N_6152);
and UO_1309 (O_1309,N_8869,N_5561);
xor UO_1310 (O_1310,N_6619,N_5967);
nand UO_1311 (O_1311,N_7794,N_6435);
nor UO_1312 (O_1312,N_9754,N_5307);
nand UO_1313 (O_1313,N_8163,N_9016);
or UO_1314 (O_1314,N_5750,N_5956);
or UO_1315 (O_1315,N_5127,N_5005);
xor UO_1316 (O_1316,N_9989,N_8827);
nand UO_1317 (O_1317,N_9422,N_6195);
and UO_1318 (O_1318,N_6148,N_9508);
nand UO_1319 (O_1319,N_6020,N_6916);
and UO_1320 (O_1320,N_9640,N_8159);
nand UO_1321 (O_1321,N_9679,N_8993);
nand UO_1322 (O_1322,N_5989,N_9852);
and UO_1323 (O_1323,N_6269,N_5162);
or UO_1324 (O_1324,N_5696,N_5698);
and UO_1325 (O_1325,N_7921,N_5239);
and UO_1326 (O_1326,N_6933,N_7582);
nand UO_1327 (O_1327,N_6874,N_8301);
nor UO_1328 (O_1328,N_6139,N_6539);
xor UO_1329 (O_1329,N_9064,N_5092);
or UO_1330 (O_1330,N_9194,N_7048);
nor UO_1331 (O_1331,N_7210,N_6547);
or UO_1332 (O_1332,N_9612,N_9880);
nor UO_1333 (O_1333,N_5909,N_7310);
nand UO_1334 (O_1334,N_8886,N_8795);
and UO_1335 (O_1335,N_6868,N_8662);
and UO_1336 (O_1336,N_7797,N_7248);
nor UO_1337 (O_1337,N_7482,N_7681);
nor UO_1338 (O_1338,N_5158,N_5355);
nand UO_1339 (O_1339,N_6888,N_5411);
nor UO_1340 (O_1340,N_6662,N_8936);
and UO_1341 (O_1341,N_8532,N_6572);
and UO_1342 (O_1342,N_9376,N_5033);
or UO_1343 (O_1343,N_9619,N_6603);
nand UO_1344 (O_1344,N_9419,N_7590);
xnor UO_1345 (O_1345,N_5404,N_5402);
and UO_1346 (O_1346,N_7172,N_9402);
xnor UO_1347 (O_1347,N_8891,N_7947);
nand UO_1348 (O_1348,N_5466,N_9460);
and UO_1349 (O_1349,N_8262,N_8888);
nand UO_1350 (O_1350,N_7876,N_8388);
or UO_1351 (O_1351,N_9680,N_6361);
and UO_1352 (O_1352,N_7763,N_8330);
or UO_1353 (O_1353,N_7174,N_5903);
nor UO_1354 (O_1354,N_7693,N_6541);
xnor UO_1355 (O_1355,N_8471,N_8903);
nor UO_1356 (O_1356,N_9056,N_9844);
nand UO_1357 (O_1357,N_5793,N_7816);
nand UO_1358 (O_1358,N_7696,N_7852);
and UO_1359 (O_1359,N_5506,N_9755);
nor UO_1360 (O_1360,N_8584,N_6801);
nor UO_1361 (O_1361,N_9104,N_9950);
or UO_1362 (O_1362,N_5502,N_8150);
xnor UO_1363 (O_1363,N_5258,N_7225);
or UO_1364 (O_1364,N_6969,N_9122);
and UO_1365 (O_1365,N_9878,N_9512);
nand UO_1366 (O_1366,N_9029,N_5374);
or UO_1367 (O_1367,N_7145,N_9209);
nand UO_1368 (O_1368,N_7056,N_6797);
xnor UO_1369 (O_1369,N_7363,N_8508);
and UO_1370 (O_1370,N_6099,N_8071);
xnor UO_1371 (O_1371,N_7849,N_8485);
nand UO_1372 (O_1372,N_6722,N_9609);
xor UO_1373 (O_1373,N_7407,N_6480);
nand UO_1374 (O_1374,N_8707,N_8635);
nand UO_1375 (O_1375,N_5868,N_8338);
or UO_1376 (O_1376,N_9620,N_8750);
or UO_1377 (O_1377,N_7377,N_8177);
nor UO_1378 (O_1378,N_8114,N_7612);
or UO_1379 (O_1379,N_6930,N_5070);
nand UO_1380 (O_1380,N_9299,N_8151);
or UO_1381 (O_1381,N_9289,N_5515);
or UO_1382 (O_1382,N_5391,N_7286);
and UO_1383 (O_1383,N_5829,N_8408);
and UO_1384 (O_1384,N_7158,N_7664);
or UO_1385 (O_1385,N_8816,N_7131);
xor UO_1386 (O_1386,N_5221,N_5815);
and UO_1387 (O_1387,N_7072,N_8329);
xnor UO_1388 (O_1388,N_9298,N_6341);
nand UO_1389 (O_1389,N_5853,N_6407);
nor UO_1390 (O_1390,N_9846,N_8796);
nor UO_1391 (O_1391,N_6826,N_8015);
nand UO_1392 (O_1392,N_6299,N_8146);
nand UO_1393 (O_1393,N_9654,N_5872);
xnor UO_1394 (O_1394,N_6655,N_7647);
nor UO_1395 (O_1395,N_6359,N_9412);
nand UO_1396 (O_1396,N_8615,N_9560);
nand UO_1397 (O_1397,N_7565,N_6294);
or UO_1398 (O_1398,N_9996,N_6786);
nand UO_1399 (O_1399,N_8537,N_5326);
nand UO_1400 (O_1400,N_8274,N_7589);
or UO_1401 (O_1401,N_8846,N_6467);
and UO_1402 (O_1402,N_8780,N_6023);
nand UO_1403 (O_1403,N_9482,N_8567);
nand UO_1404 (O_1404,N_9921,N_5603);
nand UO_1405 (O_1405,N_6605,N_6942);
nor UO_1406 (O_1406,N_6073,N_8953);
nor UO_1407 (O_1407,N_8359,N_6717);
nand UO_1408 (O_1408,N_7824,N_8872);
and UO_1409 (O_1409,N_7217,N_5879);
and UO_1410 (O_1410,N_8424,N_8474);
xnor UO_1411 (O_1411,N_7528,N_7819);
nor UO_1412 (O_1412,N_5996,N_9820);
nor UO_1413 (O_1413,N_5864,N_7855);
or UO_1414 (O_1414,N_9328,N_7574);
or UO_1415 (O_1415,N_9774,N_5532);
or UO_1416 (O_1416,N_6002,N_6557);
xor UO_1417 (O_1417,N_9395,N_5049);
and UO_1418 (O_1418,N_7831,N_7631);
and UO_1419 (O_1419,N_6106,N_8094);
or UO_1420 (O_1420,N_7698,N_6575);
nand UO_1421 (O_1421,N_8310,N_8773);
nand UO_1422 (O_1422,N_6594,N_9240);
or UO_1423 (O_1423,N_9781,N_7220);
and UO_1424 (O_1424,N_6090,N_9180);
nor UO_1425 (O_1425,N_6819,N_8868);
nand UO_1426 (O_1426,N_7660,N_9233);
nor UO_1427 (O_1427,N_9930,N_6022);
or UO_1428 (O_1428,N_5618,N_9816);
and UO_1429 (O_1429,N_7997,N_8790);
or UO_1430 (O_1430,N_8303,N_9777);
or UO_1431 (O_1431,N_8847,N_5340);
nor UO_1432 (O_1432,N_6053,N_7204);
xnor UO_1433 (O_1433,N_9617,N_5277);
or UO_1434 (O_1434,N_8517,N_8887);
and UO_1435 (O_1435,N_5609,N_6612);
xor UO_1436 (O_1436,N_7945,N_9386);
or UO_1437 (O_1437,N_8511,N_6228);
or UO_1438 (O_1438,N_8259,N_5334);
nand UO_1439 (O_1439,N_9024,N_9336);
and UO_1440 (O_1440,N_7583,N_7317);
or UO_1441 (O_1441,N_7309,N_8203);
nand UO_1442 (O_1442,N_5714,N_7435);
nor UO_1443 (O_1443,N_6056,N_5280);
nand UO_1444 (O_1444,N_9709,N_7289);
xor UO_1445 (O_1445,N_6039,N_7089);
xnor UO_1446 (O_1446,N_8559,N_9626);
and UO_1447 (O_1447,N_8713,N_5892);
and UO_1448 (O_1448,N_6744,N_5947);
or UO_1449 (O_1449,N_8478,N_6225);
xnor UO_1450 (O_1450,N_8782,N_7304);
xor UO_1451 (O_1451,N_6701,N_9265);
nor UO_1452 (O_1452,N_7186,N_6766);
or UO_1453 (O_1453,N_6367,N_7730);
nor UO_1454 (O_1454,N_8324,N_5758);
nand UO_1455 (O_1455,N_7601,N_6983);
nor UO_1456 (O_1456,N_7111,N_6025);
or UO_1457 (O_1457,N_8686,N_5577);
nand UO_1458 (O_1458,N_5354,N_8746);
nand UO_1459 (O_1459,N_9627,N_5949);
nor UO_1460 (O_1460,N_9514,N_5017);
nand UO_1461 (O_1461,N_8386,N_5330);
and UO_1462 (O_1462,N_7452,N_8044);
nand UO_1463 (O_1463,N_6095,N_5172);
and UO_1464 (O_1464,N_8229,N_6158);
and UO_1465 (O_1465,N_8088,N_6711);
and UO_1466 (O_1466,N_9206,N_6335);
or UO_1467 (O_1467,N_6473,N_9162);
nand UO_1468 (O_1468,N_5610,N_5235);
nor UO_1469 (O_1469,N_9966,N_5546);
nand UO_1470 (O_1470,N_7415,N_9801);
nand UO_1471 (O_1471,N_7962,N_9550);
and UO_1472 (O_1472,N_7917,N_8684);
xnor UO_1473 (O_1473,N_9440,N_8998);
nand UO_1474 (O_1474,N_8941,N_8181);
nor UO_1475 (O_1475,N_8947,N_7454);
or UO_1476 (O_1476,N_8945,N_9544);
and UO_1477 (O_1477,N_5036,N_8704);
nand UO_1478 (O_1478,N_7692,N_9864);
nor UO_1479 (O_1479,N_6832,N_9261);
nor UO_1480 (O_1480,N_5774,N_6640);
and UO_1481 (O_1481,N_9556,N_8841);
or UO_1482 (O_1482,N_8528,N_6636);
nand UO_1483 (O_1483,N_9970,N_5522);
nand UO_1484 (O_1484,N_5991,N_8760);
xor UO_1485 (O_1485,N_6694,N_6405);
xor UO_1486 (O_1486,N_9797,N_8101);
xnor UO_1487 (O_1487,N_9597,N_8481);
and UO_1488 (O_1488,N_5929,N_7055);
and UO_1489 (O_1489,N_9274,N_9207);
and UO_1490 (O_1490,N_6102,N_6525);
and UO_1491 (O_1491,N_7540,N_6092);
nor UO_1492 (O_1492,N_7344,N_7474);
or UO_1493 (O_1493,N_8744,N_7323);
or UO_1494 (O_1494,N_6666,N_7380);
or UO_1495 (O_1495,N_5961,N_6084);
nor UO_1496 (O_1496,N_9066,N_8800);
or UO_1497 (O_1497,N_7046,N_9454);
or UO_1498 (O_1498,N_6428,N_5454);
or UO_1499 (O_1499,N_9587,N_5942);
endmodule