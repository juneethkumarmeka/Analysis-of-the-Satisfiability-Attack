module basic_500_3000_500_6_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_221,In_189);
nor U1 (N_1,In_140,In_238);
or U2 (N_2,In_10,In_42);
or U3 (N_3,In_473,In_173);
nor U4 (N_4,In_459,In_142);
and U5 (N_5,In_145,In_39);
nor U6 (N_6,In_37,In_261);
nor U7 (N_7,In_5,In_74);
and U8 (N_8,In_301,In_223);
nor U9 (N_9,In_69,In_254);
or U10 (N_10,In_493,In_179);
nand U11 (N_11,In_81,In_316);
xnor U12 (N_12,In_488,In_117);
nand U13 (N_13,In_495,In_460);
xor U14 (N_14,In_298,In_61);
and U15 (N_15,In_129,In_426);
and U16 (N_16,In_165,In_484);
and U17 (N_17,In_198,In_480);
nor U18 (N_18,In_367,In_479);
or U19 (N_19,In_333,In_437);
nand U20 (N_20,In_359,In_497);
nand U21 (N_21,In_427,In_180);
or U22 (N_22,In_160,In_343);
nand U23 (N_23,In_197,In_88);
and U24 (N_24,In_187,In_279);
nor U25 (N_25,In_162,In_410);
and U26 (N_26,In_428,In_490);
and U27 (N_27,In_123,In_195);
xnor U28 (N_28,In_483,In_355);
nand U29 (N_29,In_85,In_40);
or U30 (N_30,In_463,In_26);
nand U31 (N_31,In_18,In_327);
or U32 (N_32,In_66,In_138);
xor U33 (N_33,In_245,In_361);
nand U34 (N_34,In_171,In_84);
and U35 (N_35,In_260,In_475);
nand U36 (N_36,In_143,In_407);
and U37 (N_37,In_275,In_309);
nand U38 (N_38,In_55,In_283);
or U39 (N_39,In_93,In_289);
or U40 (N_40,In_400,In_101);
nand U41 (N_41,In_9,In_276);
nor U42 (N_42,In_401,In_97);
or U43 (N_43,In_386,In_284);
or U44 (N_44,In_114,In_65);
or U45 (N_45,In_226,In_227);
nand U46 (N_46,In_194,In_295);
nand U47 (N_47,In_132,In_73);
or U48 (N_48,In_159,In_397);
xor U49 (N_49,In_373,In_15);
and U50 (N_50,In_371,In_71);
nand U51 (N_51,In_469,In_486);
nor U52 (N_52,In_100,In_431);
nor U53 (N_53,In_318,In_21);
nor U54 (N_54,In_24,In_322);
nor U55 (N_55,In_340,In_471);
and U56 (N_56,In_399,In_91);
nor U57 (N_57,In_476,In_262);
nor U58 (N_58,In_225,In_478);
or U59 (N_59,In_169,In_263);
and U60 (N_60,In_420,In_278);
and U61 (N_61,In_439,In_119);
nand U62 (N_62,In_308,In_383);
and U63 (N_63,In_141,In_103);
or U64 (N_64,In_115,In_163);
or U65 (N_65,In_4,In_376);
nor U66 (N_66,In_153,In_259);
and U67 (N_67,In_267,In_252);
and U68 (N_68,In_303,In_89);
nand U69 (N_69,In_216,In_498);
and U70 (N_70,In_369,In_205);
nand U71 (N_71,In_248,In_434);
nor U72 (N_72,In_315,In_464);
nand U73 (N_73,In_416,In_419);
or U74 (N_74,In_111,In_36);
nand U75 (N_75,In_19,In_20);
nand U76 (N_76,In_80,In_154);
nand U77 (N_77,In_255,In_335);
or U78 (N_78,In_177,In_213);
and U79 (N_79,In_445,In_474);
nor U80 (N_80,In_121,In_210);
nor U81 (N_81,In_362,In_294);
nor U82 (N_82,In_304,In_357);
and U83 (N_83,In_249,In_212);
xor U84 (N_84,In_417,In_29);
nor U85 (N_85,In_452,In_405);
nand U86 (N_86,In_388,In_125);
nand U87 (N_87,In_235,In_449);
and U88 (N_88,In_395,In_456);
nor U89 (N_89,In_146,In_224);
or U90 (N_90,In_257,In_51);
nor U91 (N_91,In_368,In_457);
nand U92 (N_92,In_67,In_34);
nor U93 (N_93,In_448,In_329);
nor U94 (N_94,In_482,In_70);
nand U95 (N_95,In_59,In_202);
nand U96 (N_96,In_72,In_349);
and U97 (N_97,In_491,In_82);
and U98 (N_98,In_63,In_364);
or U99 (N_99,In_323,In_351);
xnor U100 (N_100,In_46,In_353);
xnor U101 (N_101,In_320,In_326);
nor U102 (N_102,In_305,In_291);
xor U103 (N_103,In_77,In_370);
and U104 (N_104,In_172,In_50);
xnor U105 (N_105,In_130,In_219);
nor U106 (N_106,In_363,In_387);
and U107 (N_107,In_496,In_414);
xnor U108 (N_108,In_489,In_499);
nand U109 (N_109,In_60,In_433);
xor U110 (N_110,In_196,In_404);
and U111 (N_111,In_477,In_237);
nor U112 (N_112,In_211,In_185);
nor U113 (N_113,In_30,In_175);
or U114 (N_114,In_157,In_207);
and U115 (N_115,In_453,In_191);
and U116 (N_116,In_147,In_287);
or U117 (N_117,In_306,In_268);
and U118 (N_118,In_243,In_253);
nand U119 (N_119,In_347,In_168);
and U120 (N_120,In_328,In_454);
and U121 (N_121,In_150,In_311);
nor U122 (N_122,In_265,In_466);
nor U123 (N_123,In_273,In_57);
or U124 (N_124,In_461,In_403);
xnor U125 (N_125,In_319,In_22);
and U126 (N_126,In_113,In_214);
or U127 (N_127,In_174,In_470);
and U128 (N_128,In_48,In_274);
and U129 (N_129,In_2,In_421);
and U130 (N_130,In_424,In_418);
or U131 (N_131,In_487,In_124);
or U132 (N_132,In_110,In_393);
and U133 (N_133,In_94,In_133);
and U134 (N_134,In_17,In_321);
or U135 (N_135,In_348,In_256);
nand U136 (N_136,In_345,In_366);
nand U137 (N_137,In_365,In_78);
or U138 (N_138,In_352,In_167);
nand U139 (N_139,In_99,In_107);
and U140 (N_140,In_247,In_209);
or U141 (N_141,In_156,In_109);
nand U142 (N_142,In_155,In_86);
nor U143 (N_143,In_152,In_356);
nand U144 (N_144,In_242,In_6);
nand U145 (N_145,In_442,In_217);
or U146 (N_146,In_317,In_409);
and U147 (N_147,In_170,In_390);
nor U148 (N_148,In_413,In_331);
and U149 (N_149,In_98,In_446);
nand U150 (N_150,In_258,In_415);
nor U151 (N_151,In_35,In_104);
or U152 (N_152,In_151,In_408);
nand U153 (N_153,In_344,In_282);
and U154 (N_154,In_325,In_105);
nor U155 (N_155,In_465,In_389);
and U156 (N_156,In_139,In_203);
and U157 (N_157,In_87,In_447);
and U158 (N_158,In_336,In_467);
and U159 (N_159,In_451,In_128);
and U160 (N_160,In_96,In_79);
and U161 (N_161,In_443,In_38);
nand U162 (N_162,In_334,In_28);
and U163 (N_163,In_302,In_307);
nor U164 (N_164,In_206,In_0);
xor U165 (N_165,In_58,In_250);
xnor U166 (N_166,In_337,In_190);
nand U167 (N_167,In_296,In_269);
nor U168 (N_168,In_312,In_494);
and U169 (N_169,In_430,In_137);
and U170 (N_170,In_354,In_485);
and U171 (N_171,In_468,In_135);
and U172 (N_172,In_240,In_178);
xor U173 (N_173,In_8,In_49);
nor U174 (N_174,In_444,In_14);
nor U175 (N_175,In_200,In_350);
nor U176 (N_176,In_241,In_90);
and U177 (N_177,In_338,In_234);
nor U178 (N_178,In_481,In_218);
nand U179 (N_179,In_68,In_183);
or U180 (N_180,In_184,In_392);
and U181 (N_181,In_64,In_31);
and U182 (N_182,In_375,In_285);
or U183 (N_183,In_56,In_229);
or U184 (N_184,In_62,In_435);
nor U185 (N_185,In_92,In_292);
nor U186 (N_186,In_272,In_228);
or U187 (N_187,In_423,In_27);
and U188 (N_188,In_396,In_116);
or U189 (N_189,In_324,In_458);
nor U190 (N_190,In_358,In_134);
nand U191 (N_191,In_166,In_339);
or U192 (N_192,In_472,In_215);
or U193 (N_193,In_441,In_346);
nand U194 (N_194,In_384,In_300);
or U195 (N_195,In_233,In_54);
nor U196 (N_196,In_425,In_16);
nor U197 (N_197,In_264,In_83);
nor U198 (N_198,In_32,In_290);
or U199 (N_199,In_161,In_127);
or U200 (N_200,In_412,In_379);
nand U201 (N_201,In_313,In_186);
or U202 (N_202,In_158,In_251);
or U203 (N_203,In_193,In_126);
nand U204 (N_204,In_372,In_181);
and U205 (N_205,In_246,In_381);
or U206 (N_206,In_342,In_148);
nand U207 (N_207,In_25,In_402);
xnor U208 (N_208,In_394,In_332);
nor U209 (N_209,In_230,In_33);
or U210 (N_210,In_314,In_47);
nand U211 (N_211,In_108,In_45);
xnor U212 (N_212,In_75,In_231);
nor U213 (N_213,In_438,In_52);
xnor U214 (N_214,In_360,In_199);
nor U215 (N_215,In_244,In_297);
nor U216 (N_216,In_44,In_293);
and U217 (N_217,In_222,In_3);
or U218 (N_218,In_422,In_406);
and U219 (N_219,In_102,In_236);
or U220 (N_220,In_112,In_436);
or U221 (N_221,In_43,In_374);
xor U222 (N_222,In_232,In_122);
and U223 (N_223,In_7,In_398);
nor U224 (N_224,In_380,In_53);
nor U225 (N_225,In_13,In_149);
xnor U226 (N_226,In_286,In_204);
and U227 (N_227,In_385,In_377);
or U228 (N_228,In_11,In_330);
nand U229 (N_229,In_462,In_271);
and U230 (N_230,In_391,In_118);
or U231 (N_231,In_23,In_280);
and U232 (N_232,In_164,In_310);
and U233 (N_233,In_266,In_201);
or U234 (N_234,In_220,In_76);
or U235 (N_235,In_288,In_270);
or U236 (N_236,In_1,In_176);
nor U237 (N_237,In_182,In_106);
or U238 (N_238,In_192,In_382);
nand U239 (N_239,In_144,In_281);
nor U240 (N_240,In_95,In_41);
nand U241 (N_241,In_12,In_455);
nor U242 (N_242,In_299,In_188);
nand U243 (N_243,In_341,In_492);
nor U244 (N_244,In_378,In_120);
or U245 (N_245,In_432,In_136);
nor U246 (N_246,In_411,In_440);
nand U247 (N_247,In_239,In_450);
or U248 (N_248,In_277,In_429);
or U249 (N_249,In_131,In_208);
xnor U250 (N_250,In_433,In_119);
nand U251 (N_251,In_264,In_249);
nor U252 (N_252,In_281,In_363);
xnor U253 (N_253,In_78,In_268);
and U254 (N_254,In_316,In_146);
nand U255 (N_255,In_69,In_416);
nor U256 (N_256,In_424,In_474);
nand U257 (N_257,In_22,In_89);
nor U258 (N_258,In_129,In_409);
nand U259 (N_259,In_470,In_403);
or U260 (N_260,In_46,In_125);
nor U261 (N_261,In_244,In_34);
nand U262 (N_262,In_150,In_124);
and U263 (N_263,In_123,In_296);
nor U264 (N_264,In_30,In_236);
nand U265 (N_265,In_265,In_87);
nand U266 (N_266,In_427,In_266);
nor U267 (N_267,In_436,In_241);
nand U268 (N_268,In_283,In_238);
xnor U269 (N_269,In_39,In_265);
nor U270 (N_270,In_317,In_229);
nand U271 (N_271,In_471,In_255);
nor U272 (N_272,In_141,In_159);
or U273 (N_273,In_213,In_27);
nand U274 (N_274,In_466,In_404);
or U275 (N_275,In_23,In_18);
and U276 (N_276,In_350,In_485);
nor U277 (N_277,In_216,In_234);
nor U278 (N_278,In_327,In_255);
nor U279 (N_279,In_480,In_438);
or U280 (N_280,In_424,In_260);
nor U281 (N_281,In_6,In_81);
nand U282 (N_282,In_381,In_264);
nand U283 (N_283,In_118,In_162);
nand U284 (N_284,In_312,In_146);
or U285 (N_285,In_100,In_13);
and U286 (N_286,In_307,In_404);
nor U287 (N_287,In_281,In_255);
or U288 (N_288,In_337,In_93);
and U289 (N_289,In_0,In_384);
nor U290 (N_290,In_394,In_283);
or U291 (N_291,In_444,In_340);
nand U292 (N_292,In_100,In_9);
nor U293 (N_293,In_451,In_490);
nand U294 (N_294,In_147,In_208);
nand U295 (N_295,In_157,In_10);
and U296 (N_296,In_489,In_46);
nor U297 (N_297,In_66,In_309);
and U298 (N_298,In_178,In_196);
and U299 (N_299,In_438,In_396);
or U300 (N_300,In_58,In_460);
nor U301 (N_301,In_420,In_319);
nor U302 (N_302,In_302,In_300);
nor U303 (N_303,In_330,In_146);
and U304 (N_304,In_314,In_206);
and U305 (N_305,In_361,In_62);
and U306 (N_306,In_419,In_377);
nand U307 (N_307,In_467,In_32);
nand U308 (N_308,In_490,In_75);
nor U309 (N_309,In_410,In_365);
and U310 (N_310,In_477,In_396);
xor U311 (N_311,In_76,In_473);
xnor U312 (N_312,In_282,In_400);
and U313 (N_313,In_295,In_235);
xor U314 (N_314,In_381,In_166);
nand U315 (N_315,In_459,In_59);
xor U316 (N_316,In_116,In_335);
and U317 (N_317,In_432,In_312);
nand U318 (N_318,In_19,In_370);
nand U319 (N_319,In_28,In_145);
nand U320 (N_320,In_55,In_123);
or U321 (N_321,In_102,In_448);
or U322 (N_322,In_279,In_401);
xor U323 (N_323,In_161,In_124);
nor U324 (N_324,In_46,In_467);
nor U325 (N_325,In_53,In_285);
or U326 (N_326,In_202,In_449);
nor U327 (N_327,In_197,In_202);
nand U328 (N_328,In_101,In_320);
nor U329 (N_329,In_312,In_107);
and U330 (N_330,In_19,In_190);
xor U331 (N_331,In_223,In_390);
nor U332 (N_332,In_25,In_241);
and U333 (N_333,In_357,In_255);
and U334 (N_334,In_364,In_94);
or U335 (N_335,In_440,In_285);
nor U336 (N_336,In_42,In_172);
or U337 (N_337,In_199,In_384);
nor U338 (N_338,In_396,In_285);
or U339 (N_339,In_289,In_438);
or U340 (N_340,In_27,In_36);
or U341 (N_341,In_491,In_189);
and U342 (N_342,In_389,In_136);
nor U343 (N_343,In_16,In_85);
and U344 (N_344,In_287,In_246);
or U345 (N_345,In_235,In_366);
nor U346 (N_346,In_36,In_293);
and U347 (N_347,In_481,In_371);
or U348 (N_348,In_430,In_337);
and U349 (N_349,In_134,In_172);
and U350 (N_350,In_383,In_438);
and U351 (N_351,In_496,In_263);
nand U352 (N_352,In_411,In_153);
xor U353 (N_353,In_404,In_108);
and U354 (N_354,In_67,In_21);
nor U355 (N_355,In_169,In_202);
and U356 (N_356,In_317,In_101);
or U357 (N_357,In_100,In_336);
and U358 (N_358,In_464,In_313);
nor U359 (N_359,In_172,In_427);
xnor U360 (N_360,In_115,In_270);
nand U361 (N_361,In_229,In_490);
nand U362 (N_362,In_306,In_86);
or U363 (N_363,In_4,In_179);
and U364 (N_364,In_423,In_90);
xor U365 (N_365,In_227,In_388);
or U366 (N_366,In_211,In_348);
nand U367 (N_367,In_284,In_90);
or U368 (N_368,In_125,In_316);
or U369 (N_369,In_470,In_8);
and U370 (N_370,In_435,In_356);
nand U371 (N_371,In_330,In_457);
nor U372 (N_372,In_418,In_190);
and U373 (N_373,In_110,In_331);
and U374 (N_374,In_391,In_481);
nand U375 (N_375,In_181,In_262);
nand U376 (N_376,In_440,In_161);
and U377 (N_377,In_308,In_80);
nor U378 (N_378,In_78,In_415);
nor U379 (N_379,In_143,In_261);
nand U380 (N_380,In_319,In_466);
or U381 (N_381,In_386,In_394);
nor U382 (N_382,In_243,In_33);
nand U383 (N_383,In_146,In_177);
and U384 (N_384,In_275,In_357);
nand U385 (N_385,In_94,In_196);
or U386 (N_386,In_383,In_58);
nand U387 (N_387,In_381,In_210);
and U388 (N_388,In_232,In_299);
nor U389 (N_389,In_122,In_406);
or U390 (N_390,In_77,In_397);
nand U391 (N_391,In_168,In_118);
xor U392 (N_392,In_238,In_9);
xnor U393 (N_393,In_104,In_18);
nor U394 (N_394,In_125,In_298);
and U395 (N_395,In_316,In_74);
and U396 (N_396,In_25,In_195);
nor U397 (N_397,In_465,In_143);
xor U398 (N_398,In_258,In_15);
nand U399 (N_399,In_86,In_305);
nor U400 (N_400,In_493,In_242);
xor U401 (N_401,In_362,In_464);
nor U402 (N_402,In_14,In_140);
xor U403 (N_403,In_202,In_26);
nand U404 (N_404,In_19,In_475);
and U405 (N_405,In_422,In_155);
nand U406 (N_406,In_463,In_245);
or U407 (N_407,In_82,In_318);
and U408 (N_408,In_117,In_18);
and U409 (N_409,In_257,In_36);
or U410 (N_410,In_125,In_389);
nand U411 (N_411,In_178,In_359);
nand U412 (N_412,In_469,In_302);
and U413 (N_413,In_25,In_330);
nand U414 (N_414,In_465,In_339);
nor U415 (N_415,In_45,In_359);
nor U416 (N_416,In_454,In_105);
nand U417 (N_417,In_388,In_75);
and U418 (N_418,In_468,In_3);
and U419 (N_419,In_308,In_410);
nor U420 (N_420,In_229,In_53);
and U421 (N_421,In_296,In_400);
nor U422 (N_422,In_51,In_84);
or U423 (N_423,In_164,In_15);
or U424 (N_424,In_49,In_220);
and U425 (N_425,In_360,In_70);
xnor U426 (N_426,In_152,In_47);
and U427 (N_427,In_176,In_447);
nor U428 (N_428,In_207,In_452);
xnor U429 (N_429,In_289,In_491);
or U430 (N_430,In_438,In_11);
xor U431 (N_431,In_475,In_105);
nand U432 (N_432,In_164,In_329);
nand U433 (N_433,In_253,In_158);
nand U434 (N_434,In_253,In_237);
nor U435 (N_435,In_7,In_483);
nor U436 (N_436,In_129,In_158);
nand U437 (N_437,In_286,In_148);
or U438 (N_438,In_107,In_0);
and U439 (N_439,In_101,In_228);
nor U440 (N_440,In_130,In_181);
and U441 (N_441,In_19,In_382);
or U442 (N_442,In_69,In_290);
and U443 (N_443,In_404,In_441);
and U444 (N_444,In_358,In_391);
nand U445 (N_445,In_42,In_175);
nor U446 (N_446,In_447,In_246);
or U447 (N_447,In_130,In_432);
and U448 (N_448,In_49,In_254);
nor U449 (N_449,In_428,In_296);
or U450 (N_450,In_461,In_469);
nand U451 (N_451,In_141,In_452);
xnor U452 (N_452,In_120,In_313);
or U453 (N_453,In_396,In_409);
and U454 (N_454,In_287,In_414);
or U455 (N_455,In_309,In_170);
nor U456 (N_456,In_104,In_85);
nand U457 (N_457,In_307,In_443);
nand U458 (N_458,In_246,In_154);
nor U459 (N_459,In_290,In_45);
nand U460 (N_460,In_303,In_363);
nand U461 (N_461,In_27,In_129);
xor U462 (N_462,In_150,In_76);
and U463 (N_463,In_453,In_108);
nor U464 (N_464,In_148,In_197);
and U465 (N_465,In_26,In_151);
and U466 (N_466,In_91,In_193);
or U467 (N_467,In_23,In_298);
xor U468 (N_468,In_269,In_396);
nor U469 (N_469,In_41,In_141);
and U470 (N_470,In_11,In_145);
nand U471 (N_471,In_36,In_316);
xor U472 (N_472,In_405,In_294);
nor U473 (N_473,In_425,In_10);
nor U474 (N_474,In_48,In_304);
and U475 (N_475,In_206,In_128);
nor U476 (N_476,In_484,In_85);
or U477 (N_477,In_54,In_88);
nor U478 (N_478,In_400,In_248);
and U479 (N_479,In_175,In_46);
xnor U480 (N_480,In_259,In_436);
and U481 (N_481,In_207,In_468);
nor U482 (N_482,In_4,In_259);
nand U483 (N_483,In_171,In_26);
nor U484 (N_484,In_130,In_201);
and U485 (N_485,In_100,In_490);
nand U486 (N_486,In_140,In_358);
nor U487 (N_487,In_359,In_39);
or U488 (N_488,In_462,In_119);
and U489 (N_489,In_258,In_316);
nand U490 (N_490,In_252,In_309);
nor U491 (N_491,In_327,In_347);
and U492 (N_492,In_375,In_376);
nor U493 (N_493,In_264,In_472);
nand U494 (N_494,In_194,In_89);
and U495 (N_495,In_204,In_384);
and U496 (N_496,In_407,In_457);
or U497 (N_497,In_279,In_42);
nor U498 (N_498,In_177,In_32);
or U499 (N_499,In_303,In_163);
or U500 (N_500,N_175,N_440);
nor U501 (N_501,N_8,N_321);
nand U502 (N_502,N_100,N_91);
or U503 (N_503,N_383,N_307);
nor U504 (N_504,N_378,N_247);
or U505 (N_505,N_467,N_396);
or U506 (N_506,N_415,N_471);
nor U507 (N_507,N_6,N_355);
or U508 (N_508,N_33,N_296);
and U509 (N_509,N_291,N_164);
nand U510 (N_510,N_490,N_173);
or U511 (N_511,N_216,N_255);
nand U512 (N_512,N_60,N_244);
nand U513 (N_513,N_332,N_391);
nor U514 (N_514,N_305,N_446);
nand U515 (N_515,N_366,N_343);
or U516 (N_516,N_350,N_36);
nand U517 (N_517,N_417,N_299);
or U518 (N_518,N_88,N_419);
nor U519 (N_519,N_309,N_433);
nor U520 (N_520,N_435,N_287);
or U521 (N_521,N_56,N_339);
xor U522 (N_522,N_96,N_207);
and U523 (N_523,N_438,N_317);
nand U524 (N_524,N_420,N_484);
nor U525 (N_525,N_384,N_85);
nand U526 (N_526,N_374,N_155);
and U527 (N_527,N_102,N_354);
nor U528 (N_528,N_267,N_34);
and U529 (N_529,N_140,N_373);
nor U530 (N_530,N_463,N_356);
xnor U531 (N_531,N_313,N_283);
nor U532 (N_532,N_53,N_399);
nor U533 (N_533,N_365,N_495);
or U534 (N_534,N_230,N_144);
and U535 (N_535,N_375,N_326);
nand U536 (N_536,N_342,N_84);
xnor U537 (N_537,N_2,N_16);
nand U538 (N_538,N_231,N_256);
nand U539 (N_539,N_323,N_163);
nand U540 (N_540,N_398,N_178);
nor U541 (N_541,N_217,N_15);
xor U542 (N_542,N_3,N_451);
or U543 (N_543,N_371,N_331);
xnor U544 (N_544,N_314,N_90);
and U545 (N_545,N_409,N_276);
nand U546 (N_546,N_295,N_306);
nor U547 (N_547,N_42,N_477);
and U548 (N_548,N_51,N_360);
and U549 (N_549,N_361,N_447);
nor U550 (N_550,N_482,N_50);
and U551 (N_551,N_270,N_224);
and U552 (N_552,N_193,N_483);
and U553 (N_553,N_236,N_161);
and U554 (N_554,N_441,N_370);
xor U555 (N_555,N_24,N_392);
and U556 (N_556,N_376,N_214);
nand U557 (N_557,N_382,N_279);
and U558 (N_558,N_98,N_290);
or U559 (N_559,N_150,N_176);
nor U560 (N_560,N_64,N_167);
xor U561 (N_561,N_40,N_165);
or U562 (N_562,N_459,N_262);
nand U563 (N_563,N_118,N_179);
nor U564 (N_564,N_413,N_240);
and U565 (N_565,N_128,N_258);
xor U566 (N_566,N_10,N_488);
and U567 (N_567,N_431,N_257);
nand U568 (N_568,N_474,N_103);
or U569 (N_569,N_449,N_122);
or U570 (N_570,N_125,N_78);
nor U571 (N_571,N_145,N_266);
nor U572 (N_572,N_39,N_147);
and U573 (N_573,N_303,N_292);
nand U574 (N_574,N_499,N_448);
or U575 (N_575,N_212,N_472);
or U576 (N_576,N_218,N_201);
and U577 (N_577,N_221,N_202);
and U578 (N_578,N_62,N_83);
nand U579 (N_579,N_453,N_369);
and U580 (N_580,N_460,N_75);
nor U581 (N_581,N_286,N_9);
nand U582 (N_582,N_428,N_301);
nand U583 (N_583,N_473,N_385);
or U584 (N_584,N_208,N_388);
nand U585 (N_585,N_228,N_133);
and U586 (N_586,N_74,N_4);
nand U587 (N_587,N_190,N_338);
or U588 (N_588,N_426,N_436);
and U589 (N_589,N_277,N_89);
nor U590 (N_590,N_406,N_340);
and U591 (N_591,N_7,N_328);
and U592 (N_592,N_337,N_182);
nand U593 (N_593,N_159,N_5);
and U594 (N_594,N_67,N_93);
or U595 (N_595,N_14,N_380);
or U596 (N_596,N_27,N_353);
or U597 (N_597,N_11,N_273);
nand U598 (N_598,N_492,N_79);
or U599 (N_599,N_12,N_352);
nand U600 (N_600,N_403,N_478);
nand U601 (N_601,N_174,N_113);
nand U602 (N_602,N_430,N_184);
nand U603 (N_603,N_408,N_45);
nand U604 (N_604,N_17,N_181);
nor U605 (N_605,N_18,N_99);
nand U606 (N_606,N_135,N_112);
xnor U607 (N_607,N_367,N_55);
nand U608 (N_608,N_357,N_48);
nor U609 (N_609,N_358,N_316);
nand U610 (N_610,N_129,N_49);
nand U611 (N_611,N_44,N_249);
nor U612 (N_612,N_177,N_297);
or U613 (N_613,N_327,N_116);
and U614 (N_614,N_170,N_405);
or U615 (N_615,N_82,N_466);
xor U616 (N_616,N_423,N_425);
and U617 (N_617,N_481,N_268);
and U618 (N_618,N_105,N_333);
or U619 (N_619,N_265,N_136);
nand U620 (N_620,N_400,N_127);
nand U621 (N_621,N_274,N_464);
nand U622 (N_622,N_427,N_43);
nand U623 (N_623,N_293,N_227);
xor U624 (N_624,N_234,N_194);
or U625 (N_625,N_143,N_66);
and U626 (N_626,N_35,N_476);
nand U627 (N_627,N_318,N_381);
or U628 (N_628,N_245,N_465);
nor U629 (N_629,N_95,N_344);
or U630 (N_630,N_124,N_117);
or U631 (N_631,N_242,N_37);
and U632 (N_632,N_386,N_456);
or U633 (N_633,N_412,N_195);
and U634 (N_634,N_298,N_123);
and U635 (N_635,N_197,N_393);
nor U636 (N_636,N_364,N_191);
nor U637 (N_637,N_68,N_457);
nor U638 (N_638,N_437,N_302);
nor U639 (N_639,N_86,N_304);
nand U640 (N_640,N_183,N_189);
and U641 (N_641,N_402,N_429);
nand U642 (N_642,N_454,N_58);
xnor U643 (N_643,N_41,N_225);
or U644 (N_644,N_20,N_215);
xnor U645 (N_645,N_379,N_213);
or U646 (N_646,N_424,N_219);
or U647 (N_647,N_180,N_468);
nor U648 (N_648,N_196,N_233);
nor U649 (N_649,N_325,N_237);
nor U650 (N_650,N_315,N_311);
xnor U651 (N_651,N_169,N_156);
or U652 (N_652,N_132,N_461);
nor U653 (N_653,N_434,N_131);
nor U654 (N_654,N_226,N_71);
nor U655 (N_655,N_280,N_312);
or U656 (N_656,N_198,N_404);
xnor U657 (N_657,N_54,N_110);
or U658 (N_658,N_80,N_487);
nand U659 (N_659,N_469,N_25);
xor U660 (N_660,N_229,N_341);
and U661 (N_661,N_168,N_153);
nor U662 (N_662,N_101,N_232);
nor U663 (N_663,N_395,N_70);
and U664 (N_664,N_259,N_61);
and U665 (N_665,N_107,N_308);
and U666 (N_666,N_445,N_222);
or U667 (N_667,N_322,N_13);
and U668 (N_668,N_26,N_152);
nor U669 (N_669,N_238,N_462);
and U670 (N_670,N_204,N_498);
xnor U671 (N_671,N_241,N_157);
nor U672 (N_672,N_401,N_119);
or U673 (N_673,N_77,N_251);
nand U674 (N_674,N_452,N_32);
nor U675 (N_675,N_418,N_65);
nand U676 (N_676,N_23,N_319);
and U677 (N_677,N_188,N_264);
nor U678 (N_678,N_372,N_114);
or U679 (N_679,N_348,N_149);
xnor U680 (N_680,N_92,N_211);
and U681 (N_681,N_496,N_281);
and U682 (N_682,N_480,N_120);
and U683 (N_683,N_63,N_444);
or U684 (N_684,N_28,N_59);
nand U685 (N_685,N_414,N_29);
or U686 (N_686,N_253,N_141);
or U687 (N_687,N_108,N_151);
nor U688 (N_688,N_130,N_416);
xnor U689 (N_689,N_250,N_111);
or U690 (N_690,N_421,N_310);
nor U691 (N_691,N_72,N_320);
and U692 (N_692,N_21,N_494);
nor U693 (N_693,N_458,N_285);
nand U694 (N_694,N_47,N_115);
and U695 (N_695,N_289,N_200);
nor U696 (N_696,N_187,N_346);
nand U697 (N_697,N_261,N_397);
nand U698 (N_698,N_235,N_260);
nand U699 (N_699,N_347,N_186);
nor U700 (N_700,N_166,N_387);
and U701 (N_701,N_272,N_87);
and U702 (N_702,N_220,N_205);
nor U703 (N_703,N_368,N_223);
nand U704 (N_704,N_335,N_104);
nand U705 (N_705,N_109,N_172);
nand U706 (N_706,N_450,N_329);
nor U707 (N_707,N_81,N_324);
nor U708 (N_708,N_46,N_278);
nor U709 (N_709,N_410,N_282);
and U710 (N_710,N_148,N_263);
nand U711 (N_711,N_254,N_171);
nand U712 (N_712,N_390,N_439);
nor U713 (N_713,N_271,N_432);
nor U714 (N_714,N_209,N_19);
nor U715 (N_715,N_69,N_407);
or U716 (N_716,N_411,N_294);
or U717 (N_717,N_284,N_106);
and U718 (N_718,N_345,N_486);
nand U719 (N_719,N_210,N_121);
nand U720 (N_720,N_134,N_349);
nand U721 (N_721,N_475,N_73);
nor U722 (N_722,N_351,N_442);
and U723 (N_723,N_160,N_162);
or U724 (N_724,N_192,N_239);
nor U725 (N_725,N_359,N_206);
nand U726 (N_726,N_422,N_455);
nor U727 (N_727,N_0,N_269);
or U728 (N_728,N_76,N_363);
xnor U729 (N_729,N_146,N_497);
and U730 (N_730,N_491,N_362);
or U731 (N_731,N_94,N_489);
and U732 (N_732,N_185,N_139);
and U733 (N_733,N_377,N_38);
nor U734 (N_734,N_31,N_288);
nand U735 (N_735,N_1,N_330);
and U736 (N_736,N_275,N_252);
and U737 (N_737,N_300,N_479);
nor U738 (N_738,N_142,N_389);
nand U739 (N_739,N_154,N_30);
xor U740 (N_740,N_336,N_203);
nor U741 (N_741,N_158,N_248);
nor U742 (N_742,N_243,N_126);
or U743 (N_743,N_394,N_246);
nor U744 (N_744,N_199,N_485);
nor U745 (N_745,N_138,N_57);
and U746 (N_746,N_470,N_97);
nand U747 (N_747,N_137,N_52);
and U748 (N_748,N_443,N_22);
nor U749 (N_749,N_334,N_493);
nor U750 (N_750,N_36,N_485);
nor U751 (N_751,N_395,N_386);
and U752 (N_752,N_73,N_131);
or U753 (N_753,N_40,N_402);
nand U754 (N_754,N_399,N_130);
nor U755 (N_755,N_283,N_422);
or U756 (N_756,N_482,N_447);
and U757 (N_757,N_307,N_314);
or U758 (N_758,N_455,N_298);
and U759 (N_759,N_335,N_123);
nor U760 (N_760,N_295,N_386);
or U761 (N_761,N_435,N_32);
nand U762 (N_762,N_265,N_357);
or U763 (N_763,N_102,N_216);
nor U764 (N_764,N_417,N_435);
nor U765 (N_765,N_309,N_365);
and U766 (N_766,N_185,N_173);
xor U767 (N_767,N_251,N_274);
nand U768 (N_768,N_455,N_123);
and U769 (N_769,N_300,N_278);
nand U770 (N_770,N_395,N_287);
nor U771 (N_771,N_15,N_42);
nor U772 (N_772,N_124,N_495);
or U773 (N_773,N_214,N_106);
nor U774 (N_774,N_357,N_87);
xor U775 (N_775,N_471,N_14);
or U776 (N_776,N_457,N_156);
xor U777 (N_777,N_339,N_173);
nand U778 (N_778,N_5,N_17);
xnor U779 (N_779,N_450,N_226);
nor U780 (N_780,N_0,N_249);
or U781 (N_781,N_125,N_334);
nor U782 (N_782,N_215,N_9);
and U783 (N_783,N_127,N_185);
nand U784 (N_784,N_294,N_192);
nor U785 (N_785,N_180,N_266);
nor U786 (N_786,N_344,N_293);
and U787 (N_787,N_374,N_441);
nand U788 (N_788,N_287,N_154);
or U789 (N_789,N_126,N_223);
nand U790 (N_790,N_461,N_21);
or U791 (N_791,N_453,N_8);
nor U792 (N_792,N_173,N_144);
and U793 (N_793,N_400,N_48);
nand U794 (N_794,N_123,N_194);
or U795 (N_795,N_34,N_36);
nor U796 (N_796,N_468,N_241);
nor U797 (N_797,N_318,N_494);
and U798 (N_798,N_380,N_142);
xnor U799 (N_799,N_294,N_353);
nand U800 (N_800,N_310,N_369);
nor U801 (N_801,N_22,N_111);
or U802 (N_802,N_185,N_356);
or U803 (N_803,N_332,N_357);
xor U804 (N_804,N_379,N_407);
and U805 (N_805,N_223,N_290);
and U806 (N_806,N_64,N_114);
and U807 (N_807,N_464,N_185);
nor U808 (N_808,N_223,N_141);
nand U809 (N_809,N_460,N_232);
xor U810 (N_810,N_37,N_358);
and U811 (N_811,N_406,N_338);
nand U812 (N_812,N_278,N_153);
nor U813 (N_813,N_272,N_109);
and U814 (N_814,N_427,N_276);
nand U815 (N_815,N_395,N_390);
nand U816 (N_816,N_296,N_108);
xnor U817 (N_817,N_53,N_105);
nor U818 (N_818,N_4,N_139);
and U819 (N_819,N_339,N_343);
xnor U820 (N_820,N_479,N_401);
nor U821 (N_821,N_277,N_428);
or U822 (N_822,N_332,N_75);
xnor U823 (N_823,N_368,N_280);
nand U824 (N_824,N_144,N_486);
nor U825 (N_825,N_38,N_420);
and U826 (N_826,N_201,N_376);
xnor U827 (N_827,N_231,N_485);
nor U828 (N_828,N_387,N_57);
or U829 (N_829,N_127,N_274);
or U830 (N_830,N_434,N_304);
or U831 (N_831,N_385,N_175);
nand U832 (N_832,N_32,N_346);
xnor U833 (N_833,N_126,N_115);
or U834 (N_834,N_262,N_60);
nor U835 (N_835,N_283,N_292);
nand U836 (N_836,N_360,N_180);
nand U837 (N_837,N_37,N_350);
and U838 (N_838,N_99,N_374);
or U839 (N_839,N_227,N_487);
and U840 (N_840,N_260,N_445);
and U841 (N_841,N_352,N_355);
or U842 (N_842,N_432,N_464);
nor U843 (N_843,N_486,N_70);
and U844 (N_844,N_48,N_298);
nor U845 (N_845,N_335,N_331);
or U846 (N_846,N_199,N_362);
nand U847 (N_847,N_50,N_460);
nand U848 (N_848,N_174,N_124);
nor U849 (N_849,N_3,N_113);
nor U850 (N_850,N_138,N_167);
or U851 (N_851,N_461,N_369);
nor U852 (N_852,N_222,N_225);
nor U853 (N_853,N_128,N_479);
or U854 (N_854,N_272,N_40);
and U855 (N_855,N_22,N_187);
nor U856 (N_856,N_350,N_184);
nor U857 (N_857,N_288,N_41);
and U858 (N_858,N_176,N_311);
and U859 (N_859,N_434,N_471);
nor U860 (N_860,N_493,N_207);
or U861 (N_861,N_321,N_104);
xnor U862 (N_862,N_230,N_177);
nand U863 (N_863,N_37,N_484);
nor U864 (N_864,N_467,N_488);
and U865 (N_865,N_321,N_33);
nor U866 (N_866,N_387,N_161);
or U867 (N_867,N_104,N_460);
or U868 (N_868,N_436,N_200);
nor U869 (N_869,N_182,N_197);
or U870 (N_870,N_392,N_297);
or U871 (N_871,N_112,N_200);
and U872 (N_872,N_492,N_290);
nor U873 (N_873,N_230,N_184);
nand U874 (N_874,N_374,N_49);
xnor U875 (N_875,N_330,N_370);
or U876 (N_876,N_158,N_342);
nor U877 (N_877,N_214,N_322);
or U878 (N_878,N_96,N_111);
nand U879 (N_879,N_444,N_217);
nand U880 (N_880,N_467,N_398);
and U881 (N_881,N_183,N_465);
and U882 (N_882,N_119,N_104);
nand U883 (N_883,N_436,N_286);
or U884 (N_884,N_311,N_154);
or U885 (N_885,N_383,N_380);
nand U886 (N_886,N_309,N_190);
xnor U887 (N_887,N_232,N_266);
or U888 (N_888,N_267,N_363);
or U889 (N_889,N_198,N_170);
nand U890 (N_890,N_317,N_202);
nor U891 (N_891,N_365,N_156);
nand U892 (N_892,N_38,N_150);
nand U893 (N_893,N_276,N_439);
or U894 (N_894,N_43,N_238);
and U895 (N_895,N_185,N_388);
nand U896 (N_896,N_447,N_243);
nand U897 (N_897,N_209,N_266);
xor U898 (N_898,N_432,N_151);
and U899 (N_899,N_132,N_372);
and U900 (N_900,N_394,N_216);
nand U901 (N_901,N_324,N_327);
nor U902 (N_902,N_123,N_457);
or U903 (N_903,N_170,N_444);
and U904 (N_904,N_401,N_382);
nand U905 (N_905,N_303,N_286);
or U906 (N_906,N_474,N_300);
xor U907 (N_907,N_391,N_62);
and U908 (N_908,N_178,N_93);
and U909 (N_909,N_303,N_144);
or U910 (N_910,N_2,N_136);
and U911 (N_911,N_355,N_420);
nor U912 (N_912,N_473,N_376);
and U913 (N_913,N_5,N_237);
nand U914 (N_914,N_345,N_53);
or U915 (N_915,N_54,N_460);
or U916 (N_916,N_228,N_306);
nand U917 (N_917,N_375,N_208);
nor U918 (N_918,N_49,N_236);
nor U919 (N_919,N_298,N_492);
or U920 (N_920,N_276,N_152);
and U921 (N_921,N_346,N_40);
and U922 (N_922,N_405,N_148);
nand U923 (N_923,N_488,N_103);
nor U924 (N_924,N_131,N_404);
nor U925 (N_925,N_157,N_349);
nand U926 (N_926,N_253,N_38);
nor U927 (N_927,N_388,N_456);
nor U928 (N_928,N_385,N_294);
and U929 (N_929,N_168,N_444);
and U930 (N_930,N_473,N_440);
xor U931 (N_931,N_185,N_408);
or U932 (N_932,N_279,N_125);
or U933 (N_933,N_237,N_335);
or U934 (N_934,N_315,N_182);
nor U935 (N_935,N_144,N_13);
and U936 (N_936,N_412,N_68);
or U937 (N_937,N_103,N_247);
or U938 (N_938,N_200,N_333);
nor U939 (N_939,N_289,N_379);
nand U940 (N_940,N_67,N_417);
nand U941 (N_941,N_268,N_311);
nor U942 (N_942,N_97,N_111);
and U943 (N_943,N_41,N_240);
and U944 (N_944,N_75,N_95);
or U945 (N_945,N_497,N_63);
nor U946 (N_946,N_136,N_311);
nand U947 (N_947,N_12,N_231);
nor U948 (N_948,N_24,N_77);
nor U949 (N_949,N_213,N_491);
or U950 (N_950,N_147,N_216);
xnor U951 (N_951,N_131,N_132);
and U952 (N_952,N_9,N_349);
and U953 (N_953,N_99,N_140);
and U954 (N_954,N_444,N_329);
or U955 (N_955,N_407,N_170);
or U956 (N_956,N_206,N_337);
and U957 (N_957,N_296,N_345);
nor U958 (N_958,N_80,N_119);
or U959 (N_959,N_230,N_335);
nor U960 (N_960,N_322,N_308);
nor U961 (N_961,N_196,N_170);
or U962 (N_962,N_490,N_200);
nand U963 (N_963,N_499,N_462);
nand U964 (N_964,N_350,N_153);
or U965 (N_965,N_353,N_414);
nand U966 (N_966,N_427,N_65);
and U967 (N_967,N_159,N_400);
nand U968 (N_968,N_146,N_339);
nor U969 (N_969,N_52,N_320);
xor U970 (N_970,N_470,N_193);
or U971 (N_971,N_334,N_342);
or U972 (N_972,N_79,N_288);
and U973 (N_973,N_452,N_293);
and U974 (N_974,N_163,N_169);
or U975 (N_975,N_310,N_380);
nand U976 (N_976,N_38,N_250);
and U977 (N_977,N_394,N_401);
and U978 (N_978,N_361,N_39);
nor U979 (N_979,N_13,N_153);
nor U980 (N_980,N_468,N_253);
nand U981 (N_981,N_466,N_231);
and U982 (N_982,N_419,N_301);
or U983 (N_983,N_302,N_340);
or U984 (N_984,N_368,N_398);
nand U985 (N_985,N_366,N_21);
nand U986 (N_986,N_28,N_166);
nor U987 (N_987,N_277,N_249);
and U988 (N_988,N_469,N_74);
nand U989 (N_989,N_6,N_398);
nor U990 (N_990,N_85,N_359);
and U991 (N_991,N_388,N_273);
xnor U992 (N_992,N_328,N_313);
xor U993 (N_993,N_151,N_435);
xor U994 (N_994,N_301,N_283);
nand U995 (N_995,N_380,N_185);
xnor U996 (N_996,N_202,N_48);
nand U997 (N_997,N_252,N_40);
nor U998 (N_998,N_128,N_153);
nand U999 (N_999,N_64,N_344);
nand U1000 (N_1000,N_712,N_709);
nand U1001 (N_1001,N_989,N_581);
and U1002 (N_1002,N_908,N_661);
xor U1003 (N_1003,N_845,N_784);
and U1004 (N_1004,N_572,N_602);
nand U1005 (N_1005,N_974,N_592);
nand U1006 (N_1006,N_800,N_758);
nor U1007 (N_1007,N_711,N_659);
nand U1008 (N_1008,N_651,N_997);
xor U1009 (N_1009,N_623,N_621);
nor U1010 (N_1010,N_892,N_829);
and U1011 (N_1011,N_780,N_669);
or U1012 (N_1012,N_769,N_937);
nor U1013 (N_1013,N_604,N_801);
nand U1014 (N_1014,N_827,N_869);
xnor U1015 (N_1015,N_512,N_517);
nor U1016 (N_1016,N_603,N_864);
nand U1017 (N_1017,N_819,N_932);
xor U1018 (N_1018,N_676,N_835);
nor U1019 (N_1019,N_957,N_927);
nand U1020 (N_1020,N_524,N_644);
or U1021 (N_1021,N_948,N_983);
or U1022 (N_1022,N_698,N_949);
or U1023 (N_1023,N_956,N_799);
or U1024 (N_1024,N_615,N_831);
or U1025 (N_1025,N_551,N_971);
nand U1026 (N_1026,N_936,N_612);
xnor U1027 (N_1027,N_527,N_980);
or U1028 (N_1028,N_975,N_917);
nor U1029 (N_1029,N_693,N_678);
or U1030 (N_1030,N_586,N_697);
nand U1031 (N_1031,N_533,N_664);
nand U1032 (N_1032,N_738,N_787);
nor U1033 (N_1033,N_768,N_900);
nor U1034 (N_1034,N_998,N_885);
or U1035 (N_1035,N_577,N_951);
or U1036 (N_1036,N_926,N_794);
nor U1037 (N_1037,N_741,N_935);
or U1038 (N_1038,N_934,N_877);
nand U1039 (N_1039,N_876,N_857);
nand U1040 (N_1040,N_783,N_914);
or U1041 (N_1041,N_773,N_694);
and U1042 (N_1042,N_595,N_597);
nor U1043 (N_1043,N_940,N_541);
nor U1044 (N_1044,N_969,N_703);
or U1045 (N_1045,N_858,N_643);
or U1046 (N_1046,N_558,N_538);
nand U1047 (N_1047,N_728,N_886);
nand U1048 (N_1048,N_795,N_734);
xnor U1049 (N_1049,N_744,N_655);
and U1050 (N_1050,N_988,N_704);
or U1051 (N_1051,N_880,N_843);
xnor U1052 (N_1052,N_707,N_915);
nor U1053 (N_1053,N_619,N_579);
or U1054 (N_1054,N_921,N_566);
xor U1055 (N_1055,N_952,N_665);
nand U1056 (N_1056,N_777,N_640);
or U1057 (N_1057,N_739,N_755);
nor U1058 (N_1058,N_950,N_805);
and U1059 (N_1059,N_673,N_772);
or U1060 (N_1060,N_854,N_923);
or U1061 (N_1061,N_532,N_677);
nor U1062 (N_1062,N_991,N_830);
and U1063 (N_1063,N_686,N_930);
nand U1064 (N_1064,N_646,N_594);
and U1065 (N_1065,N_925,N_682);
nand U1066 (N_1066,N_961,N_587);
or U1067 (N_1067,N_607,N_641);
or U1068 (N_1068,N_993,N_903);
or U1069 (N_1069,N_902,N_836);
or U1070 (N_1070,N_723,N_815);
or U1071 (N_1071,N_844,N_508);
and U1072 (N_1072,N_807,N_504);
nand U1073 (N_1073,N_513,N_510);
nor U1074 (N_1074,N_867,N_720);
nand U1075 (N_1075,N_570,N_833);
nor U1076 (N_1076,N_992,N_946);
or U1077 (N_1077,N_618,N_786);
and U1078 (N_1078,N_528,N_825);
nor U1079 (N_1079,N_630,N_683);
or U1080 (N_1080,N_802,N_729);
or U1081 (N_1081,N_708,N_884);
and U1082 (N_1082,N_632,N_702);
xor U1083 (N_1083,N_576,N_574);
nand U1084 (N_1084,N_751,N_839);
or U1085 (N_1085,N_945,N_668);
or U1086 (N_1086,N_521,N_547);
nor U1087 (N_1087,N_593,N_943);
and U1088 (N_1088,N_778,N_753);
nor U1089 (N_1089,N_766,N_746);
nor U1090 (N_1090,N_929,N_789);
or U1091 (N_1091,N_690,N_649);
nor U1092 (N_1092,N_564,N_580);
or U1093 (N_1093,N_722,N_847);
nand U1094 (N_1094,N_964,N_660);
or U1095 (N_1095,N_796,N_792);
or U1096 (N_1096,N_529,N_743);
and U1097 (N_1097,N_507,N_501);
nand U1098 (N_1098,N_614,N_674);
or U1099 (N_1099,N_617,N_774);
nor U1100 (N_1100,N_911,N_598);
nor U1101 (N_1101,N_905,N_977);
xor U1102 (N_1102,N_539,N_613);
nor U1103 (N_1103,N_631,N_544);
nand U1104 (N_1104,N_912,N_573);
nand U1105 (N_1105,N_662,N_764);
nor U1106 (N_1106,N_752,N_653);
and U1107 (N_1107,N_756,N_578);
nor U1108 (N_1108,N_899,N_810);
xnor U1109 (N_1109,N_986,N_994);
and U1110 (N_1110,N_667,N_721);
or U1111 (N_1111,N_939,N_840);
or U1112 (N_1112,N_565,N_822);
or U1113 (N_1113,N_901,N_575);
nand U1114 (N_1114,N_505,N_629);
xnor U1115 (N_1115,N_522,N_561);
nand U1116 (N_1116,N_771,N_898);
xnor U1117 (N_1117,N_984,N_523);
nand U1118 (N_1118,N_588,N_812);
xnor U1119 (N_1119,N_941,N_955);
and U1120 (N_1120,N_890,N_556);
and U1121 (N_1121,N_832,N_973);
or U1122 (N_1122,N_874,N_979);
and U1123 (N_1123,N_928,N_972);
or U1124 (N_1124,N_820,N_685);
and U1125 (N_1125,N_608,N_616);
nand U1126 (N_1126,N_705,N_782);
xor U1127 (N_1127,N_967,N_627);
nand U1128 (N_1128,N_762,N_873);
nor U1129 (N_1129,N_846,N_828);
nand U1130 (N_1130,N_944,N_866);
nand U1131 (N_1131,N_695,N_775);
and U1132 (N_1132,N_882,N_959);
nand U1133 (N_1133,N_824,N_654);
or U1134 (N_1134,N_642,N_788);
nand U1135 (N_1135,N_813,N_860);
nor U1136 (N_1136,N_808,N_850);
nor U1137 (N_1137,N_763,N_879);
nor U1138 (N_1138,N_725,N_871);
nor U1139 (N_1139,N_680,N_715);
or U1140 (N_1140,N_981,N_918);
nor U1141 (N_1141,N_757,N_534);
nor U1142 (N_1142,N_851,N_691);
nor U1143 (N_1143,N_634,N_582);
or U1144 (N_1144,N_713,N_913);
xnor U1145 (N_1145,N_804,N_591);
xor U1146 (N_1146,N_571,N_875);
and U1147 (N_1147,N_987,N_954);
and U1148 (N_1148,N_726,N_518);
xnor U1149 (N_1149,N_754,N_790);
and U1150 (N_1150,N_520,N_910);
nand U1151 (N_1151,N_761,N_656);
nor U1152 (N_1152,N_963,N_638);
and U1153 (N_1153,N_759,N_748);
nand U1154 (N_1154,N_688,N_624);
and U1155 (N_1155,N_681,N_823);
nor U1156 (N_1156,N_793,N_610);
and U1157 (N_1157,N_826,N_855);
and U1158 (N_1158,N_803,N_600);
nand U1159 (N_1159,N_596,N_982);
nand U1160 (N_1160,N_530,N_540);
nand U1161 (N_1161,N_904,N_601);
nand U1162 (N_1162,N_809,N_853);
or U1163 (N_1163,N_666,N_732);
nor U1164 (N_1164,N_920,N_689);
nand U1165 (N_1165,N_567,N_554);
nand U1166 (N_1166,N_816,N_922);
or U1167 (N_1167,N_675,N_938);
or U1168 (N_1168,N_919,N_609);
nand U1169 (N_1169,N_657,N_933);
and U1170 (N_1170,N_650,N_856);
nand U1171 (N_1171,N_947,N_837);
or U1172 (N_1172,N_692,N_500);
nand U1173 (N_1173,N_747,N_628);
nand U1174 (N_1174,N_647,N_714);
or U1175 (N_1175,N_589,N_557);
nor U1176 (N_1176,N_701,N_716);
xnor U1177 (N_1177,N_907,N_549);
and U1178 (N_1178,N_881,N_909);
or U1179 (N_1179,N_924,N_555);
and U1180 (N_1180,N_516,N_559);
nand U1181 (N_1181,N_639,N_965);
and U1182 (N_1182,N_526,N_785);
nand U1183 (N_1183,N_821,N_684);
or U1184 (N_1184,N_888,N_672);
nand U1185 (N_1185,N_878,N_611);
and U1186 (N_1186,N_506,N_776);
and U1187 (N_1187,N_736,N_637);
xor U1188 (N_1188,N_671,N_742);
and U1189 (N_1189,N_896,N_503);
nor U1190 (N_1190,N_542,N_966);
nor U1191 (N_1191,N_731,N_553);
nand U1192 (N_1192,N_737,N_718);
or U1193 (N_1193,N_842,N_658);
nand U1194 (N_1194,N_550,N_765);
nor U1195 (N_1195,N_730,N_519);
nand U1196 (N_1196,N_648,N_872);
and U1197 (N_1197,N_625,N_895);
or U1198 (N_1198,N_968,N_568);
or U1199 (N_1199,N_841,N_515);
xor U1200 (N_1200,N_537,N_605);
or U1201 (N_1201,N_750,N_599);
nand U1202 (N_1202,N_863,N_569);
and U1203 (N_1203,N_717,N_770);
and U1204 (N_1204,N_687,N_985);
nor U1205 (N_1205,N_953,N_767);
nor U1206 (N_1206,N_719,N_699);
and U1207 (N_1207,N_727,N_663);
nand U1208 (N_1208,N_868,N_891);
or U1209 (N_1209,N_887,N_906);
nand U1210 (N_1210,N_990,N_536);
and U1211 (N_1211,N_622,N_700);
or U1212 (N_1212,N_514,N_781);
nor U1213 (N_1213,N_848,N_806);
nand U1214 (N_1214,N_552,N_916);
or U1215 (N_1215,N_735,N_779);
nor U1216 (N_1216,N_635,N_583);
or U1217 (N_1217,N_560,N_897);
nand U1218 (N_1218,N_710,N_798);
nand U1219 (N_1219,N_811,N_733);
nor U1220 (N_1220,N_760,N_861);
or U1221 (N_1221,N_724,N_942);
and U1222 (N_1222,N_652,N_525);
and U1223 (N_1223,N_562,N_585);
nand U1224 (N_1224,N_633,N_745);
nor U1225 (N_1225,N_511,N_535);
and U1226 (N_1226,N_817,N_636);
xnor U1227 (N_1227,N_889,N_706);
nand U1228 (N_1228,N_970,N_584);
and U1229 (N_1229,N_546,N_696);
or U1230 (N_1230,N_999,N_931);
nand U1231 (N_1231,N_543,N_670);
nor U1232 (N_1232,N_849,N_894);
or U1233 (N_1233,N_740,N_797);
nand U1234 (N_1234,N_996,N_814);
or U1235 (N_1235,N_995,N_834);
or U1236 (N_1236,N_852,N_978);
xnor U1237 (N_1237,N_645,N_563);
and U1238 (N_1238,N_626,N_976);
nand U1239 (N_1239,N_862,N_590);
nor U1240 (N_1240,N_679,N_893);
xor U1241 (N_1241,N_883,N_606);
xnor U1242 (N_1242,N_749,N_545);
or U1243 (N_1243,N_960,N_548);
nor U1244 (N_1244,N_818,N_958);
or U1245 (N_1245,N_531,N_859);
xnor U1246 (N_1246,N_509,N_962);
nor U1247 (N_1247,N_870,N_620);
xor U1248 (N_1248,N_865,N_838);
and U1249 (N_1249,N_502,N_791);
nor U1250 (N_1250,N_711,N_974);
nor U1251 (N_1251,N_894,N_848);
or U1252 (N_1252,N_888,N_815);
nand U1253 (N_1253,N_666,N_849);
nand U1254 (N_1254,N_557,N_754);
xor U1255 (N_1255,N_661,N_760);
or U1256 (N_1256,N_952,N_654);
xor U1257 (N_1257,N_706,N_664);
nor U1258 (N_1258,N_652,N_906);
nand U1259 (N_1259,N_813,N_537);
nand U1260 (N_1260,N_858,N_889);
and U1261 (N_1261,N_704,N_686);
nor U1262 (N_1262,N_727,N_762);
and U1263 (N_1263,N_593,N_578);
or U1264 (N_1264,N_988,N_729);
nor U1265 (N_1265,N_755,N_965);
and U1266 (N_1266,N_643,N_671);
and U1267 (N_1267,N_973,N_588);
nand U1268 (N_1268,N_942,N_989);
or U1269 (N_1269,N_681,N_568);
nand U1270 (N_1270,N_973,N_993);
or U1271 (N_1271,N_683,N_809);
nor U1272 (N_1272,N_763,N_752);
and U1273 (N_1273,N_599,N_529);
or U1274 (N_1274,N_837,N_982);
or U1275 (N_1275,N_973,N_623);
nand U1276 (N_1276,N_682,N_647);
xor U1277 (N_1277,N_731,N_629);
xnor U1278 (N_1278,N_912,N_872);
nand U1279 (N_1279,N_661,N_868);
and U1280 (N_1280,N_841,N_845);
or U1281 (N_1281,N_783,N_888);
xor U1282 (N_1282,N_663,N_808);
nor U1283 (N_1283,N_887,N_570);
nor U1284 (N_1284,N_927,N_751);
and U1285 (N_1285,N_620,N_864);
xor U1286 (N_1286,N_681,N_686);
and U1287 (N_1287,N_865,N_517);
and U1288 (N_1288,N_813,N_615);
and U1289 (N_1289,N_507,N_981);
or U1290 (N_1290,N_584,N_928);
nand U1291 (N_1291,N_838,N_648);
nor U1292 (N_1292,N_917,N_772);
and U1293 (N_1293,N_749,N_616);
or U1294 (N_1294,N_642,N_845);
and U1295 (N_1295,N_831,N_718);
or U1296 (N_1296,N_725,N_798);
nor U1297 (N_1297,N_986,N_705);
xnor U1298 (N_1298,N_632,N_737);
nor U1299 (N_1299,N_625,N_628);
xor U1300 (N_1300,N_743,N_922);
and U1301 (N_1301,N_584,N_739);
or U1302 (N_1302,N_759,N_585);
nor U1303 (N_1303,N_656,N_978);
and U1304 (N_1304,N_744,N_794);
nor U1305 (N_1305,N_585,N_909);
and U1306 (N_1306,N_569,N_571);
nand U1307 (N_1307,N_752,N_655);
nand U1308 (N_1308,N_867,N_828);
nand U1309 (N_1309,N_950,N_920);
nor U1310 (N_1310,N_698,N_969);
nand U1311 (N_1311,N_756,N_823);
or U1312 (N_1312,N_837,N_925);
nor U1313 (N_1313,N_835,N_953);
nor U1314 (N_1314,N_641,N_521);
nor U1315 (N_1315,N_938,N_702);
or U1316 (N_1316,N_909,N_658);
nand U1317 (N_1317,N_548,N_729);
nor U1318 (N_1318,N_912,N_859);
nor U1319 (N_1319,N_529,N_898);
nand U1320 (N_1320,N_958,N_952);
nor U1321 (N_1321,N_633,N_821);
xnor U1322 (N_1322,N_584,N_874);
nand U1323 (N_1323,N_599,N_545);
or U1324 (N_1324,N_754,N_623);
and U1325 (N_1325,N_557,N_652);
nor U1326 (N_1326,N_683,N_936);
and U1327 (N_1327,N_780,N_818);
nor U1328 (N_1328,N_682,N_801);
and U1329 (N_1329,N_742,N_980);
nor U1330 (N_1330,N_974,N_980);
or U1331 (N_1331,N_750,N_882);
or U1332 (N_1332,N_904,N_740);
or U1333 (N_1333,N_710,N_675);
nor U1334 (N_1334,N_693,N_674);
or U1335 (N_1335,N_998,N_688);
nand U1336 (N_1336,N_776,N_553);
or U1337 (N_1337,N_913,N_843);
nand U1338 (N_1338,N_615,N_968);
nand U1339 (N_1339,N_659,N_848);
nand U1340 (N_1340,N_723,N_525);
nor U1341 (N_1341,N_646,N_923);
nand U1342 (N_1342,N_837,N_866);
or U1343 (N_1343,N_869,N_835);
nor U1344 (N_1344,N_926,N_596);
or U1345 (N_1345,N_740,N_672);
nand U1346 (N_1346,N_974,N_843);
or U1347 (N_1347,N_706,N_847);
nor U1348 (N_1348,N_615,N_850);
or U1349 (N_1349,N_949,N_982);
or U1350 (N_1350,N_717,N_535);
and U1351 (N_1351,N_729,N_537);
and U1352 (N_1352,N_936,N_771);
nor U1353 (N_1353,N_621,N_834);
and U1354 (N_1354,N_581,N_669);
nand U1355 (N_1355,N_623,N_889);
or U1356 (N_1356,N_593,N_734);
or U1357 (N_1357,N_698,N_712);
nand U1358 (N_1358,N_969,N_640);
and U1359 (N_1359,N_676,N_974);
or U1360 (N_1360,N_831,N_736);
nand U1361 (N_1361,N_752,N_998);
and U1362 (N_1362,N_808,N_615);
and U1363 (N_1363,N_889,N_774);
nor U1364 (N_1364,N_805,N_927);
nor U1365 (N_1365,N_534,N_626);
or U1366 (N_1366,N_803,N_891);
or U1367 (N_1367,N_833,N_567);
nor U1368 (N_1368,N_634,N_555);
nand U1369 (N_1369,N_709,N_859);
nor U1370 (N_1370,N_849,N_870);
or U1371 (N_1371,N_704,N_787);
nor U1372 (N_1372,N_731,N_528);
xor U1373 (N_1373,N_806,N_574);
and U1374 (N_1374,N_671,N_818);
or U1375 (N_1375,N_821,N_573);
nor U1376 (N_1376,N_986,N_780);
nor U1377 (N_1377,N_574,N_868);
and U1378 (N_1378,N_708,N_969);
and U1379 (N_1379,N_534,N_704);
or U1380 (N_1380,N_661,N_977);
nor U1381 (N_1381,N_663,N_784);
nand U1382 (N_1382,N_712,N_669);
or U1383 (N_1383,N_574,N_553);
or U1384 (N_1384,N_833,N_636);
or U1385 (N_1385,N_928,N_878);
nor U1386 (N_1386,N_755,N_615);
nor U1387 (N_1387,N_672,N_731);
and U1388 (N_1388,N_807,N_590);
nor U1389 (N_1389,N_814,N_810);
or U1390 (N_1390,N_704,N_586);
and U1391 (N_1391,N_960,N_966);
nand U1392 (N_1392,N_650,N_652);
xnor U1393 (N_1393,N_660,N_500);
nor U1394 (N_1394,N_845,N_537);
nand U1395 (N_1395,N_866,N_699);
nor U1396 (N_1396,N_569,N_972);
xnor U1397 (N_1397,N_936,N_594);
nor U1398 (N_1398,N_979,N_684);
xnor U1399 (N_1399,N_608,N_865);
nand U1400 (N_1400,N_664,N_737);
xor U1401 (N_1401,N_799,N_500);
nor U1402 (N_1402,N_993,N_887);
nand U1403 (N_1403,N_882,N_924);
nor U1404 (N_1404,N_730,N_977);
nor U1405 (N_1405,N_618,N_714);
nor U1406 (N_1406,N_577,N_641);
nand U1407 (N_1407,N_518,N_634);
or U1408 (N_1408,N_984,N_718);
nand U1409 (N_1409,N_577,N_550);
or U1410 (N_1410,N_886,N_925);
or U1411 (N_1411,N_538,N_544);
nand U1412 (N_1412,N_572,N_910);
or U1413 (N_1413,N_941,N_533);
nor U1414 (N_1414,N_738,N_729);
and U1415 (N_1415,N_771,N_838);
and U1416 (N_1416,N_662,N_693);
nor U1417 (N_1417,N_953,N_623);
or U1418 (N_1418,N_647,N_564);
nand U1419 (N_1419,N_627,N_715);
and U1420 (N_1420,N_821,N_756);
xor U1421 (N_1421,N_593,N_753);
or U1422 (N_1422,N_844,N_789);
xnor U1423 (N_1423,N_643,N_707);
nor U1424 (N_1424,N_682,N_997);
and U1425 (N_1425,N_866,N_561);
or U1426 (N_1426,N_587,N_579);
nor U1427 (N_1427,N_645,N_877);
nand U1428 (N_1428,N_945,N_970);
xor U1429 (N_1429,N_648,N_544);
and U1430 (N_1430,N_703,N_510);
and U1431 (N_1431,N_869,N_853);
or U1432 (N_1432,N_759,N_972);
nor U1433 (N_1433,N_599,N_702);
nor U1434 (N_1434,N_708,N_815);
or U1435 (N_1435,N_770,N_794);
nor U1436 (N_1436,N_663,N_562);
or U1437 (N_1437,N_659,N_606);
nor U1438 (N_1438,N_759,N_671);
nor U1439 (N_1439,N_727,N_803);
nor U1440 (N_1440,N_642,N_817);
or U1441 (N_1441,N_844,N_606);
and U1442 (N_1442,N_843,N_951);
and U1443 (N_1443,N_769,N_873);
and U1444 (N_1444,N_587,N_631);
or U1445 (N_1445,N_561,N_830);
nand U1446 (N_1446,N_603,N_964);
or U1447 (N_1447,N_906,N_541);
xnor U1448 (N_1448,N_837,N_912);
and U1449 (N_1449,N_544,N_658);
nor U1450 (N_1450,N_659,N_738);
nor U1451 (N_1451,N_700,N_954);
nand U1452 (N_1452,N_584,N_957);
nand U1453 (N_1453,N_737,N_881);
nand U1454 (N_1454,N_987,N_652);
nor U1455 (N_1455,N_578,N_790);
nand U1456 (N_1456,N_841,N_728);
nor U1457 (N_1457,N_814,N_776);
nand U1458 (N_1458,N_790,N_625);
or U1459 (N_1459,N_629,N_632);
and U1460 (N_1460,N_510,N_937);
nor U1461 (N_1461,N_726,N_862);
nor U1462 (N_1462,N_815,N_678);
or U1463 (N_1463,N_546,N_877);
and U1464 (N_1464,N_548,N_689);
nor U1465 (N_1465,N_805,N_854);
and U1466 (N_1466,N_750,N_561);
and U1467 (N_1467,N_819,N_622);
and U1468 (N_1468,N_578,N_571);
and U1469 (N_1469,N_858,N_727);
nor U1470 (N_1470,N_569,N_589);
xnor U1471 (N_1471,N_678,N_658);
nor U1472 (N_1472,N_526,N_743);
and U1473 (N_1473,N_880,N_889);
xor U1474 (N_1474,N_887,N_704);
and U1475 (N_1475,N_647,N_905);
nor U1476 (N_1476,N_960,N_836);
or U1477 (N_1477,N_690,N_881);
or U1478 (N_1478,N_676,N_778);
nor U1479 (N_1479,N_575,N_530);
nand U1480 (N_1480,N_890,N_568);
nor U1481 (N_1481,N_508,N_634);
and U1482 (N_1482,N_698,N_766);
or U1483 (N_1483,N_584,N_546);
and U1484 (N_1484,N_566,N_856);
and U1485 (N_1485,N_610,N_824);
nor U1486 (N_1486,N_564,N_948);
nand U1487 (N_1487,N_933,N_619);
and U1488 (N_1488,N_743,N_547);
xnor U1489 (N_1489,N_585,N_781);
nor U1490 (N_1490,N_852,N_736);
nand U1491 (N_1491,N_619,N_540);
nor U1492 (N_1492,N_634,N_917);
or U1493 (N_1493,N_681,N_810);
nor U1494 (N_1494,N_879,N_545);
nand U1495 (N_1495,N_969,N_986);
nand U1496 (N_1496,N_756,N_574);
and U1497 (N_1497,N_711,N_997);
and U1498 (N_1498,N_796,N_758);
and U1499 (N_1499,N_809,N_658);
nor U1500 (N_1500,N_1045,N_1256);
xnor U1501 (N_1501,N_1396,N_1486);
nand U1502 (N_1502,N_1471,N_1296);
nor U1503 (N_1503,N_1333,N_1157);
nand U1504 (N_1504,N_1418,N_1000);
nor U1505 (N_1505,N_1320,N_1131);
or U1506 (N_1506,N_1212,N_1147);
nand U1507 (N_1507,N_1355,N_1406);
xor U1508 (N_1508,N_1439,N_1370);
nand U1509 (N_1509,N_1323,N_1059);
and U1510 (N_1510,N_1089,N_1055);
and U1511 (N_1511,N_1150,N_1160);
nand U1512 (N_1512,N_1487,N_1428);
nand U1513 (N_1513,N_1152,N_1085);
nor U1514 (N_1514,N_1291,N_1459);
or U1515 (N_1515,N_1193,N_1007);
or U1516 (N_1516,N_1113,N_1158);
nand U1517 (N_1517,N_1378,N_1096);
nor U1518 (N_1518,N_1168,N_1324);
xnor U1519 (N_1519,N_1165,N_1119);
nor U1520 (N_1520,N_1397,N_1339);
and U1521 (N_1521,N_1308,N_1376);
or U1522 (N_1522,N_1117,N_1412);
and U1523 (N_1523,N_1473,N_1340);
nor U1524 (N_1524,N_1024,N_1088);
nand U1525 (N_1525,N_1057,N_1006);
and U1526 (N_1526,N_1315,N_1034);
or U1527 (N_1527,N_1084,N_1095);
nor U1528 (N_1528,N_1071,N_1419);
and U1529 (N_1529,N_1164,N_1438);
nor U1530 (N_1530,N_1031,N_1103);
xnor U1531 (N_1531,N_1224,N_1003);
and U1532 (N_1532,N_1026,N_1306);
nor U1533 (N_1533,N_1145,N_1101);
xor U1534 (N_1534,N_1138,N_1227);
nor U1535 (N_1535,N_1022,N_1070);
nor U1536 (N_1536,N_1363,N_1077);
or U1537 (N_1537,N_1275,N_1097);
nand U1538 (N_1538,N_1192,N_1060);
nand U1539 (N_1539,N_1043,N_1407);
xor U1540 (N_1540,N_1260,N_1016);
xnor U1541 (N_1541,N_1146,N_1350);
nand U1542 (N_1542,N_1116,N_1468);
nor U1543 (N_1543,N_1074,N_1231);
and U1544 (N_1544,N_1232,N_1008);
and U1545 (N_1545,N_1399,N_1432);
or U1546 (N_1546,N_1206,N_1137);
xnor U1547 (N_1547,N_1421,N_1237);
or U1548 (N_1548,N_1234,N_1174);
xnor U1549 (N_1549,N_1049,N_1255);
nand U1550 (N_1550,N_1222,N_1081);
xor U1551 (N_1551,N_1243,N_1281);
nor U1552 (N_1552,N_1358,N_1374);
or U1553 (N_1553,N_1056,N_1280);
or U1554 (N_1554,N_1114,N_1394);
nor U1555 (N_1555,N_1038,N_1429);
nor U1556 (N_1556,N_1175,N_1140);
nor U1557 (N_1557,N_1162,N_1261);
or U1558 (N_1558,N_1287,N_1381);
and U1559 (N_1559,N_1303,N_1445);
and U1560 (N_1560,N_1436,N_1037);
and U1561 (N_1561,N_1390,N_1493);
and U1562 (N_1562,N_1442,N_1076);
and U1563 (N_1563,N_1298,N_1029);
or U1564 (N_1564,N_1182,N_1460);
nor U1565 (N_1565,N_1082,N_1433);
or U1566 (N_1566,N_1475,N_1434);
nand U1567 (N_1567,N_1293,N_1110);
nor U1568 (N_1568,N_1209,N_1127);
and U1569 (N_1569,N_1310,N_1373);
nand U1570 (N_1570,N_1080,N_1416);
and U1571 (N_1571,N_1353,N_1242);
or U1572 (N_1572,N_1249,N_1004);
nand U1573 (N_1573,N_1297,N_1120);
and U1574 (N_1574,N_1498,N_1229);
or U1575 (N_1575,N_1349,N_1267);
nor U1576 (N_1576,N_1451,N_1033);
nor U1577 (N_1577,N_1216,N_1424);
nor U1578 (N_1578,N_1321,N_1359);
xor U1579 (N_1579,N_1420,N_1448);
or U1580 (N_1580,N_1210,N_1257);
nand U1581 (N_1581,N_1200,N_1361);
or U1582 (N_1582,N_1090,N_1472);
or U1583 (N_1583,N_1148,N_1091);
and U1584 (N_1584,N_1213,N_1154);
xor U1585 (N_1585,N_1235,N_1379);
and U1586 (N_1586,N_1012,N_1130);
and U1587 (N_1587,N_1479,N_1447);
and U1588 (N_1588,N_1063,N_1017);
nor U1589 (N_1589,N_1273,N_1204);
nand U1590 (N_1590,N_1300,N_1496);
and U1591 (N_1591,N_1069,N_1041);
nor U1592 (N_1592,N_1302,N_1356);
and U1593 (N_1593,N_1129,N_1292);
xor U1594 (N_1594,N_1388,N_1497);
nand U1595 (N_1595,N_1124,N_1180);
and U1596 (N_1596,N_1371,N_1485);
nand U1597 (N_1597,N_1367,N_1347);
xor U1598 (N_1598,N_1387,N_1187);
nor U1599 (N_1599,N_1128,N_1466);
or U1600 (N_1600,N_1392,N_1372);
nor U1601 (N_1601,N_1405,N_1239);
or U1602 (N_1602,N_1105,N_1036);
nand U1603 (N_1603,N_1410,N_1177);
or U1604 (N_1604,N_1430,N_1413);
and U1605 (N_1605,N_1050,N_1400);
and U1606 (N_1606,N_1126,N_1005);
or U1607 (N_1607,N_1304,N_1369);
and U1608 (N_1608,N_1285,N_1247);
xor U1609 (N_1609,N_1214,N_1348);
or U1610 (N_1610,N_1122,N_1385);
nor U1611 (N_1611,N_1440,N_1068);
nand U1612 (N_1612,N_1318,N_1377);
and U1613 (N_1613,N_1264,N_1276);
nand U1614 (N_1614,N_1020,N_1455);
and U1615 (N_1615,N_1284,N_1289);
and U1616 (N_1616,N_1015,N_1325);
or U1617 (N_1617,N_1199,N_1048);
and U1618 (N_1618,N_1389,N_1345);
nand U1619 (N_1619,N_1141,N_1228);
or U1620 (N_1620,N_1201,N_1366);
nor U1621 (N_1621,N_1453,N_1328);
nor U1622 (N_1622,N_1384,N_1317);
nor U1623 (N_1623,N_1208,N_1401);
nand U1624 (N_1624,N_1014,N_1032);
and U1625 (N_1625,N_1279,N_1272);
xnor U1626 (N_1626,N_1002,N_1258);
nand U1627 (N_1627,N_1266,N_1094);
nand U1628 (N_1628,N_1171,N_1169);
nand U1629 (N_1629,N_1277,N_1013);
nor U1630 (N_1630,N_1312,N_1018);
or U1631 (N_1631,N_1452,N_1044);
or U1632 (N_1632,N_1327,N_1435);
and U1633 (N_1633,N_1181,N_1118);
or U1634 (N_1634,N_1295,N_1437);
nor U1635 (N_1635,N_1144,N_1046);
xor U1636 (N_1636,N_1143,N_1313);
xnor U1637 (N_1637,N_1079,N_1283);
nor U1638 (N_1638,N_1065,N_1035);
nand U1639 (N_1639,N_1125,N_1001);
nor U1640 (N_1640,N_1191,N_1215);
and U1641 (N_1641,N_1030,N_1478);
xnor U1642 (N_1642,N_1104,N_1458);
or U1643 (N_1643,N_1386,N_1155);
nor U1644 (N_1644,N_1423,N_1305);
and U1645 (N_1645,N_1488,N_1480);
xnor U1646 (N_1646,N_1268,N_1221);
or U1647 (N_1647,N_1380,N_1334);
nand U1648 (N_1648,N_1178,N_1444);
or U1649 (N_1649,N_1494,N_1454);
nand U1650 (N_1650,N_1025,N_1136);
nand U1651 (N_1651,N_1106,N_1262);
and U1652 (N_1652,N_1271,N_1245);
nor U1653 (N_1653,N_1269,N_1054);
or U1654 (N_1654,N_1058,N_1462);
or U1655 (N_1655,N_1023,N_1299);
nand U1656 (N_1656,N_1248,N_1270);
or U1657 (N_1657,N_1250,N_1446);
nand U1658 (N_1658,N_1408,N_1252);
and U1659 (N_1659,N_1490,N_1461);
nand U1660 (N_1660,N_1417,N_1330);
nand U1661 (N_1661,N_1415,N_1112);
nor U1662 (N_1662,N_1307,N_1134);
nand U1663 (N_1663,N_1111,N_1259);
and U1664 (N_1664,N_1251,N_1364);
nor U1665 (N_1665,N_1205,N_1395);
nor U1666 (N_1666,N_1391,N_1335);
and U1667 (N_1667,N_1316,N_1163);
or U1668 (N_1668,N_1087,N_1477);
and U1669 (N_1669,N_1135,N_1053);
nor U1670 (N_1670,N_1166,N_1491);
nand U1671 (N_1671,N_1064,N_1198);
or U1672 (N_1672,N_1230,N_1170);
nor U1673 (N_1673,N_1139,N_1115);
xor U1674 (N_1674,N_1109,N_1010);
nor U1675 (N_1675,N_1176,N_1078);
and U1676 (N_1676,N_1073,N_1197);
nor U1677 (N_1677,N_1241,N_1337);
nor U1678 (N_1678,N_1238,N_1286);
or U1679 (N_1679,N_1301,N_1196);
nor U1680 (N_1680,N_1086,N_1021);
nand U1681 (N_1681,N_1233,N_1067);
and U1682 (N_1682,N_1311,N_1288);
or U1683 (N_1683,N_1167,N_1188);
nand U1684 (N_1684,N_1393,N_1464);
nor U1685 (N_1685,N_1414,N_1360);
or U1686 (N_1686,N_1482,N_1483);
nand U1687 (N_1687,N_1470,N_1042);
nand U1688 (N_1688,N_1052,N_1274);
or U1689 (N_1689,N_1011,N_1083);
nor U1690 (N_1690,N_1457,N_1489);
or U1691 (N_1691,N_1357,N_1290);
or U1692 (N_1692,N_1263,N_1027);
nor U1693 (N_1693,N_1309,N_1254);
and U1694 (N_1694,N_1246,N_1265);
and U1695 (N_1695,N_1329,N_1427);
nand U1696 (N_1696,N_1422,N_1338);
or U1697 (N_1697,N_1481,N_1183);
or U1698 (N_1698,N_1108,N_1240);
nor U1699 (N_1699,N_1207,N_1362);
and U1700 (N_1700,N_1411,N_1009);
nand U1701 (N_1701,N_1403,N_1039);
and U1702 (N_1702,N_1467,N_1474);
xnor U1703 (N_1703,N_1441,N_1352);
xnor U1704 (N_1704,N_1217,N_1132);
and U1705 (N_1705,N_1469,N_1019);
nand U1706 (N_1706,N_1463,N_1365);
xor U1707 (N_1707,N_1332,N_1368);
or U1708 (N_1708,N_1425,N_1495);
nand U1709 (N_1709,N_1040,N_1426);
or U1710 (N_1710,N_1195,N_1211);
xnor U1711 (N_1711,N_1066,N_1156);
nor U1712 (N_1712,N_1172,N_1189);
nor U1713 (N_1713,N_1092,N_1398);
xor U1714 (N_1714,N_1223,N_1142);
or U1715 (N_1715,N_1102,N_1153);
or U1716 (N_1716,N_1190,N_1346);
nor U1717 (N_1717,N_1319,N_1322);
or U1718 (N_1718,N_1099,N_1186);
nand U1719 (N_1719,N_1179,N_1098);
or U1720 (N_1720,N_1184,N_1382);
nand U1721 (N_1721,N_1194,N_1121);
nor U1722 (N_1722,N_1402,N_1278);
nand U1723 (N_1723,N_1443,N_1219);
or U1724 (N_1724,N_1202,N_1161);
and U1725 (N_1725,N_1149,N_1326);
nor U1726 (N_1726,N_1203,N_1342);
or U1727 (N_1727,N_1465,N_1404);
nor U1728 (N_1728,N_1351,N_1450);
nand U1729 (N_1729,N_1100,N_1354);
nor U1730 (N_1730,N_1093,N_1159);
and U1731 (N_1731,N_1051,N_1476);
xnor U1732 (N_1732,N_1236,N_1047);
xor U1733 (N_1733,N_1107,N_1253);
nand U1734 (N_1734,N_1409,N_1314);
nor U1735 (N_1735,N_1123,N_1218);
or U1736 (N_1736,N_1173,N_1341);
nand U1737 (N_1737,N_1185,N_1383);
and U1738 (N_1738,N_1331,N_1449);
or U1739 (N_1739,N_1244,N_1294);
nand U1740 (N_1740,N_1226,N_1492);
xor U1741 (N_1741,N_1282,N_1133);
xor U1742 (N_1742,N_1336,N_1225);
nor U1743 (N_1743,N_1151,N_1343);
nand U1744 (N_1744,N_1456,N_1028);
and U1745 (N_1745,N_1220,N_1062);
nand U1746 (N_1746,N_1072,N_1344);
nand U1747 (N_1747,N_1499,N_1075);
nor U1748 (N_1748,N_1375,N_1061);
xnor U1749 (N_1749,N_1431,N_1484);
and U1750 (N_1750,N_1190,N_1268);
nand U1751 (N_1751,N_1365,N_1371);
xor U1752 (N_1752,N_1230,N_1110);
and U1753 (N_1753,N_1049,N_1235);
nand U1754 (N_1754,N_1404,N_1226);
nor U1755 (N_1755,N_1121,N_1297);
nand U1756 (N_1756,N_1017,N_1495);
or U1757 (N_1757,N_1209,N_1356);
nor U1758 (N_1758,N_1123,N_1438);
xor U1759 (N_1759,N_1252,N_1092);
and U1760 (N_1760,N_1023,N_1280);
and U1761 (N_1761,N_1277,N_1090);
nor U1762 (N_1762,N_1073,N_1208);
or U1763 (N_1763,N_1152,N_1226);
and U1764 (N_1764,N_1491,N_1100);
xnor U1765 (N_1765,N_1487,N_1186);
and U1766 (N_1766,N_1475,N_1035);
nor U1767 (N_1767,N_1036,N_1111);
or U1768 (N_1768,N_1358,N_1266);
nor U1769 (N_1769,N_1316,N_1406);
nand U1770 (N_1770,N_1185,N_1291);
or U1771 (N_1771,N_1042,N_1168);
or U1772 (N_1772,N_1473,N_1131);
nor U1773 (N_1773,N_1003,N_1372);
nor U1774 (N_1774,N_1012,N_1152);
nor U1775 (N_1775,N_1104,N_1115);
nand U1776 (N_1776,N_1118,N_1015);
and U1777 (N_1777,N_1444,N_1400);
nand U1778 (N_1778,N_1306,N_1052);
nand U1779 (N_1779,N_1012,N_1347);
nor U1780 (N_1780,N_1110,N_1244);
and U1781 (N_1781,N_1469,N_1090);
xor U1782 (N_1782,N_1166,N_1014);
nand U1783 (N_1783,N_1079,N_1384);
nand U1784 (N_1784,N_1386,N_1325);
nand U1785 (N_1785,N_1218,N_1406);
nand U1786 (N_1786,N_1368,N_1355);
and U1787 (N_1787,N_1382,N_1372);
or U1788 (N_1788,N_1305,N_1199);
nand U1789 (N_1789,N_1104,N_1216);
or U1790 (N_1790,N_1247,N_1169);
xnor U1791 (N_1791,N_1355,N_1153);
and U1792 (N_1792,N_1359,N_1492);
xnor U1793 (N_1793,N_1454,N_1026);
or U1794 (N_1794,N_1418,N_1446);
nor U1795 (N_1795,N_1366,N_1301);
and U1796 (N_1796,N_1127,N_1277);
nor U1797 (N_1797,N_1030,N_1092);
nor U1798 (N_1798,N_1345,N_1201);
nor U1799 (N_1799,N_1251,N_1158);
nand U1800 (N_1800,N_1005,N_1372);
or U1801 (N_1801,N_1171,N_1375);
or U1802 (N_1802,N_1187,N_1277);
and U1803 (N_1803,N_1255,N_1139);
or U1804 (N_1804,N_1480,N_1412);
nand U1805 (N_1805,N_1015,N_1243);
or U1806 (N_1806,N_1340,N_1155);
xor U1807 (N_1807,N_1171,N_1360);
and U1808 (N_1808,N_1415,N_1270);
or U1809 (N_1809,N_1389,N_1072);
nor U1810 (N_1810,N_1172,N_1483);
or U1811 (N_1811,N_1123,N_1382);
and U1812 (N_1812,N_1179,N_1137);
and U1813 (N_1813,N_1099,N_1181);
xnor U1814 (N_1814,N_1185,N_1303);
nor U1815 (N_1815,N_1290,N_1188);
and U1816 (N_1816,N_1392,N_1055);
and U1817 (N_1817,N_1147,N_1084);
xor U1818 (N_1818,N_1133,N_1116);
xnor U1819 (N_1819,N_1149,N_1129);
nand U1820 (N_1820,N_1041,N_1204);
nor U1821 (N_1821,N_1477,N_1377);
or U1822 (N_1822,N_1491,N_1253);
nand U1823 (N_1823,N_1303,N_1092);
and U1824 (N_1824,N_1241,N_1021);
or U1825 (N_1825,N_1489,N_1171);
and U1826 (N_1826,N_1414,N_1397);
or U1827 (N_1827,N_1031,N_1052);
and U1828 (N_1828,N_1251,N_1000);
nand U1829 (N_1829,N_1104,N_1442);
nor U1830 (N_1830,N_1054,N_1469);
nor U1831 (N_1831,N_1231,N_1098);
and U1832 (N_1832,N_1308,N_1216);
or U1833 (N_1833,N_1156,N_1201);
or U1834 (N_1834,N_1279,N_1318);
or U1835 (N_1835,N_1398,N_1307);
nand U1836 (N_1836,N_1004,N_1259);
and U1837 (N_1837,N_1357,N_1117);
nor U1838 (N_1838,N_1401,N_1037);
nor U1839 (N_1839,N_1355,N_1470);
nand U1840 (N_1840,N_1012,N_1030);
and U1841 (N_1841,N_1217,N_1108);
and U1842 (N_1842,N_1112,N_1420);
and U1843 (N_1843,N_1340,N_1422);
nand U1844 (N_1844,N_1023,N_1294);
nand U1845 (N_1845,N_1082,N_1033);
nand U1846 (N_1846,N_1121,N_1345);
nand U1847 (N_1847,N_1196,N_1019);
nand U1848 (N_1848,N_1424,N_1270);
nand U1849 (N_1849,N_1431,N_1237);
and U1850 (N_1850,N_1149,N_1248);
or U1851 (N_1851,N_1220,N_1131);
nand U1852 (N_1852,N_1391,N_1317);
nor U1853 (N_1853,N_1311,N_1227);
nor U1854 (N_1854,N_1384,N_1040);
and U1855 (N_1855,N_1378,N_1432);
or U1856 (N_1856,N_1037,N_1418);
or U1857 (N_1857,N_1052,N_1035);
and U1858 (N_1858,N_1172,N_1425);
nor U1859 (N_1859,N_1357,N_1490);
nand U1860 (N_1860,N_1206,N_1490);
xor U1861 (N_1861,N_1176,N_1084);
nor U1862 (N_1862,N_1419,N_1261);
nor U1863 (N_1863,N_1188,N_1018);
xnor U1864 (N_1864,N_1083,N_1036);
nand U1865 (N_1865,N_1080,N_1383);
nand U1866 (N_1866,N_1456,N_1049);
nand U1867 (N_1867,N_1146,N_1066);
xor U1868 (N_1868,N_1486,N_1134);
xor U1869 (N_1869,N_1250,N_1347);
nor U1870 (N_1870,N_1374,N_1217);
and U1871 (N_1871,N_1159,N_1456);
or U1872 (N_1872,N_1342,N_1006);
nand U1873 (N_1873,N_1221,N_1190);
and U1874 (N_1874,N_1497,N_1082);
or U1875 (N_1875,N_1119,N_1370);
and U1876 (N_1876,N_1201,N_1173);
and U1877 (N_1877,N_1365,N_1092);
xnor U1878 (N_1878,N_1324,N_1416);
nor U1879 (N_1879,N_1391,N_1378);
xnor U1880 (N_1880,N_1452,N_1082);
nand U1881 (N_1881,N_1393,N_1222);
nand U1882 (N_1882,N_1204,N_1047);
nor U1883 (N_1883,N_1225,N_1496);
nor U1884 (N_1884,N_1069,N_1064);
nor U1885 (N_1885,N_1061,N_1365);
nand U1886 (N_1886,N_1387,N_1076);
or U1887 (N_1887,N_1174,N_1388);
nor U1888 (N_1888,N_1497,N_1390);
or U1889 (N_1889,N_1235,N_1473);
nand U1890 (N_1890,N_1362,N_1429);
or U1891 (N_1891,N_1263,N_1178);
and U1892 (N_1892,N_1344,N_1076);
and U1893 (N_1893,N_1168,N_1200);
or U1894 (N_1894,N_1402,N_1133);
and U1895 (N_1895,N_1260,N_1297);
nor U1896 (N_1896,N_1072,N_1275);
xnor U1897 (N_1897,N_1334,N_1283);
nand U1898 (N_1898,N_1388,N_1177);
nor U1899 (N_1899,N_1146,N_1329);
and U1900 (N_1900,N_1491,N_1475);
nand U1901 (N_1901,N_1139,N_1261);
nand U1902 (N_1902,N_1417,N_1359);
and U1903 (N_1903,N_1219,N_1245);
or U1904 (N_1904,N_1277,N_1280);
nand U1905 (N_1905,N_1356,N_1090);
xor U1906 (N_1906,N_1046,N_1270);
nor U1907 (N_1907,N_1280,N_1040);
nand U1908 (N_1908,N_1131,N_1480);
or U1909 (N_1909,N_1458,N_1358);
xor U1910 (N_1910,N_1198,N_1182);
nand U1911 (N_1911,N_1404,N_1227);
nand U1912 (N_1912,N_1197,N_1414);
nand U1913 (N_1913,N_1109,N_1096);
nand U1914 (N_1914,N_1325,N_1492);
xnor U1915 (N_1915,N_1468,N_1452);
nand U1916 (N_1916,N_1062,N_1264);
and U1917 (N_1917,N_1035,N_1331);
and U1918 (N_1918,N_1215,N_1218);
and U1919 (N_1919,N_1407,N_1174);
or U1920 (N_1920,N_1185,N_1070);
nand U1921 (N_1921,N_1072,N_1295);
or U1922 (N_1922,N_1088,N_1195);
and U1923 (N_1923,N_1406,N_1343);
nor U1924 (N_1924,N_1489,N_1407);
nand U1925 (N_1925,N_1166,N_1267);
or U1926 (N_1926,N_1440,N_1080);
or U1927 (N_1927,N_1241,N_1362);
or U1928 (N_1928,N_1023,N_1115);
or U1929 (N_1929,N_1342,N_1140);
xor U1930 (N_1930,N_1470,N_1052);
or U1931 (N_1931,N_1107,N_1119);
nand U1932 (N_1932,N_1111,N_1137);
nand U1933 (N_1933,N_1095,N_1202);
nand U1934 (N_1934,N_1449,N_1339);
nand U1935 (N_1935,N_1197,N_1393);
xnor U1936 (N_1936,N_1120,N_1098);
or U1937 (N_1937,N_1280,N_1237);
nand U1938 (N_1938,N_1098,N_1201);
and U1939 (N_1939,N_1065,N_1326);
nor U1940 (N_1940,N_1363,N_1321);
nor U1941 (N_1941,N_1440,N_1178);
nor U1942 (N_1942,N_1342,N_1452);
or U1943 (N_1943,N_1143,N_1281);
or U1944 (N_1944,N_1165,N_1361);
or U1945 (N_1945,N_1290,N_1275);
xor U1946 (N_1946,N_1289,N_1392);
or U1947 (N_1947,N_1095,N_1387);
or U1948 (N_1948,N_1276,N_1488);
nor U1949 (N_1949,N_1034,N_1015);
and U1950 (N_1950,N_1202,N_1060);
or U1951 (N_1951,N_1283,N_1354);
nor U1952 (N_1952,N_1378,N_1419);
nor U1953 (N_1953,N_1359,N_1427);
nand U1954 (N_1954,N_1383,N_1062);
and U1955 (N_1955,N_1020,N_1223);
or U1956 (N_1956,N_1103,N_1404);
nand U1957 (N_1957,N_1197,N_1155);
nor U1958 (N_1958,N_1214,N_1409);
nand U1959 (N_1959,N_1199,N_1250);
nand U1960 (N_1960,N_1298,N_1270);
or U1961 (N_1961,N_1061,N_1398);
nand U1962 (N_1962,N_1251,N_1060);
or U1963 (N_1963,N_1390,N_1487);
nand U1964 (N_1964,N_1350,N_1172);
and U1965 (N_1965,N_1415,N_1057);
and U1966 (N_1966,N_1129,N_1029);
nand U1967 (N_1967,N_1210,N_1108);
nor U1968 (N_1968,N_1377,N_1089);
nor U1969 (N_1969,N_1043,N_1290);
nor U1970 (N_1970,N_1042,N_1082);
and U1971 (N_1971,N_1427,N_1057);
and U1972 (N_1972,N_1238,N_1162);
and U1973 (N_1973,N_1422,N_1448);
and U1974 (N_1974,N_1216,N_1183);
or U1975 (N_1975,N_1287,N_1454);
xnor U1976 (N_1976,N_1265,N_1104);
nand U1977 (N_1977,N_1424,N_1291);
and U1978 (N_1978,N_1446,N_1414);
nand U1979 (N_1979,N_1192,N_1047);
nor U1980 (N_1980,N_1107,N_1332);
nand U1981 (N_1981,N_1241,N_1126);
xor U1982 (N_1982,N_1001,N_1304);
and U1983 (N_1983,N_1079,N_1007);
and U1984 (N_1984,N_1075,N_1185);
nand U1985 (N_1985,N_1374,N_1123);
and U1986 (N_1986,N_1367,N_1377);
nor U1987 (N_1987,N_1437,N_1155);
nand U1988 (N_1988,N_1184,N_1289);
nand U1989 (N_1989,N_1042,N_1062);
nor U1990 (N_1990,N_1493,N_1324);
and U1991 (N_1991,N_1026,N_1080);
or U1992 (N_1992,N_1137,N_1065);
nand U1993 (N_1993,N_1038,N_1061);
nand U1994 (N_1994,N_1001,N_1108);
or U1995 (N_1995,N_1411,N_1475);
or U1996 (N_1996,N_1086,N_1380);
or U1997 (N_1997,N_1144,N_1159);
nand U1998 (N_1998,N_1387,N_1253);
nor U1999 (N_1999,N_1254,N_1390);
and U2000 (N_2000,N_1967,N_1953);
and U2001 (N_2001,N_1971,N_1812);
xor U2002 (N_2002,N_1979,N_1550);
or U2003 (N_2003,N_1770,N_1689);
or U2004 (N_2004,N_1831,N_1938);
xnor U2005 (N_2005,N_1843,N_1538);
xor U2006 (N_2006,N_1574,N_1524);
nor U2007 (N_2007,N_1792,N_1936);
and U2008 (N_2008,N_1886,N_1963);
or U2009 (N_2009,N_1521,N_1987);
and U2010 (N_2010,N_1684,N_1997);
nor U2011 (N_2011,N_1601,N_1836);
or U2012 (N_2012,N_1702,N_1691);
nor U2013 (N_2013,N_1632,N_1756);
or U2014 (N_2014,N_1842,N_1719);
nand U2015 (N_2015,N_1977,N_1942);
or U2016 (N_2016,N_1563,N_1533);
nand U2017 (N_2017,N_1976,N_1951);
or U2018 (N_2018,N_1730,N_1864);
nand U2019 (N_2019,N_1749,N_1620);
nor U2020 (N_2020,N_1784,N_1532);
nor U2021 (N_2021,N_1595,N_1518);
or U2022 (N_2022,N_1813,N_1718);
and U2023 (N_2023,N_1991,N_1782);
or U2024 (N_2024,N_1899,N_1654);
nor U2025 (N_2025,N_1698,N_1885);
nand U2026 (N_2026,N_1776,N_1858);
or U2027 (N_2027,N_1923,N_1531);
nand U2028 (N_2028,N_1775,N_1765);
and U2029 (N_2029,N_1935,N_1860);
nand U2030 (N_2030,N_1818,N_1608);
and U2031 (N_2031,N_1824,N_1832);
and U2032 (N_2032,N_1551,N_1525);
and U2033 (N_2033,N_1980,N_1777);
and U2034 (N_2034,N_1728,N_1635);
nand U2035 (N_2035,N_1580,N_1946);
nor U2036 (N_2036,N_1652,N_1578);
nor U2037 (N_2037,N_1708,N_1514);
or U2038 (N_2038,N_1859,N_1581);
and U2039 (N_2039,N_1767,N_1788);
xor U2040 (N_2040,N_1850,N_1806);
or U2041 (N_2041,N_1755,N_1695);
nor U2042 (N_2042,N_1693,N_1814);
nand U2043 (N_2043,N_1631,N_1570);
and U2044 (N_2044,N_1547,N_1764);
or U2045 (N_2045,N_1627,N_1732);
or U2046 (N_2046,N_1740,N_1862);
nor U2047 (N_2047,N_1848,N_1981);
nor U2048 (N_2048,N_1930,N_1648);
nand U2049 (N_2049,N_1807,N_1865);
nor U2050 (N_2050,N_1944,N_1681);
nor U2051 (N_2051,N_1513,N_1863);
and U2052 (N_2052,N_1828,N_1887);
nand U2053 (N_2053,N_1901,N_1933);
and U2054 (N_2054,N_1639,N_1522);
xor U2055 (N_2055,N_1705,N_1622);
and U2056 (N_2056,N_1750,N_1778);
nor U2057 (N_2057,N_1841,N_1539);
nand U2058 (N_2058,N_1616,N_1955);
and U2059 (N_2059,N_1893,N_1896);
nor U2060 (N_2060,N_1706,N_1854);
nand U2061 (N_2061,N_1676,N_1633);
nor U2062 (N_2062,N_1895,N_1736);
nor U2063 (N_2063,N_1663,N_1723);
nor U2064 (N_2064,N_1928,N_1826);
or U2065 (N_2065,N_1754,N_1875);
nor U2066 (N_2066,N_1978,N_1867);
or U2067 (N_2067,N_1996,N_1985);
nor U2068 (N_2068,N_1834,N_1903);
or U2069 (N_2069,N_1602,N_1528);
nor U2070 (N_2070,N_1894,N_1948);
xor U2071 (N_2071,N_1964,N_1805);
and U2072 (N_2072,N_1808,N_1556);
nand U2073 (N_2073,N_1995,N_1697);
and U2074 (N_2074,N_1596,N_1509);
nor U2075 (N_2075,N_1512,N_1820);
or U2076 (N_2076,N_1751,N_1900);
and U2077 (N_2077,N_1594,N_1579);
and U2078 (N_2078,N_1529,N_1816);
nand U2079 (N_2079,N_1994,N_1891);
and U2080 (N_2080,N_1604,N_1536);
and U2081 (N_2081,N_1888,N_1607);
xnor U2082 (N_2082,N_1611,N_1866);
xor U2083 (N_2083,N_1612,N_1873);
nor U2084 (N_2084,N_1999,N_1815);
nand U2085 (N_2085,N_1658,N_1629);
xnor U2086 (N_2086,N_1742,N_1564);
nor U2087 (N_2087,N_1537,N_1932);
nor U2088 (N_2088,N_1837,N_1712);
and U2089 (N_2089,N_1506,N_1647);
nor U2090 (N_2090,N_1857,N_1660);
nor U2091 (N_2091,N_1950,N_1700);
and U2092 (N_2092,N_1910,N_1990);
nand U2093 (N_2093,N_1982,N_1984);
nand U2094 (N_2094,N_1656,N_1729);
nor U2095 (N_2095,N_1657,N_1746);
nand U2096 (N_2096,N_1502,N_1825);
or U2097 (N_2097,N_1558,N_1527);
or U2098 (N_2098,N_1956,N_1752);
or U2099 (N_2099,N_1599,N_1553);
or U2100 (N_2100,N_1905,N_1795);
and U2101 (N_2101,N_1793,N_1501);
or U2102 (N_2102,N_1758,N_1572);
and U2103 (N_2103,N_1645,N_1701);
nand U2104 (N_2104,N_1710,N_1517);
or U2105 (N_2105,N_1582,N_1821);
or U2106 (N_2106,N_1716,N_1717);
and U2107 (N_2107,N_1802,N_1743);
and U2108 (N_2108,N_1630,N_1714);
or U2109 (N_2109,N_1926,N_1500);
or U2110 (N_2110,N_1838,N_1817);
or U2111 (N_2111,N_1542,N_1762);
xor U2112 (N_2112,N_1646,N_1929);
and U2113 (N_2113,N_1911,N_1739);
and U2114 (N_2114,N_1679,N_1909);
nor U2115 (N_2115,N_1849,N_1733);
or U2116 (N_2116,N_1561,N_1803);
nor U2117 (N_2117,N_1968,N_1827);
xor U2118 (N_2118,N_1884,N_1810);
xor U2119 (N_2119,N_1851,N_1941);
nand U2120 (N_2120,N_1880,N_1940);
or U2121 (N_2121,N_1721,N_1567);
or U2122 (N_2122,N_1907,N_1575);
xnor U2123 (N_2123,N_1715,N_1516);
and U2124 (N_2124,N_1783,N_1625);
or U2125 (N_2125,N_1829,N_1993);
nand U2126 (N_2126,N_1510,N_1962);
nand U2127 (N_2127,N_1677,N_1919);
and U2128 (N_2128,N_1945,N_1785);
nand U2129 (N_2129,N_1643,N_1922);
nor U2130 (N_2130,N_1641,N_1548);
nor U2131 (N_2131,N_1515,N_1722);
and U2132 (N_2132,N_1526,N_1613);
nor U2133 (N_2133,N_1519,N_1947);
nand U2134 (N_2134,N_1667,N_1690);
and U2135 (N_2135,N_1789,N_1724);
nand U2136 (N_2136,N_1560,N_1753);
nor U2137 (N_2137,N_1839,N_1897);
and U2138 (N_2138,N_1786,N_1668);
and U2139 (N_2139,N_1606,N_1798);
and U2140 (N_2140,N_1852,N_1794);
or U2141 (N_2141,N_1686,N_1954);
and U2142 (N_2142,N_1585,N_1823);
or U2143 (N_2143,N_1682,N_1576);
and U2144 (N_2144,N_1735,N_1586);
xnor U2145 (N_2145,N_1549,N_1869);
or U2146 (N_2146,N_1874,N_1559);
nor U2147 (N_2147,N_1592,N_1711);
nand U2148 (N_2148,N_1505,N_1726);
or U2149 (N_2149,N_1796,N_1797);
nor U2150 (N_2150,N_1638,N_1543);
and U2151 (N_2151,N_1904,N_1757);
or U2152 (N_2152,N_1661,N_1998);
nor U2153 (N_2153,N_1666,N_1988);
nor U2154 (N_2154,N_1844,N_1769);
and U2155 (N_2155,N_1653,N_1552);
and U2156 (N_2156,N_1876,N_1872);
nor U2157 (N_2157,N_1680,N_1508);
and U2158 (N_2158,N_1649,N_1861);
nand U2159 (N_2159,N_1881,N_1809);
nor U2160 (N_2160,N_1921,N_1853);
and U2161 (N_2161,N_1744,N_1618);
nor U2162 (N_2162,N_1833,N_1605);
nand U2163 (N_2163,N_1617,N_1745);
nor U2164 (N_2164,N_1709,N_1925);
nor U2165 (N_2165,N_1628,N_1889);
or U2166 (N_2166,N_1966,N_1882);
or U2167 (N_2167,N_1734,N_1610);
nand U2168 (N_2168,N_1912,N_1662);
nand U2169 (N_2169,N_1771,N_1787);
xor U2170 (N_2170,N_1692,N_1615);
nor U2171 (N_2171,N_1520,N_1800);
and U2172 (N_2172,N_1636,N_1665);
nand U2173 (N_2173,N_1598,N_1623);
nand U2174 (N_2174,N_1694,N_1688);
and U2175 (N_2175,N_1727,N_1687);
nand U2176 (N_2176,N_1699,N_1544);
nand U2177 (N_2177,N_1624,N_1642);
and U2178 (N_2178,N_1914,N_1673);
nand U2179 (N_2179,N_1975,N_1822);
nand U2180 (N_2180,N_1918,N_1507);
or U2181 (N_2181,N_1906,N_1614);
nand U2182 (N_2182,N_1801,N_1748);
and U2183 (N_2183,N_1591,N_1915);
xnor U2184 (N_2184,N_1637,N_1603);
nor U2185 (N_2185,N_1671,N_1983);
or U2186 (N_2186,N_1768,N_1703);
or U2187 (N_2187,N_1811,N_1685);
and U2188 (N_2188,N_1588,N_1626);
nand U2189 (N_2189,N_1713,N_1504);
xnor U2190 (N_2190,N_1846,N_1773);
or U2191 (N_2191,N_1707,N_1759);
nand U2192 (N_2192,N_1761,N_1835);
and U2193 (N_2193,N_1927,N_1651);
or U2194 (N_2194,N_1781,N_1924);
nand U2195 (N_2195,N_1961,N_1541);
and U2196 (N_2196,N_1763,N_1879);
nor U2197 (N_2197,N_1696,N_1819);
or U2198 (N_2198,N_1720,N_1779);
nor U2199 (N_2199,N_1577,N_1619);
xnor U2200 (N_2200,N_1943,N_1934);
or U2201 (N_2201,N_1937,N_1878);
and U2202 (N_2202,N_1640,N_1957);
or U2203 (N_2203,N_1949,N_1986);
and U2204 (N_2204,N_1554,N_1974);
nor U2205 (N_2205,N_1890,N_1959);
and U2206 (N_2206,N_1569,N_1659);
and U2207 (N_2207,N_1609,N_1675);
and U2208 (N_2208,N_1593,N_1568);
or U2209 (N_2209,N_1939,N_1965);
and U2210 (N_2210,N_1650,N_1562);
or U2211 (N_2211,N_1678,N_1573);
nand U2212 (N_2212,N_1672,N_1902);
or U2213 (N_2213,N_1664,N_1584);
xor U2214 (N_2214,N_1589,N_1683);
and U2215 (N_2215,N_1670,N_1540);
nand U2216 (N_2216,N_1600,N_1870);
and U2217 (N_2217,N_1908,N_1760);
nor U2218 (N_2218,N_1655,N_1621);
xor U2219 (N_2219,N_1931,N_1969);
nand U2220 (N_2220,N_1534,N_1566);
nand U2221 (N_2221,N_1503,N_1644);
and U2222 (N_2222,N_1790,N_1960);
or U2223 (N_2223,N_1546,N_1731);
or U2224 (N_2224,N_1583,N_1772);
nor U2225 (N_2225,N_1992,N_1916);
or U2226 (N_2226,N_1898,N_1725);
and U2227 (N_2227,N_1511,N_1737);
nor U2228 (N_2228,N_1883,N_1545);
xnor U2229 (N_2229,N_1970,N_1845);
or U2230 (N_2230,N_1571,N_1868);
and U2231 (N_2231,N_1840,N_1557);
nor U2232 (N_2232,N_1669,N_1856);
nand U2233 (N_2233,N_1913,N_1535);
and U2234 (N_2234,N_1791,N_1555);
xor U2235 (N_2235,N_1917,N_1920);
nor U2236 (N_2236,N_1871,N_1747);
or U2237 (N_2237,N_1877,N_1590);
and U2238 (N_2238,N_1587,N_1799);
nand U2239 (N_2239,N_1766,N_1674);
nor U2240 (N_2240,N_1774,N_1804);
nand U2241 (N_2241,N_1597,N_1738);
nor U2242 (N_2242,N_1989,N_1972);
and U2243 (N_2243,N_1634,N_1855);
or U2244 (N_2244,N_1523,N_1847);
or U2245 (N_2245,N_1741,N_1958);
or U2246 (N_2246,N_1892,N_1565);
or U2247 (N_2247,N_1780,N_1704);
or U2248 (N_2248,N_1530,N_1952);
nor U2249 (N_2249,N_1830,N_1973);
nor U2250 (N_2250,N_1936,N_1917);
and U2251 (N_2251,N_1914,N_1595);
nor U2252 (N_2252,N_1853,N_1718);
and U2253 (N_2253,N_1634,N_1644);
and U2254 (N_2254,N_1725,N_1737);
nand U2255 (N_2255,N_1525,N_1712);
nand U2256 (N_2256,N_1748,N_1997);
nand U2257 (N_2257,N_1561,N_1797);
nor U2258 (N_2258,N_1918,N_1631);
nand U2259 (N_2259,N_1837,N_1938);
or U2260 (N_2260,N_1688,N_1820);
nand U2261 (N_2261,N_1852,N_1631);
xor U2262 (N_2262,N_1504,N_1537);
and U2263 (N_2263,N_1632,N_1827);
nor U2264 (N_2264,N_1599,N_1555);
or U2265 (N_2265,N_1746,N_1813);
and U2266 (N_2266,N_1973,N_1773);
and U2267 (N_2267,N_1893,N_1621);
or U2268 (N_2268,N_1622,N_1765);
nand U2269 (N_2269,N_1715,N_1745);
nand U2270 (N_2270,N_1761,N_1795);
nand U2271 (N_2271,N_1966,N_1818);
and U2272 (N_2272,N_1884,N_1541);
xor U2273 (N_2273,N_1910,N_1710);
xnor U2274 (N_2274,N_1721,N_1572);
and U2275 (N_2275,N_1942,N_1933);
or U2276 (N_2276,N_1994,N_1873);
and U2277 (N_2277,N_1643,N_1613);
or U2278 (N_2278,N_1976,N_1738);
xor U2279 (N_2279,N_1859,N_1663);
and U2280 (N_2280,N_1686,N_1612);
and U2281 (N_2281,N_1683,N_1884);
nor U2282 (N_2282,N_1842,N_1724);
nor U2283 (N_2283,N_1782,N_1745);
nor U2284 (N_2284,N_1962,N_1855);
nor U2285 (N_2285,N_1929,N_1802);
nor U2286 (N_2286,N_1878,N_1989);
xor U2287 (N_2287,N_1863,N_1592);
and U2288 (N_2288,N_1801,N_1723);
xor U2289 (N_2289,N_1921,N_1793);
xnor U2290 (N_2290,N_1905,N_1953);
nor U2291 (N_2291,N_1786,N_1972);
and U2292 (N_2292,N_1524,N_1931);
nand U2293 (N_2293,N_1695,N_1588);
or U2294 (N_2294,N_1824,N_1831);
or U2295 (N_2295,N_1651,N_1654);
and U2296 (N_2296,N_1594,N_1996);
nor U2297 (N_2297,N_1819,N_1668);
nand U2298 (N_2298,N_1872,N_1940);
nand U2299 (N_2299,N_1544,N_1601);
nand U2300 (N_2300,N_1999,N_1809);
xor U2301 (N_2301,N_1575,N_1602);
and U2302 (N_2302,N_1983,N_1511);
nand U2303 (N_2303,N_1839,N_1761);
nor U2304 (N_2304,N_1644,N_1930);
or U2305 (N_2305,N_1597,N_1895);
or U2306 (N_2306,N_1859,N_1687);
nand U2307 (N_2307,N_1769,N_1840);
nand U2308 (N_2308,N_1882,N_1648);
nand U2309 (N_2309,N_1872,N_1970);
or U2310 (N_2310,N_1519,N_1946);
and U2311 (N_2311,N_1645,N_1896);
or U2312 (N_2312,N_1966,N_1979);
nor U2313 (N_2313,N_1519,N_1634);
nand U2314 (N_2314,N_1634,N_1569);
nand U2315 (N_2315,N_1770,N_1757);
and U2316 (N_2316,N_1844,N_1563);
nor U2317 (N_2317,N_1768,N_1578);
and U2318 (N_2318,N_1695,N_1522);
or U2319 (N_2319,N_1664,N_1546);
or U2320 (N_2320,N_1763,N_1639);
nand U2321 (N_2321,N_1646,N_1727);
or U2322 (N_2322,N_1859,N_1841);
nor U2323 (N_2323,N_1594,N_1927);
or U2324 (N_2324,N_1811,N_1901);
and U2325 (N_2325,N_1575,N_1993);
and U2326 (N_2326,N_1942,N_1909);
nand U2327 (N_2327,N_1925,N_1729);
nor U2328 (N_2328,N_1824,N_1926);
nand U2329 (N_2329,N_1963,N_1528);
or U2330 (N_2330,N_1997,N_1563);
nor U2331 (N_2331,N_1767,N_1994);
xnor U2332 (N_2332,N_1738,N_1675);
or U2333 (N_2333,N_1768,N_1819);
or U2334 (N_2334,N_1578,N_1631);
and U2335 (N_2335,N_1587,N_1610);
and U2336 (N_2336,N_1705,N_1567);
nor U2337 (N_2337,N_1976,N_1946);
nor U2338 (N_2338,N_1762,N_1609);
xnor U2339 (N_2339,N_1578,N_1975);
and U2340 (N_2340,N_1539,N_1763);
or U2341 (N_2341,N_1725,N_1994);
or U2342 (N_2342,N_1929,N_1554);
nand U2343 (N_2343,N_1821,N_1947);
nand U2344 (N_2344,N_1834,N_1545);
xor U2345 (N_2345,N_1917,N_1816);
nor U2346 (N_2346,N_1589,N_1805);
nor U2347 (N_2347,N_1550,N_1782);
or U2348 (N_2348,N_1857,N_1880);
or U2349 (N_2349,N_1971,N_1641);
nand U2350 (N_2350,N_1823,N_1605);
and U2351 (N_2351,N_1536,N_1575);
or U2352 (N_2352,N_1816,N_1932);
and U2353 (N_2353,N_1583,N_1885);
or U2354 (N_2354,N_1796,N_1710);
nor U2355 (N_2355,N_1958,N_1705);
and U2356 (N_2356,N_1654,N_1848);
or U2357 (N_2357,N_1626,N_1957);
or U2358 (N_2358,N_1844,N_1897);
xor U2359 (N_2359,N_1626,N_1625);
and U2360 (N_2360,N_1652,N_1832);
nor U2361 (N_2361,N_1640,N_1816);
or U2362 (N_2362,N_1785,N_1763);
nor U2363 (N_2363,N_1736,N_1516);
and U2364 (N_2364,N_1899,N_1980);
or U2365 (N_2365,N_1622,N_1842);
nand U2366 (N_2366,N_1560,N_1557);
nor U2367 (N_2367,N_1682,N_1892);
nor U2368 (N_2368,N_1548,N_1808);
or U2369 (N_2369,N_1737,N_1907);
nand U2370 (N_2370,N_1620,N_1766);
and U2371 (N_2371,N_1587,N_1940);
and U2372 (N_2372,N_1950,N_1681);
nor U2373 (N_2373,N_1500,N_1578);
or U2374 (N_2374,N_1935,N_1575);
or U2375 (N_2375,N_1570,N_1577);
or U2376 (N_2376,N_1759,N_1965);
or U2377 (N_2377,N_1969,N_1997);
nand U2378 (N_2378,N_1528,N_1536);
and U2379 (N_2379,N_1613,N_1518);
and U2380 (N_2380,N_1953,N_1920);
nor U2381 (N_2381,N_1580,N_1789);
nor U2382 (N_2382,N_1772,N_1519);
nand U2383 (N_2383,N_1962,N_1568);
and U2384 (N_2384,N_1667,N_1614);
and U2385 (N_2385,N_1669,N_1509);
and U2386 (N_2386,N_1647,N_1771);
nor U2387 (N_2387,N_1990,N_1521);
nor U2388 (N_2388,N_1697,N_1943);
nor U2389 (N_2389,N_1641,N_1700);
and U2390 (N_2390,N_1954,N_1861);
and U2391 (N_2391,N_1510,N_1583);
nor U2392 (N_2392,N_1556,N_1902);
nor U2393 (N_2393,N_1849,N_1935);
and U2394 (N_2394,N_1689,N_1896);
nor U2395 (N_2395,N_1567,N_1548);
or U2396 (N_2396,N_1803,N_1511);
or U2397 (N_2397,N_1645,N_1588);
nor U2398 (N_2398,N_1696,N_1763);
nand U2399 (N_2399,N_1938,N_1733);
nor U2400 (N_2400,N_1525,N_1547);
and U2401 (N_2401,N_1849,N_1572);
or U2402 (N_2402,N_1876,N_1852);
or U2403 (N_2403,N_1770,N_1873);
nand U2404 (N_2404,N_1866,N_1569);
nand U2405 (N_2405,N_1725,N_1646);
and U2406 (N_2406,N_1809,N_1681);
xor U2407 (N_2407,N_1605,N_1922);
nand U2408 (N_2408,N_1705,N_1853);
nor U2409 (N_2409,N_1714,N_1855);
and U2410 (N_2410,N_1786,N_1570);
and U2411 (N_2411,N_1530,N_1596);
nor U2412 (N_2412,N_1577,N_1574);
nor U2413 (N_2413,N_1910,N_1720);
or U2414 (N_2414,N_1883,N_1966);
nor U2415 (N_2415,N_1867,N_1635);
xnor U2416 (N_2416,N_1703,N_1684);
and U2417 (N_2417,N_1705,N_1964);
nand U2418 (N_2418,N_1908,N_1634);
nand U2419 (N_2419,N_1780,N_1618);
nor U2420 (N_2420,N_1622,N_1674);
nand U2421 (N_2421,N_1868,N_1997);
nor U2422 (N_2422,N_1876,N_1626);
nor U2423 (N_2423,N_1794,N_1861);
nor U2424 (N_2424,N_1969,N_1955);
or U2425 (N_2425,N_1556,N_1654);
xor U2426 (N_2426,N_1663,N_1651);
xnor U2427 (N_2427,N_1564,N_1984);
nor U2428 (N_2428,N_1509,N_1759);
nand U2429 (N_2429,N_1812,N_1591);
nand U2430 (N_2430,N_1781,N_1543);
or U2431 (N_2431,N_1675,N_1971);
and U2432 (N_2432,N_1540,N_1773);
nor U2433 (N_2433,N_1806,N_1641);
and U2434 (N_2434,N_1889,N_1726);
nor U2435 (N_2435,N_1984,N_1814);
nor U2436 (N_2436,N_1655,N_1809);
and U2437 (N_2437,N_1817,N_1690);
or U2438 (N_2438,N_1537,N_1721);
and U2439 (N_2439,N_1636,N_1992);
nor U2440 (N_2440,N_1929,N_1884);
nand U2441 (N_2441,N_1712,N_1816);
and U2442 (N_2442,N_1836,N_1678);
and U2443 (N_2443,N_1632,N_1644);
nor U2444 (N_2444,N_1674,N_1619);
xor U2445 (N_2445,N_1627,N_1976);
nor U2446 (N_2446,N_1837,N_1874);
and U2447 (N_2447,N_1957,N_1981);
xnor U2448 (N_2448,N_1759,N_1601);
and U2449 (N_2449,N_1683,N_1987);
or U2450 (N_2450,N_1793,N_1934);
or U2451 (N_2451,N_1682,N_1530);
nor U2452 (N_2452,N_1869,N_1963);
xor U2453 (N_2453,N_1766,N_1915);
and U2454 (N_2454,N_1946,N_1935);
nand U2455 (N_2455,N_1608,N_1568);
nand U2456 (N_2456,N_1506,N_1545);
nor U2457 (N_2457,N_1773,N_1944);
or U2458 (N_2458,N_1921,N_1705);
xnor U2459 (N_2459,N_1748,N_1777);
and U2460 (N_2460,N_1594,N_1753);
nand U2461 (N_2461,N_1691,N_1657);
nor U2462 (N_2462,N_1852,N_1702);
xor U2463 (N_2463,N_1848,N_1593);
nand U2464 (N_2464,N_1653,N_1576);
and U2465 (N_2465,N_1820,N_1656);
nand U2466 (N_2466,N_1611,N_1983);
and U2467 (N_2467,N_1783,N_1576);
and U2468 (N_2468,N_1581,N_1901);
and U2469 (N_2469,N_1816,N_1505);
nor U2470 (N_2470,N_1521,N_1687);
or U2471 (N_2471,N_1925,N_1970);
nand U2472 (N_2472,N_1866,N_1832);
nand U2473 (N_2473,N_1588,N_1825);
nor U2474 (N_2474,N_1787,N_1600);
and U2475 (N_2475,N_1655,N_1845);
and U2476 (N_2476,N_1911,N_1661);
or U2477 (N_2477,N_1905,N_1787);
nand U2478 (N_2478,N_1772,N_1639);
xor U2479 (N_2479,N_1876,N_1947);
xnor U2480 (N_2480,N_1917,N_1615);
nor U2481 (N_2481,N_1887,N_1991);
nand U2482 (N_2482,N_1690,N_1694);
and U2483 (N_2483,N_1555,N_1673);
nor U2484 (N_2484,N_1616,N_1897);
nand U2485 (N_2485,N_1747,N_1803);
and U2486 (N_2486,N_1712,N_1739);
xor U2487 (N_2487,N_1753,N_1730);
and U2488 (N_2488,N_1881,N_1602);
and U2489 (N_2489,N_1932,N_1703);
and U2490 (N_2490,N_1804,N_1665);
nand U2491 (N_2491,N_1788,N_1947);
or U2492 (N_2492,N_1783,N_1583);
nor U2493 (N_2493,N_1855,N_1836);
or U2494 (N_2494,N_1859,N_1588);
xnor U2495 (N_2495,N_1804,N_1980);
and U2496 (N_2496,N_1916,N_1675);
or U2497 (N_2497,N_1522,N_1871);
nor U2498 (N_2498,N_1519,N_1919);
nor U2499 (N_2499,N_1539,N_1835);
nand U2500 (N_2500,N_2157,N_2235);
nor U2501 (N_2501,N_2376,N_2102);
xnor U2502 (N_2502,N_2252,N_2399);
xnor U2503 (N_2503,N_2363,N_2429);
and U2504 (N_2504,N_2345,N_2439);
nand U2505 (N_2505,N_2036,N_2428);
xnor U2506 (N_2506,N_2336,N_2198);
and U2507 (N_2507,N_2007,N_2237);
xnor U2508 (N_2508,N_2201,N_2280);
or U2509 (N_2509,N_2440,N_2159);
nor U2510 (N_2510,N_2480,N_2306);
or U2511 (N_2511,N_2355,N_2431);
or U2512 (N_2512,N_2165,N_2340);
nand U2513 (N_2513,N_2073,N_2040);
nand U2514 (N_2514,N_2298,N_2289);
or U2515 (N_2515,N_2461,N_2080);
nor U2516 (N_2516,N_2259,N_2184);
nor U2517 (N_2517,N_2315,N_2227);
nand U2518 (N_2518,N_2197,N_2240);
nand U2519 (N_2519,N_2326,N_2425);
nor U2520 (N_2520,N_2027,N_2116);
or U2521 (N_2521,N_2256,N_2296);
nor U2522 (N_2522,N_2267,N_2416);
or U2523 (N_2523,N_2149,N_2087);
or U2524 (N_2524,N_2152,N_2292);
nor U2525 (N_2525,N_2190,N_2469);
and U2526 (N_2526,N_2049,N_2285);
nor U2527 (N_2527,N_2387,N_2344);
nand U2528 (N_2528,N_2166,N_2290);
or U2529 (N_2529,N_2308,N_2169);
or U2530 (N_2530,N_2111,N_2490);
nor U2531 (N_2531,N_2096,N_2451);
nand U2532 (N_2532,N_2121,N_2449);
or U2533 (N_2533,N_2066,N_2412);
nand U2534 (N_2534,N_2013,N_2448);
nor U2535 (N_2535,N_2444,N_2124);
nor U2536 (N_2536,N_2362,N_2187);
or U2537 (N_2537,N_2372,N_2337);
and U2538 (N_2538,N_2251,N_2052);
xor U2539 (N_2539,N_2411,N_2246);
and U2540 (N_2540,N_2200,N_2413);
or U2541 (N_2541,N_2402,N_2095);
or U2542 (N_2542,N_2309,N_2434);
or U2543 (N_2543,N_2163,N_2433);
and U2544 (N_2544,N_2179,N_2270);
nor U2545 (N_2545,N_2437,N_2488);
nor U2546 (N_2546,N_2286,N_2225);
nor U2547 (N_2547,N_2057,N_2368);
nand U2548 (N_2548,N_2078,N_2325);
nor U2549 (N_2549,N_2247,N_2205);
and U2550 (N_2550,N_2384,N_2317);
nand U2551 (N_2551,N_2091,N_2410);
and U2552 (N_2552,N_2193,N_2024);
nand U2553 (N_2553,N_2349,N_2082);
nor U2554 (N_2554,N_2129,N_2123);
xnor U2555 (N_2555,N_2154,N_2185);
and U2556 (N_2556,N_2168,N_2261);
or U2557 (N_2557,N_2061,N_2011);
nor U2558 (N_2558,N_2138,N_2126);
or U2559 (N_2559,N_2474,N_2183);
nand U2560 (N_2560,N_2253,N_2120);
or U2561 (N_2561,N_2456,N_2357);
and U2562 (N_2562,N_2075,N_2209);
or U2563 (N_2563,N_2400,N_2090);
and U2564 (N_2564,N_2332,N_2142);
and U2565 (N_2565,N_2125,N_2043);
and U2566 (N_2566,N_2093,N_2039);
or U2567 (N_2567,N_2343,N_2374);
xor U2568 (N_2568,N_2471,N_2419);
xnor U2569 (N_2569,N_2486,N_2021);
nand U2570 (N_2570,N_2468,N_2104);
and U2571 (N_2571,N_2359,N_2300);
nor U2572 (N_2572,N_2284,N_2484);
nand U2573 (N_2573,N_2231,N_2063);
nor U2574 (N_2574,N_2318,N_2426);
nand U2575 (N_2575,N_2348,N_2230);
or U2576 (N_2576,N_2312,N_2307);
and U2577 (N_2577,N_2353,N_2242);
or U2578 (N_2578,N_2055,N_2195);
xor U2579 (N_2579,N_2221,N_2268);
and U2580 (N_2580,N_2477,N_2015);
and U2581 (N_2581,N_2208,N_2377);
nand U2582 (N_2582,N_2141,N_2176);
or U2583 (N_2583,N_2281,N_2361);
or U2584 (N_2584,N_2446,N_2432);
nor U2585 (N_2585,N_2178,N_2465);
nand U2586 (N_2586,N_2119,N_2016);
nor U2587 (N_2587,N_2438,N_2406);
or U2588 (N_2588,N_2401,N_2450);
nand U2589 (N_2589,N_2322,N_2459);
or U2590 (N_2590,N_2464,N_2072);
nor U2591 (N_2591,N_2112,N_2238);
or U2592 (N_2592,N_2070,N_2143);
and U2593 (N_2593,N_2354,N_2350);
or U2594 (N_2594,N_2455,N_2042);
nand U2595 (N_2595,N_2222,N_2033);
and U2596 (N_2596,N_2127,N_2422);
xnor U2597 (N_2597,N_2279,N_2475);
nand U2598 (N_2598,N_2321,N_2050);
nand U2599 (N_2599,N_2071,N_2229);
or U2600 (N_2600,N_2458,N_2180);
nand U2601 (N_2601,N_2232,N_2145);
or U2602 (N_2602,N_2482,N_2099);
xor U2603 (N_2603,N_2473,N_2053);
or U2604 (N_2604,N_2398,N_2162);
and U2605 (N_2605,N_2092,N_2012);
and U2606 (N_2606,N_2217,N_2058);
or U2607 (N_2607,N_2498,N_2020);
nor U2608 (N_2608,N_2276,N_2283);
xnor U2609 (N_2609,N_2008,N_2316);
nor U2610 (N_2610,N_2250,N_2172);
and U2611 (N_2611,N_2088,N_2311);
or U2612 (N_2612,N_2103,N_2329);
and U2613 (N_2613,N_2424,N_2136);
and U2614 (N_2614,N_2206,N_2351);
xor U2615 (N_2615,N_2454,N_2463);
or U2616 (N_2616,N_2364,N_2192);
nor U2617 (N_2617,N_2175,N_2441);
nor U2618 (N_2618,N_2202,N_2327);
or U2619 (N_2619,N_2241,N_2009);
nor U2620 (N_2620,N_2499,N_2305);
nor U2621 (N_2621,N_2028,N_2097);
and U2622 (N_2622,N_2489,N_2153);
and U2623 (N_2623,N_2100,N_2128);
nor U2624 (N_2624,N_2245,N_2224);
nand U2625 (N_2625,N_2436,N_2487);
nor U2626 (N_2626,N_2442,N_2274);
xor U2627 (N_2627,N_2101,N_2333);
nand U2628 (N_2628,N_2000,N_2233);
nand U2629 (N_2629,N_2265,N_2358);
and U2630 (N_2630,N_2134,N_2151);
nand U2631 (N_2631,N_2094,N_2470);
or U2632 (N_2632,N_2135,N_2110);
or U2633 (N_2633,N_2453,N_2220);
nand U2634 (N_2634,N_2388,N_2271);
or U2635 (N_2635,N_2383,N_2079);
and U2636 (N_2636,N_2435,N_2034);
and U2637 (N_2637,N_2059,N_2223);
nor U2638 (N_2638,N_2288,N_2177);
or U2639 (N_2639,N_2334,N_2244);
nor U2640 (N_2640,N_2207,N_2031);
and U2641 (N_2641,N_2338,N_2320);
nor U2642 (N_2642,N_2018,N_2356);
nand U2643 (N_2643,N_2483,N_2109);
nand U2644 (N_2644,N_2047,N_2467);
and U2645 (N_2645,N_2065,N_2133);
or U2646 (N_2646,N_2239,N_2131);
nor U2647 (N_2647,N_2216,N_2466);
nor U2648 (N_2648,N_2485,N_2328);
xnor U2649 (N_2649,N_2452,N_2081);
or U2650 (N_2650,N_2367,N_2346);
nand U2651 (N_2651,N_2254,N_2460);
and U2652 (N_2652,N_2404,N_2248);
or U2653 (N_2653,N_2150,N_2076);
and U2654 (N_2654,N_2130,N_2392);
nor U2655 (N_2655,N_2017,N_2067);
or U2656 (N_2656,N_2215,N_2226);
or U2657 (N_2657,N_2045,N_2107);
xnor U2658 (N_2658,N_2415,N_2194);
or U2659 (N_2659,N_2046,N_2409);
nand U2660 (N_2660,N_2375,N_2331);
or U2661 (N_2661,N_2382,N_2385);
nor U2662 (N_2662,N_2196,N_2472);
nand U2663 (N_2663,N_2118,N_2029);
and U2664 (N_2664,N_2041,N_2405);
or U2665 (N_2665,N_2077,N_2211);
or U2666 (N_2666,N_2089,N_2443);
and U2667 (N_2667,N_2051,N_2064);
nor U2668 (N_2668,N_2407,N_2295);
nand U2669 (N_2669,N_2114,N_2257);
and U2670 (N_2670,N_2294,N_2023);
and U2671 (N_2671,N_2156,N_2003);
nor U2672 (N_2672,N_2174,N_2117);
nand U2673 (N_2673,N_2098,N_2005);
nor U2674 (N_2674,N_2026,N_2319);
and U2675 (N_2675,N_2113,N_2234);
xor U2676 (N_2676,N_2173,N_2379);
nor U2677 (N_2677,N_2418,N_2054);
nor U2678 (N_2678,N_2373,N_2275);
or U2679 (N_2679,N_2105,N_2293);
or U2680 (N_2680,N_2161,N_2074);
nor U2681 (N_2681,N_2203,N_2006);
nor U2682 (N_2682,N_2277,N_2212);
nor U2683 (N_2683,N_2427,N_2370);
or U2684 (N_2684,N_2144,N_2030);
or U2685 (N_2685,N_2365,N_2420);
nor U2686 (N_2686,N_2236,N_2210);
nand U2687 (N_2687,N_2085,N_2323);
or U2688 (N_2688,N_2299,N_2360);
and U2689 (N_2689,N_2214,N_2164);
nand U2690 (N_2690,N_2313,N_2297);
or U2691 (N_2691,N_2056,N_2430);
nor U2692 (N_2692,N_2394,N_2494);
or U2693 (N_2693,N_2260,N_2403);
and U2694 (N_2694,N_2019,N_2417);
and U2695 (N_2695,N_2495,N_2032);
nor U2696 (N_2696,N_2335,N_2038);
and U2697 (N_2697,N_2068,N_2170);
and U2698 (N_2698,N_2330,N_2457);
or U2699 (N_2699,N_2423,N_2002);
or U2700 (N_2700,N_2035,N_2263);
xnor U2701 (N_2701,N_2395,N_2025);
nor U2702 (N_2702,N_2083,N_2266);
and U2703 (N_2703,N_2369,N_2218);
nand U2704 (N_2704,N_2269,N_2122);
nand U2705 (N_2705,N_2302,N_2462);
xor U2706 (N_2706,N_2160,N_2137);
nand U2707 (N_2707,N_2132,N_2347);
and U2708 (N_2708,N_2243,N_2479);
or U2709 (N_2709,N_2037,N_2140);
or U2710 (N_2710,N_2199,N_2148);
xnor U2711 (N_2711,N_2108,N_2167);
nor U2712 (N_2712,N_2010,N_2291);
nor U2713 (N_2713,N_2155,N_2146);
xor U2714 (N_2714,N_2397,N_2278);
xor U2715 (N_2715,N_2171,N_2393);
nand U2716 (N_2716,N_2492,N_2390);
and U2717 (N_2717,N_2062,N_2342);
nand U2718 (N_2718,N_2371,N_2408);
xnor U2719 (N_2719,N_2249,N_2158);
or U2720 (N_2720,N_2022,N_2228);
or U2721 (N_2721,N_2421,N_2324);
and U2722 (N_2722,N_2389,N_2447);
or U2723 (N_2723,N_2380,N_2476);
and U2724 (N_2724,N_2004,N_2219);
or U2725 (N_2725,N_2414,N_2304);
nor U2726 (N_2726,N_2341,N_2491);
or U2727 (N_2727,N_2381,N_2272);
xnor U2728 (N_2728,N_2181,N_2314);
or U2729 (N_2729,N_2106,N_2001);
nand U2730 (N_2730,N_2255,N_2396);
and U2731 (N_2731,N_2115,N_2258);
and U2732 (N_2732,N_2182,N_2014);
nand U2733 (N_2733,N_2386,N_2497);
nand U2734 (N_2734,N_2044,N_2352);
nand U2735 (N_2735,N_2264,N_2084);
nor U2736 (N_2736,N_2478,N_2282);
nand U2737 (N_2737,N_2189,N_2391);
nand U2738 (N_2738,N_2191,N_2139);
nor U2739 (N_2739,N_2186,N_2287);
and U2740 (N_2740,N_2496,N_2366);
xor U2741 (N_2741,N_2481,N_2048);
and U2742 (N_2742,N_2213,N_2069);
and U2743 (N_2743,N_2188,N_2378);
nor U2744 (N_2744,N_2310,N_2204);
and U2745 (N_2745,N_2339,N_2147);
nand U2746 (N_2746,N_2262,N_2445);
nor U2747 (N_2747,N_2060,N_2493);
or U2748 (N_2748,N_2086,N_2273);
and U2749 (N_2749,N_2303,N_2301);
xor U2750 (N_2750,N_2261,N_2039);
nand U2751 (N_2751,N_2419,N_2279);
xor U2752 (N_2752,N_2329,N_2391);
or U2753 (N_2753,N_2256,N_2272);
nor U2754 (N_2754,N_2276,N_2105);
nor U2755 (N_2755,N_2191,N_2315);
xnor U2756 (N_2756,N_2132,N_2454);
nand U2757 (N_2757,N_2116,N_2445);
xor U2758 (N_2758,N_2450,N_2274);
or U2759 (N_2759,N_2304,N_2352);
nor U2760 (N_2760,N_2424,N_2161);
nor U2761 (N_2761,N_2181,N_2329);
nor U2762 (N_2762,N_2032,N_2390);
or U2763 (N_2763,N_2060,N_2348);
nor U2764 (N_2764,N_2374,N_2331);
or U2765 (N_2765,N_2115,N_2068);
or U2766 (N_2766,N_2483,N_2267);
nor U2767 (N_2767,N_2017,N_2088);
and U2768 (N_2768,N_2200,N_2092);
and U2769 (N_2769,N_2091,N_2011);
nand U2770 (N_2770,N_2051,N_2445);
nor U2771 (N_2771,N_2449,N_2358);
or U2772 (N_2772,N_2154,N_2359);
xnor U2773 (N_2773,N_2216,N_2256);
and U2774 (N_2774,N_2340,N_2287);
or U2775 (N_2775,N_2081,N_2113);
nand U2776 (N_2776,N_2180,N_2173);
or U2777 (N_2777,N_2084,N_2353);
nand U2778 (N_2778,N_2099,N_2421);
xnor U2779 (N_2779,N_2392,N_2136);
nand U2780 (N_2780,N_2149,N_2335);
xor U2781 (N_2781,N_2445,N_2490);
nor U2782 (N_2782,N_2020,N_2142);
or U2783 (N_2783,N_2187,N_2320);
nor U2784 (N_2784,N_2015,N_2455);
nand U2785 (N_2785,N_2002,N_2097);
nor U2786 (N_2786,N_2398,N_2419);
nand U2787 (N_2787,N_2375,N_2002);
or U2788 (N_2788,N_2038,N_2276);
nand U2789 (N_2789,N_2030,N_2452);
nor U2790 (N_2790,N_2193,N_2492);
nand U2791 (N_2791,N_2362,N_2307);
and U2792 (N_2792,N_2183,N_2493);
nand U2793 (N_2793,N_2025,N_2086);
nor U2794 (N_2794,N_2260,N_2208);
and U2795 (N_2795,N_2491,N_2261);
nor U2796 (N_2796,N_2292,N_2169);
nor U2797 (N_2797,N_2391,N_2468);
or U2798 (N_2798,N_2421,N_2299);
nor U2799 (N_2799,N_2301,N_2014);
nor U2800 (N_2800,N_2350,N_2340);
xor U2801 (N_2801,N_2394,N_2345);
or U2802 (N_2802,N_2289,N_2045);
and U2803 (N_2803,N_2011,N_2268);
or U2804 (N_2804,N_2352,N_2238);
nor U2805 (N_2805,N_2395,N_2157);
and U2806 (N_2806,N_2151,N_2150);
or U2807 (N_2807,N_2056,N_2103);
or U2808 (N_2808,N_2253,N_2143);
nand U2809 (N_2809,N_2486,N_2459);
nor U2810 (N_2810,N_2479,N_2330);
nor U2811 (N_2811,N_2046,N_2429);
xor U2812 (N_2812,N_2277,N_2297);
nand U2813 (N_2813,N_2420,N_2142);
nor U2814 (N_2814,N_2268,N_2316);
and U2815 (N_2815,N_2126,N_2345);
nand U2816 (N_2816,N_2441,N_2404);
nand U2817 (N_2817,N_2016,N_2401);
nand U2818 (N_2818,N_2297,N_2453);
nor U2819 (N_2819,N_2243,N_2304);
nand U2820 (N_2820,N_2147,N_2493);
and U2821 (N_2821,N_2064,N_2467);
nor U2822 (N_2822,N_2360,N_2289);
and U2823 (N_2823,N_2353,N_2339);
nand U2824 (N_2824,N_2098,N_2266);
nand U2825 (N_2825,N_2280,N_2271);
nor U2826 (N_2826,N_2132,N_2155);
nand U2827 (N_2827,N_2360,N_2140);
nor U2828 (N_2828,N_2084,N_2109);
nor U2829 (N_2829,N_2020,N_2051);
nand U2830 (N_2830,N_2430,N_2493);
nand U2831 (N_2831,N_2330,N_2360);
nand U2832 (N_2832,N_2184,N_2461);
or U2833 (N_2833,N_2060,N_2186);
or U2834 (N_2834,N_2346,N_2393);
nor U2835 (N_2835,N_2149,N_2294);
nand U2836 (N_2836,N_2102,N_2094);
nor U2837 (N_2837,N_2231,N_2492);
and U2838 (N_2838,N_2101,N_2487);
or U2839 (N_2839,N_2370,N_2130);
and U2840 (N_2840,N_2291,N_2495);
nand U2841 (N_2841,N_2248,N_2026);
and U2842 (N_2842,N_2403,N_2473);
xnor U2843 (N_2843,N_2470,N_2271);
nor U2844 (N_2844,N_2211,N_2285);
nor U2845 (N_2845,N_2050,N_2478);
nand U2846 (N_2846,N_2316,N_2431);
nor U2847 (N_2847,N_2180,N_2165);
and U2848 (N_2848,N_2031,N_2465);
and U2849 (N_2849,N_2266,N_2323);
nand U2850 (N_2850,N_2002,N_2213);
or U2851 (N_2851,N_2022,N_2447);
or U2852 (N_2852,N_2252,N_2456);
nand U2853 (N_2853,N_2243,N_2199);
nor U2854 (N_2854,N_2453,N_2022);
nand U2855 (N_2855,N_2247,N_2307);
or U2856 (N_2856,N_2178,N_2065);
nand U2857 (N_2857,N_2093,N_2476);
nor U2858 (N_2858,N_2091,N_2157);
nor U2859 (N_2859,N_2423,N_2201);
nor U2860 (N_2860,N_2290,N_2486);
and U2861 (N_2861,N_2209,N_2316);
and U2862 (N_2862,N_2296,N_2365);
nand U2863 (N_2863,N_2453,N_2145);
or U2864 (N_2864,N_2136,N_2404);
nand U2865 (N_2865,N_2185,N_2125);
nor U2866 (N_2866,N_2059,N_2347);
nand U2867 (N_2867,N_2262,N_2347);
nand U2868 (N_2868,N_2340,N_2086);
or U2869 (N_2869,N_2495,N_2473);
or U2870 (N_2870,N_2418,N_2238);
nor U2871 (N_2871,N_2109,N_2195);
or U2872 (N_2872,N_2090,N_2073);
and U2873 (N_2873,N_2140,N_2163);
nor U2874 (N_2874,N_2274,N_2000);
and U2875 (N_2875,N_2346,N_2279);
and U2876 (N_2876,N_2480,N_2213);
xor U2877 (N_2877,N_2178,N_2125);
nor U2878 (N_2878,N_2385,N_2208);
or U2879 (N_2879,N_2248,N_2282);
nor U2880 (N_2880,N_2098,N_2398);
nand U2881 (N_2881,N_2471,N_2079);
nor U2882 (N_2882,N_2369,N_2197);
and U2883 (N_2883,N_2073,N_2048);
nand U2884 (N_2884,N_2488,N_2481);
or U2885 (N_2885,N_2048,N_2071);
nand U2886 (N_2886,N_2201,N_2246);
nor U2887 (N_2887,N_2067,N_2499);
nor U2888 (N_2888,N_2030,N_2312);
or U2889 (N_2889,N_2077,N_2494);
or U2890 (N_2890,N_2050,N_2253);
or U2891 (N_2891,N_2329,N_2485);
nor U2892 (N_2892,N_2274,N_2191);
nand U2893 (N_2893,N_2001,N_2032);
nor U2894 (N_2894,N_2283,N_2446);
xor U2895 (N_2895,N_2273,N_2061);
xnor U2896 (N_2896,N_2223,N_2277);
or U2897 (N_2897,N_2433,N_2360);
nand U2898 (N_2898,N_2009,N_2276);
xor U2899 (N_2899,N_2431,N_2058);
xnor U2900 (N_2900,N_2218,N_2239);
nand U2901 (N_2901,N_2073,N_2468);
nand U2902 (N_2902,N_2170,N_2317);
nor U2903 (N_2903,N_2085,N_2083);
nor U2904 (N_2904,N_2187,N_2218);
and U2905 (N_2905,N_2314,N_2367);
or U2906 (N_2906,N_2485,N_2389);
nand U2907 (N_2907,N_2453,N_2304);
or U2908 (N_2908,N_2393,N_2326);
nand U2909 (N_2909,N_2347,N_2062);
and U2910 (N_2910,N_2087,N_2384);
and U2911 (N_2911,N_2161,N_2433);
and U2912 (N_2912,N_2402,N_2335);
nand U2913 (N_2913,N_2144,N_2443);
xnor U2914 (N_2914,N_2128,N_2211);
and U2915 (N_2915,N_2499,N_2450);
nand U2916 (N_2916,N_2000,N_2117);
or U2917 (N_2917,N_2101,N_2370);
and U2918 (N_2918,N_2048,N_2197);
and U2919 (N_2919,N_2196,N_2056);
and U2920 (N_2920,N_2408,N_2283);
nor U2921 (N_2921,N_2311,N_2182);
nor U2922 (N_2922,N_2400,N_2083);
and U2923 (N_2923,N_2041,N_2039);
or U2924 (N_2924,N_2440,N_2040);
nor U2925 (N_2925,N_2397,N_2107);
nor U2926 (N_2926,N_2294,N_2107);
or U2927 (N_2927,N_2462,N_2230);
xor U2928 (N_2928,N_2126,N_2144);
nor U2929 (N_2929,N_2069,N_2470);
nand U2930 (N_2930,N_2361,N_2079);
or U2931 (N_2931,N_2354,N_2424);
and U2932 (N_2932,N_2356,N_2350);
and U2933 (N_2933,N_2292,N_2223);
nand U2934 (N_2934,N_2134,N_2479);
nand U2935 (N_2935,N_2072,N_2121);
xor U2936 (N_2936,N_2130,N_2090);
nor U2937 (N_2937,N_2451,N_2075);
and U2938 (N_2938,N_2063,N_2460);
nor U2939 (N_2939,N_2217,N_2462);
nor U2940 (N_2940,N_2226,N_2484);
and U2941 (N_2941,N_2317,N_2040);
nor U2942 (N_2942,N_2257,N_2211);
and U2943 (N_2943,N_2062,N_2202);
and U2944 (N_2944,N_2370,N_2335);
nand U2945 (N_2945,N_2433,N_2007);
and U2946 (N_2946,N_2085,N_2112);
nor U2947 (N_2947,N_2309,N_2112);
nand U2948 (N_2948,N_2494,N_2191);
xnor U2949 (N_2949,N_2461,N_2031);
nor U2950 (N_2950,N_2317,N_2061);
and U2951 (N_2951,N_2347,N_2310);
and U2952 (N_2952,N_2236,N_2459);
and U2953 (N_2953,N_2398,N_2139);
and U2954 (N_2954,N_2488,N_2429);
xor U2955 (N_2955,N_2167,N_2078);
or U2956 (N_2956,N_2332,N_2467);
and U2957 (N_2957,N_2164,N_2216);
nor U2958 (N_2958,N_2332,N_2263);
xor U2959 (N_2959,N_2209,N_2438);
nand U2960 (N_2960,N_2433,N_2119);
or U2961 (N_2961,N_2013,N_2154);
nand U2962 (N_2962,N_2031,N_2170);
nand U2963 (N_2963,N_2136,N_2360);
nand U2964 (N_2964,N_2495,N_2188);
nor U2965 (N_2965,N_2164,N_2273);
and U2966 (N_2966,N_2343,N_2353);
or U2967 (N_2967,N_2465,N_2421);
or U2968 (N_2968,N_2404,N_2436);
nor U2969 (N_2969,N_2451,N_2192);
xor U2970 (N_2970,N_2025,N_2413);
or U2971 (N_2971,N_2285,N_2411);
nand U2972 (N_2972,N_2090,N_2196);
xnor U2973 (N_2973,N_2063,N_2005);
nor U2974 (N_2974,N_2097,N_2324);
nor U2975 (N_2975,N_2394,N_2471);
and U2976 (N_2976,N_2029,N_2115);
and U2977 (N_2977,N_2054,N_2437);
and U2978 (N_2978,N_2180,N_2050);
nor U2979 (N_2979,N_2148,N_2376);
and U2980 (N_2980,N_2342,N_2335);
and U2981 (N_2981,N_2184,N_2110);
xor U2982 (N_2982,N_2387,N_2040);
and U2983 (N_2983,N_2030,N_2371);
nand U2984 (N_2984,N_2336,N_2234);
nand U2985 (N_2985,N_2274,N_2323);
and U2986 (N_2986,N_2020,N_2266);
or U2987 (N_2987,N_2404,N_2323);
or U2988 (N_2988,N_2442,N_2456);
or U2989 (N_2989,N_2245,N_2153);
nand U2990 (N_2990,N_2420,N_2239);
or U2991 (N_2991,N_2076,N_2352);
nor U2992 (N_2992,N_2243,N_2458);
and U2993 (N_2993,N_2305,N_2282);
nor U2994 (N_2994,N_2467,N_2096);
nor U2995 (N_2995,N_2449,N_2205);
or U2996 (N_2996,N_2140,N_2227);
nand U2997 (N_2997,N_2199,N_2086);
or U2998 (N_2998,N_2363,N_2477);
nand U2999 (N_2999,N_2257,N_2197);
and UO_0 (O_0,N_2788,N_2904);
and UO_1 (O_1,N_2551,N_2623);
or UO_2 (O_2,N_2800,N_2545);
nand UO_3 (O_3,N_2794,N_2726);
nand UO_4 (O_4,N_2635,N_2677);
nand UO_5 (O_5,N_2956,N_2928);
or UO_6 (O_6,N_2652,N_2695);
nand UO_7 (O_7,N_2768,N_2560);
nand UO_8 (O_8,N_2508,N_2621);
or UO_9 (O_9,N_2611,N_2507);
nor UO_10 (O_10,N_2633,N_2616);
nor UO_11 (O_11,N_2741,N_2592);
nand UO_12 (O_12,N_2893,N_2841);
nor UO_13 (O_13,N_2713,N_2853);
or UO_14 (O_14,N_2737,N_2645);
nor UO_15 (O_15,N_2825,N_2564);
nor UO_16 (O_16,N_2784,N_2979);
and UO_17 (O_17,N_2786,N_2872);
nand UO_18 (O_18,N_2743,N_2546);
nor UO_19 (O_19,N_2550,N_2969);
or UO_20 (O_20,N_2992,N_2984);
nor UO_21 (O_21,N_2803,N_2535);
nor UO_22 (O_22,N_2547,N_2703);
nand UO_23 (O_23,N_2888,N_2603);
nand UO_24 (O_24,N_2601,N_2589);
xnor UO_25 (O_25,N_2859,N_2763);
nand UO_26 (O_26,N_2765,N_2752);
or UO_27 (O_27,N_2674,N_2529);
or UO_28 (O_28,N_2938,N_2689);
nand UO_29 (O_29,N_2697,N_2530);
xnor UO_30 (O_30,N_2563,N_2663);
and UO_31 (O_31,N_2681,N_2837);
nor UO_32 (O_32,N_2577,N_2821);
xor UO_33 (O_33,N_2540,N_2990);
nand UO_34 (O_34,N_2570,N_2690);
and UO_35 (O_35,N_2785,N_2501);
or UO_36 (O_36,N_2658,N_2636);
xor UO_37 (O_37,N_2933,N_2682);
and UO_38 (O_38,N_2554,N_2917);
nand UO_39 (O_39,N_2744,N_2526);
nor UO_40 (O_40,N_2583,N_2850);
nor UO_41 (O_41,N_2802,N_2897);
or UO_42 (O_42,N_2811,N_2885);
or UO_43 (O_43,N_2804,N_2653);
nor UO_44 (O_44,N_2980,N_2909);
nor UO_45 (O_45,N_2707,N_2659);
and UO_46 (O_46,N_2826,N_2597);
nand UO_47 (O_47,N_2721,N_2698);
and UO_48 (O_48,N_2945,N_2940);
nand UO_49 (O_49,N_2637,N_2534);
nand UO_50 (O_50,N_2762,N_2555);
nor UO_51 (O_51,N_2858,N_2617);
nand UO_52 (O_52,N_2848,N_2830);
nand UO_53 (O_53,N_2694,N_2873);
xor UO_54 (O_54,N_2751,N_2502);
nor UO_55 (O_55,N_2731,N_2774);
and UO_56 (O_56,N_2632,N_2947);
nor UO_57 (O_57,N_2609,N_2553);
nor UO_58 (O_58,N_2884,N_2516);
nor UO_59 (O_59,N_2571,N_2683);
nand UO_60 (O_60,N_2651,N_2576);
nor UO_61 (O_61,N_2913,N_2871);
nand UO_62 (O_62,N_2930,N_2996);
xor UO_63 (O_63,N_2522,N_2919);
or UO_64 (O_64,N_2720,N_2728);
nand UO_65 (O_65,N_2900,N_2886);
or UO_66 (O_66,N_2775,N_2590);
nor UO_67 (O_67,N_2839,N_2523);
and UO_68 (O_68,N_2738,N_2657);
or UO_69 (O_69,N_2916,N_2567);
or UO_70 (O_70,N_2787,N_2876);
nor UO_71 (O_71,N_2833,N_2898);
or UO_72 (O_72,N_2953,N_2532);
and UO_73 (O_73,N_2753,N_2899);
xor UO_74 (O_74,N_2520,N_2745);
nor UO_75 (O_75,N_2505,N_2757);
or UO_76 (O_76,N_2875,N_2754);
nor UO_77 (O_77,N_2701,N_2895);
or UO_78 (O_78,N_2602,N_2974);
and UO_79 (O_79,N_2951,N_2747);
nor UO_80 (O_80,N_2691,N_2963);
nand UO_81 (O_81,N_2678,N_2870);
nand UO_82 (O_82,N_2783,N_2869);
nor UO_83 (O_83,N_2629,N_2882);
or UO_84 (O_84,N_2912,N_2740);
nor UO_85 (O_85,N_2539,N_2574);
nor UO_86 (O_86,N_2982,N_2842);
and UO_87 (O_87,N_2634,N_2997);
nand UO_88 (O_88,N_2661,N_2920);
nand UO_89 (O_89,N_2662,N_2665);
and UO_90 (O_90,N_2906,N_2795);
or UO_91 (O_91,N_2509,N_2939);
or UO_92 (O_92,N_2999,N_2816);
or UO_93 (O_93,N_2558,N_2927);
or UO_94 (O_94,N_2926,N_2705);
and UO_95 (O_95,N_2618,N_2518);
and UO_96 (O_96,N_2855,N_2950);
xnor UO_97 (O_97,N_2668,N_2856);
and UO_98 (O_98,N_2536,N_2552);
or UO_99 (O_99,N_2820,N_2852);
or UO_100 (O_100,N_2638,N_2865);
nor UO_101 (O_101,N_2966,N_2500);
nand UO_102 (O_102,N_2646,N_2687);
nor UO_103 (O_103,N_2866,N_2727);
nor UO_104 (O_104,N_2828,N_2702);
nand UO_105 (O_105,N_2660,N_2595);
or UO_106 (O_106,N_2860,N_2610);
xnor UO_107 (O_107,N_2991,N_2798);
nand UO_108 (O_108,N_2769,N_2766);
or UO_109 (O_109,N_2801,N_2868);
xor UO_110 (O_110,N_2511,N_2676);
nor UO_111 (O_111,N_2575,N_2749);
nor UO_112 (O_112,N_2598,N_2704);
nor UO_113 (O_113,N_2708,N_2722);
or UO_114 (O_114,N_2932,N_2929);
and UO_115 (O_115,N_2957,N_2877);
or UO_116 (O_116,N_2515,N_2620);
xor UO_117 (O_117,N_2983,N_2504);
and UO_118 (O_118,N_2524,N_2993);
and UO_119 (O_119,N_2847,N_2773);
nand UO_120 (O_120,N_2883,N_2572);
nor UO_121 (O_121,N_2867,N_2619);
nor UO_122 (O_122,N_2580,N_2594);
nand UO_123 (O_123,N_2541,N_2622);
or UO_124 (O_124,N_2650,N_2914);
nand UO_125 (O_125,N_2792,N_2759);
or UO_126 (O_126,N_2832,N_2890);
nand UO_127 (O_127,N_2767,N_2606);
and UO_128 (O_128,N_2835,N_2559);
and UO_129 (O_129,N_2735,N_2994);
or UO_130 (O_130,N_2600,N_2986);
xnor UO_131 (O_131,N_2964,N_2975);
and UO_132 (O_132,N_2605,N_2686);
xor UO_133 (O_133,N_2840,N_2946);
nor UO_134 (O_134,N_2521,N_2542);
nand UO_135 (O_135,N_2718,N_2874);
and UO_136 (O_136,N_2760,N_2985);
xnor UO_137 (O_137,N_2781,N_2723);
nor UO_138 (O_138,N_2626,N_2696);
xor UO_139 (O_139,N_2584,N_2528);
nand UO_140 (O_140,N_2503,N_2931);
nor UO_141 (O_141,N_2711,N_2815);
xnor UO_142 (O_142,N_2981,N_2758);
or UO_143 (O_143,N_2812,N_2608);
and UO_144 (O_144,N_2565,N_2965);
nor UO_145 (O_145,N_2648,N_2878);
nand UO_146 (O_146,N_2976,N_2544);
or UO_147 (O_147,N_2789,N_2513);
or UO_148 (O_148,N_2892,N_2586);
or UO_149 (O_149,N_2908,N_2556);
xnor UO_150 (O_150,N_2714,N_2710);
nand UO_151 (O_151,N_2799,N_2607);
or UO_152 (O_152,N_2669,N_2829);
nand UO_153 (O_153,N_2962,N_2693);
nand UO_154 (O_154,N_2822,N_2922);
and UO_155 (O_155,N_2948,N_2771);
nand UO_156 (O_156,N_2548,N_2814);
nor UO_157 (O_157,N_2543,N_2639);
nand UO_158 (O_158,N_2666,N_2562);
nor UO_159 (O_159,N_2902,N_2649);
xnor UO_160 (O_160,N_2664,N_2973);
nor UO_161 (O_161,N_2712,N_2887);
and UO_162 (O_162,N_2818,N_2627);
and UO_163 (O_163,N_2844,N_2671);
and UO_164 (O_164,N_2889,N_2823);
and UO_165 (O_165,N_2700,N_2717);
or UO_166 (O_166,N_2755,N_2612);
xor UO_167 (O_167,N_2961,N_2578);
or UO_168 (O_168,N_2864,N_2734);
nor UO_169 (O_169,N_2863,N_2851);
or UO_170 (O_170,N_2761,N_2949);
or UO_171 (O_171,N_2924,N_2512);
or UO_172 (O_172,N_2831,N_2777);
and UO_173 (O_173,N_2579,N_2959);
xor UO_174 (O_174,N_2903,N_2624);
and UO_175 (O_175,N_2819,N_2506);
or UO_176 (O_176,N_2538,N_2631);
and UO_177 (O_177,N_2736,N_2834);
or UO_178 (O_178,N_2960,N_2625);
or UO_179 (O_179,N_2921,N_2630);
and UO_180 (O_180,N_2937,N_2925);
nand UO_181 (O_181,N_2673,N_2778);
nand UO_182 (O_182,N_2549,N_2854);
and UO_183 (O_183,N_2881,N_2656);
nand UO_184 (O_184,N_2644,N_2750);
nor UO_185 (O_185,N_2796,N_2846);
and UO_186 (O_186,N_2880,N_2699);
or UO_187 (O_187,N_2776,N_2813);
xor UO_188 (O_188,N_2911,N_2510);
and UO_189 (O_189,N_2587,N_2978);
xor UO_190 (O_190,N_2581,N_2967);
and UO_191 (O_191,N_2954,N_2805);
and UO_192 (O_192,N_2514,N_2614);
nor UO_193 (O_193,N_2655,N_2977);
and UO_194 (O_194,N_2642,N_2680);
and UO_195 (O_195,N_2790,N_2843);
nand UO_196 (O_196,N_2585,N_2599);
and UO_197 (O_197,N_2596,N_2810);
nand UO_198 (O_198,N_2739,N_2780);
or UO_199 (O_199,N_2910,N_2593);
nor UO_200 (O_200,N_2943,N_2688);
xnor UO_201 (O_201,N_2641,N_2746);
nor UO_202 (O_202,N_2557,N_2517);
nand UO_203 (O_203,N_2952,N_2849);
nand UO_204 (O_204,N_2807,N_2838);
and UO_205 (O_205,N_2706,N_2654);
nand UO_206 (O_206,N_2845,N_2782);
nor UO_207 (O_207,N_2923,N_2742);
or UO_208 (O_208,N_2675,N_2817);
nand UO_209 (O_209,N_2729,N_2685);
nand UO_210 (O_210,N_2862,N_2941);
or UO_211 (O_211,N_2779,N_2566);
or UO_212 (O_212,N_2915,N_2748);
nor UO_213 (O_213,N_2894,N_2809);
nand UO_214 (O_214,N_2667,N_2568);
nand UO_215 (O_215,N_2525,N_2679);
or UO_216 (O_216,N_2861,N_2643);
nand UO_217 (O_217,N_2537,N_2907);
nor UO_218 (O_218,N_2519,N_2733);
nand UO_219 (O_219,N_2808,N_2716);
or UO_220 (O_220,N_2527,N_2971);
nand UO_221 (O_221,N_2955,N_2857);
and UO_222 (O_222,N_2756,N_2934);
nor UO_223 (O_223,N_2824,N_2588);
nor UO_224 (O_224,N_2942,N_2918);
nor UO_225 (O_225,N_2647,N_2640);
nor UO_226 (O_226,N_2604,N_2561);
or UO_227 (O_227,N_2970,N_2998);
nand UO_228 (O_228,N_2901,N_2732);
or UO_229 (O_229,N_2772,N_2531);
or UO_230 (O_230,N_2672,N_2715);
nand UO_231 (O_231,N_2764,N_2944);
and UO_232 (O_232,N_2972,N_2935);
nand UO_233 (O_233,N_2724,N_2770);
nor UO_234 (O_234,N_2896,N_2573);
nor UO_235 (O_235,N_2827,N_2879);
or UO_236 (O_236,N_2615,N_2793);
and UO_237 (O_237,N_2936,N_2989);
nor UO_238 (O_238,N_2968,N_2613);
xnor UO_239 (O_239,N_2836,N_2958);
and UO_240 (O_240,N_2905,N_2891);
nand UO_241 (O_241,N_2709,N_2725);
nor UO_242 (O_242,N_2995,N_2791);
xor UO_243 (O_243,N_2670,N_2987);
and UO_244 (O_244,N_2684,N_2797);
or UO_245 (O_245,N_2591,N_2628);
and UO_246 (O_246,N_2988,N_2719);
nor UO_247 (O_247,N_2692,N_2730);
xnor UO_248 (O_248,N_2569,N_2533);
nor UO_249 (O_249,N_2582,N_2806);
xnor UO_250 (O_250,N_2754,N_2963);
or UO_251 (O_251,N_2781,N_2567);
or UO_252 (O_252,N_2593,N_2718);
or UO_253 (O_253,N_2975,N_2929);
or UO_254 (O_254,N_2725,N_2720);
nor UO_255 (O_255,N_2783,N_2786);
and UO_256 (O_256,N_2767,N_2600);
and UO_257 (O_257,N_2737,N_2812);
xor UO_258 (O_258,N_2986,N_2524);
and UO_259 (O_259,N_2599,N_2834);
nor UO_260 (O_260,N_2993,N_2569);
nor UO_261 (O_261,N_2704,N_2784);
nor UO_262 (O_262,N_2558,N_2671);
xor UO_263 (O_263,N_2634,N_2649);
nand UO_264 (O_264,N_2877,N_2926);
or UO_265 (O_265,N_2588,N_2548);
and UO_266 (O_266,N_2888,N_2667);
nand UO_267 (O_267,N_2726,N_2946);
nand UO_268 (O_268,N_2637,N_2570);
nor UO_269 (O_269,N_2889,N_2566);
nor UO_270 (O_270,N_2547,N_2822);
and UO_271 (O_271,N_2751,N_2844);
nor UO_272 (O_272,N_2632,N_2914);
or UO_273 (O_273,N_2590,N_2536);
nor UO_274 (O_274,N_2934,N_2923);
xnor UO_275 (O_275,N_2583,N_2547);
nor UO_276 (O_276,N_2760,N_2784);
and UO_277 (O_277,N_2682,N_2563);
nand UO_278 (O_278,N_2828,N_2987);
xnor UO_279 (O_279,N_2635,N_2799);
or UO_280 (O_280,N_2597,N_2689);
and UO_281 (O_281,N_2806,N_2842);
nand UO_282 (O_282,N_2765,N_2563);
xor UO_283 (O_283,N_2887,N_2665);
or UO_284 (O_284,N_2712,N_2612);
nor UO_285 (O_285,N_2824,N_2902);
or UO_286 (O_286,N_2502,N_2730);
nand UO_287 (O_287,N_2601,N_2881);
and UO_288 (O_288,N_2586,N_2833);
or UO_289 (O_289,N_2736,N_2684);
nor UO_290 (O_290,N_2827,N_2685);
nand UO_291 (O_291,N_2983,N_2672);
nor UO_292 (O_292,N_2833,N_2636);
nand UO_293 (O_293,N_2972,N_2916);
nor UO_294 (O_294,N_2628,N_2615);
nand UO_295 (O_295,N_2625,N_2871);
or UO_296 (O_296,N_2802,N_2850);
and UO_297 (O_297,N_2580,N_2798);
xor UO_298 (O_298,N_2507,N_2811);
nand UO_299 (O_299,N_2908,N_2829);
or UO_300 (O_300,N_2879,N_2668);
or UO_301 (O_301,N_2615,N_2900);
or UO_302 (O_302,N_2802,N_2789);
xor UO_303 (O_303,N_2811,N_2762);
nor UO_304 (O_304,N_2691,N_2657);
nor UO_305 (O_305,N_2536,N_2609);
or UO_306 (O_306,N_2579,N_2862);
nand UO_307 (O_307,N_2680,N_2670);
nand UO_308 (O_308,N_2763,N_2740);
nor UO_309 (O_309,N_2698,N_2788);
nand UO_310 (O_310,N_2938,N_2877);
nor UO_311 (O_311,N_2570,N_2673);
nand UO_312 (O_312,N_2695,N_2584);
xnor UO_313 (O_313,N_2739,N_2518);
nor UO_314 (O_314,N_2934,N_2627);
nor UO_315 (O_315,N_2969,N_2713);
nand UO_316 (O_316,N_2952,N_2500);
and UO_317 (O_317,N_2645,N_2558);
and UO_318 (O_318,N_2906,N_2598);
or UO_319 (O_319,N_2921,N_2777);
nand UO_320 (O_320,N_2570,N_2789);
and UO_321 (O_321,N_2705,N_2699);
or UO_322 (O_322,N_2834,N_2576);
or UO_323 (O_323,N_2840,N_2948);
nand UO_324 (O_324,N_2944,N_2627);
and UO_325 (O_325,N_2617,N_2823);
xor UO_326 (O_326,N_2911,N_2749);
nor UO_327 (O_327,N_2627,N_2687);
or UO_328 (O_328,N_2812,N_2742);
or UO_329 (O_329,N_2791,N_2699);
xor UO_330 (O_330,N_2646,N_2995);
and UO_331 (O_331,N_2939,N_2627);
and UO_332 (O_332,N_2604,N_2684);
and UO_333 (O_333,N_2612,N_2971);
and UO_334 (O_334,N_2857,N_2999);
and UO_335 (O_335,N_2898,N_2574);
nor UO_336 (O_336,N_2859,N_2641);
or UO_337 (O_337,N_2619,N_2747);
nand UO_338 (O_338,N_2732,N_2597);
and UO_339 (O_339,N_2948,N_2672);
nand UO_340 (O_340,N_2940,N_2631);
or UO_341 (O_341,N_2661,N_2562);
nor UO_342 (O_342,N_2859,N_2510);
and UO_343 (O_343,N_2835,N_2912);
nor UO_344 (O_344,N_2562,N_2603);
and UO_345 (O_345,N_2969,N_2688);
xor UO_346 (O_346,N_2930,N_2594);
nor UO_347 (O_347,N_2984,N_2608);
or UO_348 (O_348,N_2728,N_2749);
and UO_349 (O_349,N_2718,N_2568);
nand UO_350 (O_350,N_2803,N_2851);
nor UO_351 (O_351,N_2522,N_2686);
nor UO_352 (O_352,N_2769,N_2866);
xor UO_353 (O_353,N_2651,N_2706);
nand UO_354 (O_354,N_2860,N_2925);
xor UO_355 (O_355,N_2642,N_2987);
nor UO_356 (O_356,N_2972,N_2853);
and UO_357 (O_357,N_2859,N_2724);
and UO_358 (O_358,N_2896,N_2707);
and UO_359 (O_359,N_2580,N_2502);
nor UO_360 (O_360,N_2708,N_2683);
nor UO_361 (O_361,N_2522,N_2861);
and UO_362 (O_362,N_2599,N_2869);
or UO_363 (O_363,N_2744,N_2666);
and UO_364 (O_364,N_2874,N_2776);
and UO_365 (O_365,N_2864,N_2570);
and UO_366 (O_366,N_2559,N_2545);
or UO_367 (O_367,N_2574,N_2505);
or UO_368 (O_368,N_2502,N_2789);
or UO_369 (O_369,N_2923,N_2660);
or UO_370 (O_370,N_2817,N_2904);
nand UO_371 (O_371,N_2747,N_2552);
nor UO_372 (O_372,N_2778,N_2671);
xnor UO_373 (O_373,N_2676,N_2600);
xor UO_374 (O_374,N_2768,N_2578);
or UO_375 (O_375,N_2810,N_2931);
xnor UO_376 (O_376,N_2656,N_2869);
nand UO_377 (O_377,N_2616,N_2870);
nor UO_378 (O_378,N_2764,N_2501);
nand UO_379 (O_379,N_2829,N_2699);
xor UO_380 (O_380,N_2898,N_2532);
nor UO_381 (O_381,N_2653,N_2896);
nor UO_382 (O_382,N_2664,N_2694);
and UO_383 (O_383,N_2606,N_2630);
and UO_384 (O_384,N_2651,N_2550);
or UO_385 (O_385,N_2603,N_2654);
xnor UO_386 (O_386,N_2738,N_2863);
nor UO_387 (O_387,N_2968,N_2845);
or UO_388 (O_388,N_2642,N_2633);
nand UO_389 (O_389,N_2551,N_2813);
nand UO_390 (O_390,N_2629,N_2960);
and UO_391 (O_391,N_2735,N_2964);
xnor UO_392 (O_392,N_2723,N_2759);
nand UO_393 (O_393,N_2566,N_2546);
and UO_394 (O_394,N_2654,N_2898);
and UO_395 (O_395,N_2873,N_2669);
or UO_396 (O_396,N_2985,N_2686);
nand UO_397 (O_397,N_2535,N_2880);
and UO_398 (O_398,N_2565,N_2651);
nand UO_399 (O_399,N_2730,N_2817);
or UO_400 (O_400,N_2742,N_2547);
nor UO_401 (O_401,N_2759,N_2859);
or UO_402 (O_402,N_2921,N_2605);
or UO_403 (O_403,N_2531,N_2622);
nand UO_404 (O_404,N_2563,N_2824);
nor UO_405 (O_405,N_2564,N_2590);
nor UO_406 (O_406,N_2542,N_2654);
or UO_407 (O_407,N_2940,N_2975);
and UO_408 (O_408,N_2991,N_2944);
or UO_409 (O_409,N_2588,N_2885);
nand UO_410 (O_410,N_2531,N_2797);
nand UO_411 (O_411,N_2952,N_2854);
nor UO_412 (O_412,N_2961,N_2554);
nand UO_413 (O_413,N_2970,N_2939);
or UO_414 (O_414,N_2887,N_2738);
nor UO_415 (O_415,N_2896,N_2797);
nor UO_416 (O_416,N_2856,N_2836);
nand UO_417 (O_417,N_2674,N_2522);
nor UO_418 (O_418,N_2634,N_2823);
and UO_419 (O_419,N_2960,N_2783);
nor UO_420 (O_420,N_2972,N_2941);
nand UO_421 (O_421,N_2931,N_2782);
nand UO_422 (O_422,N_2674,N_2683);
nand UO_423 (O_423,N_2907,N_2887);
nand UO_424 (O_424,N_2582,N_2828);
xor UO_425 (O_425,N_2859,N_2715);
or UO_426 (O_426,N_2628,N_2724);
nor UO_427 (O_427,N_2619,N_2545);
nand UO_428 (O_428,N_2729,N_2960);
or UO_429 (O_429,N_2959,N_2845);
and UO_430 (O_430,N_2771,N_2958);
xor UO_431 (O_431,N_2760,N_2544);
and UO_432 (O_432,N_2556,N_2781);
and UO_433 (O_433,N_2776,N_2807);
and UO_434 (O_434,N_2998,N_2842);
nand UO_435 (O_435,N_2535,N_2810);
xnor UO_436 (O_436,N_2607,N_2575);
nor UO_437 (O_437,N_2915,N_2886);
nor UO_438 (O_438,N_2576,N_2745);
nand UO_439 (O_439,N_2692,N_2652);
nor UO_440 (O_440,N_2631,N_2679);
or UO_441 (O_441,N_2526,N_2589);
nand UO_442 (O_442,N_2590,N_2799);
nor UO_443 (O_443,N_2502,N_2757);
nand UO_444 (O_444,N_2639,N_2911);
and UO_445 (O_445,N_2661,N_2969);
xnor UO_446 (O_446,N_2529,N_2726);
nor UO_447 (O_447,N_2582,N_2814);
or UO_448 (O_448,N_2752,N_2512);
nand UO_449 (O_449,N_2756,N_2602);
nor UO_450 (O_450,N_2997,N_2958);
or UO_451 (O_451,N_2701,N_2707);
nor UO_452 (O_452,N_2657,N_2968);
xnor UO_453 (O_453,N_2575,N_2658);
xor UO_454 (O_454,N_2670,N_2547);
and UO_455 (O_455,N_2601,N_2722);
nand UO_456 (O_456,N_2937,N_2951);
nand UO_457 (O_457,N_2995,N_2635);
or UO_458 (O_458,N_2734,N_2838);
xnor UO_459 (O_459,N_2971,N_2624);
nor UO_460 (O_460,N_2741,N_2556);
or UO_461 (O_461,N_2617,N_2961);
nor UO_462 (O_462,N_2960,N_2560);
xnor UO_463 (O_463,N_2524,N_2776);
nand UO_464 (O_464,N_2850,N_2615);
nor UO_465 (O_465,N_2755,N_2691);
or UO_466 (O_466,N_2946,N_2683);
nand UO_467 (O_467,N_2683,N_2942);
nor UO_468 (O_468,N_2675,N_2538);
nand UO_469 (O_469,N_2920,N_2871);
or UO_470 (O_470,N_2726,N_2720);
xnor UO_471 (O_471,N_2800,N_2599);
and UO_472 (O_472,N_2570,N_2945);
nor UO_473 (O_473,N_2689,N_2873);
or UO_474 (O_474,N_2880,N_2567);
or UO_475 (O_475,N_2587,N_2765);
and UO_476 (O_476,N_2597,N_2575);
or UO_477 (O_477,N_2767,N_2719);
and UO_478 (O_478,N_2664,N_2905);
nand UO_479 (O_479,N_2606,N_2762);
or UO_480 (O_480,N_2991,N_2973);
and UO_481 (O_481,N_2652,N_2873);
or UO_482 (O_482,N_2786,N_2551);
or UO_483 (O_483,N_2627,N_2533);
nor UO_484 (O_484,N_2939,N_2596);
nor UO_485 (O_485,N_2695,N_2741);
xor UO_486 (O_486,N_2715,N_2735);
or UO_487 (O_487,N_2624,N_2811);
or UO_488 (O_488,N_2804,N_2918);
nor UO_489 (O_489,N_2897,N_2879);
nand UO_490 (O_490,N_2866,N_2634);
nand UO_491 (O_491,N_2899,N_2962);
and UO_492 (O_492,N_2701,N_2550);
nand UO_493 (O_493,N_2612,N_2862);
nor UO_494 (O_494,N_2783,N_2752);
and UO_495 (O_495,N_2794,N_2967);
xnor UO_496 (O_496,N_2822,N_2597);
nand UO_497 (O_497,N_2908,N_2997);
xor UO_498 (O_498,N_2636,N_2773);
or UO_499 (O_499,N_2557,N_2947);
endmodule