module basic_500_3000_500_60_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_127,In_458);
or U1 (N_1,In_487,In_89);
nand U2 (N_2,In_237,In_201);
nor U3 (N_3,In_153,In_62);
nor U4 (N_4,In_199,In_366);
nor U5 (N_5,In_336,In_297);
or U6 (N_6,In_410,In_350);
nor U7 (N_7,In_359,In_49);
and U8 (N_8,In_453,In_29);
nor U9 (N_9,In_322,In_79);
or U10 (N_10,In_399,In_1);
nor U11 (N_11,In_324,In_149);
xor U12 (N_12,In_284,In_92);
nor U13 (N_13,In_100,In_242);
and U14 (N_14,In_99,In_270);
or U15 (N_15,In_415,In_150);
and U16 (N_16,In_185,In_22);
nand U17 (N_17,In_42,In_264);
and U18 (N_18,In_274,In_216);
nor U19 (N_19,In_381,In_280);
nand U20 (N_20,In_391,In_132);
nor U21 (N_21,In_262,In_94);
or U22 (N_22,In_311,In_442);
nor U23 (N_23,In_183,In_301);
nand U24 (N_24,In_379,In_427);
nor U25 (N_25,In_470,In_20);
nor U26 (N_26,In_107,In_471);
nand U27 (N_27,In_226,In_74);
nor U28 (N_28,In_479,In_174);
or U29 (N_29,In_388,In_243);
nor U30 (N_30,In_346,In_239);
nand U31 (N_31,In_90,In_402);
or U32 (N_32,In_56,In_141);
and U33 (N_33,In_302,In_455);
xnor U34 (N_34,In_133,In_58);
or U35 (N_35,In_358,In_469);
or U36 (N_36,In_236,In_326);
or U37 (N_37,In_123,In_308);
nand U38 (N_38,In_317,In_215);
and U39 (N_39,In_283,In_66);
or U40 (N_40,In_34,In_116);
nor U41 (N_41,In_265,In_76);
and U42 (N_42,In_357,In_443);
xnor U43 (N_43,In_347,In_281);
and U44 (N_44,In_300,In_447);
and U45 (N_45,In_148,In_329);
xnor U46 (N_46,In_178,In_200);
xor U47 (N_47,In_436,In_320);
nand U48 (N_48,In_495,In_9);
or U49 (N_49,In_491,In_333);
xnor U50 (N_50,N_34,In_253);
and U51 (N_51,In_108,In_38);
nor U52 (N_52,In_59,In_371);
xnor U53 (N_53,N_45,In_356);
and U54 (N_54,N_21,In_23);
xnor U55 (N_55,In_298,In_287);
xnor U56 (N_56,In_225,In_407);
xnor U57 (N_57,In_106,In_383);
nor U58 (N_58,In_212,In_286);
and U59 (N_59,In_273,In_21);
xnor U60 (N_60,N_26,In_478);
and U61 (N_61,In_248,In_77);
and U62 (N_62,In_257,In_485);
xnor U63 (N_63,N_18,In_91);
nand U64 (N_64,In_52,In_192);
nand U65 (N_65,N_46,In_84);
and U66 (N_66,In_306,In_65);
nand U67 (N_67,N_2,In_271);
nor U68 (N_68,In_196,In_187);
nand U69 (N_69,In_457,In_335);
and U70 (N_70,In_426,In_2);
xor U71 (N_71,In_289,In_213);
nand U72 (N_72,In_223,In_0);
nand U73 (N_73,In_362,In_327);
nor U74 (N_74,In_250,In_206);
or U75 (N_75,In_450,In_54);
xnor U76 (N_76,In_365,In_285);
nand U77 (N_77,N_7,In_130);
or U78 (N_78,In_499,In_463);
nand U79 (N_79,In_377,In_343);
xor U80 (N_80,In_345,In_230);
xnor U81 (N_81,N_23,N_41);
nor U82 (N_82,In_131,In_303);
nor U83 (N_83,In_494,In_218);
nand U84 (N_84,In_44,In_97);
and U85 (N_85,N_25,In_87);
nand U86 (N_86,In_184,In_15);
xor U87 (N_87,In_168,In_35);
and U88 (N_88,In_451,In_98);
nor U89 (N_89,In_288,In_423);
nor U90 (N_90,In_181,In_466);
and U91 (N_91,In_293,In_46);
or U92 (N_92,In_432,In_24);
nand U93 (N_93,In_63,In_348);
nor U94 (N_94,In_119,In_269);
nand U95 (N_95,N_31,In_373);
and U96 (N_96,In_17,In_31);
nand U97 (N_97,In_454,In_53);
and U98 (N_98,In_41,In_331);
or U99 (N_99,In_96,In_268);
xnor U100 (N_100,N_27,In_80);
or U101 (N_101,In_395,In_481);
nand U102 (N_102,In_165,In_10);
or U103 (N_103,In_477,In_382);
nor U104 (N_104,In_173,N_95);
or U105 (N_105,N_69,In_144);
nor U106 (N_106,In_456,In_368);
nand U107 (N_107,In_352,In_85);
and U108 (N_108,In_459,In_472);
or U109 (N_109,In_69,In_191);
nor U110 (N_110,In_386,N_83);
and U111 (N_111,In_138,In_78);
or U112 (N_112,In_344,N_89);
or U113 (N_113,In_205,In_460);
or U114 (N_114,In_228,In_401);
xor U115 (N_115,In_290,In_145);
xor U116 (N_116,In_369,In_384);
nor U117 (N_117,N_73,N_29);
xor U118 (N_118,In_473,In_146);
nand U119 (N_119,In_406,In_476);
nor U120 (N_120,In_13,N_4);
nand U121 (N_121,In_431,In_439);
xnor U122 (N_122,In_118,In_93);
nand U123 (N_123,In_489,In_323);
nor U124 (N_124,In_313,In_207);
and U125 (N_125,In_414,In_259);
or U126 (N_126,N_43,In_389);
or U127 (N_127,In_341,In_75);
and U128 (N_128,In_251,N_48);
or U129 (N_129,In_68,In_231);
and U130 (N_130,N_62,In_304);
nand U131 (N_131,N_64,In_88);
nand U132 (N_132,N_90,In_449);
nand U133 (N_133,In_355,In_428);
and U134 (N_134,In_433,In_12);
nand U135 (N_135,In_444,In_486);
nor U136 (N_136,In_14,N_87);
nor U137 (N_137,In_394,In_480);
or U138 (N_138,In_310,In_227);
nand U139 (N_139,In_50,In_246);
nor U140 (N_140,N_13,N_10);
nand U141 (N_141,N_16,In_339);
nand U142 (N_142,In_134,N_53);
or U143 (N_143,In_167,In_363);
or U144 (N_144,In_3,In_198);
or U145 (N_145,In_390,In_28);
or U146 (N_146,N_51,In_400);
nor U147 (N_147,In_140,In_376);
and U148 (N_148,N_74,In_27);
xnor U149 (N_149,N_55,In_222);
xor U150 (N_150,In_364,In_81);
nand U151 (N_151,In_424,In_435);
nor U152 (N_152,In_135,In_67);
nand U153 (N_153,In_186,N_114);
nand U154 (N_154,N_134,In_385);
xor U155 (N_155,In_163,In_448);
nand U156 (N_156,N_57,In_147);
or U157 (N_157,N_35,N_120);
or U158 (N_158,In_217,In_263);
nor U159 (N_159,In_137,N_141);
and U160 (N_160,N_118,In_421);
or U161 (N_161,In_255,In_397);
xnor U162 (N_162,In_374,In_55);
xor U163 (N_163,N_15,In_387);
or U164 (N_164,In_72,In_316);
nor U165 (N_165,In_151,In_408);
and U166 (N_166,In_484,In_398);
and U167 (N_167,N_94,In_474);
nor U168 (N_168,N_30,In_482);
nor U169 (N_169,N_88,N_37);
or U170 (N_170,In_214,In_156);
xor U171 (N_171,In_493,In_354);
nand U172 (N_172,In_249,N_54);
xor U173 (N_173,N_119,In_48);
and U174 (N_174,N_96,In_170);
xnor U175 (N_175,In_171,In_372);
nand U176 (N_176,In_220,N_52);
xnor U177 (N_177,In_464,In_16);
xor U178 (N_178,In_202,In_315);
and U179 (N_179,In_26,N_132);
nor U180 (N_180,In_112,In_61);
nand U181 (N_181,In_221,N_136);
and U182 (N_182,In_244,In_351);
and U183 (N_183,In_124,In_497);
nor U184 (N_184,In_47,In_73);
and U185 (N_185,In_83,In_430);
xnor U186 (N_186,In_314,In_419);
or U187 (N_187,In_349,N_49);
nand U188 (N_188,In_71,In_177);
xnor U189 (N_189,In_115,In_294);
nand U190 (N_190,In_256,In_321);
nand U191 (N_191,N_84,N_60);
or U192 (N_192,In_405,In_169);
and U193 (N_193,In_162,In_440);
or U194 (N_194,In_6,N_28);
xnor U195 (N_195,N_99,In_155);
or U196 (N_196,In_332,In_43);
or U197 (N_197,N_130,N_97);
and U198 (N_198,In_411,In_412);
nand U199 (N_199,N_40,N_127);
and U200 (N_200,N_33,In_370);
nand U201 (N_201,In_319,N_11);
xnor U202 (N_202,In_292,N_72);
or U203 (N_203,In_445,N_151);
or U204 (N_204,N_100,N_169);
nor U205 (N_205,In_245,In_465);
or U206 (N_206,In_438,In_160);
nand U207 (N_207,N_63,N_184);
or U208 (N_208,In_70,N_101);
and U209 (N_209,In_60,N_106);
or U210 (N_210,In_299,In_429);
nand U211 (N_211,In_241,In_224);
and U212 (N_212,In_434,In_64);
and U213 (N_213,In_158,N_135);
nand U214 (N_214,In_125,In_11);
xnor U215 (N_215,N_108,In_483);
nand U216 (N_216,In_232,N_162);
or U217 (N_217,N_155,In_203);
nand U218 (N_218,N_22,N_12);
or U219 (N_219,N_153,In_254);
nor U220 (N_220,N_111,In_238);
and U221 (N_221,N_197,In_95);
xor U222 (N_222,N_193,N_5);
nor U223 (N_223,N_50,In_101);
xor U224 (N_224,In_325,N_138);
xor U225 (N_225,In_4,N_107);
nand U226 (N_226,N_112,N_170);
or U227 (N_227,N_36,In_361);
and U228 (N_228,In_404,In_114);
or U229 (N_229,N_152,N_14);
xor U230 (N_230,In_139,In_417);
nor U231 (N_231,In_25,In_413);
and U232 (N_232,In_425,N_188);
nor U233 (N_233,N_104,N_32);
or U234 (N_234,In_33,N_123);
and U235 (N_235,In_111,In_109);
xnor U236 (N_236,In_378,In_266);
and U237 (N_237,In_154,N_82);
xor U238 (N_238,N_144,N_113);
nand U239 (N_239,N_44,In_211);
nand U240 (N_240,In_157,N_176);
nor U241 (N_241,N_20,N_187);
nand U242 (N_242,In_267,N_8);
or U243 (N_243,N_189,N_180);
or U244 (N_244,N_105,N_124);
and U245 (N_245,In_209,N_70);
or U246 (N_246,N_93,In_5);
nand U247 (N_247,N_142,N_3);
xor U248 (N_248,N_81,In_403);
xor U249 (N_249,In_260,In_420);
xor U250 (N_250,In_338,N_206);
nand U251 (N_251,In_190,In_82);
and U252 (N_252,In_467,In_296);
nand U253 (N_253,N_211,In_104);
xnor U254 (N_254,N_241,N_65);
xor U255 (N_255,N_232,In_129);
nor U256 (N_256,N_171,In_8);
or U257 (N_257,In_117,In_353);
nor U258 (N_258,N_209,In_152);
nand U259 (N_259,In_105,N_131);
and U260 (N_260,N_156,In_240);
and U261 (N_261,N_76,In_103);
and U262 (N_262,In_380,In_18);
nand U263 (N_263,In_307,In_312);
nor U264 (N_264,N_208,N_129);
and U265 (N_265,N_58,N_215);
nand U266 (N_266,N_239,In_488);
or U267 (N_267,N_174,In_126);
or U268 (N_268,In_45,N_240);
nor U269 (N_269,N_143,N_212);
nand U270 (N_270,In_277,In_143);
xor U271 (N_271,N_178,N_230);
xor U272 (N_272,N_61,In_121);
xor U273 (N_273,N_39,N_228);
nor U274 (N_274,In_110,In_36);
or U275 (N_275,In_360,N_223);
nand U276 (N_276,In_30,In_330);
or U277 (N_277,In_490,N_1);
nor U278 (N_278,In_461,In_416);
and U279 (N_279,N_56,In_172);
nor U280 (N_280,N_150,N_139);
and U281 (N_281,N_166,N_9);
nand U282 (N_282,In_462,In_441);
xor U283 (N_283,N_148,In_37);
and U284 (N_284,N_231,In_193);
xnor U285 (N_285,N_24,In_409);
or U286 (N_286,N_92,In_234);
xnor U287 (N_287,In_142,In_102);
nor U288 (N_288,In_342,In_496);
nor U289 (N_289,N_186,N_19);
nand U290 (N_290,N_137,In_175);
nand U291 (N_291,In_279,N_17);
or U292 (N_292,N_182,N_217);
nor U293 (N_293,In_468,In_452);
nand U294 (N_294,In_51,N_219);
xnor U295 (N_295,N_225,In_235);
and U296 (N_296,In_437,In_328);
xnor U297 (N_297,N_203,In_39);
and U298 (N_298,N_172,N_126);
and U299 (N_299,N_201,In_446);
or U300 (N_300,N_165,N_133);
xor U301 (N_301,N_159,N_244);
and U302 (N_302,N_85,N_255);
and U303 (N_303,N_121,N_214);
nand U304 (N_304,In_278,In_375);
nor U305 (N_305,N_229,N_233);
nor U306 (N_306,In_204,N_270);
or U307 (N_307,N_249,N_195);
nor U308 (N_308,N_200,N_274);
and U309 (N_309,N_252,N_79);
nor U310 (N_310,N_279,N_245);
or U311 (N_311,In_258,In_194);
or U312 (N_312,N_247,N_80);
nand U313 (N_313,In_337,N_190);
nor U314 (N_314,N_294,N_102);
nand U315 (N_315,N_6,In_7);
nor U316 (N_316,N_277,N_295);
and U317 (N_317,In_367,N_261);
and U318 (N_318,N_145,N_196);
nor U319 (N_319,N_213,N_289);
or U320 (N_320,In_291,In_166);
and U321 (N_321,N_287,N_86);
nand U322 (N_322,N_71,N_297);
xor U323 (N_323,N_236,N_282);
nor U324 (N_324,N_181,N_299);
xor U325 (N_325,N_291,N_183);
nand U326 (N_326,N_226,N_167);
nand U327 (N_327,N_163,In_261);
or U328 (N_328,N_161,N_227);
nor U329 (N_329,In_40,In_418);
nor U330 (N_330,In_179,N_234);
nand U331 (N_331,N_125,In_86);
or U332 (N_332,N_68,In_396);
nor U333 (N_333,N_204,N_248);
nand U334 (N_334,In_318,N_168);
xor U335 (N_335,N_238,N_272);
xor U336 (N_336,N_254,N_285);
xor U337 (N_337,N_264,N_115);
nand U338 (N_338,N_250,N_91);
or U339 (N_339,In_164,N_205);
nand U340 (N_340,In_159,N_198);
and U341 (N_341,N_164,N_271);
nor U342 (N_342,N_260,In_32);
nor U343 (N_343,N_38,N_157);
xor U344 (N_344,In_334,N_276);
xor U345 (N_345,N_207,N_283);
nor U346 (N_346,N_173,N_0);
nand U347 (N_347,N_177,In_161);
nor U348 (N_348,N_222,N_175);
xnor U349 (N_349,In_422,N_59);
nor U350 (N_350,N_147,N_327);
nor U351 (N_351,N_321,N_317);
or U352 (N_352,N_324,N_312);
nand U353 (N_353,N_251,N_339);
or U354 (N_354,N_140,N_47);
nor U355 (N_355,N_330,N_154);
and U356 (N_356,In_393,N_146);
or U357 (N_357,N_149,In_189);
nand U358 (N_358,In_176,N_336);
and U359 (N_359,N_243,In_392);
xor U360 (N_360,N_216,In_210);
xnor U361 (N_361,N_109,N_300);
or U362 (N_362,N_242,N_284);
nor U363 (N_363,N_309,N_292);
and U364 (N_364,N_306,N_110);
xnor U365 (N_365,N_314,In_282);
xor U366 (N_366,In_197,N_256);
and U367 (N_367,N_340,N_349);
nand U368 (N_368,N_335,N_286);
xnor U369 (N_369,N_311,In_247);
xnor U370 (N_370,In_276,In_219);
xor U371 (N_371,N_237,N_246);
and U372 (N_372,N_308,N_266);
nor U373 (N_373,N_262,N_265);
or U374 (N_374,N_128,N_75);
or U375 (N_375,N_273,N_191);
nand U376 (N_376,In_19,N_103);
nand U377 (N_377,N_199,N_268);
xor U378 (N_378,N_98,N_342);
and U379 (N_379,N_345,In_188);
and U380 (N_380,N_258,N_160);
or U381 (N_381,N_185,N_334);
or U382 (N_382,N_303,In_275);
nand U383 (N_383,N_331,N_158);
nor U384 (N_384,N_310,N_179);
nor U385 (N_385,N_307,In_122);
xnor U386 (N_386,N_320,In_182);
xnor U387 (N_387,N_269,N_42);
and U388 (N_388,N_301,N_333);
nand U389 (N_389,In_136,N_263);
xor U390 (N_390,N_325,N_332);
or U391 (N_391,N_117,N_122);
nor U392 (N_392,N_77,In_295);
and U393 (N_393,N_341,N_288);
nand U394 (N_394,In_113,N_323);
nor U395 (N_395,N_290,N_296);
and U396 (N_396,N_78,In_309);
and U397 (N_397,N_259,N_329);
and U398 (N_398,In_272,N_319);
nand U399 (N_399,N_338,In_475);
xor U400 (N_400,In_229,N_370);
and U401 (N_401,N_384,N_348);
xor U402 (N_402,N_218,N_389);
and U403 (N_403,In_252,N_391);
nand U404 (N_404,N_318,N_379);
xnor U405 (N_405,In_340,In_498);
nor U406 (N_406,N_378,N_281);
nand U407 (N_407,N_363,N_360);
nand U408 (N_408,N_374,N_396);
nand U409 (N_409,N_390,N_386);
nand U410 (N_410,N_344,N_221);
and U411 (N_411,N_383,N_395);
and U412 (N_412,N_356,N_367);
nand U413 (N_413,N_355,N_359);
nor U414 (N_414,N_365,In_305);
or U415 (N_415,N_398,N_328);
or U416 (N_416,N_381,N_368);
or U417 (N_417,N_369,N_202);
or U418 (N_418,N_394,N_371);
xor U419 (N_419,N_343,N_346);
or U420 (N_420,In_208,In_128);
nor U421 (N_421,N_192,N_375);
or U422 (N_422,N_278,N_366);
and U423 (N_423,N_235,N_116);
nand U424 (N_424,N_354,In_120);
or U425 (N_425,N_267,N_322);
nand U426 (N_426,N_337,N_392);
nor U427 (N_427,N_380,N_66);
or U428 (N_428,In_233,In_180);
nor U429 (N_429,N_302,N_351);
and U430 (N_430,N_67,N_280);
or U431 (N_431,N_347,N_373);
nand U432 (N_432,In_195,N_358);
and U433 (N_433,N_353,N_385);
xor U434 (N_434,N_315,N_361);
nand U435 (N_435,N_220,N_364);
xnor U436 (N_436,N_298,N_388);
nor U437 (N_437,N_382,N_393);
xor U438 (N_438,N_316,N_194);
nor U439 (N_439,N_304,N_397);
nor U440 (N_440,N_387,In_492);
nand U441 (N_441,In_57,N_352);
and U442 (N_442,N_372,N_399);
and U443 (N_443,N_377,N_376);
nand U444 (N_444,N_293,N_326);
nand U445 (N_445,N_313,N_362);
nand U446 (N_446,N_210,N_275);
and U447 (N_447,N_350,N_257);
and U448 (N_448,N_224,N_357);
and U449 (N_449,N_253,N_305);
nor U450 (N_450,N_405,N_446);
and U451 (N_451,N_433,N_407);
and U452 (N_452,N_449,N_424);
xor U453 (N_453,N_414,N_430);
and U454 (N_454,N_438,N_419);
and U455 (N_455,N_439,N_427);
and U456 (N_456,N_425,N_400);
nand U457 (N_457,N_443,N_413);
nand U458 (N_458,N_448,N_435);
nor U459 (N_459,N_423,N_437);
nor U460 (N_460,N_429,N_406);
xor U461 (N_461,N_428,N_434);
or U462 (N_462,N_410,N_404);
nor U463 (N_463,N_442,N_412);
nand U464 (N_464,N_418,N_402);
or U465 (N_465,N_420,N_409);
xnor U466 (N_466,N_447,N_421);
nand U467 (N_467,N_441,N_440);
nor U468 (N_468,N_431,N_426);
xnor U469 (N_469,N_444,N_401);
and U470 (N_470,N_408,N_403);
xnor U471 (N_471,N_432,N_416);
nand U472 (N_472,N_422,N_445);
and U473 (N_473,N_436,N_415);
and U474 (N_474,N_411,N_417);
nor U475 (N_475,N_413,N_407);
nand U476 (N_476,N_446,N_429);
xor U477 (N_477,N_435,N_400);
xnor U478 (N_478,N_446,N_411);
nand U479 (N_479,N_449,N_427);
nand U480 (N_480,N_421,N_430);
nor U481 (N_481,N_408,N_423);
xor U482 (N_482,N_406,N_418);
and U483 (N_483,N_408,N_429);
nor U484 (N_484,N_423,N_401);
or U485 (N_485,N_447,N_428);
and U486 (N_486,N_405,N_442);
nor U487 (N_487,N_435,N_438);
xor U488 (N_488,N_442,N_432);
xor U489 (N_489,N_413,N_435);
or U490 (N_490,N_444,N_440);
nand U491 (N_491,N_437,N_412);
xor U492 (N_492,N_432,N_431);
xor U493 (N_493,N_401,N_414);
nor U494 (N_494,N_432,N_441);
and U495 (N_495,N_422,N_425);
and U496 (N_496,N_445,N_403);
xnor U497 (N_497,N_441,N_419);
nand U498 (N_498,N_439,N_434);
or U499 (N_499,N_413,N_421);
xor U500 (N_500,N_488,N_483);
nand U501 (N_501,N_495,N_459);
or U502 (N_502,N_487,N_450);
or U503 (N_503,N_491,N_461);
or U504 (N_504,N_484,N_462);
nor U505 (N_505,N_481,N_485);
nand U506 (N_506,N_463,N_466);
and U507 (N_507,N_474,N_452);
nor U508 (N_508,N_473,N_475);
or U509 (N_509,N_458,N_453);
nor U510 (N_510,N_489,N_457);
nor U511 (N_511,N_456,N_460);
nor U512 (N_512,N_492,N_494);
xor U513 (N_513,N_477,N_496);
nor U514 (N_514,N_498,N_469);
nand U515 (N_515,N_471,N_476);
xnor U516 (N_516,N_478,N_480);
or U517 (N_517,N_499,N_479);
xor U518 (N_518,N_467,N_493);
nor U519 (N_519,N_490,N_486);
and U520 (N_520,N_455,N_451);
nand U521 (N_521,N_464,N_497);
nor U522 (N_522,N_470,N_468);
and U523 (N_523,N_472,N_482);
and U524 (N_524,N_454,N_465);
nand U525 (N_525,N_499,N_456);
nor U526 (N_526,N_483,N_476);
and U527 (N_527,N_479,N_472);
nor U528 (N_528,N_460,N_474);
or U529 (N_529,N_486,N_493);
xor U530 (N_530,N_463,N_454);
xor U531 (N_531,N_482,N_469);
nand U532 (N_532,N_469,N_491);
xor U533 (N_533,N_471,N_460);
xor U534 (N_534,N_480,N_466);
and U535 (N_535,N_451,N_469);
and U536 (N_536,N_465,N_471);
or U537 (N_537,N_492,N_467);
xor U538 (N_538,N_484,N_492);
or U539 (N_539,N_460,N_488);
nand U540 (N_540,N_451,N_483);
nor U541 (N_541,N_470,N_475);
nand U542 (N_542,N_480,N_489);
or U543 (N_543,N_484,N_460);
or U544 (N_544,N_483,N_481);
nand U545 (N_545,N_479,N_460);
xnor U546 (N_546,N_481,N_463);
nor U547 (N_547,N_489,N_467);
and U548 (N_548,N_472,N_456);
xnor U549 (N_549,N_453,N_462);
or U550 (N_550,N_532,N_548);
nor U551 (N_551,N_518,N_543);
xor U552 (N_552,N_533,N_524);
nor U553 (N_553,N_516,N_501);
nand U554 (N_554,N_508,N_520);
nand U555 (N_555,N_535,N_502);
nand U556 (N_556,N_546,N_514);
or U557 (N_557,N_529,N_505);
nor U558 (N_558,N_525,N_517);
and U559 (N_559,N_521,N_542);
nor U560 (N_560,N_504,N_540);
nor U561 (N_561,N_507,N_523);
nand U562 (N_562,N_544,N_519);
and U563 (N_563,N_531,N_549);
nand U564 (N_564,N_522,N_537);
nand U565 (N_565,N_510,N_534);
xor U566 (N_566,N_547,N_536);
nand U567 (N_567,N_512,N_503);
nand U568 (N_568,N_509,N_500);
xor U569 (N_569,N_530,N_541);
xnor U570 (N_570,N_527,N_528);
xor U571 (N_571,N_538,N_539);
xor U572 (N_572,N_526,N_506);
and U573 (N_573,N_515,N_511);
or U574 (N_574,N_513,N_545);
nand U575 (N_575,N_512,N_506);
nor U576 (N_576,N_540,N_546);
nor U577 (N_577,N_533,N_510);
nand U578 (N_578,N_542,N_505);
nand U579 (N_579,N_505,N_526);
or U580 (N_580,N_532,N_502);
nor U581 (N_581,N_505,N_530);
or U582 (N_582,N_547,N_541);
and U583 (N_583,N_530,N_524);
or U584 (N_584,N_529,N_548);
nor U585 (N_585,N_525,N_510);
xor U586 (N_586,N_522,N_545);
nor U587 (N_587,N_518,N_507);
or U588 (N_588,N_538,N_521);
xnor U589 (N_589,N_525,N_523);
nand U590 (N_590,N_519,N_526);
nor U591 (N_591,N_508,N_530);
and U592 (N_592,N_548,N_508);
nor U593 (N_593,N_517,N_522);
nor U594 (N_594,N_521,N_513);
or U595 (N_595,N_542,N_509);
and U596 (N_596,N_539,N_544);
xor U597 (N_597,N_540,N_517);
nor U598 (N_598,N_506,N_503);
nand U599 (N_599,N_523,N_540);
and U600 (N_600,N_584,N_556);
or U601 (N_601,N_571,N_582);
and U602 (N_602,N_561,N_558);
nand U603 (N_603,N_575,N_579);
or U604 (N_604,N_596,N_580);
nand U605 (N_605,N_593,N_559);
nor U606 (N_606,N_589,N_594);
or U607 (N_607,N_550,N_554);
or U608 (N_608,N_557,N_578);
nor U609 (N_609,N_565,N_574);
nand U610 (N_610,N_599,N_592);
xnor U611 (N_611,N_590,N_585);
xnor U612 (N_612,N_562,N_586);
and U613 (N_613,N_595,N_583);
xor U614 (N_614,N_568,N_581);
or U615 (N_615,N_577,N_564);
or U616 (N_616,N_560,N_552);
nor U617 (N_617,N_551,N_563);
nor U618 (N_618,N_569,N_591);
nor U619 (N_619,N_566,N_567);
xnor U620 (N_620,N_597,N_573);
or U621 (N_621,N_572,N_553);
nor U622 (N_622,N_588,N_587);
or U623 (N_623,N_555,N_598);
nor U624 (N_624,N_576,N_570);
nor U625 (N_625,N_576,N_557);
nor U626 (N_626,N_573,N_575);
xnor U627 (N_627,N_567,N_575);
or U628 (N_628,N_556,N_598);
xnor U629 (N_629,N_565,N_571);
nor U630 (N_630,N_574,N_588);
and U631 (N_631,N_569,N_584);
or U632 (N_632,N_550,N_567);
and U633 (N_633,N_568,N_565);
or U634 (N_634,N_568,N_597);
nor U635 (N_635,N_596,N_563);
or U636 (N_636,N_569,N_597);
or U637 (N_637,N_569,N_562);
nand U638 (N_638,N_550,N_590);
nor U639 (N_639,N_589,N_572);
or U640 (N_640,N_564,N_561);
or U641 (N_641,N_554,N_593);
nor U642 (N_642,N_566,N_558);
nor U643 (N_643,N_566,N_552);
nand U644 (N_644,N_570,N_586);
nor U645 (N_645,N_591,N_586);
xnor U646 (N_646,N_564,N_586);
nand U647 (N_647,N_580,N_579);
nor U648 (N_648,N_573,N_586);
and U649 (N_649,N_582,N_575);
xnor U650 (N_650,N_649,N_646);
and U651 (N_651,N_619,N_605);
or U652 (N_652,N_638,N_606);
and U653 (N_653,N_622,N_600);
xnor U654 (N_654,N_633,N_640);
or U655 (N_655,N_642,N_621);
xnor U656 (N_656,N_611,N_625);
nor U657 (N_657,N_624,N_614);
or U658 (N_658,N_603,N_618);
nor U659 (N_659,N_636,N_617);
or U660 (N_660,N_647,N_616);
or U661 (N_661,N_612,N_645);
or U662 (N_662,N_602,N_644);
or U663 (N_663,N_628,N_626);
nor U664 (N_664,N_627,N_630);
nor U665 (N_665,N_607,N_631);
and U666 (N_666,N_637,N_609);
and U667 (N_667,N_629,N_641);
and U668 (N_668,N_610,N_620);
xor U669 (N_669,N_613,N_643);
xor U670 (N_670,N_601,N_648);
nor U671 (N_671,N_635,N_639);
nand U672 (N_672,N_608,N_623);
nand U673 (N_673,N_604,N_634);
and U674 (N_674,N_632,N_615);
xnor U675 (N_675,N_628,N_642);
or U676 (N_676,N_613,N_600);
or U677 (N_677,N_649,N_633);
nand U678 (N_678,N_645,N_603);
or U679 (N_679,N_639,N_636);
xnor U680 (N_680,N_601,N_631);
xnor U681 (N_681,N_618,N_609);
xor U682 (N_682,N_606,N_635);
xnor U683 (N_683,N_610,N_638);
xor U684 (N_684,N_630,N_633);
nand U685 (N_685,N_649,N_644);
or U686 (N_686,N_629,N_605);
nand U687 (N_687,N_612,N_614);
nor U688 (N_688,N_642,N_646);
nand U689 (N_689,N_605,N_640);
or U690 (N_690,N_606,N_613);
xor U691 (N_691,N_649,N_601);
and U692 (N_692,N_617,N_618);
or U693 (N_693,N_634,N_633);
and U694 (N_694,N_605,N_616);
nand U695 (N_695,N_649,N_630);
or U696 (N_696,N_614,N_606);
xnor U697 (N_697,N_632,N_621);
nor U698 (N_698,N_621,N_610);
nor U699 (N_699,N_636,N_612);
xnor U700 (N_700,N_660,N_657);
nand U701 (N_701,N_666,N_676);
and U702 (N_702,N_695,N_699);
nor U703 (N_703,N_694,N_656);
or U704 (N_704,N_692,N_658);
xor U705 (N_705,N_669,N_685);
nand U706 (N_706,N_682,N_668);
nor U707 (N_707,N_677,N_696);
nand U708 (N_708,N_691,N_663);
xor U709 (N_709,N_654,N_698);
nand U710 (N_710,N_665,N_675);
or U711 (N_711,N_672,N_650);
or U712 (N_712,N_693,N_683);
xnor U713 (N_713,N_671,N_659);
nand U714 (N_714,N_653,N_689);
xor U715 (N_715,N_664,N_652);
and U716 (N_716,N_651,N_679);
or U717 (N_717,N_670,N_655);
and U718 (N_718,N_681,N_667);
nor U719 (N_719,N_690,N_687);
nor U720 (N_720,N_684,N_686);
or U721 (N_721,N_678,N_688);
and U722 (N_722,N_673,N_674);
nand U723 (N_723,N_662,N_680);
and U724 (N_724,N_697,N_661);
nand U725 (N_725,N_659,N_666);
xnor U726 (N_726,N_667,N_698);
or U727 (N_727,N_687,N_677);
xnor U728 (N_728,N_675,N_685);
nor U729 (N_729,N_669,N_689);
nand U730 (N_730,N_690,N_654);
nand U731 (N_731,N_680,N_656);
nand U732 (N_732,N_650,N_674);
or U733 (N_733,N_661,N_682);
nand U734 (N_734,N_656,N_689);
nor U735 (N_735,N_661,N_666);
nor U736 (N_736,N_669,N_696);
nor U737 (N_737,N_662,N_661);
xor U738 (N_738,N_668,N_684);
xor U739 (N_739,N_682,N_657);
nand U740 (N_740,N_688,N_680);
or U741 (N_741,N_655,N_658);
nor U742 (N_742,N_682,N_651);
xnor U743 (N_743,N_683,N_686);
nand U744 (N_744,N_657,N_674);
xnor U745 (N_745,N_659,N_673);
or U746 (N_746,N_668,N_653);
and U747 (N_747,N_659,N_688);
or U748 (N_748,N_682,N_679);
nor U749 (N_749,N_653,N_661);
xor U750 (N_750,N_734,N_718);
nor U751 (N_751,N_720,N_708);
nor U752 (N_752,N_703,N_709);
nand U753 (N_753,N_740,N_701);
and U754 (N_754,N_742,N_702);
and U755 (N_755,N_739,N_719);
nand U756 (N_756,N_745,N_711);
nor U757 (N_757,N_733,N_746);
or U758 (N_758,N_744,N_724);
xor U759 (N_759,N_706,N_715);
nor U760 (N_760,N_714,N_712);
or U761 (N_761,N_704,N_747);
nor U762 (N_762,N_723,N_722);
or U763 (N_763,N_748,N_749);
or U764 (N_764,N_705,N_700);
nor U765 (N_765,N_741,N_713);
nand U766 (N_766,N_730,N_710);
nand U767 (N_767,N_727,N_728);
xnor U768 (N_768,N_721,N_737);
nand U769 (N_769,N_743,N_738);
or U770 (N_770,N_731,N_732);
or U771 (N_771,N_716,N_735);
nor U772 (N_772,N_725,N_729);
or U773 (N_773,N_717,N_736);
xnor U774 (N_774,N_726,N_707);
nor U775 (N_775,N_703,N_704);
and U776 (N_776,N_712,N_737);
and U777 (N_777,N_707,N_736);
xnor U778 (N_778,N_743,N_742);
nand U779 (N_779,N_728,N_703);
nor U780 (N_780,N_726,N_703);
nand U781 (N_781,N_731,N_746);
nor U782 (N_782,N_704,N_741);
nor U783 (N_783,N_723,N_708);
nand U784 (N_784,N_719,N_742);
nor U785 (N_785,N_708,N_727);
nor U786 (N_786,N_709,N_726);
nand U787 (N_787,N_740,N_725);
xnor U788 (N_788,N_734,N_706);
and U789 (N_789,N_721,N_712);
and U790 (N_790,N_748,N_713);
xnor U791 (N_791,N_749,N_707);
xnor U792 (N_792,N_745,N_738);
nor U793 (N_793,N_708,N_714);
or U794 (N_794,N_736,N_714);
or U795 (N_795,N_720,N_710);
nor U796 (N_796,N_707,N_740);
and U797 (N_797,N_728,N_724);
xnor U798 (N_798,N_734,N_724);
nand U799 (N_799,N_715,N_749);
and U800 (N_800,N_770,N_764);
and U801 (N_801,N_782,N_791);
or U802 (N_802,N_761,N_778);
nor U803 (N_803,N_787,N_771);
xnor U804 (N_804,N_779,N_757);
or U805 (N_805,N_773,N_774);
and U806 (N_806,N_754,N_793);
nand U807 (N_807,N_756,N_799);
xor U808 (N_808,N_762,N_777);
and U809 (N_809,N_755,N_796);
and U810 (N_810,N_784,N_775);
or U811 (N_811,N_772,N_767);
and U812 (N_812,N_783,N_769);
nand U813 (N_813,N_763,N_758);
xor U814 (N_814,N_753,N_794);
and U815 (N_815,N_759,N_781);
and U816 (N_816,N_795,N_751);
and U817 (N_817,N_766,N_768);
or U818 (N_818,N_786,N_789);
xor U819 (N_819,N_765,N_797);
nand U820 (N_820,N_798,N_790);
nand U821 (N_821,N_788,N_785);
xnor U822 (N_822,N_750,N_752);
xor U823 (N_823,N_780,N_776);
or U824 (N_824,N_760,N_792);
xnor U825 (N_825,N_776,N_764);
nand U826 (N_826,N_780,N_790);
xnor U827 (N_827,N_758,N_776);
nor U828 (N_828,N_782,N_760);
or U829 (N_829,N_768,N_777);
xnor U830 (N_830,N_773,N_785);
or U831 (N_831,N_759,N_750);
and U832 (N_832,N_771,N_795);
or U833 (N_833,N_758,N_762);
xnor U834 (N_834,N_780,N_786);
or U835 (N_835,N_793,N_779);
nand U836 (N_836,N_754,N_768);
and U837 (N_837,N_767,N_796);
nor U838 (N_838,N_771,N_797);
or U839 (N_839,N_756,N_764);
nand U840 (N_840,N_755,N_782);
and U841 (N_841,N_782,N_754);
nor U842 (N_842,N_776,N_777);
nand U843 (N_843,N_796,N_776);
xor U844 (N_844,N_787,N_785);
or U845 (N_845,N_794,N_793);
nand U846 (N_846,N_784,N_774);
nor U847 (N_847,N_765,N_766);
nor U848 (N_848,N_781,N_772);
nand U849 (N_849,N_752,N_762);
or U850 (N_850,N_839,N_817);
nor U851 (N_851,N_807,N_800);
xnor U852 (N_852,N_810,N_801);
and U853 (N_853,N_835,N_804);
and U854 (N_854,N_844,N_823);
or U855 (N_855,N_811,N_816);
and U856 (N_856,N_829,N_820);
or U857 (N_857,N_821,N_843);
nor U858 (N_858,N_848,N_803);
nor U859 (N_859,N_827,N_849);
and U860 (N_860,N_826,N_841);
xor U861 (N_861,N_813,N_824);
and U862 (N_862,N_833,N_842);
xnor U863 (N_863,N_808,N_814);
nand U864 (N_864,N_845,N_840);
xor U865 (N_865,N_847,N_809);
or U866 (N_866,N_830,N_802);
nor U867 (N_867,N_825,N_836);
or U868 (N_868,N_846,N_818);
and U869 (N_869,N_832,N_806);
nor U870 (N_870,N_831,N_805);
and U871 (N_871,N_828,N_838);
nand U872 (N_872,N_815,N_819);
nor U873 (N_873,N_834,N_812);
and U874 (N_874,N_822,N_837);
nand U875 (N_875,N_838,N_814);
nand U876 (N_876,N_845,N_838);
or U877 (N_877,N_800,N_846);
or U878 (N_878,N_841,N_806);
nor U879 (N_879,N_829,N_825);
nor U880 (N_880,N_807,N_823);
nor U881 (N_881,N_810,N_812);
or U882 (N_882,N_825,N_841);
and U883 (N_883,N_825,N_839);
and U884 (N_884,N_808,N_848);
xnor U885 (N_885,N_802,N_818);
nand U886 (N_886,N_834,N_800);
xor U887 (N_887,N_832,N_822);
nand U888 (N_888,N_818,N_848);
or U889 (N_889,N_811,N_830);
or U890 (N_890,N_847,N_805);
nand U891 (N_891,N_846,N_810);
and U892 (N_892,N_819,N_825);
and U893 (N_893,N_840,N_818);
nor U894 (N_894,N_818,N_842);
nand U895 (N_895,N_822,N_812);
or U896 (N_896,N_819,N_842);
xor U897 (N_897,N_822,N_805);
and U898 (N_898,N_813,N_827);
and U899 (N_899,N_840,N_806);
or U900 (N_900,N_875,N_879);
and U901 (N_901,N_882,N_892);
nand U902 (N_902,N_884,N_888);
xor U903 (N_903,N_886,N_872);
nand U904 (N_904,N_895,N_880);
xor U905 (N_905,N_851,N_866);
or U906 (N_906,N_896,N_877);
nand U907 (N_907,N_857,N_852);
or U908 (N_908,N_850,N_863);
and U909 (N_909,N_862,N_893);
nor U910 (N_910,N_854,N_874);
nand U911 (N_911,N_897,N_870);
or U912 (N_912,N_890,N_894);
nor U913 (N_913,N_867,N_899);
nor U914 (N_914,N_859,N_883);
or U915 (N_915,N_860,N_881);
xnor U916 (N_916,N_868,N_898);
nand U917 (N_917,N_871,N_855);
or U918 (N_918,N_887,N_856);
and U919 (N_919,N_853,N_878);
nor U920 (N_920,N_858,N_885);
xor U921 (N_921,N_869,N_864);
nand U922 (N_922,N_861,N_873);
nor U923 (N_923,N_865,N_876);
and U924 (N_924,N_891,N_889);
xnor U925 (N_925,N_880,N_889);
or U926 (N_926,N_854,N_883);
or U927 (N_927,N_889,N_852);
xor U928 (N_928,N_896,N_889);
nor U929 (N_929,N_853,N_867);
nor U930 (N_930,N_891,N_861);
and U931 (N_931,N_873,N_898);
and U932 (N_932,N_877,N_899);
nor U933 (N_933,N_895,N_860);
and U934 (N_934,N_888,N_850);
xor U935 (N_935,N_866,N_871);
nand U936 (N_936,N_884,N_873);
and U937 (N_937,N_866,N_888);
xor U938 (N_938,N_862,N_886);
nand U939 (N_939,N_868,N_866);
nor U940 (N_940,N_890,N_878);
xor U941 (N_941,N_883,N_856);
or U942 (N_942,N_881,N_893);
xnor U943 (N_943,N_866,N_897);
nor U944 (N_944,N_871,N_885);
or U945 (N_945,N_866,N_859);
xnor U946 (N_946,N_881,N_884);
nand U947 (N_947,N_888,N_854);
nand U948 (N_948,N_862,N_880);
nor U949 (N_949,N_889,N_855);
nor U950 (N_950,N_934,N_926);
nor U951 (N_951,N_909,N_946);
and U952 (N_952,N_931,N_938);
nand U953 (N_953,N_928,N_906);
or U954 (N_954,N_941,N_945);
nor U955 (N_955,N_922,N_901);
or U956 (N_956,N_924,N_903);
or U957 (N_957,N_907,N_911);
nand U958 (N_958,N_915,N_916);
nor U959 (N_959,N_905,N_933);
and U960 (N_960,N_939,N_947);
xnor U961 (N_961,N_925,N_923);
nand U962 (N_962,N_949,N_921);
nand U963 (N_963,N_910,N_904);
or U964 (N_964,N_927,N_932);
and U965 (N_965,N_929,N_900);
nor U966 (N_966,N_920,N_944);
nor U967 (N_967,N_937,N_919);
and U968 (N_968,N_930,N_913);
or U969 (N_969,N_914,N_917);
xnor U970 (N_970,N_936,N_942);
nor U971 (N_971,N_935,N_902);
or U972 (N_972,N_943,N_912);
xor U973 (N_973,N_908,N_940);
xnor U974 (N_974,N_948,N_918);
nand U975 (N_975,N_925,N_907);
nand U976 (N_976,N_911,N_939);
xnor U977 (N_977,N_913,N_941);
xnor U978 (N_978,N_945,N_931);
xnor U979 (N_979,N_916,N_910);
nand U980 (N_980,N_934,N_933);
nand U981 (N_981,N_924,N_948);
nand U982 (N_982,N_937,N_949);
xnor U983 (N_983,N_909,N_942);
nor U984 (N_984,N_910,N_924);
or U985 (N_985,N_927,N_918);
nand U986 (N_986,N_938,N_908);
or U987 (N_987,N_912,N_927);
or U988 (N_988,N_925,N_924);
nand U989 (N_989,N_908,N_945);
or U990 (N_990,N_919,N_944);
nand U991 (N_991,N_907,N_916);
nand U992 (N_992,N_948,N_939);
nor U993 (N_993,N_923,N_933);
or U994 (N_994,N_921,N_910);
or U995 (N_995,N_941,N_930);
nand U996 (N_996,N_943,N_916);
xor U997 (N_997,N_922,N_913);
and U998 (N_998,N_906,N_914);
and U999 (N_999,N_903,N_907);
nor U1000 (N_1000,N_969,N_973);
or U1001 (N_1001,N_977,N_975);
xor U1002 (N_1002,N_970,N_990);
or U1003 (N_1003,N_991,N_966);
and U1004 (N_1004,N_999,N_952);
or U1005 (N_1005,N_996,N_980);
xor U1006 (N_1006,N_961,N_972);
nor U1007 (N_1007,N_987,N_957);
and U1008 (N_1008,N_974,N_953);
xnor U1009 (N_1009,N_959,N_958);
nand U1010 (N_1010,N_982,N_956);
nor U1011 (N_1011,N_976,N_981);
xor U1012 (N_1012,N_984,N_962);
xnor U1013 (N_1013,N_971,N_978);
nor U1014 (N_1014,N_998,N_951);
nor U1015 (N_1015,N_960,N_979);
nor U1016 (N_1016,N_950,N_986);
xor U1017 (N_1017,N_994,N_989);
and U1018 (N_1018,N_988,N_995);
xnor U1019 (N_1019,N_997,N_983);
nor U1020 (N_1020,N_965,N_993);
nand U1021 (N_1021,N_968,N_985);
or U1022 (N_1022,N_992,N_954);
and U1023 (N_1023,N_967,N_964);
or U1024 (N_1024,N_955,N_963);
nor U1025 (N_1025,N_972,N_986);
and U1026 (N_1026,N_986,N_976);
xor U1027 (N_1027,N_965,N_979);
or U1028 (N_1028,N_993,N_976);
or U1029 (N_1029,N_999,N_983);
nor U1030 (N_1030,N_954,N_997);
xor U1031 (N_1031,N_950,N_961);
nor U1032 (N_1032,N_963,N_999);
nand U1033 (N_1033,N_967,N_966);
nand U1034 (N_1034,N_994,N_987);
xnor U1035 (N_1035,N_971,N_962);
or U1036 (N_1036,N_967,N_969);
xor U1037 (N_1037,N_984,N_977);
and U1038 (N_1038,N_959,N_966);
xnor U1039 (N_1039,N_994,N_996);
xnor U1040 (N_1040,N_971,N_977);
and U1041 (N_1041,N_952,N_990);
and U1042 (N_1042,N_985,N_952);
or U1043 (N_1043,N_961,N_969);
or U1044 (N_1044,N_982,N_974);
nor U1045 (N_1045,N_999,N_988);
and U1046 (N_1046,N_987,N_975);
xnor U1047 (N_1047,N_956,N_999);
nand U1048 (N_1048,N_974,N_997);
xnor U1049 (N_1049,N_952,N_983);
xor U1050 (N_1050,N_1003,N_1047);
nand U1051 (N_1051,N_1027,N_1008);
xnor U1052 (N_1052,N_1033,N_1007);
xnor U1053 (N_1053,N_1042,N_1022);
xor U1054 (N_1054,N_1005,N_1001);
xor U1055 (N_1055,N_1045,N_1006);
xnor U1056 (N_1056,N_1012,N_1018);
nand U1057 (N_1057,N_1028,N_1040);
or U1058 (N_1058,N_1020,N_1048);
nor U1059 (N_1059,N_1019,N_1016);
nor U1060 (N_1060,N_1049,N_1034);
xnor U1061 (N_1061,N_1002,N_1000);
and U1062 (N_1062,N_1041,N_1038);
xnor U1063 (N_1063,N_1031,N_1043);
and U1064 (N_1064,N_1037,N_1011);
nand U1065 (N_1065,N_1023,N_1039);
nand U1066 (N_1066,N_1009,N_1004);
or U1067 (N_1067,N_1036,N_1014);
nor U1068 (N_1068,N_1044,N_1032);
nand U1069 (N_1069,N_1026,N_1013);
nand U1070 (N_1070,N_1024,N_1015);
or U1071 (N_1071,N_1017,N_1030);
nand U1072 (N_1072,N_1029,N_1010);
nor U1073 (N_1073,N_1035,N_1021);
or U1074 (N_1074,N_1025,N_1046);
nand U1075 (N_1075,N_1002,N_1003);
xor U1076 (N_1076,N_1005,N_1041);
xor U1077 (N_1077,N_1044,N_1043);
xor U1078 (N_1078,N_1038,N_1007);
and U1079 (N_1079,N_1030,N_1020);
or U1080 (N_1080,N_1029,N_1003);
nor U1081 (N_1081,N_1038,N_1036);
or U1082 (N_1082,N_1010,N_1036);
nand U1083 (N_1083,N_1038,N_1015);
or U1084 (N_1084,N_1000,N_1028);
nor U1085 (N_1085,N_1028,N_1013);
nand U1086 (N_1086,N_1027,N_1029);
nor U1087 (N_1087,N_1040,N_1018);
or U1088 (N_1088,N_1026,N_1030);
or U1089 (N_1089,N_1022,N_1005);
xnor U1090 (N_1090,N_1042,N_1018);
nor U1091 (N_1091,N_1017,N_1033);
xnor U1092 (N_1092,N_1017,N_1048);
nand U1093 (N_1093,N_1029,N_1011);
nor U1094 (N_1094,N_1047,N_1037);
or U1095 (N_1095,N_1024,N_1046);
nand U1096 (N_1096,N_1009,N_1013);
or U1097 (N_1097,N_1038,N_1022);
or U1098 (N_1098,N_1041,N_1010);
and U1099 (N_1099,N_1021,N_1045);
xor U1100 (N_1100,N_1089,N_1087);
nor U1101 (N_1101,N_1061,N_1059);
nor U1102 (N_1102,N_1070,N_1062);
or U1103 (N_1103,N_1068,N_1057);
nand U1104 (N_1104,N_1065,N_1095);
nand U1105 (N_1105,N_1071,N_1096);
or U1106 (N_1106,N_1066,N_1054);
nor U1107 (N_1107,N_1067,N_1053);
nand U1108 (N_1108,N_1097,N_1099);
nand U1109 (N_1109,N_1055,N_1098);
nand U1110 (N_1110,N_1084,N_1076);
nand U1111 (N_1111,N_1069,N_1074);
and U1112 (N_1112,N_1051,N_1092);
nor U1113 (N_1113,N_1064,N_1050);
or U1114 (N_1114,N_1063,N_1080);
nor U1115 (N_1115,N_1082,N_1085);
nor U1116 (N_1116,N_1052,N_1078);
nand U1117 (N_1117,N_1079,N_1083);
and U1118 (N_1118,N_1058,N_1075);
and U1119 (N_1119,N_1081,N_1086);
xor U1120 (N_1120,N_1056,N_1093);
and U1121 (N_1121,N_1072,N_1060);
nand U1122 (N_1122,N_1088,N_1094);
nand U1123 (N_1123,N_1091,N_1073);
xnor U1124 (N_1124,N_1090,N_1077);
or U1125 (N_1125,N_1072,N_1064);
and U1126 (N_1126,N_1079,N_1063);
nand U1127 (N_1127,N_1054,N_1052);
or U1128 (N_1128,N_1054,N_1060);
nand U1129 (N_1129,N_1060,N_1092);
nor U1130 (N_1130,N_1066,N_1057);
nor U1131 (N_1131,N_1063,N_1078);
nand U1132 (N_1132,N_1072,N_1071);
nand U1133 (N_1133,N_1084,N_1083);
and U1134 (N_1134,N_1069,N_1078);
xnor U1135 (N_1135,N_1091,N_1053);
nand U1136 (N_1136,N_1076,N_1062);
nand U1137 (N_1137,N_1081,N_1064);
nor U1138 (N_1138,N_1080,N_1097);
nand U1139 (N_1139,N_1094,N_1055);
nor U1140 (N_1140,N_1082,N_1075);
nand U1141 (N_1141,N_1083,N_1065);
nand U1142 (N_1142,N_1050,N_1059);
or U1143 (N_1143,N_1057,N_1099);
or U1144 (N_1144,N_1082,N_1094);
nor U1145 (N_1145,N_1091,N_1092);
nor U1146 (N_1146,N_1083,N_1050);
nor U1147 (N_1147,N_1060,N_1069);
xnor U1148 (N_1148,N_1096,N_1089);
xor U1149 (N_1149,N_1094,N_1068);
and U1150 (N_1150,N_1108,N_1147);
and U1151 (N_1151,N_1131,N_1149);
xor U1152 (N_1152,N_1140,N_1136);
and U1153 (N_1153,N_1104,N_1100);
nand U1154 (N_1154,N_1121,N_1106);
xnor U1155 (N_1155,N_1115,N_1137);
nor U1156 (N_1156,N_1135,N_1112);
or U1157 (N_1157,N_1117,N_1142);
or U1158 (N_1158,N_1130,N_1129);
and U1159 (N_1159,N_1114,N_1110);
xnor U1160 (N_1160,N_1124,N_1143);
nand U1161 (N_1161,N_1141,N_1146);
xor U1162 (N_1162,N_1138,N_1123);
and U1163 (N_1163,N_1111,N_1109);
xor U1164 (N_1164,N_1120,N_1105);
nand U1165 (N_1165,N_1116,N_1139);
nor U1166 (N_1166,N_1118,N_1127);
nor U1167 (N_1167,N_1145,N_1126);
xor U1168 (N_1168,N_1128,N_1148);
xor U1169 (N_1169,N_1107,N_1125);
nor U1170 (N_1170,N_1134,N_1144);
or U1171 (N_1171,N_1122,N_1101);
nor U1172 (N_1172,N_1133,N_1113);
nand U1173 (N_1173,N_1103,N_1102);
or U1174 (N_1174,N_1132,N_1119);
xor U1175 (N_1175,N_1122,N_1139);
nor U1176 (N_1176,N_1129,N_1137);
or U1177 (N_1177,N_1145,N_1133);
nand U1178 (N_1178,N_1115,N_1107);
xnor U1179 (N_1179,N_1120,N_1139);
nor U1180 (N_1180,N_1146,N_1102);
or U1181 (N_1181,N_1133,N_1142);
xor U1182 (N_1182,N_1126,N_1116);
xnor U1183 (N_1183,N_1124,N_1132);
and U1184 (N_1184,N_1145,N_1110);
xnor U1185 (N_1185,N_1134,N_1148);
or U1186 (N_1186,N_1122,N_1118);
xnor U1187 (N_1187,N_1132,N_1127);
xor U1188 (N_1188,N_1123,N_1106);
or U1189 (N_1189,N_1136,N_1117);
nand U1190 (N_1190,N_1101,N_1109);
and U1191 (N_1191,N_1108,N_1100);
xnor U1192 (N_1192,N_1136,N_1122);
nor U1193 (N_1193,N_1127,N_1129);
xnor U1194 (N_1194,N_1129,N_1138);
and U1195 (N_1195,N_1101,N_1110);
xnor U1196 (N_1196,N_1109,N_1113);
nand U1197 (N_1197,N_1110,N_1134);
nand U1198 (N_1198,N_1144,N_1129);
nor U1199 (N_1199,N_1122,N_1138);
xor U1200 (N_1200,N_1192,N_1150);
nor U1201 (N_1201,N_1179,N_1153);
nand U1202 (N_1202,N_1166,N_1173);
nand U1203 (N_1203,N_1171,N_1154);
and U1204 (N_1204,N_1180,N_1177);
and U1205 (N_1205,N_1167,N_1157);
and U1206 (N_1206,N_1182,N_1174);
and U1207 (N_1207,N_1160,N_1194);
or U1208 (N_1208,N_1198,N_1151);
xnor U1209 (N_1209,N_1175,N_1159);
and U1210 (N_1210,N_1176,N_1185);
nand U1211 (N_1211,N_1152,N_1170);
nand U1212 (N_1212,N_1158,N_1156);
nor U1213 (N_1213,N_1163,N_1186);
or U1214 (N_1214,N_1168,N_1188);
nand U1215 (N_1215,N_1199,N_1190);
nand U1216 (N_1216,N_1191,N_1161);
nand U1217 (N_1217,N_1195,N_1184);
nor U1218 (N_1218,N_1183,N_1165);
and U1219 (N_1219,N_1172,N_1162);
xor U1220 (N_1220,N_1178,N_1187);
xnor U1221 (N_1221,N_1169,N_1155);
xnor U1222 (N_1222,N_1181,N_1189);
xnor U1223 (N_1223,N_1196,N_1193);
and U1224 (N_1224,N_1197,N_1164);
xnor U1225 (N_1225,N_1182,N_1188);
nor U1226 (N_1226,N_1183,N_1151);
or U1227 (N_1227,N_1151,N_1194);
nor U1228 (N_1228,N_1194,N_1170);
or U1229 (N_1229,N_1194,N_1197);
and U1230 (N_1230,N_1193,N_1168);
nand U1231 (N_1231,N_1189,N_1163);
xor U1232 (N_1232,N_1172,N_1180);
and U1233 (N_1233,N_1175,N_1165);
or U1234 (N_1234,N_1192,N_1183);
and U1235 (N_1235,N_1157,N_1178);
and U1236 (N_1236,N_1196,N_1186);
nor U1237 (N_1237,N_1186,N_1184);
or U1238 (N_1238,N_1159,N_1192);
or U1239 (N_1239,N_1193,N_1167);
xor U1240 (N_1240,N_1166,N_1162);
nand U1241 (N_1241,N_1196,N_1154);
or U1242 (N_1242,N_1156,N_1161);
or U1243 (N_1243,N_1173,N_1177);
nand U1244 (N_1244,N_1161,N_1150);
or U1245 (N_1245,N_1159,N_1158);
and U1246 (N_1246,N_1154,N_1157);
or U1247 (N_1247,N_1193,N_1197);
xnor U1248 (N_1248,N_1152,N_1158);
and U1249 (N_1249,N_1180,N_1192);
or U1250 (N_1250,N_1213,N_1201);
or U1251 (N_1251,N_1215,N_1218);
nor U1252 (N_1252,N_1222,N_1203);
nand U1253 (N_1253,N_1230,N_1227);
nand U1254 (N_1254,N_1236,N_1235);
nor U1255 (N_1255,N_1209,N_1233);
or U1256 (N_1256,N_1206,N_1216);
nor U1257 (N_1257,N_1231,N_1229);
xor U1258 (N_1258,N_1220,N_1238);
xnor U1259 (N_1259,N_1239,N_1244);
or U1260 (N_1260,N_1232,N_1225);
nand U1261 (N_1261,N_1249,N_1214);
nor U1262 (N_1262,N_1240,N_1241);
xnor U1263 (N_1263,N_1207,N_1246);
and U1264 (N_1264,N_1210,N_1202);
nor U1265 (N_1265,N_1212,N_1224);
or U1266 (N_1266,N_1243,N_1217);
xnor U1267 (N_1267,N_1242,N_1234);
or U1268 (N_1268,N_1219,N_1223);
and U1269 (N_1269,N_1245,N_1205);
xnor U1270 (N_1270,N_1211,N_1247);
nand U1271 (N_1271,N_1237,N_1204);
nor U1272 (N_1272,N_1228,N_1221);
nor U1273 (N_1273,N_1208,N_1248);
nand U1274 (N_1274,N_1200,N_1226);
nand U1275 (N_1275,N_1204,N_1210);
nor U1276 (N_1276,N_1214,N_1219);
and U1277 (N_1277,N_1214,N_1241);
and U1278 (N_1278,N_1223,N_1241);
xor U1279 (N_1279,N_1215,N_1204);
xnor U1280 (N_1280,N_1243,N_1211);
or U1281 (N_1281,N_1209,N_1205);
or U1282 (N_1282,N_1236,N_1239);
xor U1283 (N_1283,N_1216,N_1211);
xor U1284 (N_1284,N_1221,N_1233);
or U1285 (N_1285,N_1248,N_1200);
or U1286 (N_1286,N_1205,N_1204);
nor U1287 (N_1287,N_1200,N_1236);
and U1288 (N_1288,N_1246,N_1241);
and U1289 (N_1289,N_1241,N_1211);
xnor U1290 (N_1290,N_1215,N_1234);
and U1291 (N_1291,N_1204,N_1213);
nor U1292 (N_1292,N_1243,N_1221);
nand U1293 (N_1293,N_1216,N_1220);
and U1294 (N_1294,N_1243,N_1237);
nor U1295 (N_1295,N_1245,N_1216);
xnor U1296 (N_1296,N_1240,N_1229);
nand U1297 (N_1297,N_1229,N_1214);
and U1298 (N_1298,N_1222,N_1234);
or U1299 (N_1299,N_1237,N_1221);
nand U1300 (N_1300,N_1294,N_1291);
nand U1301 (N_1301,N_1286,N_1262);
or U1302 (N_1302,N_1255,N_1284);
or U1303 (N_1303,N_1274,N_1281);
nand U1304 (N_1304,N_1293,N_1264);
and U1305 (N_1305,N_1283,N_1258);
nand U1306 (N_1306,N_1271,N_1280);
nor U1307 (N_1307,N_1275,N_1259);
xnor U1308 (N_1308,N_1266,N_1298);
xor U1309 (N_1309,N_1277,N_1287);
nand U1310 (N_1310,N_1297,N_1289);
xor U1311 (N_1311,N_1285,N_1252);
and U1312 (N_1312,N_1288,N_1290);
xor U1313 (N_1313,N_1263,N_1251);
or U1314 (N_1314,N_1278,N_1295);
and U1315 (N_1315,N_1299,N_1270);
nand U1316 (N_1316,N_1296,N_1254);
and U1317 (N_1317,N_1261,N_1250);
nor U1318 (N_1318,N_1292,N_1279);
xor U1319 (N_1319,N_1267,N_1265);
nand U1320 (N_1320,N_1268,N_1282);
nor U1321 (N_1321,N_1253,N_1256);
nor U1322 (N_1322,N_1260,N_1273);
xor U1323 (N_1323,N_1269,N_1272);
nor U1324 (N_1324,N_1257,N_1276);
nor U1325 (N_1325,N_1278,N_1261);
xnor U1326 (N_1326,N_1260,N_1284);
nand U1327 (N_1327,N_1274,N_1269);
nand U1328 (N_1328,N_1298,N_1294);
nor U1329 (N_1329,N_1257,N_1296);
xnor U1330 (N_1330,N_1299,N_1281);
xor U1331 (N_1331,N_1298,N_1250);
or U1332 (N_1332,N_1272,N_1290);
xnor U1333 (N_1333,N_1271,N_1257);
xor U1334 (N_1334,N_1289,N_1253);
nor U1335 (N_1335,N_1277,N_1251);
nor U1336 (N_1336,N_1284,N_1281);
xnor U1337 (N_1337,N_1251,N_1259);
and U1338 (N_1338,N_1296,N_1297);
nor U1339 (N_1339,N_1269,N_1295);
nand U1340 (N_1340,N_1275,N_1263);
or U1341 (N_1341,N_1269,N_1268);
nor U1342 (N_1342,N_1268,N_1294);
xnor U1343 (N_1343,N_1269,N_1252);
and U1344 (N_1344,N_1284,N_1280);
xnor U1345 (N_1345,N_1285,N_1257);
and U1346 (N_1346,N_1261,N_1251);
or U1347 (N_1347,N_1267,N_1264);
nand U1348 (N_1348,N_1290,N_1285);
nor U1349 (N_1349,N_1294,N_1287);
nand U1350 (N_1350,N_1310,N_1343);
and U1351 (N_1351,N_1301,N_1319);
xnor U1352 (N_1352,N_1303,N_1312);
or U1353 (N_1353,N_1306,N_1320);
nor U1354 (N_1354,N_1349,N_1326);
nor U1355 (N_1355,N_1347,N_1333);
and U1356 (N_1356,N_1328,N_1332);
or U1357 (N_1357,N_1314,N_1327);
nand U1358 (N_1358,N_1302,N_1313);
nor U1359 (N_1359,N_1308,N_1331);
and U1360 (N_1360,N_1344,N_1321);
or U1361 (N_1361,N_1300,N_1336);
and U1362 (N_1362,N_1335,N_1339);
nand U1363 (N_1363,N_1329,N_1323);
nand U1364 (N_1364,N_1318,N_1304);
nand U1365 (N_1365,N_1340,N_1311);
and U1366 (N_1366,N_1317,N_1346);
nor U1367 (N_1367,N_1338,N_1309);
nor U1368 (N_1368,N_1322,N_1341);
or U1369 (N_1369,N_1348,N_1330);
or U1370 (N_1370,N_1316,N_1334);
xnor U1371 (N_1371,N_1315,N_1342);
or U1372 (N_1372,N_1307,N_1324);
nand U1373 (N_1373,N_1305,N_1325);
nand U1374 (N_1374,N_1337,N_1345);
nand U1375 (N_1375,N_1302,N_1319);
nor U1376 (N_1376,N_1323,N_1345);
nor U1377 (N_1377,N_1322,N_1308);
nand U1378 (N_1378,N_1316,N_1301);
and U1379 (N_1379,N_1347,N_1305);
or U1380 (N_1380,N_1334,N_1349);
and U1381 (N_1381,N_1314,N_1325);
nor U1382 (N_1382,N_1329,N_1309);
xor U1383 (N_1383,N_1311,N_1314);
xnor U1384 (N_1384,N_1305,N_1327);
xnor U1385 (N_1385,N_1331,N_1347);
nand U1386 (N_1386,N_1308,N_1349);
nand U1387 (N_1387,N_1337,N_1331);
nand U1388 (N_1388,N_1312,N_1329);
or U1389 (N_1389,N_1319,N_1318);
xnor U1390 (N_1390,N_1345,N_1331);
nor U1391 (N_1391,N_1309,N_1308);
xnor U1392 (N_1392,N_1343,N_1327);
nand U1393 (N_1393,N_1329,N_1306);
nand U1394 (N_1394,N_1333,N_1316);
nand U1395 (N_1395,N_1318,N_1300);
and U1396 (N_1396,N_1306,N_1338);
nand U1397 (N_1397,N_1318,N_1306);
and U1398 (N_1398,N_1340,N_1327);
nor U1399 (N_1399,N_1323,N_1340);
and U1400 (N_1400,N_1377,N_1370);
nor U1401 (N_1401,N_1399,N_1391);
nand U1402 (N_1402,N_1379,N_1394);
xnor U1403 (N_1403,N_1381,N_1393);
nand U1404 (N_1404,N_1350,N_1383);
and U1405 (N_1405,N_1363,N_1373);
or U1406 (N_1406,N_1390,N_1388);
nor U1407 (N_1407,N_1369,N_1365);
or U1408 (N_1408,N_1368,N_1359);
xor U1409 (N_1409,N_1355,N_1395);
nand U1410 (N_1410,N_1382,N_1392);
nand U1411 (N_1411,N_1396,N_1361);
nor U1412 (N_1412,N_1375,N_1374);
nor U1413 (N_1413,N_1367,N_1352);
or U1414 (N_1414,N_1385,N_1357);
xnor U1415 (N_1415,N_1371,N_1380);
nand U1416 (N_1416,N_1366,N_1351);
nand U1417 (N_1417,N_1364,N_1389);
xor U1418 (N_1418,N_1360,N_1362);
xor U1419 (N_1419,N_1372,N_1356);
nand U1420 (N_1420,N_1378,N_1353);
nand U1421 (N_1421,N_1387,N_1398);
nor U1422 (N_1422,N_1397,N_1386);
and U1423 (N_1423,N_1376,N_1354);
or U1424 (N_1424,N_1358,N_1384);
nor U1425 (N_1425,N_1364,N_1370);
and U1426 (N_1426,N_1390,N_1385);
nand U1427 (N_1427,N_1358,N_1391);
and U1428 (N_1428,N_1350,N_1382);
nor U1429 (N_1429,N_1388,N_1394);
nor U1430 (N_1430,N_1367,N_1386);
or U1431 (N_1431,N_1387,N_1394);
or U1432 (N_1432,N_1373,N_1354);
xor U1433 (N_1433,N_1379,N_1364);
nand U1434 (N_1434,N_1367,N_1363);
nand U1435 (N_1435,N_1368,N_1397);
xor U1436 (N_1436,N_1365,N_1360);
xor U1437 (N_1437,N_1350,N_1378);
nand U1438 (N_1438,N_1355,N_1352);
nor U1439 (N_1439,N_1363,N_1353);
nor U1440 (N_1440,N_1359,N_1374);
nor U1441 (N_1441,N_1356,N_1376);
and U1442 (N_1442,N_1387,N_1355);
and U1443 (N_1443,N_1387,N_1360);
and U1444 (N_1444,N_1351,N_1388);
nor U1445 (N_1445,N_1376,N_1398);
nor U1446 (N_1446,N_1395,N_1368);
nor U1447 (N_1447,N_1394,N_1354);
and U1448 (N_1448,N_1394,N_1364);
or U1449 (N_1449,N_1378,N_1360);
or U1450 (N_1450,N_1420,N_1409);
nand U1451 (N_1451,N_1408,N_1400);
nand U1452 (N_1452,N_1427,N_1412);
nor U1453 (N_1453,N_1431,N_1401);
nor U1454 (N_1454,N_1443,N_1419);
and U1455 (N_1455,N_1434,N_1441);
nor U1456 (N_1456,N_1444,N_1445);
nor U1457 (N_1457,N_1426,N_1403);
or U1458 (N_1458,N_1423,N_1447);
and U1459 (N_1459,N_1424,N_1416);
or U1460 (N_1460,N_1421,N_1407);
xnor U1461 (N_1461,N_1402,N_1428);
nor U1462 (N_1462,N_1429,N_1430);
nand U1463 (N_1463,N_1418,N_1405);
nor U1464 (N_1464,N_1417,N_1425);
nand U1465 (N_1465,N_1446,N_1439);
and U1466 (N_1466,N_1411,N_1435);
nand U1467 (N_1467,N_1406,N_1436);
nand U1468 (N_1468,N_1410,N_1440);
nor U1469 (N_1469,N_1404,N_1442);
xor U1470 (N_1470,N_1414,N_1438);
xor U1471 (N_1471,N_1433,N_1422);
or U1472 (N_1472,N_1449,N_1415);
xor U1473 (N_1473,N_1413,N_1432);
and U1474 (N_1474,N_1448,N_1437);
nand U1475 (N_1475,N_1408,N_1426);
and U1476 (N_1476,N_1418,N_1413);
and U1477 (N_1477,N_1409,N_1415);
nand U1478 (N_1478,N_1404,N_1449);
xor U1479 (N_1479,N_1419,N_1428);
nand U1480 (N_1480,N_1422,N_1400);
nand U1481 (N_1481,N_1421,N_1430);
nand U1482 (N_1482,N_1410,N_1430);
nor U1483 (N_1483,N_1420,N_1417);
xor U1484 (N_1484,N_1442,N_1426);
xnor U1485 (N_1485,N_1438,N_1433);
xor U1486 (N_1486,N_1431,N_1404);
nor U1487 (N_1487,N_1414,N_1442);
xnor U1488 (N_1488,N_1425,N_1446);
or U1489 (N_1489,N_1420,N_1418);
nand U1490 (N_1490,N_1413,N_1449);
nand U1491 (N_1491,N_1432,N_1433);
nor U1492 (N_1492,N_1435,N_1415);
xnor U1493 (N_1493,N_1428,N_1444);
nand U1494 (N_1494,N_1425,N_1424);
or U1495 (N_1495,N_1426,N_1432);
xnor U1496 (N_1496,N_1449,N_1420);
and U1497 (N_1497,N_1402,N_1415);
nand U1498 (N_1498,N_1438,N_1422);
and U1499 (N_1499,N_1437,N_1433);
xor U1500 (N_1500,N_1489,N_1461);
or U1501 (N_1501,N_1490,N_1473);
xor U1502 (N_1502,N_1472,N_1462);
nand U1503 (N_1503,N_1451,N_1465);
xor U1504 (N_1504,N_1458,N_1466);
and U1505 (N_1505,N_1474,N_1498);
nor U1506 (N_1506,N_1467,N_1450);
nand U1507 (N_1507,N_1469,N_1495);
and U1508 (N_1508,N_1483,N_1491);
xnor U1509 (N_1509,N_1493,N_1499);
nor U1510 (N_1510,N_1480,N_1496);
nor U1511 (N_1511,N_1479,N_1471);
or U1512 (N_1512,N_1454,N_1494);
xnor U1513 (N_1513,N_1485,N_1455);
nor U1514 (N_1514,N_1452,N_1463);
nor U1515 (N_1515,N_1453,N_1497);
or U1516 (N_1516,N_1484,N_1478);
nand U1517 (N_1517,N_1459,N_1464);
or U1518 (N_1518,N_1456,N_1470);
or U1519 (N_1519,N_1475,N_1468);
nor U1520 (N_1520,N_1477,N_1487);
and U1521 (N_1521,N_1492,N_1460);
xor U1522 (N_1522,N_1476,N_1481);
xnor U1523 (N_1523,N_1457,N_1482);
and U1524 (N_1524,N_1486,N_1488);
nor U1525 (N_1525,N_1463,N_1482);
or U1526 (N_1526,N_1490,N_1482);
and U1527 (N_1527,N_1455,N_1457);
nand U1528 (N_1528,N_1475,N_1454);
nand U1529 (N_1529,N_1478,N_1473);
nor U1530 (N_1530,N_1477,N_1456);
or U1531 (N_1531,N_1474,N_1483);
nand U1532 (N_1532,N_1496,N_1450);
nor U1533 (N_1533,N_1453,N_1482);
or U1534 (N_1534,N_1459,N_1456);
and U1535 (N_1535,N_1471,N_1478);
or U1536 (N_1536,N_1463,N_1455);
nor U1537 (N_1537,N_1464,N_1481);
nand U1538 (N_1538,N_1484,N_1464);
nand U1539 (N_1539,N_1466,N_1484);
xor U1540 (N_1540,N_1476,N_1451);
nand U1541 (N_1541,N_1456,N_1469);
nor U1542 (N_1542,N_1484,N_1460);
or U1543 (N_1543,N_1479,N_1456);
or U1544 (N_1544,N_1493,N_1466);
nor U1545 (N_1545,N_1464,N_1475);
and U1546 (N_1546,N_1468,N_1467);
and U1547 (N_1547,N_1467,N_1487);
or U1548 (N_1548,N_1490,N_1452);
and U1549 (N_1549,N_1463,N_1457);
and U1550 (N_1550,N_1533,N_1500);
xor U1551 (N_1551,N_1545,N_1509);
nand U1552 (N_1552,N_1538,N_1511);
xor U1553 (N_1553,N_1528,N_1544);
or U1554 (N_1554,N_1539,N_1512);
or U1555 (N_1555,N_1526,N_1530);
or U1556 (N_1556,N_1531,N_1521);
and U1557 (N_1557,N_1527,N_1516);
or U1558 (N_1558,N_1517,N_1543);
xnor U1559 (N_1559,N_1524,N_1541);
xnor U1560 (N_1560,N_1506,N_1534);
nand U1561 (N_1561,N_1515,N_1501);
and U1562 (N_1562,N_1535,N_1523);
xnor U1563 (N_1563,N_1548,N_1504);
or U1564 (N_1564,N_1508,N_1513);
nand U1565 (N_1565,N_1514,N_1503);
nand U1566 (N_1566,N_1542,N_1546);
nor U1567 (N_1567,N_1532,N_1520);
nand U1568 (N_1568,N_1525,N_1510);
nand U1569 (N_1569,N_1549,N_1529);
nor U1570 (N_1570,N_1540,N_1522);
or U1571 (N_1571,N_1519,N_1507);
and U1572 (N_1572,N_1502,N_1536);
or U1573 (N_1573,N_1518,N_1547);
nand U1574 (N_1574,N_1537,N_1505);
nor U1575 (N_1575,N_1531,N_1524);
nor U1576 (N_1576,N_1534,N_1533);
xnor U1577 (N_1577,N_1542,N_1510);
or U1578 (N_1578,N_1515,N_1530);
and U1579 (N_1579,N_1535,N_1530);
nor U1580 (N_1580,N_1507,N_1500);
nor U1581 (N_1581,N_1528,N_1543);
and U1582 (N_1582,N_1501,N_1532);
xnor U1583 (N_1583,N_1506,N_1511);
nand U1584 (N_1584,N_1540,N_1521);
and U1585 (N_1585,N_1540,N_1507);
or U1586 (N_1586,N_1524,N_1547);
and U1587 (N_1587,N_1512,N_1507);
xnor U1588 (N_1588,N_1538,N_1523);
xnor U1589 (N_1589,N_1541,N_1502);
nand U1590 (N_1590,N_1539,N_1514);
or U1591 (N_1591,N_1534,N_1544);
xor U1592 (N_1592,N_1517,N_1534);
nor U1593 (N_1593,N_1508,N_1521);
nand U1594 (N_1594,N_1525,N_1545);
and U1595 (N_1595,N_1537,N_1538);
nand U1596 (N_1596,N_1501,N_1530);
xnor U1597 (N_1597,N_1508,N_1545);
and U1598 (N_1598,N_1502,N_1518);
nor U1599 (N_1599,N_1525,N_1548);
nor U1600 (N_1600,N_1590,N_1584);
or U1601 (N_1601,N_1598,N_1579);
or U1602 (N_1602,N_1566,N_1555);
nor U1603 (N_1603,N_1550,N_1594);
or U1604 (N_1604,N_1571,N_1589);
xnor U1605 (N_1605,N_1573,N_1596);
nor U1606 (N_1606,N_1578,N_1552);
nor U1607 (N_1607,N_1556,N_1560);
or U1608 (N_1608,N_1581,N_1572);
and U1609 (N_1609,N_1554,N_1564);
nor U1610 (N_1610,N_1585,N_1559);
or U1611 (N_1611,N_1595,N_1586);
nor U1612 (N_1612,N_1582,N_1562);
nor U1613 (N_1613,N_1563,N_1587);
xnor U1614 (N_1614,N_1553,N_1576);
nand U1615 (N_1615,N_1591,N_1575);
nand U1616 (N_1616,N_1565,N_1599);
and U1617 (N_1617,N_1580,N_1558);
and U1618 (N_1618,N_1561,N_1583);
xnor U1619 (N_1619,N_1592,N_1570);
nor U1620 (N_1620,N_1588,N_1597);
or U1621 (N_1621,N_1557,N_1551);
nand U1622 (N_1622,N_1574,N_1568);
nand U1623 (N_1623,N_1577,N_1593);
and U1624 (N_1624,N_1569,N_1567);
xor U1625 (N_1625,N_1550,N_1572);
xnor U1626 (N_1626,N_1568,N_1595);
xnor U1627 (N_1627,N_1597,N_1576);
nor U1628 (N_1628,N_1582,N_1552);
xnor U1629 (N_1629,N_1579,N_1593);
nor U1630 (N_1630,N_1553,N_1582);
nor U1631 (N_1631,N_1550,N_1554);
or U1632 (N_1632,N_1591,N_1598);
or U1633 (N_1633,N_1589,N_1594);
nor U1634 (N_1634,N_1594,N_1557);
and U1635 (N_1635,N_1570,N_1551);
nand U1636 (N_1636,N_1567,N_1575);
nand U1637 (N_1637,N_1576,N_1590);
nand U1638 (N_1638,N_1558,N_1557);
xor U1639 (N_1639,N_1553,N_1587);
nand U1640 (N_1640,N_1579,N_1554);
nand U1641 (N_1641,N_1587,N_1552);
nand U1642 (N_1642,N_1552,N_1551);
or U1643 (N_1643,N_1551,N_1592);
nand U1644 (N_1644,N_1552,N_1568);
nand U1645 (N_1645,N_1578,N_1577);
or U1646 (N_1646,N_1583,N_1595);
nor U1647 (N_1647,N_1557,N_1588);
xnor U1648 (N_1648,N_1558,N_1588);
or U1649 (N_1649,N_1559,N_1582);
nand U1650 (N_1650,N_1646,N_1619);
nor U1651 (N_1651,N_1611,N_1630);
nor U1652 (N_1652,N_1644,N_1626);
or U1653 (N_1653,N_1628,N_1636);
or U1654 (N_1654,N_1618,N_1607);
or U1655 (N_1655,N_1609,N_1601);
nand U1656 (N_1656,N_1627,N_1649);
nand U1657 (N_1657,N_1606,N_1638);
xor U1658 (N_1658,N_1645,N_1617);
nand U1659 (N_1659,N_1640,N_1600);
and U1660 (N_1660,N_1639,N_1610);
nand U1661 (N_1661,N_1631,N_1625);
xor U1662 (N_1662,N_1608,N_1616);
nand U1663 (N_1663,N_1604,N_1647);
nor U1664 (N_1664,N_1642,N_1614);
nor U1665 (N_1665,N_1603,N_1635);
nor U1666 (N_1666,N_1615,N_1622);
or U1667 (N_1667,N_1641,N_1629);
nand U1668 (N_1668,N_1623,N_1602);
xnor U1669 (N_1669,N_1633,N_1632);
nand U1670 (N_1670,N_1613,N_1624);
or U1671 (N_1671,N_1620,N_1634);
or U1672 (N_1672,N_1621,N_1648);
nand U1673 (N_1673,N_1612,N_1643);
or U1674 (N_1674,N_1605,N_1637);
xor U1675 (N_1675,N_1635,N_1623);
nor U1676 (N_1676,N_1643,N_1608);
nor U1677 (N_1677,N_1620,N_1640);
nor U1678 (N_1678,N_1617,N_1632);
or U1679 (N_1679,N_1624,N_1622);
and U1680 (N_1680,N_1619,N_1621);
nor U1681 (N_1681,N_1616,N_1629);
or U1682 (N_1682,N_1601,N_1629);
nand U1683 (N_1683,N_1605,N_1616);
or U1684 (N_1684,N_1637,N_1602);
xnor U1685 (N_1685,N_1606,N_1635);
or U1686 (N_1686,N_1646,N_1644);
or U1687 (N_1687,N_1626,N_1635);
or U1688 (N_1688,N_1640,N_1642);
xor U1689 (N_1689,N_1617,N_1649);
nor U1690 (N_1690,N_1633,N_1620);
or U1691 (N_1691,N_1606,N_1619);
xor U1692 (N_1692,N_1604,N_1625);
nand U1693 (N_1693,N_1616,N_1636);
nor U1694 (N_1694,N_1630,N_1602);
nand U1695 (N_1695,N_1643,N_1629);
and U1696 (N_1696,N_1607,N_1604);
nor U1697 (N_1697,N_1618,N_1601);
nand U1698 (N_1698,N_1603,N_1627);
nand U1699 (N_1699,N_1638,N_1602);
xor U1700 (N_1700,N_1656,N_1673);
and U1701 (N_1701,N_1668,N_1698);
nand U1702 (N_1702,N_1663,N_1684);
and U1703 (N_1703,N_1677,N_1694);
and U1704 (N_1704,N_1667,N_1699);
nor U1705 (N_1705,N_1666,N_1652);
and U1706 (N_1706,N_1665,N_1669);
xnor U1707 (N_1707,N_1670,N_1664);
nand U1708 (N_1708,N_1686,N_1676);
xor U1709 (N_1709,N_1688,N_1679);
nand U1710 (N_1710,N_1662,N_1654);
and U1711 (N_1711,N_1680,N_1657);
and U1712 (N_1712,N_1689,N_1650);
nand U1713 (N_1713,N_1687,N_1674);
nor U1714 (N_1714,N_1682,N_1678);
nand U1715 (N_1715,N_1683,N_1691);
and U1716 (N_1716,N_1660,N_1697);
or U1717 (N_1717,N_1693,N_1653);
nor U1718 (N_1718,N_1672,N_1655);
or U1719 (N_1719,N_1692,N_1659);
xor U1720 (N_1720,N_1696,N_1695);
xor U1721 (N_1721,N_1671,N_1681);
nand U1722 (N_1722,N_1690,N_1661);
xor U1723 (N_1723,N_1658,N_1685);
and U1724 (N_1724,N_1675,N_1651);
nand U1725 (N_1725,N_1677,N_1697);
or U1726 (N_1726,N_1670,N_1698);
and U1727 (N_1727,N_1692,N_1695);
and U1728 (N_1728,N_1678,N_1680);
nand U1729 (N_1729,N_1674,N_1650);
nand U1730 (N_1730,N_1655,N_1674);
nor U1731 (N_1731,N_1670,N_1676);
or U1732 (N_1732,N_1675,N_1662);
nand U1733 (N_1733,N_1672,N_1667);
and U1734 (N_1734,N_1688,N_1654);
and U1735 (N_1735,N_1689,N_1664);
xor U1736 (N_1736,N_1668,N_1685);
xor U1737 (N_1737,N_1661,N_1695);
xor U1738 (N_1738,N_1658,N_1692);
nand U1739 (N_1739,N_1662,N_1697);
or U1740 (N_1740,N_1650,N_1667);
or U1741 (N_1741,N_1684,N_1676);
nor U1742 (N_1742,N_1652,N_1679);
nor U1743 (N_1743,N_1655,N_1673);
nand U1744 (N_1744,N_1689,N_1672);
xnor U1745 (N_1745,N_1650,N_1695);
and U1746 (N_1746,N_1674,N_1675);
and U1747 (N_1747,N_1658,N_1688);
nand U1748 (N_1748,N_1679,N_1666);
nor U1749 (N_1749,N_1694,N_1654);
xnor U1750 (N_1750,N_1708,N_1728);
nand U1751 (N_1751,N_1735,N_1725);
nor U1752 (N_1752,N_1746,N_1737);
nor U1753 (N_1753,N_1740,N_1702);
and U1754 (N_1754,N_1700,N_1720);
nand U1755 (N_1755,N_1729,N_1748);
and U1756 (N_1756,N_1741,N_1713);
xnor U1757 (N_1757,N_1704,N_1747);
nand U1758 (N_1758,N_1743,N_1721);
nand U1759 (N_1759,N_1705,N_1712);
nand U1760 (N_1760,N_1707,N_1749);
xor U1761 (N_1761,N_1717,N_1716);
nor U1762 (N_1762,N_1719,N_1711);
or U1763 (N_1763,N_1727,N_1738);
or U1764 (N_1764,N_1742,N_1714);
and U1765 (N_1765,N_1745,N_1736);
xnor U1766 (N_1766,N_1744,N_1706);
or U1767 (N_1767,N_1703,N_1732);
and U1768 (N_1768,N_1718,N_1731);
nor U1769 (N_1769,N_1733,N_1730);
and U1770 (N_1770,N_1723,N_1709);
nor U1771 (N_1771,N_1739,N_1710);
xnor U1772 (N_1772,N_1701,N_1734);
xnor U1773 (N_1773,N_1726,N_1724);
and U1774 (N_1774,N_1722,N_1715);
or U1775 (N_1775,N_1709,N_1712);
and U1776 (N_1776,N_1741,N_1735);
xnor U1777 (N_1777,N_1701,N_1716);
xor U1778 (N_1778,N_1732,N_1749);
and U1779 (N_1779,N_1708,N_1746);
nor U1780 (N_1780,N_1729,N_1725);
nand U1781 (N_1781,N_1748,N_1713);
nor U1782 (N_1782,N_1709,N_1703);
nand U1783 (N_1783,N_1734,N_1736);
nand U1784 (N_1784,N_1743,N_1742);
nand U1785 (N_1785,N_1728,N_1749);
nand U1786 (N_1786,N_1717,N_1707);
or U1787 (N_1787,N_1734,N_1702);
or U1788 (N_1788,N_1731,N_1726);
or U1789 (N_1789,N_1702,N_1721);
and U1790 (N_1790,N_1737,N_1719);
xor U1791 (N_1791,N_1732,N_1709);
xor U1792 (N_1792,N_1714,N_1747);
xor U1793 (N_1793,N_1719,N_1745);
nand U1794 (N_1794,N_1741,N_1731);
xnor U1795 (N_1795,N_1742,N_1745);
xor U1796 (N_1796,N_1723,N_1728);
or U1797 (N_1797,N_1736,N_1737);
xnor U1798 (N_1798,N_1717,N_1703);
nand U1799 (N_1799,N_1742,N_1725);
and U1800 (N_1800,N_1798,N_1759);
nand U1801 (N_1801,N_1770,N_1793);
xnor U1802 (N_1802,N_1750,N_1767);
xor U1803 (N_1803,N_1751,N_1781);
nor U1804 (N_1804,N_1765,N_1790);
xnor U1805 (N_1805,N_1796,N_1771);
and U1806 (N_1806,N_1774,N_1787);
and U1807 (N_1807,N_1789,N_1777);
nor U1808 (N_1808,N_1757,N_1786);
xor U1809 (N_1809,N_1756,N_1760);
nand U1810 (N_1810,N_1794,N_1755);
xor U1811 (N_1811,N_1773,N_1758);
and U1812 (N_1812,N_1754,N_1785);
or U1813 (N_1813,N_1753,N_1766);
nor U1814 (N_1814,N_1799,N_1764);
and U1815 (N_1815,N_1769,N_1776);
xnor U1816 (N_1816,N_1768,N_1788);
nor U1817 (N_1817,N_1797,N_1782);
nand U1818 (N_1818,N_1775,N_1762);
xor U1819 (N_1819,N_1791,N_1779);
or U1820 (N_1820,N_1792,N_1772);
nand U1821 (N_1821,N_1784,N_1780);
or U1822 (N_1822,N_1783,N_1778);
or U1823 (N_1823,N_1752,N_1795);
nand U1824 (N_1824,N_1763,N_1761);
xor U1825 (N_1825,N_1751,N_1755);
nand U1826 (N_1826,N_1768,N_1787);
nor U1827 (N_1827,N_1798,N_1758);
and U1828 (N_1828,N_1781,N_1772);
nor U1829 (N_1829,N_1798,N_1750);
nor U1830 (N_1830,N_1768,N_1790);
nand U1831 (N_1831,N_1775,N_1760);
nor U1832 (N_1832,N_1794,N_1774);
or U1833 (N_1833,N_1767,N_1766);
xnor U1834 (N_1834,N_1763,N_1777);
xor U1835 (N_1835,N_1794,N_1785);
and U1836 (N_1836,N_1762,N_1758);
or U1837 (N_1837,N_1770,N_1779);
or U1838 (N_1838,N_1789,N_1757);
nand U1839 (N_1839,N_1759,N_1765);
and U1840 (N_1840,N_1789,N_1778);
and U1841 (N_1841,N_1769,N_1784);
or U1842 (N_1842,N_1780,N_1788);
and U1843 (N_1843,N_1792,N_1757);
or U1844 (N_1844,N_1785,N_1789);
or U1845 (N_1845,N_1780,N_1750);
or U1846 (N_1846,N_1771,N_1792);
nand U1847 (N_1847,N_1789,N_1772);
or U1848 (N_1848,N_1781,N_1793);
xor U1849 (N_1849,N_1755,N_1778);
and U1850 (N_1850,N_1806,N_1804);
or U1851 (N_1851,N_1824,N_1830);
nand U1852 (N_1852,N_1808,N_1839);
or U1853 (N_1853,N_1812,N_1843);
xor U1854 (N_1854,N_1840,N_1834);
or U1855 (N_1855,N_1813,N_1842);
nor U1856 (N_1856,N_1846,N_1833);
xor U1857 (N_1857,N_1809,N_1811);
or U1858 (N_1858,N_1823,N_1828);
and U1859 (N_1859,N_1837,N_1803);
nor U1860 (N_1860,N_1819,N_1820);
nor U1861 (N_1861,N_1827,N_1838);
xor U1862 (N_1862,N_1822,N_1831);
nor U1863 (N_1863,N_1845,N_1818);
nand U1864 (N_1864,N_1814,N_1805);
or U1865 (N_1865,N_1817,N_1844);
xor U1866 (N_1866,N_1826,N_1815);
xor U1867 (N_1867,N_1816,N_1836);
nor U1868 (N_1868,N_1800,N_1848);
xor U1869 (N_1869,N_1849,N_1825);
or U1870 (N_1870,N_1801,N_1829);
xnor U1871 (N_1871,N_1835,N_1821);
xor U1872 (N_1872,N_1832,N_1841);
xor U1873 (N_1873,N_1802,N_1810);
xor U1874 (N_1874,N_1847,N_1807);
nor U1875 (N_1875,N_1823,N_1804);
xor U1876 (N_1876,N_1839,N_1807);
nor U1877 (N_1877,N_1848,N_1804);
nor U1878 (N_1878,N_1814,N_1844);
or U1879 (N_1879,N_1829,N_1819);
and U1880 (N_1880,N_1815,N_1831);
xnor U1881 (N_1881,N_1838,N_1813);
and U1882 (N_1882,N_1811,N_1843);
xnor U1883 (N_1883,N_1812,N_1801);
or U1884 (N_1884,N_1801,N_1807);
nand U1885 (N_1885,N_1838,N_1815);
and U1886 (N_1886,N_1839,N_1826);
nor U1887 (N_1887,N_1816,N_1830);
nor U1888 (N_1888,N_1805,N_1820);
or U1889 (N_1889,N_1847,N_1821);
nand U1890 (N_1890,N_1837,N_1820);
xnor U1891 (N_1891,N_1833,N_1815);
or U1892 (N_1892,N_1847,N_1811);
nand U1893 (N_1893,N_1840,N_1818);
and U1894 (N_1894,N_1835,N_1843);
and U1895 (N_1895,N_1800,N_1807);
nor U1896 (N_1896,N_1808,N_1809);
and U1897 (N_1897,N_1815,N_1806);
or U1898 (N_1898,N_1819,N_1827);
xor U1899 (N_1899,N_1820,N_1804);
and U1900 (N_1900,N_1869,N_1856);
or U1901 (N_1901,N_1899,N_1873);
and U1902 (N_1902,N_1876,N_1877);
nor U1903 (N_1903,N_1853,N_1882);
xnor U1904 (N_1904,N_1888,N_1870);
or U1905 (N_1905,N_1896,N_1887);
nand U1906 (N_1906,N_1892,N_1855);
or U1907 (N_1907,N_1861,N_1857);
or U1908 (N_1908,N_1864,N_1891);
nand U1909 (N_1909,N_1859,N_1889);
or U1910 (N_1910,N_1854,N_1868);
and U1911 (N_1911,N_1884,N_1894);
xnor U1912 (N_1912,N_1874,N_1872);
nor U1913 (N_1913,N_1881,N_1878);
xnor U1914 (N_1914,N_1850,N_1886);
or U1915 (N_1915,N_1860,N_1866);
nand U1916 (N_1916,N_1867,N_1865);
nor U1917 (N_1917,N_1883,N_1871);
or U1918 (N_1918,N_1890,N_1875);
xor U1919 (N_1919,N_1897,N_1879);
and U1920 (N_1920,N_1885,N_1851);
and U1921 (N_1921,N_1898,N_1862);
and U1922 (N_1922,N_1895,N_1893);
nand U1923 (N_1923,N_1852,N_1880);
nor U1924 (N_1924,N_1863,N_1858);
xnor U1925 (N_1925,N_1886,N_1887);
nand U1926 (N_1926,N_1884,N_1855);
and U1927 (N_1927,N_1890,N_1889);
or U1928 (N_1928,N_1860,N_1850);
xor U1929 (N_1929,N_1897,N_1859);
or U1930 (N_1930,N_1850,N_1869);
and U1931 (N_1931,N_1874,N_1861);
or U1932 (N_1932,N_1888,N_1889);
nor U1933 (N_1933,N_1869,N_1885);
or U1934 (N_1934,N_1871,N_1881);
or U1935 (N_1935,N_1870,N_1853);
nor U1936 (N_1936,N_1869,N_1859);
xnor U1937 (N_1937,N_1857,N_1881);
nor U1938 (N_1938,N_1877,N_1867);
and U1939 (N_1939,N_1863,N_1874);
nand U1940 (N_1940,N_1870,N_1862);
nand U1941 (N_1941,N_1874,N_1853);
xnor U1942 (N_1942,N_1873,N_1863);
and U1943 (N_1943,N_1866,N_1875);
xnor U1944 (N_1944,N_1851,N_1892);
nor U1945 (N_1945,N_1886,N_1874);
nor U1946 (N_1946,N_1856,N_1863);
or U1947 (N_1947,N_1868,N_1867);
and U1948 (N_1948,N_1887,N_1889);
and U1949 (N_1949,N_1867,N_1888);
xor U1950 (N_1950,N_1907,N_1920);
xnor U1951 (N_1951,N_1913,N_1924);
and U1952 (N_1952,N_1940,N_1906);
or U1953 (N_1953,N_1902,N_1930);
nand U1954 (N_1954,N_1908,N_1926);
or U1955 (N_1955,N_1919,N_1916);
and U1956 (N_1956,N_1914,N_1933);
nand U1957 (N_1957,N_1939,N_1918);
or U1958 (N_1958,N_1943,N_1903);
or U1959 (N_1959,N_1905,N_1912);
and U1960 (N_1960,N_1921,N_1931);
nor U1961 (N_1961,N_1937,N_1934);
or U1962 (N_1962,N_1947,N_1948);
and U1963 (N_1963,N_1946,N_1917);
and U1964 (N_1964,N_1925,N_1932);
nor U1965 (N_1965,N_1942,N_1929);
and U1966 (N_1966,N_1938,N_1936);
xor U1967 (N_1967,N_1945,N_1909);
and U1968 (N_1968,N_1927,N_1900);
nand U1969 (N_1969,N_1901,N_1922);
xor U1970 (N_1970,N_1910,N_1928);
nand U1971 (N_1971,N_1904,N_1923);
nand U1972 (N_1972,N_1941,N_1915);
nor U1973 (N_1973,N_1935,N_1911);
xnor U1974 (N_1974,N_1949,N_1944);
nand U1975 (N_1975,N_1939,N_1919);
nand U1976 (N_1976,N_1938,N_1921);
nor U1977 (N_1977,N_1936,N_1914);
nand U1978 (N_1978,N_1921,N_1930);
nor U1979 (N_1979,N_1934,N_1922);
or U1980 (N_1980,N_1921,N_1936);
xnor U1981 (N_1981,N_1944,N_1919);
xnor U1982 (N_1982,N_1920,N_1932);
or U1983 (N_1983,N_1905,N_1940);
and U1984 (N_1984,N_1924,N_1935);
nor U1985 (N_1985,N_1908,N_1941);
nor U1986 (N_1986,N_1910,N_1935);
or U1987 (N_1987,N_1939,N_1937);
nor U1988 (N_1988,N_1931,N_1946);
or U1989 (N_1989,N_1939,N_1942);
or U1990 (N_1990,N_1913,N_1915);
nand U1991 (N_1991,N_1911,N_1929);
nor U1992 (N_1992,N_1908,N_1945);
or U1993 (N_1993,N_1940,N_1949);
and U1994 (N_1994,N_1904,N_1933);
xnor U1995 (N_1995,N_1930,N_1919);
nand U1996 (N_1996,N_1936,N_1904);
nand U1997 (N_1997,N_1920,N_1930);
nor U1998 (N_1998,N_1902,N_1949);
xor U1999 (N_1999,N_1945,N_1932);
xnor U2000 (N_2000,N_1979,N_1955);
nor U2001 (N_2001,N_1968,N_1965);
xor U2002 (N_2002,N_1954,N_1959);
xnor U2003 (N_2003,N_1952,N_1978);
and U2004 (N_2004,N_1969,N_1985);
nand U2005 (N_2005,N_1977,N_1964);
or U2006 (N_2006,N_1972,N_1951);
and U2007 (N_2007,N_1988,N_1989);
xnor U2008 (N_2008,N_1990,N_1962);
or U2009 (N_2009,N_1986,N_1974);
nor U2010 (N_2010,N_1963,N_1994);
nor U2011 (N_2011,N_1982,N_1970);
nor U2012 (N_2012,N_1980,N_1987);
nor U2013 (N_2013,N_1976,N_1960);
nor U2014 (N_2014,N_1981,N_1975);
or U2015 (N_2015,N_1957,N_1995);
xor U2016 (N_2016,N_1998,N_1967);
nor U2017 (N_2017,N_1971,N_1953);
nor U2018 (N_2018,N_1996,N_1961);
nor U2019 (N_2019,N_1966,N_1956);
nor U2020 (N_2020,N_1958,N_1991);
and U2021 (N_2021,N_1950,N_1993);
xor U2022 (N_2022,N_1997,N_1983);
or U2023 (N_2023,N_1999,N_1984);
nand U2024 (N_2024,N_1992,N_1973);
xor U2025 (N_2025,N_1993,N_1984);
nand U2026 (N_2026,N_1995,N_1967);
or U2027 (N_2027,N_1997,N_1952);
xnor U2028 (N_2028,N_1992,N_1981);
nand U2029 (N_2029,N_1977,N_1984);
nor U2030 (N_2030,N_1967,N_1989);
xor U2031 (N_2031,N_1953,N_1982);
nand U2032 (N_2032,N_1963,N_1961);
and U2033 (N_2033,N_1999,N_1968);
nand U2034 (N_2034,N_1978,N_1970);
nor U2035 (N_2035,N_1959,N_1964);
xnor U2036 (N_2036,N_1980,N_1976);
xnor U2037 (N_2037,N_1972,N_1956);
nand U2038 (N_2038,N_1984,N_1991);
nand U2039 (N_2039,N_1958,N_1984);
nand U2040 (N_2040,N_1989,N_1998);
nor U2041 (N_2041,N_1972,N_1996);
nor U2042 (N_2042,N_1995,N_1993);
nor U2043 (N_2043,N_1991,N_1974);
nor U2044 (N_2044,N_1963,N_1971);
and U2045 (N_2045,N_1963,N_1995);
and U2046 (N_2046,N_1950,N_1997);
or U2047 (N_2047,N_1998,N_1969);
nand U2048 (N_2048,N_1952,N_1981);
or U2049 (N_2049,N_1961,N_1992);
nor U2050 (N_2050,N_2038,N_2027);
nor U2051 (N_2051,N_2028,N_2034);
nor U2052 (N_2052,N_2020,N_2019);
and U2053 (N_2053,N_2049,N_2018);
nand U2054 (N_2054,N_2024,N_2001);
nor U2055 (N_2055,N_2013,N_2007);
xor U2056 (N_2056,N_2039,N_2022);
or U2057 (N_2057,N_2031,N_2033);
nor U2058 (N_2058,N_2045,N_2014);
nor U2059 (N_2059,N_2015,N_2040);
xor U2060 (N_2060,N_2012,N_2037);
xor U2061 (N_2061,N_2004,N_2016);
or U2062 (N_2062,N_2000,N_2047);
nand U2063 (N_2063,N_2009,N_2029);
and U2064 (N_2064,N_2006,N_2002);
nor U2065 (N_2065,N_2008,N_2042);
or U2066 (N_2066,N_2005,N_2030);
or U2067 (N_2067,N_2041,N_2044);
or U2068 (N_2068,N_2011,N_2026);
xnor U2069 (N_2069,N_2032,N_2048);
or U2070 (N_2070,N_2025,N_2036);
and U2071 (N_2071,N_2043,N_2035);
nor U2072 (N_2072,N_2017,N_2021);
or U2073 (N_2073,N_2003,N_2046);
and U2074 (N_2074,N_2023,N_2010);
xor U2075 (N_2075,N_2033,N_2010);
or U2076 (N_2076,N_2039,N_2005);
and U2077 (N_2077,N_2043,N_2019);
and U2078 (N_2078,N_2025,N_2027);
xor U2079 (N_2079,N_2009,N_2019);
or U2080 (N_2080,N_2006,N_2012);
xor U2081 (N_2081,N_2030,N_2019);
nor U2082 (N_2082,N_2010,N_2047);
and U2083 (N_2083,N_2028,N_2027);
xnor U2084 (N_2084,N_2020,N_2033);
or U2085 (N_2085,N_2041,N_2011);
or U2086 (N_2086,N_2005,N_2024);
nor U2087 (N_2087,N_2028,N_2005);
or U2088 (N_2088,N_2036,N_2000);
nand U2089 (N_2089,N_2026,N_2023);
or U2090 (N_2090,N_2015,N_2025);
xor U2091 (N_2091,N_2020,N_2023);
nor U2092 (N_2092,N_2033,N_2026);
nand U2093 (N_2093,N_2018,N_2025);
xnor U2094 (N_2094,N_2020,N_2034);
xnor U2095 (N_2095,N_2034,N_2027);
and U2096 (N_2096,N_2046,N_2034);
nor U2097 (N_2097,N_2046,N_2009);
and U2098 (N_2098,N_2044,N_2024);
xnor U2099 (N_2099,N_2040,N_2048);
xnor U2100 (N_2100,N_2056,N_2057);
or U2101 (N_2101,N_2075,N_2088);
and U2102 (N_2102,N_2053,N_2062);
nand U2103 (N_2103,N_2082,N_2058);
or U2104 (N_2104,N_2095,N_2078);
nand U2105 (N_2105,N_2090,N_2083);
or U2106 (N_2106,N_2055,N_2084);
nand U2107 (N_2107,N_2070,N_2085);
nand U2108 (N_2108,N_2073,N_2081);
or U2109 (N_2109,N_2064,N_2077);
and U2110 (N_2110,N_2097,N_2091);
and U2111 (N_2111,N_2050,N_2076);
xnor U2112 (N_2112,N_2066,N_2074);
or U2113 (N_2113,N_2093,N_2052);
and U2114 (N_2114,N_2072,N_2051);
and U2115 (N_2115,N_2079,N_2094);
nor U2116 (N_2116,N_2061,N_2067);
nor U2117 (N_2117,N_2098,N_2080);
or U2118 (N_2118,N_2071,N_2089);
and U2119 (N_2119,N_2069,N_2087);
or U2120 (N_2120,N_2054,N_2060);
nand U2121 (N_2121,N_2096,N_2092);
or U2122 (N_2122,N_2086,N_2065);
or U2123 (N_2123,N_2099,N_2068);
or U2124 (N_2124,N_2059,N_2063);
or U2125 (N_2125,N_2052,N_2088);
nand U2126 (N_2126,N_2094,N_2053);
and U2127 (N_2127,N_2092,N_2097);
nor U2128 (N_2128,N_2078,N_2090);
or U2129 (N_2129,N_2055,N_2060);
nor U2130 (N_2130,N_2066,N_2059);
nand U2131 (N_2131,N_2089,N_2085);
nand U2132 (N_2132,N_2065,N_2062);
or U2133 (N_2133,N_2080,N_2069);
nor U2134 (N_2134,N_2082,N_2097);
and U2135 (N_2135,N_2068,N_2058);
and U2136 (N_2136,N_2084,N_2066);
or U2137 (N_2137,N_2093,N_2081);
nor U2138 (N_2138,N_2071,N_2096);
nor U2139 (N_2139,N_2075,N_2054);
nand U2140 (N_2140,N_2076,N_2098);
xor U2141 (N_2141,N_2069,N_2093);
or U2142 (N_2142,N_2094,N_2057);
nor U2143 (N_2143,N_2054,N_2092);
and U2144 (N_2144,N_2050,N_2090);
nor U2145 (N_2145,N_2077,N_2063);
and U2146 (N_2146,N_2082,N_2098);
or U2147 (N_2147,N_2059,N_2071);
nor U2148 (N_2148,N_2081,N_2066);
nand U2149 (N_2149,N_2081,N_2085);
nand U2150 (N_2150,N_2135,N_2148);
nor U2151 (N_2151,N_2126,N_2102);
nand U2152 (N_2152,N_2103,N_2122);
xor U2153 (N_2153,N_2133,N_2108);
and U2154 (N_2154,N_2119,N_2101);
nand U2155 (N_2155,N_2128,N_2124);
nand U2156 (N_2156,N_2120,N_2121);
nor U2157 (N_2157,N_2104,N_2114);
xor U2158 (N_2158,N_2107,N_2139);
nor U2159 (N_2159,N_2109,N_2146);
and U2160 (N_2160,N_2138,N_2137);
nand U2161 (N_2161,N_2127,N_2130);
and U2162 (N_2162,N_2147,N_2132);
xor U2163 (N_2163,N_2134,N_2129);
and U2164 (N_2164,N_2141,N_2145);
nand U2165 (N_2165,N_2110,N_2123);
nor U2166 (N_2166,N_2144,N_2125);
and U2167 (N_2167,N_2117,N_2140);
xnor U2168 (N_2168,N_2105,N_2100);
or U2169 (N_2169,N_2116,N_2149);
or U2170 (N_2170,N_2106,N_2113);
xor U2171 (N_2171,N_2112,N_2111);
xnor U2172 (N_2172,N_2136,N_2142);
nor U2173 (N_2173,N_2115,N_2118);
nor U2174 (N_2174,N_2143,N_2131);
nand U2175 (N_2175,N_2122,N_2131);
xor U2176 (N_2176,N_2148,N_2113);
nor U2177 (N_2177,N_2118,N_2139);
nand U2178 (N_2178,N_2128,N_2145);
nor U2179 (N_2179,N_2108,N_2127);
or U2180 (N_2180,N_2120,N_2106);
nand U2181 (N_2181,N_2109,N_2127);
nor U2182 (N_2182,N_2119,N_2125);
xnor U2183 (N_2183,N_2129,N_2145);
nand U2184 (N_2184,N_2122,N_2136);
nand U2185 (N_2185,N_2113,N_2126);
nand U2186 (N_2186,N_2114,N_2141);
or U2187 (N_2187,N_2121,N_2118);
xor U2188 (N_2188,N_2149,N_2140);
nor U2189 (N_2189,N_2149,N_2101);
or U2190 (N_2190,N_2100,N_2138);
nand U2191 (N_2191,N_2103,N_2120);
nor U2192 (N_2192,N_2100,N_2123);
nand U2193 (N_2193,N_2125,N_2137);
and U2194 (N_2194,N_2147,N_2130);
nand U2195 (N_2195,N_2118,N_2127);
and U2196 (N_2196,N_2102,N_2107);
and U2197 (N_2197,N_2112,N_2145);
and U2198 (N_2198,N_2120,N_2118);
or U2199 (N_2199,N_2135,N_2106);
and U2200 (N_2200,N_2193,N_2155);
xor U2201 (N_2201,N_2154,N_2153);
nor U2202 (N_2202,N_2172,N_2169);
or U2203 (N_2203,N_2176,N_2159);
nand U2204 (N_2204,N_2196,N_2164);
and U2205 (N_2205,N_2174,N_2192);
and U2206 (N_2206,N_2173,N_2167);
nand U2207 (N_2207,N_2186,N_2165);
or U2208 (N_2208,N_2199,N_2187);
and U2209 (N_2209,N_2166,N_2150);
nand U2210 (N_2210,N_2160,N_2195);
nor U2211 (N_2211,N_2191,N_2182);
and U2212 (N_2212,N_2188,N_2190);
xor U2213 (N_2213,N_2175,N_2156);
xor U2214 (N_2214,N_2177,N_2158);
xnor U2215 (N_2215,N_2185,N_2181);
and U2216 (N_2216,N_2157,N_2197);
nor U2217 (N_2217,N_2194,N_2198);
nand U2218 (N_2218,N_2178,N_2151);
or U2219 (N_2219,N_2184,N_2179);
xnor U2220 (N_2220,N_2163,N_2168);
or U2221 (N_2221,N_2161,N_2152);
or U2222 (N_2222,N_2189,N_2171);
xor U2223 (N_2223,N_2180,N_2162);
and U2224 (N_2224,N_2170,N_2183);
xor U2225 (N_2225,N_2173,N_2175);
nand U2226 (N_2226,N_2197,N_2154);
or U2227 (N_2227,N_2178,N_2162);
nand U2228 (N_2228,N_2192,N_2187);
or U2229 (N_2229,N_2185,N_2173);
or U2230 (N_2230,N_2178,N_2171);
and U2231 (N_2231,N_2166,N_2199);
and U2232 (N_2232,N_2152,N_2197);
nor U2233 (N_2233,N_2164,N_2179);
nor U2234 (N_2234,N_2182,N_2195);
xnor U2235 (N_2235,N_2194,N_2189);
nor U2236 (N_2236,N_2194,N_2170);
or U2237 (N_2237,N_2191,N_2197);
xor U2238 (N_2238,N_2152,N_2187);
xnor U2239 (N_2239,N_2157,N_2158);
xnor U2240 (N_2240,N_2191,N_2150);
or U2241 (N_2241,N_2185,N_2178);
nand U2242 (N_2242,N_2164,N_2155);
or U2243 (N_2243,N_2197,N_2193);
nor U2244 (N_2244,N_2175,N_2158);
nor U2245 (N_2245,N_2159,N_2157);
nor U2246 (N_2246,N_2154,N_2196);
nor U2247 (N_2247,N_2190,N_2151);
and U2248 (N_2248,N_2190,N_2186);
nor U2249 (N_2249,N_2164,N_2174);
and U2250 (N_2250,N_2208,N_2230);
and U2251 (N_2251,N_2221,N_2210);
nor U2252 (N_2252,N_2223,N_2243);
nor U2253 (N_2253,N_2215,N_2241);
or U2254 (N_2254,N_2237,N_2225);
and U2255 (N_2255,N_2202,N_2200);
xnor U2256 (N_2256,N_2235,N_2212);
and U2257 (N_2257,N_2232,N_2224);
nand U2258 (N_2258,N_2206,N_2244);
nand U2259 (N_2259,N_2211,N_2236);
and U2260 (N_2260,N_2227,N_2222);
nor U2261 (N_2261,N_2228,N_2203);
nor U2262 (N_2262,N_2242,N_2245);
xor U2263 (N_2263,N_2233,N_2231);
nor U2264 (N_2264,N_2234,N_2229);
and U2265 (N_2265,N_2218,N_2240);
nor U2266 (N_2266,N_2214,N_2217);
and U2267 (N_2267,N_2226,N_2201);
nand U2268 (N_2268,N_2247,N_2205);
nand U2269 (N_2269,N_2238,N_2216);
or U2270 (N_2270,N_2248,N_2249);
nor U2271 (N_2271,N_2207,N_2220);
and U2272 (N_2272,N_2219,N_2239);
nand U2273 (N_2273,N_2213,N_2204);
nand U2274 (N_2274,N_2209,N_2246);
nor U2275 (N_2275,N_2224,N_2218);
or U2276 (N_2276,N_2249,N_2202);
or U2277 (N_2277,N_2215,N_2212);
or U2278 (N_2278,N_2226,N_2204);
xnor U2279 (N_2279,N_2231,N_2249);
nand U2280 (N_2280,N_2206,N_2222);
and U2281 (N_2281,N_2240,N_2205);
nor U2282 (N_2282,N_2238,N_2242);
nor U2283 (N_2283,N_2238,N_2217);
or U2284 (N_2284,N_2224,N_2227);
or U2285 (N_2285,N_2243,N_2246);
and U2286 (N_2286,N_2200,N_2238);
or U2287 (N_2287,N_2211,N_2203);
nand U2288 (N_2288,N_2234,N_2218);
nor U2289 (N_2289,N_2212,N_2236);
and U2290 (N_2290,N_2224,N_2222);
nand U2291 (N_2291,N_2230,N_2232);
nor U2292 (N_2292,N_2215,N_2218);
xnor U2293 (N_2293,N_2240,N_2246);
nor U2294 (N_2294,N_2225,N_2235);
and U2295 (N_2295,N_2214,N_2247);
nand U2296 (N_2296,N_2223,N_2225);
or U2297 (N_2297,N_2225,N_2243);
or U2298 (N_2298,N_2213,N_2245);
and U2299 (N_2299,N_2208,N_2233);
and U2300 (N_2300,N_2260,N_2297);
nor U2301 (N_2301,N_2291,N_2298);
or U2302 (N_2302,N_2255,N_2266);
or U2303 (N_2303,N_2268,N_2271);
nand U2304 (N_2304,N_2261,N_2286);
nor U2305 (N_2305,N_2272,N_2253);
or U2306 (N_2306,N_2277,N_2264);
nor U2307 (N_2307,N_2282,N_2284);
and U2308 (N_2308,N_2273,N_2270);
nor U2309 (N_2309,N_2258,N_2252);
nand U2310 (N_2310,N_2254,N_2278);
nor U2311 (N_2311,N_2285,N_2294);
or U2312 (N_2312,N_2257,N_2299);
and U2313 (N_2313,N_2288,N_2262);
nand U2314 (N_2314,N_2274,N_2293);
and U2315 (N_2315,N_2259,N_2265);
or U2316 (N_2316,N_2251,N_2256);
xor U2317 (N_2317,N_2267,N_2279);
nand U2318 (N_2318,N_2275,N_2287);
and U2319 (N_2319,N_2280,N_2263);
nor U2320 (N_2320,N_2283,N_2290);
nand U2321 (N_2321,N_2250,N_2296);
nand U2322 (N_2322,N_2289,N_2295);
xnor U2323 (N_2323,N_2269,N_2276);
nor U2324 (N_2324,N_2281,N_2292);
nand U2325 (N_2325,N_2293,N_2285);
and U2326 (N_2326,N_2289,N_2270);
or U2327 (N_2327,N_2286,N_2291);
and U2328 (N_2328,N_2273,N_2290);
or U2329 (N_2329,N_2271,N_2262);
nand U2330 (N_2330,N_2270,N_2274);
nor U2331 (N_2331,N_2281,N_2287);
and U2332 (N_2332,N_2295,N_2274);
or U2333 (N_2333,N_2274,N_2275);
or U2334 (N_2334,N_2281,N_2299);
and U2335 (N_2335,N_2296,N_2254);
or U2336 (N_2336,N_2295,N_2256);
or U2337 (N_2337,N_2290,N_2252);
and U2338 (N_2338,N_2285,N_2262);
nand U2339 (N_2339,N_2287,N_2268);
xnor U2340 (N_2340,N_2271,N_2256);
and U2341 (N_2341,N_2281,N_2275);
nor U2342 (N_2342,N_2275,N_2261);
and U2343 (N_2343,N_2284,N_2255);
nand U2344 (N_2344,N_2284,N_2265);
nor U2345 (N_2345,N_2289,N_2278);
nand U2346 (N_2346,N_2295,N_2250);
nor U2347 (N_2347,N_2287,N_2291);
and U2348 (N_2348,N_2292,N_2276);
and U2349 (N_2349,N_2260,N_2288);
nand U2350 (N_2350,N_2314,N_2316);
nand U2351 (N_2351,N_2304,N_2338);
nor U2352 (N_2352,N_2300,N_2306);
nand U2353 (N_2353,N_2332,N_2323);
xnor U2354 (N_2354,N_2309,N_2325);
xor U2355 (N_2355,N_2326,N_2318);
nor U2356 (N_2356,N_2343,N_2337);
nand U2357 (N_2357,N_2319,N_2349);
nor U2358 (N_2358,N_2315,N_2305);
nor U2359 (N_2359,N_2339,N_2340);
and U2360 (N_2360,N_2335,N_2322);
xor U2361 (N_2361,N_2330,N_2331);
or U2362 (N_2362,N_2336,N_2311);
xor U2363 (N_2363,N_2303,N_2345);
xnor U2364 (N_2364,N_2348,N_2333);
nor U2365 (N_2365,N_2327,N_2346);
nor U2366 (N_2366,N_2341,N_2301);
nand U2367 (N_2367,N_2320,N_2302);
xor U2368 (N_2368,N_2334,N_2328);
xnor U2369 (N_2369,N_2307,N_2310);
nand U2370 (N_2370,N_2321,N_2308);
or U2371 (N_2371,N_2342,N_2324);
xnor U2372 (N_2372,N_2317,N_2329);
nand U2373 (N_2373,N_2347,N_2312);
xnor U2374 (N_2374,N_2344,N_2313);
and U2375 (N_2375,N_2306,N_2322);
or U2376 (N_2376,N_2314,N_2313);
nand U2377 (N_2377,N_2304,N_2320);
and U2378 (N_2378,N_2342,N_2306);
xnor U2379 (N_2379,N_2305,N_2314);
xnor U2380 (N_2380,N_2340,N_2306);
and U2381 (N_2381,N_2349,N_2347);
nor U2382 (N_2382,N_2307,N_2347);
xnor U2383 (N_2383,N_2328,N_2338);
nor U2384 (N_2384,N_2301,N_2324);
and U2385 (N_2385,N_2307,N_2321);
or U2386 (N_2386,N_2328,N_2341);
xor U2387 (N_2387,N_2324,N_2345);
and U2388 (N_2388,N_2306,N_2326);
and U2389 (N_2389,N_2303,N_2337);
nand U2390 (N_2390,N_2346,N_2315);
and U2391 (N_2391,N_2312,N_2304);
or U2392 (N_2392,N_2307,N_2327);
and U2393 (N_2393,N_2306,N_2343);
xnor U2394 (N_2394,N_2321,N_2316);
or U2395 (N_2395,N_2319,N_2331);
and U2396 (N_2396,N_2325,N_2313);
nand U2397 (N_2397,N_2308,N_2345);
nor U2398 (N_2398,N_2325,N_2349);
and U2399 (N_2399,N_2341,N_2327);
nor U2400 (N_2400,N_2398,N_2374);
nor U2401 (N_2401,N_2371,N_2373);
or U2402 (N_2402,N_2395,N_2356);
and U2403 (N_2403,N_2382,N_2361);
nor U2404 (N_2404,N_2378,N_2377);
and U2405 (N_2405,N_2365,N_2391);
xor U2406 (N_2406,N_2364,N_2397);
nor U2407 (N_2407,N_2376,N_2390);
nand U2408 (N_2408,N_2392,N_2358);
nand U2409 (N_2409,N_2396,N_2366);
nor U2410 (N_2410,N_2363,N_2352);
and U2411 (N_2411,N_2379,N_2394);
nand U2412 (N_2412,N_2369,N_2355);
nor U2413 (N_2413,N_2350,N_2384);
or U2414 (N_2414,N_2399,N_2383);
nor U2415 (N_2415,N_2368,N_2388);
or U2416 (N_2416,N_2385,N_2367);
nand U2417 (N_2417,N_2353,N_2393);
xnor U2418 (N_2418,N_2360,N_2370);
nor U2419 (N_2419,N_2389,N_2375);
or U2420 (N_2420,N_2362,N_2387);
nand U2421 (N_2421,N_2357,N_2380);
nand U2422 (N_2422,N_2386,N_2372);
or U2423 (N_2423,N_2359,N_2381);
nor U2424 (N_2424,N_2351,N_2354);
or U2425 (N_2425,N_2356,N_2367);
and U2426 (N_2426,N_2369,N_2394);
or U2427 (N_2427,N_2364,N_2363);
or U2428 (N_2428,N_2362,N_2357);
and U2429 (N_2429,N_2393,N_2376);
xnor U2430 (N_2430,N_2355,N_2391);
and U2431 (N_2431,N_2360,N_2371);
or U2432 (N_2432,N_2394,N_2393);
xnor U2433 (N_2433,N_2354,N_2396);
xor U2434 (N_2434,N_2382,N_2391);
nand U2435 (N_2435,N_2375,N_2386);
nor U2436 (N_2436,N_2367,N_2387);
xnor U2437 (N_2437,N_2394,N_2381);
or U2438 (N_2438,N_2374,N_2390);
nor U2439 (N_2439,N_2373,N_2356);
nand U2440 (N_2440,N_2372,N_2382);
nor U2441 (N_2441,N_2376,N_2366);
nor U2442 (N_2442,N_2391,N_2396);
and U2443 (N_2443,N_2371,N_2369);
or U2444 (N_2444,N_2370,N_2371);
or U2445 (N_2445,N_2393,N_2364);
nand U2446 (N_2446,N_2375,N_2394);
or U2447 (N_2447,N_2378,N_2383);
nand U2448 (N_2448,N_2398,N_2397);
nand U2449 (N_2449,N_2351,N_2384);
and U2450 (N_2450,N_2440,N_2404);
or U2451 (N_2451,N_2438,N_2408);
nor U2452 (N_2452,N_2422,N_2432);
nor U2453 (N_2453,N_2416,N_2439);
and U2454 (N_2454,N_2401,N_2447);
xor U2455 (N_2455,N_2412,N_2429);
and U2456 (N_2456,N_2413,N_2410);
nand U2457 (N_2457,N_2402,N_2419);
or U2458 (N_2458,N_2443,N_2418);
xor U2459 (N_2459,N_2434,N_2445);
nor U2460 (N_2460,N_2400,N_2421);
nor U2461 (N_2461,N_2430,N_2426);
or U2462 (N_2462,N_2441,N_2409);
xor U2463 (N_2463,N_2425,N_2436);
nand U2464 (N_2464,N_2446,N_2437);
and U2465 (N_2465,N_2411,N_2449);
or U2466 (N_2466,N_2417,N_2405);
nand U2467 (N_2467,N_2435,N_2444);
nor U2468 (N_2468,N_2442,N_2433);
or U2469 (N_2469,N_2424,N_2448);
nor U2470 (N_2470,N_2427,N_2403);
nand U2471 (N_2471,N_2407,N_2428);
and U2472 (N_2472,N_2420,N_2415);
nand U2473 (N_2473,N_2414,N_2423);
and U2474 (N_2474,N_2431,N_2406);
and U2475 (N_2475,N_2422,N_2427);
or U2476 (N_2476,N_2433,N_2445);
xor U2477 (N_2477,N_2401,N_2400);
nor U2478 (N_2478,N_2404,N_2405);
nor U2479 (N_2479,N_2411,N_2417);
nand U2480 (N_2480,N_2401,N_2405);
and U2481 (N_2481,N_2408,N_2427);
xnor U2482 (N_2482,N_2435,N_2421);
nor U2483 (N_2483,N_2443,N_2434);
or U2484 (N_2484,N_2402,N_2413);
nand U2485 (N_2485,N_2440,N_2442);
nand U2486 (N_2486,N_2439,N_2414);
and U2487 (N_2487,N_2447,N_2412);
nor U2488 (N_2488,N_2414,N_2431);
or U2489 (N_2489,N_2447,N_2414);
and U2490 (N_2490,N_2415,N_2405);
and U2491 (N_2491,N_2430,N_2432);
or U2492 (N_2492,N_2449,N_2404);
nand U2493 (N_2493,N_2443,N_2441);
or U2494 (N_2494,N_2427,N_2435);
and U2495 (N_2495,N_2448,N_2443);
xnor U2496 (N_2496,N_2427,N_2420);
xor U2497 (N_2497,N_2414,N_2444);
nor U2498 (N_2498,N_2434,N_2442);
and U2499 (N_2499,N_2410,N_2436);
nor U2500 (N_2500,N_2487,N_2469);
and U2501 (N_2501,N_2453,N_2459);
nand U2502 (N_2502,N_2486,N_2464);
and U2503 (N_2503,N_2498,N_2491);
nor U2504 (N_2504,N_2489,N_2455);
nor U2505 (N_2505,N_2492,N_2493);
nor U2506 (N_2506,N_2497,N_2466);
xor U2507 (N_2507,N_2495,N_2468);
or U2508 (N_2508,N_2470,N_2457);
or U2509 (N_2509,N_2490,N_2471);
nor U2510 (N_2510,N_2477,N_2460);
and U2511 (N_2511,N_2483,N_2475);
and U2512 (N_2512,N_2485,N_2467);
or U2513 (N_2513,N_2499,N_2484);
xor U2514 (N_2514,N_2458,N_2496);
xnor U2515 (N_2515,N_2456,N_2474);
nand U2516 (N_2516,N_2463,N_2482);
and U2517 (N_2517,N_2452,N_2472);
nand U2518 (N_2518,N_2473,N_2494);
nand U2519 (N_2519,N_2488,N_2465);
nor U2520 (N_2520,N_2450,N_2462);
and U2521 (N_2521,N_2454,N_2480);
xnor U2522 (N_2522,N_2478,N_2479);
or U2523 (N_2523,N_2476,N_2451);
and U2524 (N_2524,N_2481,N_2461);
xnor U2525 (N_2525,N_2457,N_2478);
xor U2526 (N_2526,N_2469,N_2498);
or U2527 (N_2527,N_2493,N_2479);
and U2528 (N_2528,N_2487,N_2471);
nor U2529 (N_2529,N_2461,N_2457);
xor U2530 (N_2530,N_2476,N_2489);
or U2531 (N_2531,N_2486,N_2495);
or U2532 (N_2532,N_2452,N_2464);
nor U2533 (N_2533,N_2480,N_2491);
or U2534 (N_2534,N_2492,N_2499);
xor U2535 (N_2535,N_2459,N_2496);
nand U2536 (N_2536,N_2450,N_2484);
nand U2537 (N_2537,N_2476,N_2467);
and U2538 (N_2538,N_2480,N_2494);
or U2539 (N_2539,N_2484,N_2471);
xnor U2540 (N_2540,N_2490,N_2474);
and U2541 (N_2541,N_2486,N_2494);
nor U2542 (N_2542,N_2460,N_2483);
and U2543 (N_2543,N_2466,N_2473);
and U2544 (N_2544,N_2484,N_2474);
or U2545 (N_2545,N_2456,N_2473);
nand U2546 (N_2546,N_2453,N_2492);
and U2547 (N_2547,N_2470,N_2455);
nor U2548 (N_2548,N_2480,N_2482);
xor U2549 (N_2549,N_2461,N_2460);
nor U2550 (N_2550,N_2517,N_2505);
xor U2551 (N_2551,N_2534,N_2547);
or U2552 (N_2552,N_2524,N_2533);
xnor U2553 (N_2553,N_2541,N_2539);
and U2554 (N_2554,N_2501,N_2523);
nor U2555 (N_2555,N_2500,N_2529);
and U2556 (N_2556,N_2509,N_2521);
nand U2557 (N_2557,N_2525,N_2548);
and U2558 (N_2558,N_2522,N_2519);
nand U2559 (N_2559,N_2544,N_2543);
and U2560 (N_2560,N_2527,N_2512);
nand U2561 (N_2561,N_2542,N_2549);
xor U2562 (N_2562,N_2540,N_2507);
and U2563 (N_2563,N_2506,N_2531);
xor U2564 (N_2564,N_2538,N_2545);
and U2565 (N_2565,N_2514,N_2516);
xnor U2566 (N_2566,N_2530,N_2537);
xor U2567 (N_2567,N_2536,N_2520);
nor U2568 (N_2568,N_2515,N_2504);
or U2569 (N_2569,N_2513,N_2526);
and U2570 (N_2570,N_2503,N_2510);
and U2571 (N_2571,N_2535,N_2511);
and U2572 (N_2572,N_2532,N_2508);
nor U2573 (N_2573,N_2502,N_2518);
nand U2574 (N_2574,N_2528,N_2546);
xor U2575 (N_2575,N_2512,N_2537);
nor U2576 (N_2576,N_2524,N_2529);
and U2577 (N_2577,N_2503,N_2537);
and U2578 (N_2578,N_2522,N_2530);
nand U2579 (N_2579,N_2537,N_2522);
nand U2580 (N_2580,N_2548,N_2537);
or U2581 (N_2581,N_2529,N_2547);
or U2582 (N_2582,N_2536,N_2503);
xor U2583 (N_2583,N_2502,N_2527);
and U2584 (N_2584,N_2500,N_2507);
or U2585 (N_2585,N_2532,N_2534);
or U2586 (N_2586,N_2516,N_2506);
nor U2587 (N_2587,N_2508,N_2523);
nor U2588 (N_2588,N_2530,N_2511);
and U2589 (N_2589,N_2519,N_2526);
nor U2590 (N_2590,N_2540,N_2530);
nor U2591 (N_2591,N_2529,N_2534);
and U2592 (N_2592,N_2512,N_2548);
nor U2593 (N_2593,N_2526,N_2512);
nand U2594 (N_2594,N_2511,N_2506);
or U2595 (N_2595,N_2512,N_2531);
or U2596 (N_2596,N_2544,N_2503);
xor U2597 (N_2597,N_2549,N_2548);
or U2598 (N_2598,N_2518,N_2520);
and U2599 (N_2599,N_2508,N_2504);
and U2600 (N_2600,N_2567,N_2590);
nor U2601 (N_2601,N_2555,N_2566);
xnor U2602 (N_2602,N_2597,N_2574);
or U2603 (N_2603,N_2573,N_2554);
or U2604 (N_2604,N_2579,N_2576);
nor U2605 (N_2605,N_2553,N_2570);
or U2606 (N_2606,N_2588,N_2558);
and U2607 (N_2607,N_2561,N_2552);
nor U2608 (N_2608,N_2565,N_2563);
or U2609 (N_2609,N_2596,N_2583);
nand U2610 (N_2610,N_2556,N_2568);
xnor U2611 (N_2611,N_2562,N_2572);
nor U2612 (N_2612,N_2586,N_2580);
xor U2613 (N_2613,N_2559,N_2564);
xor U2614 (N_2614,N_2581,N_2599);
nand U2615 (N_2615,N_2577,N_2560);
xnor U2616 (N_2616,N_2587,N_2578);
nand U2617 (N_2617,N_2598,N_2594);
xor U2618 (N_2618,N_2569,N_2595);
and U2619 (N_2619,N_2584,N_2551);
nor U2620 (N_2620,N_2557,N_2589);
and U2621 (N_2621,N_2575,N_2593);
nand U2622 (N_2622,N_2571,N_2585);
or U2623 (N_2623,N_2550,N_2582);
and U2624 (N_2624,N_2591,N_2592);
or U2625 (N_2625,N_2589,N_2568);
xnor U2626 (N_2626,N_2586,N_2557);
and U2627 (N_2627,N_2575,N_2551);
and U2628 (N_2628,N_2570,N_2574);
or U2629 (N_2629,N_2586,N_2577);
xnor U2630 (N_2630,N_2561,N_2571);
and U2631 (N_2631,N_2577,N_2597);
xnor U2632 (N_2632,N_2574,N_2584);
xor U2633 (N_2633,N_2595,N_2591);
or U2634 (N_2634,N_2556,N_2558);
and U2635 (N_2635,N_2586,N_2578);
xor U2636 (N_2636,N_2554,N_2553);
nor U2637 (N_2637,N_2596,N_2558);
nor U2638 (N_2638,N_2598,N_2550);
nand U2639 (N_2639,N_2564,N_2560);
or U2640 (N_2640,N_2556,N_2597);
nand U2641 (N_2641,N_2586,N_2596);
xor U2642 (N_2642,N_2591,N_2569);
and U2643 (N_2643,N_2593,N_2595);
nand U2644 (N_2644,N_2562,N_2550);
or U2645 (N_2645,N_2579,N_2555);
and U2646 (N_2646,N_2569,N_2597);
xor U2647 (N_2647,N_2597,N_2552);
nor U2648 (N_2648,N_2588,N_2597);
nand U2649 (N_2649,N_2585,N_2588);
xor U2650 (N_2650,N_2634,N_2608);
nor U2651 (N_2651,N_2635,N_2640);
or U2652 (N_2652,N_2626,N_2631);
nand U2653 (N_2653,N_2643,N_2638);
and U2654 (N_2654,N_2622,N_2611);
and U2655 (N_2655,N_2615,N_2609);
xor U2656 (N_2656,N_2644,N_2646);
nor U2657 (N_2657,N_2618,N_2607);
nor U2658 (N_2658,N_2604,N_2649);
or U2659 (N_2659,N_2645,N_2625);
or U2660 (N_2660,N_2614,N_2616);
and U2661 (N_2661,N_2619,N_2639);
or U2662 (N_2662,N_2610,N_2623);
nor U2663 (N_2663,N_2620,N_2605);
nand U2664 (N_2664,N_2600,N_2637);
or U2665 (N_2665,N_2630,N_2647);
and U2666 (N_2666,N_2624,N_2628);
or U2667 (N_2667,N_2621,N_2633);
nand U2668 (N_2668,N_2629,N_2602);
nand U2669 (N_2669,N_2627,N_2603);
nor U2670 (N_2670,N_2648,N_2601);
nand U2671 (N_2671,N_2606,N_2617);
or U2672 (N_2672,N_2641,N_2632);
and U2673 (N_2673,N_2636,N_2612);
xnor U2674 (N_2674,N_2642,N_2613);
xor U2675 (N_2675,N_2600,N_2602);
xnor U2676 (N_2676,N_2609,N_2604);
xnor U2677 (N_2677,N_2602,N_2621);
xnor U2678 (N_2678,N_2614,N_2639);
and U2679 (N_2679,N_2615,N_2649);
nor U2680 (N_2680,N_2646,N_2643);
and U2681 (N_2681,N_2609,N_2630);
nor U2682 (N_2682,N_2631,N_2630);
and U2683 (N_2683,N_2612,N_2649);
nor U2684 (N_2684,N_2637,N_2645);
xor U2685 (N_2685,N_2629,N_2600);
or U2686 (N_2686,N_2610,N_2611);
and U2687 (N_2687,N_2620,N_2648);
nand U2688 (N_2688,N_2649,N_2645);
nor U2689 (N_2689,N_2620,N_2602);
nor U2690 (N_2690,N_2648,N_2646);
xnor U2691 (N_2691,N_2629,N_2618);
or U2692 (N_2692,N_2645,N_2629);
or U2693 (N_2693,N_2618,N_2616);
xor U2694 (N_2694,N_2639,N_2615);
nand U2695 (N_2695,N_2620,N_2603);
and U2696 (N_2696,N_2603,N_2649);
xnor U2697 (N_2697,N_2635,N_2633);
or U2698 (N_2698,N_2647,N_2643);
and U2699 (N_2699,N_2647,N_2611);
and U2700 (N_2700,N_2658,N_2655);
or U2701 (N_2701,N_2667,N_2663);
and U2702 (N_2702,N_2673,N_2678);
nor U2703 (N_2703,N_2698,N_2659);
and U2704 (N_2704,N_2681,N_2664);
nor U2705 (N_2705,N_2675,N_2690);
or U2706 (N_2706,N_2680,N_2669);
nor U2707 (N_2707,N_2686,N_2666);
xnor U2708 (N_2708,N_2682,N_2679);
nor U2709 (N_2709,N_2657,N_2651);
and U2710 (N_2710,N_2662,N_2670);
xnor U2711 (N_2711,N_2696,N_2665);
xnor U2712 (N_2712,N_2656,N_2683);
and U2713 (N_2713,N_2687,N_2685);
nor U2714 (N_2714,N_2697,N_2660);
nor U2715 (N_2715,N_2674,N_2695);
or U2716 (N_2716,N_2650,N_2677);
and U2717 (N_2717,N_2654,N_2652);
nor U2718 (N_2718,N_2694,N_2692);
and U2719 (N_2719,N_2668,N_2689);
or U2720 (N_2720,N_2661,N_2684);
nor U2721 (N_2721,N_2653,N_2676);
and U2722 (N_2722,N_2672,N_2699);
nand U2723 (N_2723,N_2691,N_2688);
xor U2724 (N_2724,N_2693,N_2671);
xnor U2725 (N_2725,N_2653,N_2690);
xnor U2726 (N_2726,N_2671,N_2659);
nand U2727 (N_2727,N_2685,N_2694);
and U2728 (N_2728,N_2656,N_2662);
or U2729 (N_2729,N_2655,N_2657);
and U2730 (N_2730,N_2671,N_2683);
or U2731 (N_2731,N_2695,N_2687);
nand U2732 (N_2732,N_2676,N_2651);
nor U2733 (N_2733,N_2681,N_2687);
xnor U2734 (N_2734,N_2675,N_2659);
and U2735 (N_2735,N_2666,N_2688);
nor U2736 (N_2736,N_2650,N_2654);
and U2737 (N_2737,N_2652,N_2650);
and U2738 (N_2738,N_2686,N_2664);
nand U2739 (N_2739,N_2670,N_2696);
nor U2740 (N_2740,N_2656,N_2695);
nand U2741 (N_2741,N_2686,N_2672);
nor U2742 (N_2742,N_2672,N_2652);
and U2743 (N_2743,N_2675,N_2660);
nand U2744 (N_2744,N_2672,N_2690);
nor U2745 (N_2745,N_2690,N_2668);
nor U2746 (N_2746,N_2689,N_2662);
xor U2747 (N_2747,N_2655,N_2676);
xor U2748 (N_2748,N_2687,N_2674);
nor U2749 (N_2749,N_2692,N_2696);
and U2750 (N_2750,N_2729,N_2711);
nand U2751 (N_2751,N_2701,N_2703);
or U2752 (N_2752,N_2726,N_2731);
xnor U2753 (N_2753,N_2709,N_2744);
nor U2754 (N_2754,N_2745,N_2721);
nor U2755 (N_2755,N_2738,N_2718);
or U2756 (N_2756,N_2747,N_2713);
nor U2757 (N_2757,N_2715,N_2741);
nand U2758 (N_2758,N_2730,N_2728);
xnor U2759 (N_2759,N_2720,N_2727);
xor U2760 (N_2760,N_2714,N_2725);
or U2761 (N_2761,N_2716,N_2735);
nor U2762 (N_2762,N_2737,N_2740);
nand U2763 (N_2763,N_2707,N_2700);
and U2764 (N_2764,N_2736,N_2708);
or U2765 (N_2765,N_2743,N_2717);
xor U2766 (N_2766,N_2722,N_2719);
or U2767 (N_2767,N_2712,N_2746);
nand U2768 (N_2768,N_2734,N_2710);
and U2769 (N_2769,N_2749,N_2706);
xnor U2770 (N_2770,N_2742,N_2732);
nand U2771 (N_2771,N_2739,N_2748);
nand U2772 (N_2772,N_2724,N_2704);
nor U2773 (N_2773,N_2733,N_2702);
nand U2774 (N_2774,N_2723,N_2705);
and U2775 (N_2775,N_2731,N_2733);
nand U2776 (N_2776,N_2737,N_2712);
nor U2777 (N_2777,N_2702,N_2731);
or U2778 (N_2778,N_2738,N_2747);
or U2779 (N_2779,N_2708,N_2743);
nor U2780 (N_2780,N_2730,N_2703);
xnor U2781 (N_2781,N_2739,N_2719);
or U2782 (N_2782,N_2739,N_2737);
and U2783 (N_2783,N_2722,N_2730);
and U2784 (N_2784,N_2742,N_2725);
xnor U2785 (N_2785,N_2706,N_2713);
nand U2786 (N_2786,N_2717,N_2746);
and U2787 (N_2787,N_2746,N_2704);
xor U2788 (N_2788,N_2718,N_2708);
nand U2789 (N_2789,N_2714,N_2746);
or U2790 (N_2790,N_2735,N_2728);
nor U2791 (N_2791,N_2724,N_2708);
xor U2792 (N_2792,N_2700,N_2740);
xor U2793 (N_2793,N_2710,N_2721);
xor U2794 (N_2794,N_2720,N_2715);
and U2795 (N_2795,N_2724,N_2713);
nand U2796 (N_2796,N_2734,N_2724);
nand U2797 (N_2797,N_2713,N_2701);
nor U2798 (N_2798,N_2734,N_2744);
nor U2799 (N_2799,N_2748,N_2743);
nand U2800 (N_2800,N_2767,N_2789);
xnor U2801 (N_2801,N_2774,N_2754);
and U2802 (N_2802,N_2775,N_2785);
nand U2803 (N_2803,N_2773,N_2757);
xnor U2804 (N_2804,N_2788,N_2759);
nor U2805 (N_2805,N_2758,N_2764);
or U2806 (N_2806,N_2783,N_2790);
or U2807 (N_2807,N_2784,N_2768);
or U2808 (N_2808,N_2752,N_2794);
xor U2809 (N_2809,N_2756,N_2770);
nor U2810 (N_2810,N_2763,N_2753);
or U2811 (N_2811,N_2797,N_2792);
nor U2812 (N_2812,N_2786,N_2782);
and U2813 (N_2813,N_2791,N_2796);
nor U2814 (N_2814,N_2777,N_2781);
or U2815 (N_2815,N_2787,N_2793);
nor U2816 (N_2816,N_2750,N_2798);
nor U2817 (N_2817,N_2799,N_2762);
xor U2818 (N_2818,N_2771,N_2776);
or U2819 (N_2819,N_2795,N_2760);
nor U2820 (N_2820,N_2761,N_2769);
nor U2821 (N_2821,N_2779,N_2765);
nand U2822 (N_2822,N_2780,N_2755);
xor U2823 (N_2823,N_2766,N_2751);
nor U2824 (N_2824,N_2778,N_2772);
and U2825 (N_2825,N_2750,N_2788);
or U2826 (N_2826,N_2786,N_2799);
and U2827 (N_2827,N_2766,N_2790);
xor U2828 (N_2828,N_2783,N_2789);
nor U2829 (N_2829,N_2775,N_2768);
xnor U2830 (N_2830,N_2774,N_2773);
and U2831 (N_2831,N_2763,N_2794);
or U2832 (N_2832,N_2794,N_2790);
and U2833 (N_2833,N_2779,N_2754);
nor U2834 (N_2834,N_2788,N_2790);
or U2835 (N_2835,N_2768,N_2781);
nand U2836 (N_2836,N_2768,N_2776);
nor U2837 (N_2837,N_2756,N_2797);
nand U2838 (N_2838,N_2775,N_2756);
nor U2839 (N_2839,N_2757,N_2755);
nand U2840 (N_2840,N_2750,N_2764);
nor U2841 (N_2841,N_2766,N_2755);
or U2842 (N_2842,N_2769,N_2789);
nor U2843 (N_2843,N_2783,N_2759);
and U2844 (N_2844,N_2773,N_2798);
nor U2845 (N_2845,N_2764,N_2771);
nor U2846 (N_2846,N_2754,N_2791);
or U2847 (N_2847,N_2795,N_2761);
and U2848 (N_2848,N_2766,N_2759);
xnor U2849 (N_2849,N_2769,N_2751);
nand U2850 (N_2850,N_2837,N_2848);
xor U2851 (N_2851,N_2832,N_2815);
or U2852 (N_2852,N_2814,N_2821);
nand U2853 (N_2853,N_2824,N_2820);
xor U2854 (N_2854,N_2841,N_2845);
nand U2855 (N_2855,N_2829,N_2849);
or U2856 (N_2856,N_2805,N_2827);
nor U2857 (N_2857,N_2804,N_2833);
or U2858 (N_2858,N_2818,N_2819);
nand U2859 (N_2859,N_2811,N_2806);
or U2860 (N_2860,N_2840,N_2803);
xor U2861 (N_2861,N_2822,N_2802);
or U2862 (N_2862,N_2843,N_2844);
nand U2863 (N_2863,N_2826,N_2816);
nand U2864 (N_2864,N_2830,N_2836);
nand U2865 (N_2865,N_2808,N_2800);
xnor U2866 (N_2866,N_2823,N_2842);
nand U2867 (N_2867,N_2812,N_2834);
xor U2868 (N_2868,N_2801,N_2817);
nor U2869 (N_2869,N_2825,N_2831);
or U2870 (N_2870,N_2835,N_2810);
nand U2871 (N_2871,N_2828,N_2813);
nand U2872 (N_2872,N_2846,N_2838);
and U2873 (N_2873,N_2809,N_2839);
or U2874 (N_2874,N_2807,N_2847);
xnor U2875 (N_2875,N_2846,N_2844);
xor U2876 (N_2876,N_2821,N_2834);
nor U2877 (N_2877,N_2828,N_2849);
nand U2878 (N_2878,N_2808,N_2814);
xor U2879 (N_2879,N_2813,N_2827);
xnor U2880 (N_2880,N_2834,N_2801);
xnor U2881 (N_2881,N_2814,N_2845);
nand U2882 (N_2882,N_2813,N_2821);
nor U2883 (N_2883,N_2808,N_2806);
nor U2884 (N_2884,N_2825,N_2802);
or U2885 (N_2885,N_2809,N_2811);
nor U2886 (N_2886,N_2819,N_2805);
nor U2887 (N_2887,N_2802,N_2831);
nand U2888 (N_2888,N_2817,N_2816);
nand U2889 (N_2889,N_2844,N_2827);
nor U2890 (N_2890,N_2804,N_2821);
and U2891 (N_2891,N_2803,N_2846);
nor U2892 (N_2892,N_2802,N_2849);
xnor U2893 (N_2893,N_2807,N_2818);
nand U2894 (N_2894,N_2843,N_2818);
and U2895 (N_2895,N_2809,N_2821);
nor U2896 (N_2896,N_2823,N_2810);
nand U2897 (N_2897,N_2816,N_2834);
or U2898 (N_2898,N_2835,N_2825);
nand U2899 (N_2899,N_2807,N_2830);
and U2900 (N_2900,N_2897,N_2850);
nor U2901 (N_2901,N_2871,N_2885);
xnor U2902 (N_2902,N_2886,N_2894);
nor U2903 (N_2903,N_2898,N_2887);
or U2904 (N_2904,N_2870,N_2884);
nand U2905 (N_2905,N_2891,N_2855);
nor U2906 (N_2906,N_2876,N_2878);
nor U2907 (N_2907,N_2888,N_2873);
and U2908 (N_2908,N_2899,N_2893);
or U2909 (N_2909,N_2857,N_2877);
and U2910 (N_2910,N_2856,N_2896);
nor U2911 (N_2911,N_2881,N_2890);
nand U2912 (N_2912,N_2853,N_2862);
or U2913 (N_2913,N_2892,N_2852);
nor U2914 (N_2914,N_2851,N_2863);
nor U2915 (N_2915,N_2860,N_2879);
or U2916 (N_2916,N_2865,N_2889);
nor U2917 (N_2917,N_2859,N_2875);
or U2918 (N_2918,N_2868,N_2864);
or U2919 (N_2919,N_2883,N_2880);
or U2920 (N_2920,N_2869,N_2858);
nand U2921 (N_2921,N_2867,N_2866);
xor U2922 (N_2922,N_2874,N_2872);
and U2923 (N_2923,N_2854,N_2861);
nand U2924 (N_2924,N_2882,N_2895);
or U2925 (N_2925,N_2850,N_2885);
nor U2926 (N_2926,N_2870,N_2876);
nand U2927 (N_2927,N_2867,N_2888);
xor U2928 (N_2928,N_2897,N_2863);
or U2929 (N_2929,N_2870,N_2861);
nand U2930 (N_2930,N_2850,N_2877);
or U2931 (N_2931,N_2880,N_2882);
or U2932 (N_2932,N_2855,N_2889);
or U2933 (N_2933,N_2863,N_2880);
or U2934 (N_2934,N_2889,N_2881);
nand U2935 (N_2935,N_2897,N_2858);
and U2936 (N_2936,N_2857,N_2896);
nor U2937 (N_2937,N_2889,N_2884);
nand U2938 (N_2938,N_2891,N_2866);
nand U2939 (N_2939,N_2877,N_2869);
nor U2940 (N_2940,N_2858,N_2895);
nand U2941 (N_2941,N_2885,N_2865);
or U2942 (N_2942,N_2887,N_2862);
nor U2943 (N_2943,N_2890,N_2898);
nor U2944 (N_2944,N_2893,N_2870);
nand U2945 (N_2945,N_2865,N_2856);
and U2946 (N_2946,N_2887,N_2854);
nor U2947 (N_2947,N_2877,N_2891);
nor U2948 (N_2948,N_2867,N_2871);
or U2949 (N_2949,N_2889,N_2874);
or U2950 (N_2950,N_2933,N_2930);
or U2951 (N_2951,N_2919,N_2939);
xnor U2952 (N_2952,N_2929,N_2945);
nand U2953 (N_2953,N_2902,N_2910);
nand U2954 (N_2954,N_2927,N_2926);
and U2955 (N_2955,N_2936,N_2903);
nor U2956 (N_2956,N_2906,N_2904);
xnor U2957 (N_2957,N_2916,N_2900);
nor U2958 (N_2958,N_2922,N_2920);
nand U2959 (N_2959,N_2944,N_2924);
nor U2960 (N_2960,N_2928,N_2923);
nand U2961 (N_2961,N_2914,N_2940);
nor U2962 (N_2962,N_2948,N_2921);
or U2963 (N_2963,N_2943,N_2905);
or U2964 (N_2964,N_2918,N_2912);
xnor U2965 (N_2965,N_2937,N_2938);
nand U2966 (N_2966,N_2935,N_2925);
and U2967 (N_2967,N_2915,N_2907);
nor U2968 (N_2968,N_2913,N_2931);
nand U2969 (N_2969,N_2917,N_2908);
and U2970 (N_2970,N_2909,N_2947);
nor U2971 (N_2971,N_2901,N_2911);
xor U2972 (N_2972,N_2942,N_2934);
or U2973 (N_2973,N_2932,N_2941);
or U2974 (N_2974,N_2946,N_2949);
nor U2975 (N_2975,N_2944,N_2914);
and U2976 (N_2976,N_2923,N_2913);
nor U2977 (N_2977,N_2936,N_2929);
xor U2978 (N_2978,N_2903,N_2948);
nor U2979 (N_2979,N_2919,N_2921);
xor U2980 (N_2980,N_2905,N_2930);
xor U2981 (N_2981,N_2925,N_2931);
xnor U2982 (N_2982,N_2907,N_2931);
or U2983 (N_2983,N_2902,N_2930);
nand U2984 (N_2984,N_2932,N_2945);
xor U2985 (N_2985,N_2908,N_2909);
nor U2986 (N_2986,N_2914,N_2923);
xnor U2987 (N_2987,N_2919,N_2947);
or U2988 (N_2988,N_2942,N_2929);
nand U2989 (N_2989,N_2936,N_2902);
nand U2990 (N_2990,N_2917,N_2932);
and U2991 (N_2991,N_2921,N_2903);
xnor U2992 (N_2992,N_2916,N_2930);
or U2993 (N_2993,N_2926,N_2943);
and U2994 (N_2994,N_2948,N_2900);
nor U2995 (N_2995,N_2918,N_2929);
xor U2996 (N_2996,N_2918,N_2927);
and U2997 (N_2997,N_2934,N_2921);
xnor U2998 (N_2998,N_2909,N_2910);
or U2999 (N_2999,N_2907,N_2914);
and UO_0 (O_0,N_2998,N_2991);
or UO_1 (O_1,N_2967,N_2955);
xnor UO_2 (O_2,N_2992,N_2950);
nand UO_3 (O_3,N_2989,N_2976);
nor UO_4 (O_4,N_2995,N_2978);
and UO_5 (O_5,N_2990,N_2988);
or UO_6 (O_6,N_2973,N_2979);
xnor UO_7 (O_7,N_2969,N_2974);
nand UO_8 (O_8,N_2985,N_2965);
and UO_9 (O_9,N_2980,N_2957);
nor UO_10 (O_10,N_2962,N_2981);
nor UO_11 (O_11,N_2987,N_2963);
xor UO_12 (O_12,N_2971,N_2954);
or UO_13 (O_13,N_2959,N_2996);
nand UO_14 (O_14,N_2952,N_2951);
nand UO_15 (O_15,N_2999,N_2958);
or UO_16 (O_16,N_2982,N_2986);
nand UO_17 (O_17,N_2972,N_2977);
and UO_18 (O_18,N_2975,N_2984);
nor UO_19 (O_19,N_2993,N_2983);
xor UO_20 (O_20,N_2968,N_2960);
and UO_21 (O_21,N_2994,N_2966);
nor UO_22 (O_22,N_2970,N_2961);
or UO_23 (O_23,N_2964,N_2956);
nand UO_24 (O_24,N_2997,N_2953);
or UO_25 (O_25,N_2984,N_2965);
nor UO_26 (O_26,N_2989,N_2987);
or UO_27 (O_27,N_2975,N_2967);
or UO_28 (O_28,N_2979,N_2989);
and UO_29 (O_29,N_2989,N_2960);
nor UO_30 (O_30,N_2990,N_2985);
nand UO_31 (O_31,N_2955,N_2969);
xnor UO_32 (O_32,N_2995,N_2963);
xor UO_33 (O_33,N_2963,N_2970);
and UO_34 (O_34,N_2973,N_2996);
and UO_35 (O_35,N_2957,N_2993);
or UO_36 (O_36,N_2992,N_2965);
xor UO_37 (O_37,N_2979,N_2963);
nor UO_38 (O_38,N_2955,N_2991);
xnor UO_39 (O_39,N_2992,N_2987);
or UO_40 (O_40,N_2977,N_2967);
and UO_41 (O_41,N_2960,N_2985);
xor UO_42 (O_42,N_2984,N_2992);
and UO_43 (O_43,N_2953,N_2979);
and UO_44 (O_44,N_2979,N_2968);
nor UO_45 (O_45,N_2988,N_2976);
or UO_46 (O_46,N_2996,N_2977);
and UO_47 (O_47,N_2960,N_2996);
and UO_48 (O_48,N_2980,N_2959);
nand UO_49 (O_49,N_2954,N_2956);
nor UO_50 (O_50,N_2979,N_2993);
or UO_51 (O_51,N_2985,N_2977);
nor UO_52 (O_52,N_2976,N_2954);
nor UO_53 (O_53,N_2960,N_2993);
xnor UO_54 (O_54,N_2991,N_2959);
nor UO_55 (O_55,N_2986,N_2981);
or UO_56 (O_56,N_2963,N_2994);
nand UO_57 (O_57,N_2976,N_2994);
nand UO_58 (O_58,N_2962,N_2968);
xor UO_59 (O_59,N_2988,N_2999);
nand UO_60 (O_60,N_2987,N_2964);
nand UO_61 (O_61,N_2987,N_2974);
xor UO_62 (O_62,N_2979,N_2959);
or UO_63 (O_63,N_2970,N_2991);
and UO_64 (O_64,N_2993,N_2964);
xnor UO_65 (O_65,N_2984,N_2958);
nor UO_66 (O_66,N_2959,N_2974);
nor UO_67 (O_67,N_2979,N_2969);
xnor UO_68 (O_68,N_2986,N_2961);
nand UO_69 (O_69,N_2955,N_2950);
nor UO_70 (O_70,N_2975,N_2997);
nor UO_71 (O_71,N_2959,N_2957);
and UO_72 (O_72,N_2960,N_2963);
nand UO_73 (O_73,N_2961,N_2998);
nand UO_74 (O_74,N_2970,N_2972);
nand UO_75 (O_75,N_2950,N_2962);
xnor UO_76 (O_76,N_2990,N_2982);
nand UO_77 (O_77,N_2999,N_2973);
nand UO_78 (O_78,N_2996,N_2980);
and UO_79 (O_79,N_2975,N_2970);
or UO_80 (O_80,N_2969,N_2954);
nand UO_81 (O_81,N_2956,N_2994);
nand UO_82 (O_82,N_2985,N_2992);
nand UO_83 (O_83,N_2978,N_2996);
nor UO_84 (O_84,N_2972,N_2996);
nand UO_85 (O_85,N_2982,N_2985);
nor UO_86 (O_86,N_2992,N_2954);
and UO_87 (O_87,N_2971,N_2980);
nor UO_88 (O_88,N_2966,N_2968);
or UO_89 (O_89,N_2997,N_2986);
xor UO_90 (O_90,N_2993,N_2980);
nor UO_91 (O_91,N_2961,N_2964);
nand UO_92 (O_92,N_2972,N_2965);
and UO_93 (O_93,N_2997,N_2998);
or UO_94 (O_94,N_2982,N_2995);
nor UO_95 (O_95,N_2984,N_2986);
xor UO_96 (O_96,N_2968,N_2982);
nand UO_97 (O_97,N_2991,N_2956);
xnor UO_98 (O_98,N_2988,N_2958);
nand UO_99 (O_99,N_2953,N_2988);
or UO_100 (O_100,N_2954,N_2982);
xor UO_101 (O_101,N_2952,N_2963);
nand UO_102 (O_102,N_2986,N_2991);
and UO_103 (O_103,N_2994,N_2980);
nor UO_104 (O_104,N_2987,N_2976);
xnor UO_105 (O_105,N_2975,N_2999);
xnor UO_106 (O_106,N_2970,N_2986);
nor UO_107 (O_107,N_2999,N_2972);
nand UO_108 (O_108,N_2989,N_2988);
nand UO_109 (O_109,N_2954,N_2968);
nand UO_110 (O_110,N_2980,N_2987);
xnor UO_111 (O_111,N_2971,N_2996);
or UO_112 (O_112,N_2996,N_2988);
xor UO_113 (O_113,N_2959,N_2966);
and UO_114 (O_114,N_2972,N_2959);
and UO_115 (O_115,N_2985,N_2952);
nand UO_116 (O_116,N_2986,N_2957);
and UO_117 (O_117,N_2980,N_2999);
nand UO_118 (O_118,N_2950,N_2953);
and UO_119 (O_119,N_2996,N_2990);
and UO_120 (O_120,N_2981,N_2953);
nand UO_121 (O_121,N_2999,N_2982);
xor UO_122 (O_122,N_2976,N_2952);
or UO_123 (O_123,N_2968,N_2967);
nand UO_124 (O_124,N_2995,N_2985);
nand UO_125 (O_125,N_2971,N_2984);
xor UO_126 (O_126,N_2963,N_2958);
nor UO_127 (O_127,N_2992,N_2976);
nand UO_128 (O_128,N_2991,N_2974);
or UO_129 (O_129,N_2989,N_2982);
xnor UO_130 (O_130,N_2994,N_2955);
nor UO_131 (O_131,N_2992,N_2967);
nor UO_132 (O_132,N_2993,N_2981);
or UO_133 (O_133,N_2987,N_2971);
and UO_134 (O_134,N_2968,N_2992);
xnor UO_135 (O_135,N_2971,N_2976);
or UO_136 (O_136,N_2962,N_2952);
or UO_137 (O_137,N_2971,N_2995);
or UO_138 (O_138,N_2991,N_2979);
and UO_139 (O_139,N_2986,N_2973);
nor UO_140 (O_140,N_2989,N_2998);
nand UO_141 (O_141,N_2971,N_2978);
nor UO_142 (O_142,N_2992,N_2995);
nand UO_143 (O_143,N_2978,N_2998);
xor UO_144 (O_144,N_2967,N_2998);
xor UO_145 (O_145,N_2997,N_2979);
and UO_146 (O_146,N_2967,N_2978);
or UO_147 (O_147,N_2987,N_2986);
and UO_148 (O_148,N_2988,N_2983);
xnor UO_149 (O_149,N_2962,N_2979);
nand UO_150 (O_150,N_2989,N_2954);
xor UO_151 (O_151,N_2970,N_2992);
nor UO_152 (O_152,N_2979,N_2966);
xor UO_153 (O_153,N_2950,N_2973);
nand UO_154 (O_154,N_2980,N_2970);
xnor UO_155 (O_155,N_2963,N_2976);
nor UO_156 (O_156,N_2950,N_2981);
and UO_157 (O_157,N_2960,N_2966);
nand UO_158 (O_158,N_2951,N_2984);
nand UO_159 (O_159,N_2964,N_2967);
xnor UO_160 (O_160,N_2998,N_2952);
nor UO_161 (O_161,N_2964,N_2960);
nor UO_162 (O_162,N_2997,N_2990);
nor UO_163 (O_163,N_2959,N_2986);
and UO_164 (O_164,N_2969,N_2992);
nor UO_165 (O_165,N_2980,N_2978);
nand UO_166 (O_166,N_2961,N_2969);
nor UO_167 (O_167,N_2975,N_2983);
xnor UO_168 (O_168,N_2963,N_2991);
and UO_169 (O_169,N_2990,N_2971);
xnor UO_170 (O_170,N_2966,N_2990);
xor UO_171 (O_171,N_2967,N_2958);
xnor UO_172 (O_172,N_2951,N_2983);
nor UO_173 (O_173,N_2952,N_2977);
nand UO_174 (O_174,N_2972,N_2971);
xnor UO_175 (O_175,N_2965,N_2959);
or UO_176 (O_176,N_2958,N_2952);
or UO_177 (O_177,N_2998,N_2994);
and UO_178 (O_178,N_2974,N_2978);
xnor UO_179 (O_179,N_2962,N_2966);
and UO_180 (O_180,N_2994,N_2996);
xor UO_181 (O_181,N_2957,N_2955);
xnor UO_182 (O_182,N_2991,N_2981);
nand UO_183 (O_183,N_2999,N_2993);
nor UO_184 (O_184,N_2952,N_2972);
nor UO_185 (O_185,N_2980,N_2982);
or UO_186 (O_186,N_2968,N_2957);
and UO_187 (O_187,N_2988,N_2951);
xnor UO_188 (O_188,N_2996,N_2986);
nand UO_189 (O_189,N_2960,N_2994);
and UO_190 (O_190,N_2965,N_2962);
xnor UO_191 (O_191,N_2974,N_2961);
and UO_192 (O_192,N_2970,N_2965);
and UO_193 (O_193,N_2987,N_2977);
nand UO_194 (O_194,N_2976,N_2984);
or UO_195 (O_195,N_2979,N_2998);
nor UO_196 (O_196,N_2960,N_2997);
and UO_197 (O_197,N_2973,N_2984);
xor UO_198 (O_198,N_2957,N_2982);
nor UO_199 (O_199,N_2999,N_2989);
nor UO_200 (O_200,N_2964,N_2983);
nor UO_201 (O_201,N_2958,N_2973);
and UO_202 (O_202,N_2972,N_2961);
nand UO_203 (O_203,N_2980,N_2979);
or UO_204 (O_204,N_2963,N_2973);
xor UO_205 (O_205,N_2960,N_2965);
nand UO_206 (O_206,N_2950,N_2959);
xnor UO_207 (O_207,N_2975,N_2969);
and UO_208 (O_208,N_2972,N_2963);
nand UO_209 (O_209,N_2985,N_2999);
xor UO_210 (O_210,N_2980,N_2984);
and UO_211 (O_211,N_2975,N_2991);
or UO_212 (O_212,N_2980,N_2977);
nor UO_213 (O_213,N_2973,N_2971);
and UO_214 (O_214,N_2992,N_2980);
xnor UO_215 (O_215,N_2992,N_2952);
nor UO_216 (O_216,N_2983,N_2952);
nor UO_217 (O_217,N_2972,N_2960);
nor UO_218 (O_218,N_2970,N_2956);
or UO_219 (O_219,N_2981,N_2961);
nand UO_220 (O_220,N_2964,N_2999);
or UO_221 (O_221,N_2984,N_2966);
and UO_222 (O_222,N_2989,N_2985);
nand UO_223 (O_223,N_2963,N_2982);
nand UO_224 (O_224,N_2957,N_2956);
nand UO_225 (O_225,N_2965,N_2968);
and UO_226 (O_226,N_2957,N_2978);
nand UO_227 (O_227,N_2997,N_2971);
and UO_228 (O_228,N_2952,N_2956);
nor UO_229 (O_229,N_2999,N_2967);
nand UO_230 (O_230,N_2967,N_2957);
xor UO_231 (O_231,N_2994,N_2967);
or UO_232 (O_232,N_2955,N_2998);
or UO_233 (O_233,N_2980,N_2950);
nor UO_234 (O_234,N_2987,N_2982);
nor UO_235 (O_235,N_2957,N_2981);
xnor UO_236 (O_236,N_2998,N_2972);
xor UO_237 (O_237,N_2987,N_2956);
xnor UO_238 (O_238,N_2979,N_2950);
nor UO_239 (O_239,N_2950,N_2976);
xnor UO_240 (O_240,N_2991,N_2964);
and UO_241 (O_241,N_2955,N_2995);
nand UO_242 (O_242,N_2965,N_2971);
nand UO_243 (O_243,N_2990,N_2963);
nand UO_244 (O_244,N_2987,N_2993);
xnor UO_245 (O_245,N_2979,N_2974);
nor UO_246 (O_246,N_2970,N_2993);
nand UO_247 (O_247,N_2991,N_2958);
nor UO_248 (O_248,N_2981,N_2978);
nor UO_249 (O_249,N_2964,N_2963);
xor UO_250 (O_250,N_2960,N_2984);
xnor UO_251 (O_251,N_2973,N_2982);
nor UO_252 (O_252,N_2950,N_2986);
nand UO_253 (O_253,N_2967,N_2976);
and UO_254 (O_254,N_2998,N_2987);
and UO_255 (O_255,N_2969,N_2998);
and UO_256 (O_256,N_2995,N_2972);
nor UO_257 (O_257,N_2991,N_2992);
xor UO_258 (O_258,N_2982,N_2952);
nor UO_259 (O_259,N_2959,N_2989);
nand UO_260 (O_260,N_2990,N_2998);
xor UO_261 (O_261,N_2972,N_2954);
nor UO_262 (O_262,N_2962,N_2987);
xor UO_263 (O_263,N_2994,N_2981);
nand UO_264 (O_264,N_2956,N_2981);
nand UO_265 (O_265,N_2975,N_2988);
nor UO_266 (O_266,N_2980,N_2965);
nor UO_267 (O_267,N_2984,N_2952);
xnor UO_268 (O_268,N_2964,N_2954);
nor UO_269 (O_269,N_2980,N_2966);
or UO_270 (O_270,N_2997,N_2983);
nand UO_271 (O_271,N_2956,N_2986);
or UO_272 (O_272,N_2965,N_2974);
xor UO_273 (O_273,N_2983,N_2979);
and UO_274 (O_274,N_2983,N_2957);
nand UO_275 (O_275,N_2968,N_2958);
nand UO_276 (O_276,N_2965,N_2998);
and UO_277 (O_277,N_2969,N_2965);
nor UO_278 (O_278,N_2994,N_2997);
nor UO_279 (O_279,N_2955,N_2968);
or UO_280 (O_280,N_2997,N_2992);
nand UO_281 (O_281,N_2951,N_2969);
nor UO_282 (O_282,N_2990,N_2967);
xnor UO_283 (O_283,N_2958,N_2962);
nand UO_284 (O_284,N_2961,N_2988);
xnor UO_285 (O_285,N_2995,N_2959);
nor UO_286 (O_286,N_2952,N_2960);
xor UO_287 (O_287,N_2982,N_2975);
and UO_288 (O_288,N_2953,N_2962);
nand UO_289 (O_289,N_2976,N_2956);
and UO_290 (O_290,N_2958,N_2981);
or UO_291 (O_291,N_2967,N_2988);
nor UO_292 (O_292,N_2959,N_2999);
nand UO_293 (O_293,N_2967,N_2970);
or UO_294 (O_294,N_2953,N_2999);
xor UO_295 (O_295,N_2971,N_2975);
nand UO_296 (O_296,N_2958,N_2992);
or UO_297 (O_297,N_2974,N_2993);
xnor UO_298 (O_298,N_2996,N_2995);
and UO_299 (O_299,N_2962,N_2999);
or UO_300 (O_300,N_2960,N_2976);
and UO_301 (O_301,N_2986,N_2980);
or UO_302 (O_302,N_2951,N_2955);
or UO_303 (O_303,N_2951,N_2995);
and UO_304 (O_304,N_2966,N_2998);
or UO_305 (O_305,N_2991,N_2983);
nand UO_306 (O_306,N_2962,N_2956);
and UO_307 (O_307,N_2966,N_2956);
or UO_308 (O_308,N_2974,N_2963);
nor UO_309 (O_309,N_2984,N_2950);
nor UO_310 (O_310,N_2971,N_2993);
or UO_311 (O_311,N_2983,N_2969);
xor UO_312 (O_312,N_2964,N_2992);
nand UO_313 (O_313,N_2993,N_2973);
nand UO_314 (O_314,N_2994,N_2984);
and UO_315 (O_315,N_2997,N_2958);
and UO_316 (O_316,N_2962,N_2972);
nor UO_317 (O_317,N_2978,N_2972);
or UO_318 (O_318,N_2974,N_2954);
xnor UO_319 (O_319,N_2966,N_2995);
nor UO_320 (O_320,N_2967,N_2972);
and UO_321 (O_321,N_2973,N_2988);
xor UO_322 (O_322,N_2991,N_2951);
nor UO_323 (O_323,N_2989,N_2991);
nor UO_324 (O_324,N_2995,N_2952);
xor UO_325 (O_325,N_2987,N_2996);
nor UO_326 (O_326,N_2981,N_2983);
or UO_327 (O_327,N_2965,N_2978);
and UO_328 (O_328,N_2977,N_2956);
or UO_329 (O_329,N_2985,N_2961);
nand UO_330 (O_330,N_2984,N_2967);
nor UO_331 (O_331,N_2998,N_2975);
and UO_332 (O_332,N_2956,N_2995);
nor UO_333 (O_333,N_2959,N_2975);
or UO_334 (O_334,N_2988,N_2993);
nand UO_335 (O_335,N_2989,N_2972);
nand UO_336 (O_336,N_2976,N_2961);
nor UO_337 (O_337,N_2958,N_2980);
and UO_338 (O_338,N_2975,N_2966);
xor UO_339 (O_339,N_2990,N_2968);
nand UO_340 (O_340,N_2980,N_2960);
xnor UO_341 (O_341,N_2978,N_2993);
nand UO_342 (O_342,N_2959,N_2990);
nor UO_343 (O_343,N_2953,N_2958);
nand UO_344 (O_344,N_2976,N_2990);
or UO_345 (O_345,N_2982,N_2967);
xor UO_346 (O_346,N_2972,N_2950);
xnor UO_347 (O_347,N_2989,N_2975);
and UO_348 (O_348,N_2965,N_2999);
nand UO_349 (O_349,N_2958,N_2961);
xnor UO_350 (O_350,N_2971,N_2992);
nor UO_351 (O_351,N_2971,N_2967);
nor UO_352 (O_352,N_2990,N_2954);
and UO_353 (O_353,N_2974,N_2967);
nand UO_354 (O_354,N_2988,N_2950);
and UO_355 (O_355,N_2992,N_2957);
xor UO_356 (O_356,N_2999,N_2961);
nor UO_357 (O_357,N_2982,N_2961);
nand UO_358 (O_358,N_2977,N_2984);
xor UO_359 (O_359,N_2967,N_2960);
nor UO_360 (O_360,N_2956,N_2996);
and UO_361 (O_361,N_2990,N_2983);
nand UO_362 (O_362,N_2998,N_2959);
and UO_363 (O_363,N_2994,N_2962);
nor UO_364 (O_364,N_2952,N_2961);
nor UO_365 (O_365,N_2972,N_2973);
xnor UO_366 (O_366,N_2952,N_2954);
and UO_367 (O_367,N_2997,N_2965);
and UO_368 (O_368,N_2970,N_2976);
xnor UO_369 (O_369,N_2961,N_2955);
or UO_370 (O_370,N_2997,N_2968);
or UO_371 (O_371,N_2957,N_2985);
nand UO_372 (O_372,N_2965,N_2986);
xor UO_373 (O_373,N_2996,N_2992);
or UO_374 (O_374,N_2994,N_2979);
and UO_375 (O_375,N_2990,N_2970);
nand UO_376 (O_376,N_2960,N_2981);
and UO_377 (O_377,N_2975,N_2994);
and UO_378 (O_378,N_2951,N_2998);
xnor UO_379 (O_379,N_2978,N_2961);
or UO_380 (O_380,N_2975,N_2976);
nand UO_381 (O_381,N_2961,N_2962);
nor UO_382 (O_382,N_2983,N_2950);
xor UO_383 (O_383,N_2991,N_2995);
and UO_384 (O_384,N_2987,N_2991);
nand UO_385 (O_385,N_2970,N_2988);
xnor UO_386 (O_386,N_2971,N_2989);
nor UO_387 (O_387,N_2976,N_2978);
xnor UO_388 (O_388,N_2981,N_2996);
and UO_389 (O_389,N_2957,N_2958);
nand UO_390 (O_390,N_2982,N_2988);
and UO_391 (O_391,N_2962,N_2977);
nor UO_392 (O_392,N_2977,N_2958);
nor UO_393 (O_393,N_2976,N_2991);
nand UO_394 (O_394,N_2982,N_2981);
nor UO_395 (O_395,N_2985,N_2980);
xnor UO_396 (O_396,N_2963,N_2968);
nor UO_397 (O_397,N_2976,N_2999);
nor UO_398 (O_398,N_2957,N_2951);
and UO_399 (O_399,N_2970,N_2983);
nand UO_400 (O_400,N_2954,N_2979);
nor UO_401 (O_401,N_2992,N_2956);
xnor UO_402 (O_402,N_2965,N_2973);
nor UO_403 (O_403,N_2970,N_2999);
nor UO_404 (O_404,N_2951,N_2954);
nor UO_405 (O_405,N_2982,N_2997);
or UO_406 (O_406,N_2966,N_2996);
nor UO_407 (O_407,N_2973,N_2992);
nand UO_408 (O_408,N_2991,N_2962);
nor UO_409 (O_409,N_2977,N_2981);
nor UO_410 (O_410,N_2980,N_2956);
nor UO_411 (O_411,N_2987,N_2957);
nand UO_412 (O_412,N_2971,N_2999);
and UO_413 (O_413,N_2950,N_2954);
and UO_414 (O_414,N_2955,N_2999);
and UO_415 (O_415,N_2984,N_2996);
xor UO_416 (O_416,N_2977,N_2965);
xnor UO_417 (O_417,N_2962,N_2955);
or UO_418 (O_418,N_2952,N_2965);
nand UO_419 (O_419,N_2987,N_2966);
or UO_420 (O_420,N_2986,N_2953);
or UO_421 (O_421,N_2989,N_2953);
and UO_422 (O_422,N_2967,N_2963);
xnor UO_423 (O_423,N_2986,N_2969);
or UO_424 (O_424,N_2964,N_2997);
nand UO_425 (O_425,N_2963,N_2998);
and UO_426 (O_426,N_2969,N_2976);
and UO_427 (O_427,N_2961,N_2997);
nand UO_428 (O_428,N_2979,N_2967);
and UO_429 (O_429,N_2990,N_2979);
xnor UO_430 (O_430,N_2959,N_2994);
or UO_431 (O_431,N_2989,N_2963);
or UO_432 (O_432,N_2960,N_2973);
nor UO_433 (O_433,N_2952,N_2973);
nor UO_434 (O_434,N_2952,N_2966);
xnor UO_435 (O_435,N_2993,N_2976);
or UO_436 (O_436,N_2981,N_2976);
nor UO_437 (O_437,N_2972,N_2985);
or UO_438 (O_438,N_2950,N_2982);
nand UO_439 (O_439,N_2963,N_2962);
nor UO_440 (O_440,N_2993,N_2992);
nand UO_441 (O_441,N_2969,N_2967);
nand UO_442 (O_442,N_2950,N_2977);
and UO_443 (O_443,N_2975,N_2955);
and UO_444 (O_444,N_2973,N_2964);
or UO_445 (O_445,N_2997,N_2972);
nand UO_446 (O_446,N_2968,N_2973);
xnor UO_447 (O_447,N_2958,N_2959);
nor UO_448 (O_448,N_2961,N_2989);
xor UO_449 (O_449,N_2989,N_2993);
nor UO_450 (O_450,N_2982,N_2953);
xor UO_451 (O_451,N_2954,N_2981);
and UO_452 (O_452,N_2965,N_2966);
nand UO_453 (O_453,N_2969,N_2988);
nor UO_454 (O_454,N_2971,N_2953);
nand UO_455 (O_455,N_2990,N_2987);
nand UO_456 (O_456,N_2973,N_2994);
and UO_457 (O_457,N_2988,N_2974);
and UO_458 (O_458,N_2964,N_2952);
nand UO_459 (O_459,N_2964,N_2986);
nand UO_460 (O_460,N_2960,N_2958);
nor UO_461 (O_461,N_2970,N_2955);
and UO_462 (O_462,N_2992,N_2951);
nor UO_463 (O_463,N_2993,N_2950);
nand UO_464 (O_464,N_2986,N_2992);
or UO_465 (O_465,N_2990,N_2975);
nor UO_466 (O_466,N_2993,N_2956);
nor UO_467 (O_467,N_2952,N_2957);
nor UO_468 (O_468,N_2987,N_2952);
nand UO_469 (O_469,N_2979,N_2982);
nor UO_470 (O_470,N_2978,N_2988);
nand UO_471 (O_471,N_2977,N_2999);
nand UO_472 (O_472,N_2969,N_2995);
or UO_473 (O_473,N_2963,N_2985);
xnor UO_474 (O_474,N_2959,N_2982);
and UO_475 (O_475,N_2952,N_2980);
xnor UO_476 (O_476,N_2997,N_2951);
or UO_477 (O_477,N_2965,N_2979);
and UO_478 (O_478,N_2982,N_2966);
xnor UO_479 (O_479,N_2983,N_2995);
xor UO_480 (O_480,N_2958,N_2971);
nand UO_481 (O_481,N_2956,N_2972);
or UO_482 (O_482,N_2952,N_2974);
xnor UO_483 (O_483,N_2971,N_2981);
and UO_484 (O_484,N_2968,N_2969);
nor UO_485 (O_485,N_2956,N_2965);
nor UO_486 (O_486,N_2983,N_2956);
nand UO_487 (O_487,N_2978,N_2958);
xnor UO_488 (O_488,N_2991,N_2982);
xor UO_489 (O_489,N_2975,N_2961);
nand UO_490 (O_490,N_2954,N_2965);
or UO_491 (O_491,N_2982,N_2996);
nor UO_492 (O_492,N_2971,N_2988);
nor UO_493 (O_493,N_2964,N_2958);
nor UO_494 (O_494,N_2965,N_2963);
and UO_495 (O_495,N_2986,N_2988);
xor UO_496 (O_496,N_2985,N_2993);
and UO_497 (O_497,N_2996,N_2957);
or UO_498 (O_498,N_2953,N_2976);
and UO_499 (O_499,N_2955,N_2981);
endmodule